// Benchmark "voter" written by ABC on Mon Sep 11 23:36:32 2023

module voter ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] ,
    \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] ,
    \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] ,
    \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
    \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
    \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] ,
    \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] ,
    \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] ,
    \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] ,
    \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
    \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
    \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] ,
    \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] ,
    \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] ,
    \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] ,
    \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
    \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
    \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] ,
    \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] ,
    \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] ,
    \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] ,
    \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
    \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
    \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] ,
    \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] ,
    \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] ,
    \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] ,
    \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
    \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
    \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] ,
    \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] ,
    \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] ,
    \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] ,
    \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
    \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
    \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] ,
    \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] ,
    \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] ,
    \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] ,
    \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
    \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
    \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] ,
    \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] ,
    \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] ,
    \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] ,
    \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
    \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
    \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] ,
    \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] ,
    \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] ,
    \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] ,
    \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
    \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
    \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] ,
    \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] ,
    \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] ,
    \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] ,
    \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
    \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
    \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] ,
    \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] ,
    \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] ,
    \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] ,
    \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
    \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
    \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] ,
    \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] ,
    \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] ,
    \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] ,
    \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
    \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
    \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] ,
    \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] ,
    \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] ,
    \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] ,
    \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
    \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
    \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] ,
    \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] ,
    \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] ,
    \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] ,
    \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
    \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
    \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] ,
    \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] ,
    \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] ,
    \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] ,
    \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
    \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
    \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] ,
    \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] ,
    \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] ,
    \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] ,
    \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
    \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
    \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] ,
    \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] ,
    \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] ,
    \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] ,
    \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
    \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
    \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] ,
    \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] ,
    \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] ,
    \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] ,
    \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
    \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
    \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] ,
    \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] ,
    \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] ,
    \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] ,
    \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
    \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
    \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] ,
    \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] ,
    \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] ,
    \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] ,
    \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
    \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
    \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] ,
    \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] ,
    \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] ,
    \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] ,
    \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
    \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
    \A[1000] ,
    maj  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] ,
    \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] ,
    \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] ,
    \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] ,
    \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
    \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
    \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] ,
    \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] ,
    \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] ,
    \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] ,
    \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
    \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
    \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] ,
    \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] ,
    \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] ,
    \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] ,
    \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
    \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
    \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] ,
    \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] ,
    \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] ,
    \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] ,
    \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
    \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
    \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] ,
    \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] ,
    \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] ,
    \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] ,
    \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
    \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
    \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] ,
    \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] ,
    \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] ,
    \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] ,
    \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
    \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
    \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] ,
    \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] ,
    \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] ,
    \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] ,
    \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
    \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
    \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] ,
    \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] ,
    \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] ,
    \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] ,
    \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
    \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
    \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] ,
    \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] ,
    \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] ,
    \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] ,
    \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
    \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
    \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] ,
    \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] ,
    \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] ,
    \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] ,
    \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
    \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
    \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] ,
    \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] ,
    \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] ,
    \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] ,
    \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
    \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
    \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] ,
    \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] ,
    \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] ,
    \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] ,
    \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
    \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
    \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] ,
    \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] ,
    \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] ,
    \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] ,
    \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
    \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
    \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] ,
    \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] ,
    \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] ,
    \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] ,
    \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
    \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
    \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] ,
    \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] ,
    \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] ,
    \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] ,
    \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
    \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
    \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] ,
    \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] ,
    \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] ,
    \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] ,
    \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
    \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
    \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] ,
    \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] ,
    \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] ,
    \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] ,
    \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
    \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
    \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] ,
    \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] ,
    \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] ,
    \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] ,
    \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
    \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
    \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] ,
    \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] ,
    \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] ,
    \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] ,
    \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
    \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
    \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] ,
    \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] ,
    \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] ,
    \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] ,
    \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
    \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
    \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] ,
    \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] ,
    \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] ,
    \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] ,
    \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
    \A[999] , \A[1000] ;
  output maj;
  wire new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_,
    new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_,
    new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_,
    new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_,
    new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_,
    new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_,
    new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_,
    new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_,
    new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_,
    new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_,
    new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_,
    new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_,
    new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_,
    new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_,
    new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_,
    new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_,
    new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_,
    new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_,
    new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_,
    new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_,
    new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_,
    new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_,
    new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_,
    new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_,
    new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_,
    new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_,
    new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_,
    new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_,
    new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_,
    new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_,
    new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_,
    new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_,
    new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_,
    new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_,
    new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_,
    new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_,
    new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_,
    new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_,
    new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_,
    new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_,
    new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_,
    new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_,
    new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_,
    new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_,
    new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_,
    new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_,
    new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_,
    new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_,
    new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_,
    new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_,
    new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_,
    new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_,
    new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_,
    new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_,
    new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_,
    new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_,
    new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_,
    new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_,
    new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_,
    new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_,
    new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_,
    new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_,
    new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_,
    new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_,
    new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_,
    new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_,
    new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_,
    new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_,
    new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_,
    new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_,
    new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_,
    new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_,
    new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_,
    new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_,
    new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_,
    new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_,
    new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_,
    new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_,
    new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_,
    new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_,
    new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_,
    new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_,
    new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_,
    new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_,
    new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_,
    new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_,
    new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_,
    new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_,
    new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_,
    new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_,
    new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_,
    new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_,
    new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_,
    new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_,
    new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_,
    new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_,
    new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_,
    new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_,
    new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_,
    new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_,
    new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_,
    new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_,
    new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_,
    new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_,
    new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_,
    new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_,
    new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_,
    new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_,
    new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_,
    new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_,
    new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_,
    new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_,
    new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_,
    new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_,
    new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_,
    new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_,
    new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_,
    new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_,
    new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_,
    new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_,
    new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_,
    new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_,
    new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_,
    new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_,
    new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_,
    new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_,
    new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_,
    new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_,
    new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_,
    new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_,
    new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_,
    new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_,
    new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_,
    new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_,
    new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_,
    new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_,
    new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_,
    new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_,
    new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_,
    new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_,
    new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_,
    new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_,
    new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_,
    new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_,
    new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_,
    new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_,
    new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_,
    new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_,
    new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_,
    new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_,
    new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_,
    new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_,
    new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_,
    new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_,
    new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_,
    new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_,
    new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_,
    new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_,
    new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_,
    new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_,
    new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_,
    new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_,
    new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_,
    new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_,
    new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_,
    new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_,
    new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_,
    new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_,
    new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_,
    new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_,
    new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_,
    new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_,
    new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_,
    new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_,
    new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_,
    new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_,
    new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_,
    new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_,
    new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_,
    new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_,
    new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_,
    new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_,
    new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_,
    new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_,
    new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_,
    new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_,
    new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_,
    new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_,
    new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_,
    new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_,
    new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_,
    new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_,
    new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_,
    new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_,
    new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_,
    new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_,
    new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_,
    new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_,
    new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_,
    new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_,
    new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12147_, new_n12148_, new_n12149_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12333_, new_n12334_, new_n12335_,
    new_n12336_, new_n12337_, new_n12338_, new_n12339_, new_n12340_,
    new_n12341_, new_n12342_, new_n12343_, new_n12344_, new_n12345_,
    new_n12346_, new_n12347_, new_n12348_, new_n12349_, new_n12350_,
    new_n12351_, new_n12352_, new_n12353_, new_n12354_, new_n12355_,
    new_n12356_, new_n12357_, new_n12358_, new_n12359_, new_n12360_,
    new_n12361_, new_n12362_, new_n12363_, new_n12364_, new_n12365_,
    new_n12366_, new_n12367_, new_n12368_, new_n12369_, new_n12370_,
    new_n12371_, new_n12372_, new_n12373_, new_n12374_, new_n12375_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12384_, new_n12385_,
    new_n12386_, new_n12387_, new_n12388_, new_n12389_, new_n12390_,
    new_n12391_, new_n12392_, new_n12393_, new_n12394_, new_n12395_,
    new_n12396_, new_n12397_, new_n12398_, new_n12399_, new_n12400_,
    new_n12401_, new_n12402_, new_n12403_, new_n12404_, new_n12405_,
    new_n12406_, new_n12407_, new_n12408_, new_n12409_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12420_,
    new_n12421_, new_n12422_, new_n12423_, new_n12424_, new_n12425_,
    new_n12426_, new_n12427_, new_n12428_, new_n12429_, new_n12430_,
    new_n12431_, new_n12432_, new_n12433_, new_n12434_, new_n12435_,
    new_n12436_, new_n12437_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14075_,
    new_n14076_, new_n14077_, new_n14078_, new_n14079_, new_n14080_,
    new_n14081_, new_n14082_, new_n14083_, new_n14084_, new_n14085_,
    new_n14086_, new_n14087_, new_n14088_, new_n14089_, new_n14090_,
    new_n14091_, new_n14092_, new_n14093_, new_n14094_, new_n14095_,
    new_n14096_, new_n14097_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14103_, new_n14104_, new_n14105_,
    new_n14106_, new_n14107_, new_n14108_, new_n14109_, new_n14110_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14117_, new_n14118_, new_n14119_, new_n14120_,
    new_n14121_, new_n14122_, new_n14123_, new_n14124_, new_n14125_,
    new_n14126_, new_n14127_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14133_, new_n14134_, new_n14135_,
    new_n14136_, new_n14137_, new_n14138_, new_n14139_, new_n14140_,
    new_n14141_, new_n14142_, new_n14143_, new_n14144_, new_n14145_,
    new_n14146_, new_n14147_, new_n14148_, new_n14149_, new_n14150_,
    new_n14151_, new_n14152_, new_n14153_, new_n14154_, new_n14155_,
    new_n14156_, new_n14157_, new_n14158_, new_n14159_, new_n14160_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14205_,
    new_n14206_, new_n14207_, new_n14208_, new_n14209_, new_n14210_,
    new_n14211_, new_n14212_, new_n14213_, new_n14214_, new_n14215_,
    new_n14216_, new_n14217_, new_n14218_, new_n14219_, new_n14220_,
    new_n14221_, new_n14222_, new_n14223_, new_n14224_, new_n14225_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14241_, new_n14242_, new_n14243_, new_n14244_, new_n14245_,
    new_n14246_, new_n14247_, new_n14248_, new_n14249_, new_n14250_,
    new_n14251_, new_n14252_, new_n14253_, new_n14254_, new_n14255_,
    new_n14256_, new_n14257_, new_n14258_, new_n14259_, new_n14260_,
    new_n14261_, new_n14262_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14268_, new_n14269_, new_n14270_,
    new_n14271_, new_n14272_, new_n14273_, new_n14274_, new_n14275_,
    new_n14276_, new_n14277_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14284_, new_n14285_,
    new_n14286_, new_n14287_, new_n14288_, new_n14289_, new_n14290_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14342_, new_n14343_, new_n14344_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14416_, new_n14417_, new_n14418_, new_n14419_, new_n14420_,
    new_n14421_, new_n14422_, new_n14423_, new_n14424_, new_n14425_,
    new_n14426_, new_n14427_, new_n14428_, new_n14429_, new_n14430_,
    new_n14431_, new_n14432_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14465_,
    new_n14466_, new_n14467_, new_n14468_, new_n14469_, new_n14470_,
    new_n14471_, new_n14472_, new_n14473_, new_n14474_, new_n14475_,
    new_n14476_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14481_, new_n14482_, new_n14483_, new_n14484_, new_n14485_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14595_,
    new_n14596_, new_n14597_, new_n14598_, new_n14599_, new_n14600_,
    new_n14601_, new_n14602_, new_n14603_, new_n14604_, new_n14605_,
    new_n14606_, new_n14607_, new_n14608_, new_n14609_, new_n14610_,
    new_n14611_, new_n14612_, new_n14613_, new_n14614_, new_n14615_,
    new_n14616_, new_n14617_, new_n14618_, new_n14619_, new_n14620_,
    new_n14621_, new_n14622_, new_n14623_, new_n14624_, new_n14625_,
    new_n14626_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14840_,
    new_n14841_, new_n14842_, new_n14843_, new_n14844_, new_n14845_,
    new_n14846_, new_n14847_, new_n14848_, new_n14849_, new_n14850_,
    new_n14851_, new_n14852_, new_n14853_, new_n14854_, new_n14855_,
    new_n14856_, new_n14857_, new_n14858_, new_n14859_, new_n14860_,
    new_n14861_, new_n14862_, new_n14863_, new_n14864_, new_n14865_,
    new_n14866_, new_n14867_, new_n14868_, new_n14869_, new_n14870_,
    new_n14871_, new_n14872_, new_n14873_, new_n14874_, new_n14875_,
    new_n14876_, new_n14877_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14887_, new_n14888_, new_n14889_, new_n14890_,
    new_n14891_, new_n14892_, new_n14893_, new_n14894_, new_n14895_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14902_, new_n14903_, new_n14904_, new_n14905_,
    new_n14906_, new_n14907_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15328_, new_n15329_, new_n15330_,
    new_n15331_, new_n15332_, new_n15333_, new_n15334_, new_n15335_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15381_, new_n15382_, new_n15383_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15390_,
    new_n15391_, new_n15392_, new_n15393_, new_n15394_, new_n15395_,
    new_n15396_, new_n15397_, new_n15398_, new_n15399_, new_n15400_,
    new_n15401_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15438_, new_n15439_, new_n15440_,
    new_n15441_, new_n15442_, new_n15443_, new_n15444_, new_n15445_,
    new_n15446_, new_n15447_, new_n15448_, new_n15449_, new_n15450_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15494_, new_n15495_,
    new_n15496_, new_n15497_, new_n15498_, new_n15499_, new_n15500_,
    new_n15501_, new_n15502_, new_n15503_, new_n15504_, new_n15505_,
    new_n15506_, new_n15507_, new_n15508_, new_n15509_, new_n15510_,
    new_n15511_, new_n15512_, new_n15513_, new_n15514_, new_n15515_,
    new_n15516_, new_n15517_, new_n15518_, new_n15519_, new_n15520_,
    new_n15521_, new_n15522_, new_n15523_, new_n15524_, new_n15525_,
    new_n15526_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15531_, new_n15532_, new_n15533_, new_n15534_, new_n15535_,
    new_n15536_, new_n15537_, new_n15538_, new_n15539_, new_n15540_,
    new_n15541_, new_n15542_, new_n15543_, new_n15544_, new_n15545_,
    new_n15546_, new_n15547_, new_n15548_, new_n15549_, new_n15550_,
    new_n15551_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16349_, new_n16350_,
    new_n16351_, new_n16352_, new_n16353_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16361_, new_n16362_, new_n16363_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16489_, new_n16490_,
    new_n16491_, new_n16492_, new_n16493_, new_n16494_, new_n16495_,
    new_n16496_, new_n16497_, new_n16498_, new_n16499_, new_n16500_,
    new_n16501_, new_n16502_, new_n16503_, new_n16504_, new_n16505_,
    new_n16506_, new_n16507_, new_n16508_, new_n16509_, new_n16510_,
    new_n16511_, new_n16512_, new_n16513_, new_n16514_, new_n16515_,
    new_n16516_, new_n16517_, new_n16518_, new_n16519_, new_n16520_,
    new_n16521_, new_n16522_, new_n16523_, new_n16524_, new_n16525_,
    new_n16526_, new_n16527_, new_n16528_, new_n16529_, new_n16530_,
    new_n16531_, new_n16532_, new_n16533_, new_n16534_, new_n16535_,
    new_n16536_, new_n16537_, new_n16538_, new_n16539_, new_n16540_,
    new_n16541_, new_n16542_, new_n16543_, new_n16544_, new_n16545_,
    new_n16546_, new_n16547_, new_n16548_, new_n16549_, new_n16550_,
    new_n16551_, new_n16552_, new_n16553_, new_n16554_, new_n16555_,
    new_n16556_, new_n16557_, new_n16558_, new_n16559_, new_n16560_,
    new_n16561_, new_n16562_, new_n16563_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16618_, new_n16619_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16659_, new_n16660_,
    new_n16661_, new_n16662_, new_n16663_, new_n16664_, new_n16665_,
    new_n16666_, new_n16667_, new_n16668_, new_n16669_, new_n16670_,
    new_n16671_, new_n16672_, new_n16673_, new_n16674_, new_n16675_,
    new_n16676_, new_n16677_, new_n16678_, new_n16679_, new_n16680_,
    new_n16681_, new_n16682_, new_n16683_, new_n16684_, new_n16685_,
    new_n16686_, new_n16687_, new_n16688_, new_n16689_, new_n16690_,
    new_n16691_, new_n16692_, new_n16693_, new_n16694_, new_n16695_,
    new_n16696_, new_n16697_, new_n16698_, new_n16699_, new_n16700_,
    new_n16701_, new_n16702_, new_n16703_, new_n16704_, new_n16705_,
    new_n16706_, new_n16707_, new_n16708_, new_n16709_, new_n16710_,
    new_n16711_, new_n16712_, new_n16713_, new_n16714_, new_n16715_,
    new_n16716_, new_n16717_, new_n16718_, new_n16719_, new_n16720_,
    new_n16721_, new_n16722_, new_n16723_, new_n16724_, new_n16725_,
    new_n16726_, new_n16727_, new_n16728_, new_n16729_, new_n16730_,
    new_n16731_, new_n16732_, new_n16733_, new_n16734_, new_n16735_,
    new_n16736_, new_n16737_, new_n16738_, new_n16739_, new_n16740_,
    new_n16741_, new_n16742_, new_n16743_, new_n16744_, new_n16745_,
    new_n16746_, new_n16747_, new_n16748_, new_n16749_, new_n16750_,
    new_n16751_, new_n16752_, new_n16753_, new_n16754_, new_n16755_,
    new_n16756_, new_n16757_, new_n16758_, new_n16759_, new_n16760_,
    new_n16761_, new_n16762_, new_n16763_, new_n16764_, new_n16765_,
    new_n16766_, new_n16767_, new_n16768_, new_n16769_, new_n16770_,
    new_n16771_, new_n16772_, new_n16773_, new_n16774_, new_n16775_,
    new_n16776_, new_n16777_, new_n16778_, new_n16779_, new_n16780_,
    new_n16781_, new_n16782_, new_n16783_, new_n16784_, new_n16785_,
    new_n16786_, new_n16787_, new_n16788_, new_n16789_, new_n16790_,
    new_n16791_, new_n16792_, new_n16793_, new_n16794_, new_n16795_,
    new_n16796_, new_n16797_, new_n16798_, new_n16799_, new_n16800_,
    new_n16801_, new_n16802_, new_n16803_, new_n16804_, new_n16805_,
    new_n16806_, new_n16807_, new_n16808_, new_n16809_, new_n16810_,
    new_n16811_, new_n16812_, new_n16813_, new_n16814_, new_n16815_,
    new_n16816_, new_n16817_, new_n16818_, new_n16819_, new_n16820_,
    new_n16821_, new_n16822_, new_n16823_, new_n16824_, new_n16825_,
    new_n16826_, new_n16827_, new_n16828_, new_n16829_, new_n16830_,
    new_n16831_, new_n16832_, new_n16833_, new_n16834_, new_n16835_,
    new_n16836_, new_n16837_, new_n16838_, new_n16839_, new_n16840_,
    new_n16841_, new_n16842_, new_n16843_, new_n16844_, new_n16845_,
    new_n16846_, new_n16847_, new_n16848_, new_n16849_, new_n16850_,
    new_n16851_, new_n16852_, new_n16853_, new_n16854_, new_n16855_,
    new_n16856_, new_n16857_, new_n16858_, new_n16859_, new_n16860_,
    new_n16861_, new_n16862_, new_n16863_, new_n16864_, new_n16865_,
    new_n16866_, new_n16867_, new_n16868_, new_n16869_, new_n16870_,
    new_n16871_, new_n16872_, new_n16873_, new_n16874_, new_n16875_,
    new_n16876_, new_n16877_, new_n16878_, new_n16879_, new_n16880_,
    new_n16881_, new_n16882_, new_n16883_, new_n16884_, new_n16885_,
    new_n16886_, new_n16887_, new_n16888_, new_n16889_, new_n16890_,
    new_n16891_, new_n16892_, new_n16893_, new_n16894_, new_n16895_,
    new_n16896_, new_n16897_, new_n16898_, new_n16899_, new_n16900_,
    new_n16901_, new_n16902_, new_n16903_, new_n16904_, new_n16905_,
    new_n16906_, new_n16907_, new_n16908_, new_n16909_, new_n16910_,
    new_n16911_, new_n16912_, new_n16913_, new_n16914_, new_n16915_,
    new_n16916_, new_n16917_, new_n16918_, new_n16919_, new_n16920_,
    new_n16921_, new_n16922_, new_n16923_, new_n16924_, new_n16925_,
    new_n16926_, new_n16927_, new_n16928_, new_n16929_, new_n16930_,
    new_n16931_, new_n16932_, new_n16933_, new_n16934_, new_n16935_,
    new_n16936_, new_n16937_, new_n16938_, new_n16939_, new_n16940_,
    new_n16941_, new_n16942_, new_n16943_, new_n16944_, new_n16945_,
    new_n16946_, new_n16947_, new_n16948_, new_n16949_, new_n16950_,
    new_n16951_, new_n16952_, new_n16953_, new_n16954_, new_n16955_,
    new_n16956_, new_n16957_, new_n16958_, new_n16959_, new_n16960_,
    new_n16961_, new_n16962_, new_n16963_, new_n16964_, new_n16965_,
    new_n16966_, new_n16967_, new_n16968_, new_n16969_, new_n16970_,
    new_n16971_, new_n16972_, new_n16973_, new_n16974_, new_n16975_,
    new_n16976_, new_n16977_, new_n16978_, new_n16979_, new_n16980_,
    new_n16981_, new_n16982_, new_n16983_, new_n16984_, new_n16985_,
    new_n16986_, new_n16987_, new_n16988_, new_n16989_, new_n16990_,
    new_n16991_, new_n16992_, new_n16993_, new_n16994_, new_n16995_,
    new_n16996_, new_n16997_, new_n16998_, new_n16999_, new_n17000_,
    new_n17001_, new_n17002_, new_n17003_, new_n17004_, new_n17005_,
    new_n17006_, new_n17007_, new_n17008_, new_n17009_, new_n17010_,
    new_n17011_, new_n17012_, new_n17013_, new_n17014_, new_n17015_,
    new_n17016_, new_n17017_, new_n17018_, new_n17019_, new_n17020_,
    new_n17021_, new_n17022_, new_n17023_, new_n17024_, new_n17025_,
    new_n17026_, new_n17027_, new_n17028_, new_n17029_, new_n17030_,
    new_n17031_, new_n17032_, new_n17033_, new_n17034_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17039_, new_n17040_,
    new_n17041_, new_n17042_, new_n17043_, new_n17044_, new_n17045_,
    new_n17046_, new_n17047_, new_n17048_, new_n17049_, new_n17050_,
    new_n17051_, new_n17052_, new_n17053_, new_n17054_, new_n17055_,
    new_n17056_, new_n17057_, new_n17058_, new_n17059_, new_n17060_,
    new_n17061_, new_n17062_, new_n17063_, new_n17064_, new_n17065_,
    new_n17066_, new_n17067_, new_n17068_, new_n17069_, new_n17070_,
    new_n17071_, new_n17072_, new_n17073_, new_n17074_, new_n17075_,
    new_n17076_, new_n17077_, new_n17078_, new_n17079_, new_n17080_,
    new_n17081_, new_n17082_, new_n17083_, new_n17084_, new_n17085_,
    new_n17086_, new_n17087_, new_n17088_, new_n17089_, new_n17090_,
    new_n17091_, new_n17092_, new_n17093_, new_n17094_, new_n17095_,
    new_n17096_, new_n17097_, new_n17098_, new_n17099_, new_n17100_,
    new_n17101_, new_n17102_, new_n17103_, new_n17104_, new_n17105_,
    new_n17106_, new_n17107_, new_n17108_, new_n17109_, new_n17110_,
    new_n17111_, new_n17112_, new_n17113_, new_n17114_, new_n17115_,
    new_n17116_, new_n17117_, new_n17118_, new_n17119_, new_n17120_,
    new_n17121_, new_n17122_, new_n17123_, new_n17124_, new_n17125_,
    new_n17126_, new_n17127_, new_n17128_, new_n17129_, new_n17130_,
    new_n17131_, new_n17132_, new_n17133_, new_n17134_, new_n17135_,
    new_n17136_, new_n17137_, new_n17138_, new_n17139_, new_n17140_,
    new_n17141_, new_n17142_, new_n17143_, new_n17144_, new_n17145_,
    new_n17146_, new_n17147_, new_n17148_, new_n17149_, new_n17150_,
    new_n17151_, new_n17152_, new_n17153_, new_n17154_, new_n17155_,
    new_n17156_, new_n17157_, new_n17158_, new_n17159_, new_n17160_,
    new_n17161_, new_n17162_, new_n17163_, new_n17164_, new_n17165_,
    new_n17166_, new_n17167_, new_n17168_, new_n17169_, new_n17170_,
    new_n17171_, new_n17172_, new_n17173_, new_n17174_, new_n17175_,
    new_n17176_, new_n17177_, new_n17178_, new_n17179_, new_n17180_,
    new_n17181_, new_n17182_, new_n17183_, new_n17184_, new_n17185_,
    new_n17186_, new_n17187_, new_n17188_, new_n17189_, new_n17190_,
    new_n17191_, new_n17192_, new_n17193_, new_n17194_, new_n17195_,
    new_n17196_, new_n17197_, new_n17198_, new_n17199_, new_n17200_,
    new_n17201_, new_n17202_, new_n17203_, new_n17204_, new_n17205_,
    new_n17206_, new_n17207_, new_n17208_, new_n17209_, new_n17210_,
    new_n17211_, new_n17212_, new_n17213_, new_n17214_, new_n17215_,
    new_n17216_, new_n17217_, new_n17218_, new_n17219_, new_n17220_,
    new_n17221_, new_n17222_, new_n17223_, new_n17224_, new_n17225_,
    new_n17226_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17233_, new_n17234_, new_n17235_,
    new_n17236_, new_n17237_, new_n17238_, new_n17239_, new_n17240_,
    new_n17241_, new_n17242_, new_n17243_, new_n17244_, new_n17245_,
    new_n17246_, new_n17247_, new_n17248_, new_n17249_, new_n17250_,
    new_n17251_, new_n17252_, new_n17253_, new_n17254_, new_n17255_,
    new_n17256_, new_n17257_, new_n17258_, new_n17259_, new_n17260_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17283_, new_n17284_, new_n17285_,
    new_n17286_, new_n17287_, new_n17288_, new_n17289_, new_n17290_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17345_,
    new_n17346_, new_n17347_, new_n17348_, new_n17349_, new_n17350_,
    new_n17351_, new_n17352_, new_n17353_, new_n17354_, new_n17355_,
    new_n17356_, new_n17357_, new_n17358_, new_n17359_, new_n17360_,
    new_n17361_, new_n17362_, new_n17363_, new_n17364_, new_n17365_,
    new_n17366_, new_n17367_, new_n17368_, new_n17369_, new_n17370_,
    new_n17371_, new_n17372_, new_n17373_, new_n17374_, new_n17375_,
    new_n17376_, new_n17377_, new_n17378_, new_n17379_, new_n17380_,
    new_n17381_, new_n17382_, new_n17383_, new_n17384_, new_n17385_,
    new_n17386_, new_n17387_, new_n17388_, new_n17389_, new_n17390_,
    new_n17391_, new_n17392_, new_n17393_, new_n17394_, new_n17395_,
    new_n17396_, new_n17397_, new_n17398_, new_n17399_, new_n17400_,
    new_n17401_, new_n17402_, new_n17403_, new_n17404_, new_n17405_,
    new_n17406_, new_n17407_, new_n17408_, new_n17409_, new_n17410_,
    new_n17411_, new_n17412_, new_n17413_, new_n17414_, new_n17415_,
    new_n17416_, new_n17417_, new_n17418_, new_n17419_, new_n17420_,
    new_n17421_, new_n17422_, new_n17423_, new_n17424_, new_n17425_,
    new_n17426_, new_n17427_, new_n17428_, new_n17429_, new_n17430_,
    new_n17431_, new_n17432_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17438_, new_n17439_, new_n17440_,
    new_n17441_, new_n17442_, new_n17443_, new_n17444_, new_n17445_,
    new_n17446_, new_n17447_, new_n17448_, new_n17449_, new_n17450_,
    new_n17451_, new_n17452_, new_n17453_, new_n17454_, new_n17455_,
    new_n17456_, new_n17457_, new_n17458_, new_n17459_, new_n17460_,
    new_n17461_, new_n17462_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17468_, new_n17469_, new_n17470_,
    new_n17471_, new_n17472_, new_n17473_, new_n17474_, new_n17475_,
    new_n17476_, new_n17477_, new_n17478_, new_n17479_, new_n17480_,
    new_n17481_, new_n17482_, new_n17483_, new_n17484_, new_n17485_,
    new_n17486_, new_n17487_, new_n17488_, new_n17489_, new_n17490_,
    new_n17491_, new_n17492_, new_n17493_, new_n17494_, new_n17495_,
    new_n17496_, new_n17497_, new_n17498_, new_n17499_, new_n17500_,
    new_n17501_, new_n17502_, new_n17503_, new_n17504_, new_n17505_,
    new_n17506_, new_n17507_, new_n17508_, new_n17509_, new_n17510_,
    new_n17511_, new_n17512_, new_n17513_, new_n17514_, new_n17515_,
    new_n17516_, new_n17517_, new_n17518_, new_n17519_, new_n17520_,
    new_n17521_, new_n17522_, new_n17523_, new_n17524_, new_n17525_,
    new_n17526_, new_n17527_, new_n17528_, new_n17529_, new_n17530_,
    new_n17531_, new_n17532_, new_n17533_, new_n17534_, new_n17535_,
    new_n17536_, new_n17537_, new_n17538_, new_n17539_, new_n17540_,
    new_n17541_, new_n17542_, new_n17543_, new_n17544_, new_n17545_,
    new_n17546_, new_n17547_, new_n17548_, new_n17549_, new_n17550_,
    new_n17551_, new_n17552_, new_n17553_, new_n17554_, new_n17555_,
    new_n17556_, new_n17557_, new_n17558_, new_n17559_, new_n17560_,
    new_n17561_, new_n17562_, new_n17563_, new_n17564_, new_n17565_,
    new_n17566_, new_n17567_, new_n17568_, new_n17569_, new_n17570_,
    new_n17571_, new_n17572_, new_n17573_, new_n17574_, new_n17575_,
    new_n17576_, new_n17577_, new_n17578_, new_n17579_, new_n17580_,
    new_n17581_, new_n17582_, new_n17583_, new_n17584_, new_n17585_,
    new_n17586_, new_n17587_, new_n17588_, new_n17589_, new_n17590_,
    new_n17591_, new_n17592_, new_n17593_, new_n17594_, new_n17595_,
    new_n17596_, new_n17597_, new_n17598_, new_n17599_, new_n17600_,
    new_n17601_, new_n17602_, new_n17603_, new_n17604_, new_n17605_,
    new_n17606_, new_n17607_, new_n17608_, new_n17609_, new_n17610_,
    new_n17611_, new_n17612_, new_n17613_, new_n17614_, new_n17615_,
    new_n17616_, new_n17617_, new_n17618_, new_n17619_, new_n17620_,
    new_n17621_, new_n17622_, new_n17623_, new_n17624_, new_n17625_,
    new_n17626_, new_n17627_, new_n17628_, new_n17629_, new_n17630_,
    new_n17631_, new_n17632_, new_n17633_, new_n17634_, new_n17635_,
    new_n17636_, new_n17637_, new_n17638_, new_n17639_, new_n17640_,
    new_n17641_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17667_, new_n17668_, new_n17669_, new_n17670_,
    new_n17671_, new_n17672_, new_n17673_, new_n17674_, new_n17675_,
    new_n17676_, new_n17677_, new_n17678_, new_n17679_, new_n17680_,
    new_n17681_, new_n17682_, new_n17683_, new_n17684_, new_n17685_,
    new_n17686_, new_n17687_, new_n17688_, new_n17689_, new_n17690_,
    new_n17691_, new_n17692_, new_n17693_, new_n17694_, new_n17695_,
    new_n17696_, new_n17697_, new_n17698_, new_n17699_, new_n17700_,
    new_n17701_, new_n17702_, new_n17703_, new_n17704_, new_n17705_,
    new_n17706_, new_n17707_, new_n17708_, new_n17709_, new_n17710_,
    new_n17711_, new_n17712_, new_n17713_, new_n17714_, new_n17715_,
    new_n17716_, new_n17717_, new_n17718_, new_n17719_, new_n17720_,
    new_n17721_, new_n17722_, new_n17723_, new_n17724_, new_n17725_,
    new_n17726_, new_n17727_, new_n17728_, new_n17729_, new_n17730_,
    new_n17731_, new_n17732_, new_n17733_, new_n17734_, new_n17735_,
    new_n17736_, new_n17737_, new_n17738_, new_n17739_, new_n17740_,
    new_n17741_, new_n17742_, new_n17743_, new_n17744_, new_n17745_,
    new_n17746_, new_n17747_, new_n17748_, new_n17749_, new_n17750_,
    new_n17751_, new_n17752_, new_n17753_, new_n17754_, new_n17755_,
    new_n17756_, new_n17757_, new_n17758_, new_n17759_, new_n17760_,
    new_n17761_, new_n17762_, new_n17763_, new_n17764_, new_n17765_,
    new_n17766_, new_n17767_, new_n17768_, new_n17769_, new_n17770_,
    new_n17771_, new_n17772_, new_n17773_, new_n17774_, new_n17775_,
    new_n17776_, new_n17777_, new_n17778_, new_n17779_, new_n17780_,
    new_n17781_, new_n17782_, new_n17783_, new_n17784_, new_n17785_,
    new_n17786_, new_n17787_, new_n17788_, new_n17789_, new_n17790_,
    new_n17791_, new_n17792_, new_n17793_, new_n17794_, new_n17795_,
    new_n17796_, new_n17797_, new_n17798_, new_n17799_, new_n17800_,
    new_n17801_, new_n17802_, new_n17803_, new_n17804_, new_n17805_,
    new_n17806_, new_n17807_, new_n17808_, new_n17809_, new_n17810_,
    new_n17811_, new_n17812_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17824_, new_n17825_,
    new_n17826_, new_n17827_, new_n17828_, new_n17829_, new_n17830_,
    new_n17831_, new_n17832_, new_n17833_, new_n17834_, new_n17835_,
    new_n17836_, new_n17837_, new_n17838_, new_n17839_, new_n17840_,
    new_n17841_, new_n17842_, new_n17843_, new_n17844_, new_n17845_,
    new_n17846_, new_n17847_, new_n17848_, new_n17849_, new_n17850_,
    new_n17851_, new_n17852_, new_n17853_, new_n17854_, new_n17855_,
    new_n17856_, new_n17857_, new_n17858_, new_n17859_, new_n17860_,
    new_n17861_, new_n17862_, new_n17863_, new_n17864_, new_n17865_,
    new_n17866_, new_n17867_, new_n17868_, new_n17869_, new_n17870_,
    new_n17871_, new_n17872_, new_n17873_, new_n17874_, new_n17875_,
    new_n17876_, new_n17877_, new_n17878_, new_n17879_, new_n17880_,
    new_n17881_, new_n17882_, new_n17883_, new_n17884_, new_n17885_,
    new_n17886_, new_n17887_, new_n17888_, new_n17889_, new_n17890_,
    new_n17891_, new_n17892_, new_n17893_, new_n17894_, new_n17895_,
    new_n17896_, new_n17897_, new_n17898_, new_n17899_, new_n17900_,
    new_n17901_, new_n17902_, new_n17903_, new_n17904_, new_n17905_,
    new_n17906_, new_n17907_, new_n17908_, new_n17909_, new_n17910_,
    new_n17911_, new_n17912_, new_n17913_, new_n17914_, new_n17915_,
    new_n17916_, new_n17917_, new_n17918_, new_n17919_, new_n17920_,
    new_n17921_, new_n17922_, new_n17923_, new_n17924_, new_n17925_,
    new_n17926_, new_n17927_, new_n17928_, new_n17929_, new_n17930_,
    new_n17931_, new_n17932_, new_n17933_, new_n17934_, new_n17935_,
    new_n17936_, new_n17937_, new_n17938_, new_n17939_, new_n17940_,
    new_n17941_, new_n17942_, new_n17943_, new_n17944_, new_n17945_,
    new_n17946_, new_n17947_, new_n17948_, new_n17949_, new_n17950_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17970_,
    new_n17971_, new_n17972_, new_n17973_, new_n17974_, new_n17975_,
    new_n17976_, new_n17977_, new_n17978_, new_n17979_, new_n17980_,
    new_n17981_, new_n17982_, new_n17983_, new_n17984_, new_n17985_,
    new_n17986_, new_n17987_, new_n17988_, new_n17989_, new_n17990_,
    new_n17991_, new_n17992_, new_n17993_, new_n17994_, new_n17995_,
    new_n17996_, new_n17997_, new_n17998_, new_n17999_, new_n18000_,
    new_n18001_, new_n18002_, new_n18003_, new_n18004_, new_n18005_,
    new_n18006_, new_n18007_, new_n18008_, new_n18009_, new_n18010_,
    new_n18011_, new_n18012_, new_n18013_, new_n18014_, new_n18015_,
    new_n18016_, new_n18017_, new_n18018_, new_n18019_, new_n18020_,
    new_n18021_, new_n18022_, new_n18023_, new_n18024_, new_n18025_,
    new_n18026_, new_n18027_, new_n18028_, new_n18029_, new_n18030_,
    new_n18031_, new_n18032_, new_n18033_, new_n18034_, new_n18035_,
    new_n18036_, new_n18037_, new_n18038_, new_n18039_, new_n18040_,
    new_n18041_, new_n18042_, new_n18043_, new_n18044_, new_n18045_,
    new_n18046_, new_n18047_, new_n18048_, new_n18049_, new_n18050_,
    new_n18051_, new_n18052_, new_n18053_, new_n18054_, new_n18055_,
    new_n18056_, new_n18057_, new_n18058_, new_n18059_, new_n18060_,
    new_n18061_, new_n18062_, new_n18063_, new_n18064_, new_n18065_,
    new_n18066_, new_n18067_, new_n18068_, new_n18069_, new_n18070_,
    new_n18071_, new_n18072_, new_n18073_, new_n18074_, new_n18075_,
    new_n18076_, new_n18077_, new_n18078_, new_n18079_, new_n18080_,
    new_n18081_, new_n18082_, new_n18083_, new_n18084_, new_n18085_,
    new_n18086_, new_n18087_, new_n18088_, new_n18089_, new_n18090_,
    new_n18091_, new_n18092_, new_n18093_, new_n18094_, new_n18095_,
    new_n18096_, new_n18097_, new_n18098_, new_n18099_, new_n18100_,
    new_n18101_, new_n18102_, new_n18103_, new_n18104_, new_n18105_,
    new_n18106_, new_n18107_, new_n18108_, new_n18109_, new_n18110_,
    new_n18111_, new_n18112_, new_n18113_, new_n18114_, new_n18115_,
    new_n18116_, new_n18117_, new_n18118_, new_n18119_, new_n18120_,
    new_n18121_, new_n18122_, new_n18123_, new_n18124_, new_n18125_,
    new_n18126_, new_n18127_, new_n18128_, new_n18129_, new_n18130_,
    new_n18131_, new_n18132_, new_n18133_, new_n18134_, new_n18135_,
    new_n18136_, new_n18137_, new_n18138_, new_n18139_, new_n18140_,
    new_n18141_, new_n18142_, new_n18143_, new_n18144_, new_n18145_,
    new_n18146_, new_n18147_, new_n18148_, new_n18149_, new_n18150_,
    new_n18151_, new_n18152_, new_n18153_, new_n18154_, new_n18155_,
    new_n18156_, new_n18157_, new_n18158_, new_n18159_, new_n18160_,
    new_n18161_, new_n18162_, new_n18163_, new_n18164_, new_n18165_,
    new_n18166_, new_n18167_, new_n18168_, new_n18169_, new_n18170_,
    new_n18171_, new_n18172_, new_n18173_, new_n18174_, new_n18175_,
    new_n18176_, new_n18177_, new_n18178_, new_n18179_, new_n18180_,
    new_n18181_, new_n18182_, new_n18183_, new_n18184_, new_n18185_,
    new_n18186_, new_n18187_, new_n18188_, new_n18189_, new_n18190_,
    new_n18191_, new_n18192_, new_n18193_, new_n18194_, new_n18195_,
    new_n18196_, new_n18197_, new_n18198_, new_n18199_, new_n18200_,
    new_n18201_, new_n18202_, new_n18203_, new_n18204_, new_n18205_,
    new_n18206_, new_n18207_, new_n18208_, new_n18209_, new_n18210_,
    new_n18211_, new_n18212_, new_n18213_, new_n18214_, new_n18215_,
    new_n18216_, new_n18217_, new_n18218_, new_n18219_, new_n18220_,
    new_n18221_, new_n18222_, new_n18223_, new_n18224_, new_n18225_,
    new_n18226_, new_n18227_, new_n18228_, new_n18229_, new_n18230_,
    new_n18231_, new_n18232_, new_n18233_, new_n18234_, new_n18235_,
    new_n18236_, new_n18237_, new_n18238_, new_n18239_, new_n18240_,
    new_n18241_, new_n18242_, new_n18243_, new_n18244_, new_n18245_,
    new_n18246_, new_n18247_, new_n18248_, new_n18249_, new_n18250_,
    new_n18251_, new_n18252_, new_n18253_, new_n18254_, new_n18255_,
    new_n18256_, new_n18257_, new_n18258_, new_n18259_, new_n18260_,
    new_n18261_, new_n18262_, new_n18263_, new_n18264_, new_n18265_,
    new_n18266_, new_n18267_, new_n18268_, new_n18269_, new_n18270_,
    new_n18271_, new_n18272_, new_n18273_, new_n18274_, new_n18275_,
    new_n18276_, new_n18277_, new_n18278_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18376_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18381_, new_n18382_, new_n18383_, new_n18384_, new_n18385_,
    new_n18386_, new_n18387_, new_n18388_, new_n18389_, new_n18390_,
    new_n18391_, new_n18392_, new_n18393_, new_n18394_, new_n18395_,
    new_n18396_, new_n18397_, new_n18398_, new_n18399_, new_n18400_,
    new_n18401_, new_n18402_, new_n18403_, new_n18404_, new_n18405_,
    new_n18406_, new_n18407_, new_n18408_, new_n18409_, new_n18410_,
    new_n18411_, new_n18412_, new_n18413_, new_n18414_, new_n18415_,
    new_n18416_, new_n18417_, new_n18418_, new_n18419_, new_n18420_,
    new_n18421_, new_n18422_, new_n18423_, new_n18424_, new_n18425_,
    new_n18426_, new_n18427_, new_n18428_, new_n18429_, new_n18430_,
    new_n18431_, new_n18432_, new_n18433_, new_n18434_, new_n18435_,
    new_n18436_, new_n18437_, new_n18438_, new_n18439_, new_n18440_,
    new_n18441_, new_n18442_, new_n18443_, new_n18444_, new_n18445_,
    new_n18446_, new_n18447_, new_n18448_, new_n18449_, new_n18450_,
    new_n18451_, new_n18452_, new_n18453_, new_n18454_, new_n18455_,
    new_n18456_, new_n18457_, new_n18458_, new_n18459_, new_n18460_,
    new_n18461_, new_n18462_, new_n18463_, new_n18464_, new_n18465_,
    new_n18466_, new_n18467_, new_n18468_, new_n18469_, new_n18470_,
    new_n18471_, new_n18472_, new_n18473_, new_n18474_, new_n18475_,
    new_n18476_, new_n18477_, new_n18478_, new_n18479_, new_n18480_,
    new_n18481_, new_n18482_, new_n18483_, new_n18484_, new_n18485_,
    new_n18486_, new_n18487_, new_n18488_, new_n18489_, new_n18490_,
    new_n18491_, new_n18492_, new_n18493_, new_n18494_, new_n18495_,
    new_n18496_, new_n18497_, new_n18498_, new_n18499_, new_n18500_,
    new_n18501_, new_n18502_, new_n18503_, new_n18504_, new_n18505_,
    new_n18506_, new_n18507_, new_n18508_, new_n18509_, new_n18510_,
    new_n18511_, new_n18512_, new_n18513_, new_n18514_, new_n18515_,
    new_n18516_, new_n18517_, new_n18518_, new_n18519_, new_n18520_,
    new_n18521_, new_n18522_, new_n18523_, new_n18524_, new_n18525_,
    new_n18526_, new_n18527_, new_n18528_, new_n18529_, new_n18530_,
    new_n18531_, new_n18532_, new_n18533_, new_n18534_, new_n18535_,
    new_n18536_, new_n18537_, new_n18538_, new_n18539_, new_n18540_,
    new_n18541_, new_n18542_, new_n18543_, new_n18544_, new_n18545_,
    new_n18546_, new_n18547_, new_n18548_, new_n18549_, new_n18550_,
    new_n18551_, new_n18552_, new_n18553_, new_n18554_, new_n18555_,
    new_n18556_, new_n18557_, new_n18558_, new_n18559_, new_n18560_,
    new_n18561_, new_n18562_, new_n18563_, new_n18564_, new_n18565_,
    new_n18566_, new_n18567_, new_n18568_, new_n18569_, new_n18570_,
    new_n18571_, new_n18572_, new_n18573_, new_n18574_, new_n18575_,
    new_n18576_, new_n18577_, new_n18578_, new_n18579_, new_n18580_,
    new_n18581_, new_n18582_, new_n18583_, new_n18584_, new_n18585_,
    new_n18586_, new_n18587_, new_n18588_, new_n18589_, new_n18590_,
    new_n18591_, new_n18592_, new_n18593_, new_n18594_, new_n18595_,
    new_n18596_, new_n18597_, new_n18598_, new_n18599_, new_n18600_,
    new_n18601_, new_n18602_, new_n18603_, new_n18604_, new_n18605_,
    new_n18606_, new_n18607_, new_n18608_, new_n18609_, new_n18610_,
    new_n18611_, new_n18612_, new_n18613_, new_n18614_, new_n18615_,
    new_n18616_, new_n18617_, new_n18618_, new_n18619_, new_n18620_,
    new_n18621_, new_n18622_, new_n18623_, new_n18624_, new_n18625_,
    new_n18626_, new_n18627_, new_n18628_, new_n18629_, new_n18630_,
    new_n18631_, new_n18632_, new_n18633_, new_n18634_, new_n18635_,
    new_n18636_, new_n18637_, new_n18638_, new_n18639_, new_n18640_,
    new_n18641_, new_n18642_, new_n18643_, new_n18644_, new_n18645_,
    new_n18646_, new_n18647_, new_n18648_, new_n18649_, new_n18650_,
    new_n18651_, new_n18652_, new_n18653_, new_n18654_, new_n18655_,
    new_n18656_, new_n18657_, new_n18658_, new_n18659_, new_n18660_,
    new_n18661_, new_n18662_, new_n18663_, new_n18664_, new_n18665_,
    new_n18666_, new_n18667_, new_n18668_, new_n18669_, new_n18670_,
    new_n18671_, new_n18672_, new_n18673_, new_n18674_, new_n18675_,
    new_n18676_, new_n18677_, new_n18678_, new_n18679_, new_n18680_,
    new_n18681_, new_n18682_, new_n18683_, new_n18684_, new_n18685_,
    new_n18686_, new_n18687_, new_n18688_, new_n18689_, new_n18690_,
    new_n18691_, new_n18692_, new_n18693_, new_n18694_, new_n18695_,
    new_n18696_, new_n18697_, new_n18698_, new_n18699_, new_n18700_,
    new_n18701_, new_n18702_, new_n18703_, new_n18704_, new_n18705_,
    new_n18706_, new_n18707_, new_n18708_, new_n18709_, new_n18710_,
    new_n18711_, new_n18712_, new_n18713_, new_n18714_, new_n18715_,
    new_n18716_, new_n18717_, new_n18718_, new_n18719_, new_n18720_,
    new_n18721_, new_n18722_, new_n18723_, new_n18724_, new_n18725_,
    new_n18726_, new_n18727_, new_n18728_, new_n18729_, new_n18730_,
    new_n18731_, new_n18732_, new_n18733_, new_n18734_, new_n18735_,
    new_n18736_, new_n18737_, new_n18738_, new_n18739_, new_n18740_,
    new_n18741_, new_n18742_, new_n18743_, new_n18744_, new_n18745_,
    new_n18746_, new_n18747_, new_n18748_, new_n18749_, new_n18750_,
    new_n18751_, new_n18752_, new_n18753_, new_n18754_, new_n18755_,
    new_n18756_, new_n18757_, new_n18758_, new_n18759_, new_n18760_,
    new_n18761_, new_n18762_, new_n18763_, new_n18764_, new_n18765_,
    new_n18766_, new_n18767_, new_n18768_, new_n18769_, new_n18770_,
    new_n18771_, new_n18772_, new_n18773_, new_n18774_, new_n18775_,
    new_n18776_, new_n18777_, new_n18778_, new_n18779_, new_n18780_,
    new_n18781_, new_n18782_, new_n18783_, new_n18784_, new_n18785_,
    new_n18786_, new_n18787_, new_n18788_, new_n18789_, new_n18790_,
    new_n18791_, new_n18792_, new_n18793_, new_n18794_, new_n18795_,
    new_n18796_, new_n18797_, new_n18798_, new_n18799_, new_n18800_,
    new_n18801_, new_n18802_, new_n18803_, new_n18804_, new_n18805_,
    new_n18806_, new_n18807_, new_n18808_, new_n18809_, new_n18810_,
    new_n18811_, new_n18812_, new_n18813_, new_n18814_, new_n18815_,
    new_n18816_, new_n18817_, new_n18818_, new_n18819_, new_n18820_,
    new_n18821_, new_n18822_, new_n18823_, new_n18824_, new_n18825_,
    new_n18826_, new_n18827_, new_n18828_, new_n18829_, new_n18830_,
    new_n18831_, new_n18832_, new_n18833_, new_n18834_, new_n18835_,
    new_n18836_, new_n18837_, new_n18838_, new_n18839_, new_n18840_,
    new_n18841_, new_n18842_, new_n18843_, new_n18844_, new_n18845_,
    new_n18846_, new_n18847_, new_n18848_, new_n18849_, new_n18850_,
    new_n18851_, new_n18852_, new_n18853_, new_n18854_, new_n18855_,
    new_n18856_, new_n18857_, new_n18858_, new_n18859_, new_n18860_,
    new_n18861_, new_n18862_, new_n18863_, new_n18864_, new_n18865_,
    new_n18866_, new_n18867_, new_n18868_, new_n18869_, new_n18870_,
    new_n18871_, new_n18872_, new_n18873_, new_n18874_, new_n18875_,
    new_n18876_, new_n18877_, new_n18878_, new_n18879_, new_n18880_,
    new_n18881_, new_n18882_, new_n18883_, new_n18884_, new_n18885_,
    new_n18886_, new_n18887_, new_n18888_, new_n18889_, new_n18890_,
    new_n18891_, new_n18892_, new_n18893_, new_n18894_, new_n18895_,
    new_n18896_, new_n18897_, new_n18898_, new_n18899_, new_n18900_,
    new_n18901_, new_n18902_, new_n18903_, new_n18904_, new_n18905_,
    new_n18906_, new_n18907_, new_n18908_, new_n18909_, new_n18910_,
    new_n18911_, new_n18912_, new_n18913_, new_n18914_, new_n18915_,
    new_n18916_, new_n18917_, new_n18918_, new_n18919_, new_n18920_,
    new_n18921_, new_n18922_, new_n18923_, new_n18924_, new_n18925_,
    new_n18926_, new_n18927_, new_n18928_, new_n18929_, new_n18930_,
    new_n18931_, new_n18932_, new_n18933_, new_n18934_, new_n18935_,
    new_n18936_, new_n18937_, new_n18938_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18944_, new_n18945_,
    new_n18946_, new_n18947_, new_n18948_, new_n18949_, new_n18950_,
    new_n18951_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19107_, new_n19108_, new_n19109_, new_n19110_,
    new_n19111_, new_n19112_, new_n19113_, new_n19114_, new_n19115_,
    new_n19116_, new_n19117_, new_n19118_, new_n19119_, new_n19120_,
    new_n19121_, new_n19122_, new_n19123_, new_n19124_, new_n19125_,
    new_n19126_, new_n19127_, new_n19128_, new_n19129_, new_n19130_,
    new_n19131_, new_n19132_, new_n19133_, new_n19134_, new_n19135_,
    new_n19136_, new_n19137_, new_n19138_, new_n19139_, new_n19140_,
    new_n19141_, new_n19142_, new_n19143_, new_n19144_, new_n19145_,
    new_n19146_, new_n19147_, new_n19148_, new_n19149_, new_n19150_,
    new_n19151_, new_n19152_, new_n19153_, new_n19154_, new_n19155_,
    new_n19156_, new_n19157_, new_n19158_, new_n19159_, new_n19160_,
    new_n19161_, new_n19162_, new_n19163_, new_n19164_, new_n19165_,
    new_n19166_, new_n19167_, new_n19168_, new_n19169_, new_n19170_,
    new_n19171_, new_n19172_, new_n19173_, new_n19174_, new_n19175_,
    new_n19176_, new_n19177_, new_n19178_, new_n19179_, new_n19180_,
    new_n19181_, new_n19182_, new_n19183_, new_n19184_, new_n19185_,
    new_n19186_, new_n19187_, new_n19188_, new_n19189_, new_n19190_,
    new_n19191_, new_n19192_, new_n19193_, new_n19194_, new_n19195_,
    new_n19196_, new_n19197_, new_n19198_, new_n19199_, new_n19200_,
    new_n19201_, new_n19202_, new_n19203_, new_n19204_, new_n19205_,
    new_n19206_, new_n19207_, new_n19208_, new_n19209_, new_n19210_,
    new_n19211_, new_n19212_, new_n19213_, new_n19214_, new_n19215_,
    new_n19216_, new_n19217_, new_n19218_, new_n19219_, new_n19220_,
    new_n19221_, new_n19222_, new_n19223_, new_n19224_, new_n19225_,
    new_n19226_, new_n19227_, new_n19228_, new_n19229_, new_n19230_,
    new_n19231_, new_n19232_, new_n19233_, new_n19234_, new_n19235_,
    new_n19236_, new_n19237_, new_n19238_, new_n19239_, new_n19240_,
    new_n19241_, new_n19242_, new_n19243_, new_n19244_, new_n19245_,
    new_n19246_, new_n19247_, new_n19248_, new_n19249_, new_n19250_,
    new_n19251_, new_n19252_, new_n19253_, new_n19254_, new_n19255_,
    new_n19256_, new_n19257_, new_n19258_, new_n19259_, new_n19260_,
    new_n19261_, new_n19262_, new_n19263_, new_n19264_, new_n19265_,
    new_n19266_, new_n19267_, new_n19268_, new_n19269_, new_n19270_,
    new_n19271_, new_n19272_, new_n19273_, new_n19274_, new_n19275_,
    new_n19276_, new_n19277_, new_n19278_, new_n19279_, new_n19280_,
    new_n19281_, new_n19282_, new_n19283_, new_n19284_, new_n19285_,
    new_n19286_, new_n19287_, new_n19288_, new_n19289_, new_n19290_,
    new_n19291_, new_n19292_, new_n19293_, new_n19294_, new_n19295_,
    new_n19296_, new_n19297_, new_n19298_, new_n19299_, new_n19300_,
    new_n19301_, new_n19302_, new_n19303_, new_n19304_, new_n19305_,
    new_n19306_, new_n19307_, new_n19308_, new_n19309_, new_n19310_,
    new_n19311_, new_n19312_, new_n19313_, new_n19314_, new_n19315_,
    new_n19316_, new_n19317_, new_n19318_, new_n19319_, new_n19320_,
    new_n19321_, new_n19322_, new_n19323_, new_n19324_, new_n19325_,
    new_n19326_, new_n19327_, new_n19328_, new_n19329_, new_n19330_,
    new_n19331_, new_n19332_, new_n19333_, new_n19334_, new_n19335_,
    new_n19336_, new_n19337_, new_n19338_, new_n19339_, new_n19340_,
    new_n19341_, new_n19342_, new_n19343_, new_n19344_, new_n19345_,
    new_n19346_, new_n19347_, new_n19348_, new_n19349_, new_n19350_,
    new_n19351_, new_n19352_, new_n19353_, new_n19354_, new_n19355_,
    new_n19356_, new_n19357_, new_n19358_, new_n19359_, new_n19360_,
    new_n19361_, new_n19362_, new_n19363_, new_n19364_, new_n19365_,
    new_n19366_, new_n19367_, new_n19368_, new_n19369_, new_n19370_,
    new_n19371_, new_n19372_, new_n19373_, new_n19374_, new_n19375_,
    new_n19376_, new_n19377_, new_n19378_, new_n19379_, new_n19380_,
    new_n19381_, new_n19382_, new_n19383_, new_n19384_, new_n19385_,
    new_n19386_, new_n19387_, new_n19388_, new_n19389_, new_n19390_,
    new_n19391_, new_n19392_, new_n19393_, new_n19394_, new_n19395_,
    new_n19396_, new_n19397_, new_n19398_, new_n19399_, new_n19400_,
    new_n19401_, new_n19402_, new_n19403_, new_n19404_, new_n19405_,
    new_n19406_, new_n19407_, new_n19408_, new_n19409_, new_n19410_,
    new_n19411_, new_n19412_, new_n19413_, new_n19414_, new_n19415_,
    new_n19416_, new_n19417_, new_n19418_, new_n19419_, new_n19420_,
    new_n19421_, new_n19422_, new_n19423_, new_n19424_, new_n19425_,
    new_n19426_, new_n19427_, new_n19428_, new_n19429_, new_n19430_,
    new_n19431_, new_n19432_, new_n19433_, new_n19434_, new_n19435_,
    new_n19436_, new_n19437_, new_n19438_, new_n19439_, new_n19440_,
    new_n19441_, new_n19442_, new_n19443_, new_n19444_, new_n19445_,
    new_n19446_, new_n19447_, new_n19448_, new_n19449_, new_n19450_,
    new_n19451_, new_n19452_, new_n19453_, new_n19454_, new_n19455_,
    new_n19456_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19513_, new_n19514_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19738_, new_n19739_, new_n19740_,
    new_n19741_, new_n19742_, new_n19743_, new_n19744_, new_n19745_,
    new_n19746_, new_n19747_, new_n19748_, new_n19749_, new_n19750_,
    new_n19751_, new_n19752_, new_n19753_, new_n19754_, new_n19755_,
    new_n19756_, new_n19757_, new_n19758_, new_n19759_, new_n19760_,
    new_n19761_, new_n19762_, new_n19763_, new_n19764_, new_n19765_,
    new_n19766_, new_n19767_, new_n19768_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19779_, new_n19780_, new_n19783_, new_n19787_,
    new_n19789_, new_n19790_, new_n19791_, new_n19792_, new_n19793_,
    new_n19794_, new_n19795_, new_n19796_, new_n19797_, new_n19798_;
  INV_X1     g00000(.I(\A[938] ), .ZN(new_n1003_));
  NOR2_X1    g00001(.A1(new_n1003_), .A2(\A[937] ), .ZN(new_n1004_));
  NAND2_X1   g00002(.A1(new_n1003_), .A2(\A[937] ), .ZN(new_n1005_));
  NAND2_X1   g00003(.A1(new_n1005_), .A2(\A[939] ), .ZN(new_n1006_));
  INV_X1     g00004(.I(\A[937] ), .ZN(new_n1007_));
  NOR2_X1    g00005(.A1(new_n1007_), .A2(\A[938] ), .ZN(new_n1008_));
  NOR2_X1    g00006(.A1(new_n1004_), .A2(new_n1008_), .ZN(new_n1009_));
  OAI22_X1   g00007(.A1(new_n1009_), .A2(\A[939] ), .B1(new_n1006_), .B2(new_n1004_), .ZN(new_n1010_));
  INV_X1     g00008(.I(\A[941] ), .ZN(new_n1011_));
  NOR2_X1    g00009(.A1(new_n1011_), .A2(\A[940] ), .ZN(new_n1012_));
  NAND2_X1   g00010(.A1(new_n1011_), .A2(\A[940] ), .ZN(new_n1013_));
  NAND2_X1   g00011(.A1(new_n1013_), .A2(\A[942] ), .ZN(new_n1014_));
  INV_X1     g00012(.I(\A[940] ), .ZN(new_n1015_));
  NOR2_X1    g00013(.A1(new_n1015_), .A2(\A[941] ), .ZN(new_n1016_));
  NOR2_X1    g00014(.A1(new_n1012_), .A2(new_n1016_), .ZN(new_n1017_));
  OAI22_X1   g00015(.A1(new_n1017_), .A2(\A[942] ), .B1(new_n1014_), .B2(new_n1012_), .ZN(new_n1018_));
  XOR2_X1    g00016(.A1(new_n1010_), .A2(new_n1018_), .Z(new_n1019_));
  INV_X1     g00017(.I(\A[942] ), .ZN(new_n1020_));
  NOR2_X1    g00018(.A1(new_n1015_), .A2(new_n1011_), .ZN(new_n1021_));
  INV_X1     g00019(.I(new_n1021_), .ZN(new_n1022_));
  OAI21_X1   g00020(.A1(new_n1017_), .A2(new_n1020_), .B(new_n1022_), .ZN(new_n1023_));
  INV_X1     g00021(.I(\A[939] ), .ZN(new_n1024_));
  NOR2_X1    g00022(.A1(new_n1007_), .A2(new_n1003_), .ZN(new_n1025_));
  INV_X1     g00023(.I(new_n1025_), .ZN(new_n1026_));
  OAI21_X1   g00024(.A1(new_n1009_), .A2(new_n1024_), .B(new_n1026_), .ZN(new_n1027_));
  NAND2_X1   g00025(.A1(new_n1007_), .A2(\A[938] ), .ZN(new_n1028_));
  NOR2_X1    g00026(.A1(new_n1008_), .A2(new_n1024_), .ZN(new_n1029_));
  NAND2_X1   g00027(.A1(new_n1028_), .A2(new_n1005_), .ZN(new_n1030_));
  AOI22_X1   g00028(.A1(new_n1030_), .A2(new_n1024_), .B1(new_n1029_), .B2(new_n1028_), .ZN(new_n1031_));
  NAND2_X1   g00029(.A1(new_n1015_), .A2(\A[941] ), .ZN(new_n1032_));
  NOR2_X1    g00030(.A1(new_n1016_), .A2(new_n1020_), .ZN(new_n1033_));
  NAND2_X1   g00031(.A1(new_n1032_), .A2(new_n1013_), .ZN(new_n1034_));
  AOI22_X1   g00032(.A1(new_n1034_), .A2(new_n1020_), .B1(new_n1033_), .B2(new_n1032_), .ZN(new_n1035_));
  NOR2_X1    g00033(.A1(new_n1031_), .A2(new_n1035_), .ZN(new_n1036_));
  NAND3_X1   g00034(.A1(new_n1036_), .A2(new_n1023_), .A3(new_n1027_), .ZN(new_n1037_));
  NAND2_X1   g00035(.A1(new_n1019_), .A2(new_n1037_), .ZN(new_n1038_));
  INV_X1     g00036(.I(\A[933] ), .ZN(new_n1039_));
  INV_X1     g00037(.I(\A[931] ), .ZN(new_n1040_));
  NAND2_X1   g00038(.A1(new_n1040_), .A2(\A[932] ), .ZN(new_n1041_));
  NOR2_X1    g00039(.A1(new_n1040_), .A2(\A[932] ), .ZN(new_n1042_));
  NOR2_X1    g00040(.A1(new_n1042_), .A2(new_n1039_), .ZN(new_n1043_));
  INV_X1     g00041(.I(\A[932] ), .ZN(new_n1044_));
  NAND2_X1   g00042(.A1(new_n1044_), .A2(\A[931] ), .ZN(new_n1045_));
  NAND2_X1   g00043(.A1(new_n1041_), .A2(new_n1045_), .ZN(new_n1046_));
  AOI22_X1   g00044(.A1(new_n1046_), .A2(new_n1039_), .B1(new_n1043_), .B2(new_n1041_), .ZN(new_n1047_));
  INV_X1     g00045(.I(\A[936] ), .ZN(new_n1048_));
  INV_X1     g00046(.I(\A[934] ), .ZN(new_n1049_));
  NAND2_X1   g00047(.A1(new_n1049_), .A2(\A[935] ), .ZN(new_n1050_));
  INV_X1     g00048(.I(\A[935] ), .ZN(new_n1051_));
  AOI21_X1   g00049(.A1(\A[934] ), .A2(new_n1051_), .B(new_n1048_), .ZN(new_n1052_));
  NAND2_X1   g00050(.A1(new_n1051_), .A2(\A[934] ), .ZN(new_n1053_));
  NAND2_X1   g00051(.A1(new_n1050_), .A2(new_n1053_), .ZN(new_n1054_));
  AOI22_X1   g00052(.A1(new_n1054_), .A2(new_n1048_), .B1(new_n1050_), .B2(new_n1052_), .ZN(new_n1055_));
  XOR2_X1    g00053(.A1(new_n1047_), .A2(new_n1055_), .Z(new_n1056_));
  NOR2_X1    g00054(.A1(new_n1051_), .A2(\A[934] ), .ZN(new_n1057_));
  NOR2_X1    g00055(.A1(new_n1049_), .A2(\A[935] ), .ZN(new_n1058_));
  NOR2_X1    g00056(.A1(new_n1057_), .A2(new_n1058_), .ZN(new_n1059_));
  NOR2_X1    g00057(.A1(new_n1049_), .A2(new_n1051_), .ZN(new_n1060_));
  INV_X1     g00058(.I(new_n1060_), .ZN(new_n1061_));
  OAI21_X1   g00059(.A1(new_n1059_), .A2(new_n1048_), .B(new_n1061_), .ZN(new_n1062_));
  NOR2_X1    g00060(.A1(new_n1044_), .A2(\A[931] ), .ZN(new_n1063_));
  NOR2_X1    g00061(.A1(new_n1063_), .A2(new_n1042_), .ZN(new_n1064_));
  NOR2_X1    g00062(.A1(new_n1040_), .A2(new_n1044_), .ZN(new_n1065_));
  INV_X1     g00063(.I(new_n1065_), .ZN(new_n1066_));
  OAI21_X1   g00064(.A1(new_n1064_), .A2(new_n1039_), .B(new_n1066_), .ZN(new_n1067_));
  NOR2_X1    g00065(.A1(new_n1047_), .A2(new_n1055_), .ZN(new_n1068_));
  NAND3_X1   g00066(.A1(new_n1068_), .A2(new_n1062_), .A3(new_n1067_), .ZN(new_n1069_));
  NAND2_X1   g00067(.A1(new_n1056_), .A2(new_n1069_), .ZN(new_n1070_));
  XOR2_X1    g00068(.A1(new_n1038_), .A2(new_n1070_), .Z(new_n1071_));
  INV_X1     g00069(.I(\A[927] ), .ZN(new_n1072_));
  INV_X1     g00070(.I(\A[925] ), .ZN(new_n1073_));
  NAND2_X1   g00071(.A1(new_n1073_), .A2(\A[926] ), .ZN(new_n1074_));
  NOR2_X1    g00072(.A1(new_n1073_), .A2(\A[926] ), .ZN(new_n1075_));
  NOR2_X1    g00073(.A1(new_n1075_), .A2(new_n1072_), .ZN(new_n1076_));
  INV_X1     g00074(.I(\A[926] ), .ZN(new_n1077_));
  NAND2_X1   g00075(.A1(new_n1077_), .A2(\A[925] ), .ZN(new_n1078_));
  NAND2_X1   g00076(.A1(new_n1074_), .A2(new_n1078_), .ZN(new_n1079_));
  AOI22_X1   g00077(.A1(new_n1079_), .A2(new_n1072_), .B1(new_n1076_), .B2(new_n1074_), .ZN(new_n1080_));
  INV_X1     g00078(.I(\A[930] ), .ZN(new_n1081_));
  INV_X1     g00079(.I(\A[928] ), .ZN(new_n1082_));
  NAND2_X1   g00080(.A1(new_n1082_), .A2(\A[929] ), .ZN(new_n1083_));
  INV_X1     g00081(.I(\A[929] ), .ZN(new_n1084_));
  AOI21_X1   g00082(.A1(\A[928] ), .A2(new_n1084_), .B(new_n1081_), .ZN(new_n1085_));
  NAND2_X1   g00083(.A1(new_n1084_), .A2(\A[928] ), .ZN(new_n1086_));
  NAND2_X1   g00084(.A1(new_n1083_), .A2(new_n1086_), .ZN(new_n1087_));
  AOI22_X1   g00085(.A1(new_n1087_), .A2(new_n1081_), .B1(new_n1083_), .B2(new_n1085_), .ZN(new_n1088_));
  XOR2_X1    g00086(.A1(new_n1080_), .A2(new_n1088_), .Z(new_n1089_));
  AND2_X2    g00087(.A1(new_n1083_), .A2(new_n1086_), .Z(new_n1090_));
  NOR2_X1    g00088(.A1(new_n1082_), .A2(new_n1084_), .ZN(new_n1091_));
  INV_X1     g00089(.I(new_n1091_), .ZN(new_n1092_));
  OAI21_X1   g00090(.A1(new_n1090_), .A2(new_n1081_), .B(new_n1092_), .ZN(new_n1093_));
  NOR2_X1    g00091(.A1(new_n1077_), .A2(\A[925] ), .ZN(new_n1094_));
  NOR2_X1    g00092(.A1(new_n1094_), .A2(new_n1075_), .ZN(new_n1095_));
  NOR2_X1    g00093(.A1(new_n1073_), .A2(new_n1077_), .ZN(new_n1096_));
  INV_X1     g00094(.I(new_n1096_), .ZN(new_n1097_));
  OAI21_X1   g00095(.A1(new_n1095_), .A2(new_n1072_), .B(new_n1097_), .ZN(new_n1098_));
  NOR2_X1    g00096(.A1(new_n1080_), .A2(new_n1088_), .ZN(new_n1099_));
  NAND3_X1   g00097(.A1(new_n1099_), .A2(new_n1093_), .A3(new_n1098_), .ZN(new_n1100_));
  NAND2_X1   g00098(.A1(new_n1089_), .A2(new_n1100_), .ZN(new_n1101_));
  INV_X1     g00099(.I(\A[921] ), .ZN(new_n1102_));
  INV_X1     g00100(.I(\A[919] ), .ZN(new_n1103_));
  NAND2_X1   g00101(.A1(new_n1103_), .A2(\A[920] ), .ZN(new_n1104_));
  NOR2_X1    g00102(.A1(new_n1103_), .A2(\A[920] ), .ZN(new_n1105_));
  NOR2_X1    g00103(.A1(new_n1105_), .A2(new_n1102_), .ZN(new_n1106_));
  INV_X1     g00104(.I(\A[920] ), .ZN(new_n1107_));
  NAND2_X1   g00105(.A1(new_n1107_), .A2(\A[919] ), .ZN(new_n1108_));
  NAND2_X1   g00106(.A1(new_n1104_), .A2(new_n1108_), .ZN(new_n1109_));
  AOI22_X1   g00107(.A1(new_n1109_), .A2(new_n1102_), .B1(new_n1106_), .B2(new_n1104_), .ZN(new_n1110_));
  INV_X1     g00108(.I(\A[924] ), .ZN(new_n1111_));
  INV_X1     g00109(.I(\A[922] ), .ZN(new_n1112_));
  NAND2_X1   g00110(.A1(new_n1112_), .A2(\A[923] ), .ZN(new_n1113_));
  INV_X1     g00111(.I(\A[923] ), .ZN(new_n1114_));
  AOI21_X1   g00112(.A1(\A[922] ), .A2(new_n1114_), .B(new_n1111_), .ZN(new_n1115_));
  NAND2_X1   g00113(.A1(new_n1114_), .A2(\A[922] ), .ZN(new_n1116_));
  NAND2_X1   g00114(.A1(new_n1113_), .A2(new_n1116_), .ZN(new_n1117_));
  AOI22_X1   g00115(.A1(new_n1117_), .A2(new_n1111_), .B1(new_n1113_), .B2(new_n1115_), .ZN(new_n1118_));
  XOR2_X1    g00116(.A1(new_n1110_), .A2(new_n1118_), .Z(new_n1119_));
  XNOR2_X1   g00117(.A1(\A[922] ), .A2(\A[923] ), .ZN(new_n1120_));
  NOR2_X1    g00118(.A1(new_n1112_), .A2(new_n1114_), .ZN(new_n1121_));
  INV_X1     g00119(.I(new_n1121_), .ZN(new_n1122_));
  OAI21_X1   g00120(.A1(new_n1120_), .A2(new_n1111_), .B(new_n1122_), .ZN(new_n1123_));
  NOR2_X1    g00121(.A1(new_n1107_), .A2(\A[919] ), .ZN(new_n1124_));
  NOR2_X1    g00122(.A1(new_n1124_), .A2(new_n1105_), .ZN(new_n1125_));
  NOR2_X1    g00123(.A1(new_n1103_), .A2(new_n1107_), .ZN(new_n1126_));
  INV_X1     g00124(.I(new_n1126_), .ZN(new_n1127_));
  OAI21_X1   g00125(.A1(new_n1125_), .A2(new_n1102_), .B(new_n1127_), .ZN(new_n1128_));
  NOR2_X1    g00126(.A1(new_n1110_), .A2(new_n1118_), .ZN(new_n1129_));
  NAND3_X1   g00127(.A1(new_n1129_), .A2(new_n1123_), .A3(new_n1128_), .ZN(new_n1130_));
  NAND2_X1   g00128(.A1(new_n1119_), .A2(new_n1130_), .ZN(new_n1131_));
  XOR2_X1    g00129(.A1(new_n1101_), .A2(new_n1131_), .Z(new_n1132_));
  XOR2_X1    g00130(.A1(new_n1071_), .A2(new_n1132_), .Z(new_n1133_));
  INV_X1     g00131(.I(\A[914] ), .ZN(new_n1134_));
  NOR2_X1    g00132(.A1(new_n1134_), .A2(\A[913] ), .ZN(new_n1135_));
  NAND2_X1   g00133(.A1(new_n1134_), .A2(\A[913] ), .ZN(new_n1136_));
  NAND2_X1   g00134(.A1(new_n1136_), .A2(\A[915] ), .ZN(new_n1137_));
  INV_X1     g00135(.I(\A[913] ), .ZN(new_n1138_));
  NOR2_X1    g00136(.A1(new_n1138_), .A2(\A[914] ), .ZN(new_n1139_));
  NOR2_X1    g00137(.A1(new_n1135_), .A2(new_n1139_), .ZN(new_n1140_));
  OAI22_X1   g00138(.A1(new_n1140_), .A2(\A[915] ), .B1(new_n1137_), .B2(new_n1135_), .ZN(new_n1141_));
  INV_X1     g00139(.I(\A[917] ), .ZN(new_n1142_));
  NOR2_X1    g00140(.A1(new_n1142_), .A2(\A[916] ), .ZN(new_n1143_));
  NAND2_X1   g00141(.A1(new_n1142_), .A2(\A[916] ), .ZN(new_n1144_));
  NAND2_X1   g00142(.A1(new_n1144_), .A2(\A[918] ), .ZN(new_n1145_));
  INV_X1     g00143(.I(\A[916] ), .ZN(new_n1146_));
  NOR2_X1    g00144(.A1(new_n1146_), .A2(\A[917] ), .ZN(new_n1147_));
  NOR2_X1    g00145(.A1(new_n1143_), .A2(new_n1147_), .ZN(new_n1148_));
  OAI22_X1   g00146(.A1(new_n1148_), .A2(\A[918] ), .B1(new_n1145_), .B2(new_n1143_), .ZN(new_n1149_));
  XOR2_X1    g00147(.A1(new_n1141_), .A2(new_n1149_), .Z(new_n1150_));
  INV_X1     g00148(.I(\A[918] ), .ZN(new_n1151_));
  NOR2_X1    g00149(.A1(new_n1146_), .A2(new_n1142_), .ZN(new_n1152_));
  INV_X1     g00150(.I(new_n1152_), .ZN(new_n1153_));
  OAI21_X1   g00151(.A1(new_n1148_), .A2(new_n1151_), .B(new_n1153_), .ZN(new_n1154_));
  INV_X1     g00152(.I(\A[915] ), .ZN(new_n1155_));
  NOR2_X1    g00153(.A1(new_n1138_), .A2(new_n1134_), .ZN(new_n1156_));
  INV_X1     g00154(.I(new_n1156_), .ZN(new_n1157_));
  OAI21_X1   g00155(.A1(new_n1140_), .A2(new_n1155_), .B(new_n1157_), .ZN(new_n1158_));
  NAND2_X1   g00156(.A1(new_n1138_), .A2(\A[914] ), .ZN(new_n1159_));
  NOR2_X1    g00157(.A1(new_n1139_), .A2(new_n1155_), .ZN(new_n1160_));
  NAND2_X1   g00158(.A1(new_n1159_), .A2(new_n1136_), .ZN(new_n1161_));
  AOI22_X1   g00159(.A1(new_n1161_), .A2(new_n1155_), .B1(new_n1160_), .B2(new_n1159_), .ZN(new_n1162_));
  NAND2_X1   g00160(.A1(new_n1146_), .A2(\A[917] ), .ZN(new_n1163_));
  NOR2_X1    g00161(.A1(new_n1147_), .A2(new_n1151_), .ZN(new_n1164_));
  NAND2_X1   g00162(.A1(new_n1163_), .A2(new_n1144_), .ZN(new_n1165_));
  AOI22_X1   g00163(.A1(new_n1165_), .A2(new_n1151_), .B1(new_n1164_), .B2(new_n1163_), .ZN(new_n1166_));
  NOR2_X1    g00164(.A1(new_n1162_), .A2(new_n1166_), .ZN(new_n1167_));
  NAND3_X1   g00165(.A1(new_n1167_), .A2(new_n1154_), .A3(new_n1158_), .ZN(new_n1168_));
  NAND2_X1   g00166(.A1(new_n1150_), .A2(new_n1168_), .ZN(new_n1169_));
  INV_X1     g00167(.I(\A[909] ), .ZN(new_n1170_));
  INV_X1     g00168(.I(\A[907] ), .ZN(new_n1171_));
  NAND2_X1   g00169(.A1(new_n1171_), .A2(\A[908] ), .ZN(new_n1172_));
  NOR2_X1    g00170(.A1(new_n1171_), .A2(\A[908] ), .ZN(new_n1173_));
  NOR2_X1    g00171(.A1(new_n1173_), .A2(new_n1170_), .ZN(new_n1174_));
  INV_X1     g00172(.I(\A[908] ), .ZN(new_n1175_));
  NAND2_X1   g00173(.A1(new_n1175_), .A2(\A[907] ), .ZN(new_n1176_));
  NAND2_X1   g00174(.A1(new_n1172_), .A2(new_n1176_), .ZN(new_n1177_));
  AOI22_X1   g00175(.A1(new_n1177_), .A2(new_n1170_), .B1(new_n1174_), .B2(new_n1172_), .ZN(new_n1178_));
  INV_X1     g00176(.I(\A[912] ), .ZN(new_n1179_));
  INV_X1     g00177(.I(\A[910] ), .ZN(new_n1180_));
  NAND2_X1   g00178(.A1(new_n1180_), .A2(\A[911] ), .ZN(new_n1181_));
  INV_X1     g00179(.I(\A[911] ), .ZN(new_n1182_));
  AOI21_X1   g00180(.A1(\A[910] ), .A2(new_n1182_), .B(new_n1179_), .ZN(new_n1183_));
  NAND2_X1   g00181(.A1(new_n1182_), .A2(\A[910] ), .ZN(new_n1184_));
  NAND2_X1   g00182(.A1(new_n1181_), .A2(new_n1184_), .ZN(new_n1185_));
  AOI22_X1   g00183(.A1(new_n1185_), .A2(new_n1179_), .B1(new_n1181_), .B2(new_n1183_), .ZN(new_n1186_));
  XOR2_X1    g00184(.A1(new_n1178_), .A2(new_n1186_), .Z(new_n1187_));
  AND2_X2    g00185(.A1(new_n1181_), .A2(new_n1184_), .Z(new_n1188_));
  NOR2_X1    g00186(.A1(new_n1180_), .A2(new_n1182_), .ZN(new_n1189_));
  INV_X1     g00187(.I(new_n1189_), .ZN(new_n1190_));
  OAI21_X1   g00188(.A1(new_n1188_), .A2(new_n1179_), .B(new_n1190_), .ZN(new_n1191_));
  NOR2_X1    g00189(.A1(new_n1175_), .A2(\A[907] ), .ZN(new_n1192_));
  NOR2_X1    g00190(.A1(new_n1192_), .A2(new_n1173_), .ZN(new_n1193_));
  NOR2_X1    g00191(.A1(new_n1171_), .A2(new_n1175_), .ZN(new_n1194_));
  INV_X1     g00192(.I(new_n1194_), .ZN(new_n1195_));
  OAI21_X1   g00193(.A1(new_n1193_), .A2(new_n1170_), .B(new_n1195_), .ZN(new_n1196_));
  NOR2_X1    g00194(.A1(new_n1178_), .A2(new_n1186_), .ZN(new_n1197_));
  NAND3_X1   g00195(.A1(new_n1197_), .A2(new_n1191_), .A3(new_n1196_), .ZN(new_n1198_));
  NAND2_X1   g00196(.A1(new_n1187_), .A2(new_n1198_), .ZN(new_n1199_));
  XOR2_X1    g00197(.A1(new_n1169_), .A2(new_n1199_), .Z(new_n1200_));
  INV_X1     g00198(.I(\A[903] ), .ZN(new_n1201_));
  INV_X1     g00199(.I(\A[901] ), .ZN(new_n1202_));
  NAND2_X1   g00200(.A1(new_n1202_), .A2(\A[902] ), .ZN(new_n1203_));
  NOR2_X1    g00201(.A1(new_n1202_), .A2(\A[902] ), .ZN(new_n1204_));
  NOR2_X1    g00202(.A1(new_n1204_), .A2(new_n1201_), .ZN(new_n1205_));
  INV_X1     g00203(.I(\A[902] ), .ZN(new_n1206_));
  NAND2_X1   g00204(.A1(new_n1206_), .A2(\A[901] ), .ZN(new_n1207_));
  NAND2_X1   g00205(.A1(new_n1203_), .A2(new_n1207_), .ZN(new_n1208_));
  AOI22_X1   g00206(.A1(new_n1208_), .A2(new_n1201_), .B1(new_n1205_), .B2(new_n1203_), .ZN(new_n1209_));
  INV_X1     g00207(.I(\A[906] ), .ZN(new_n1210_));
  INV_X1     g00208(.I(\A[904] ), .ZN(new_n1211_));
  NAND2_X1   g00209(.A1(new_n1211_), .A2(\A[905] ), .ZN(new_n1212_));
  NOR2_X1    g00210(.A1(new_n1211_), .A2(\A[905] ), .ZN(new_n1213_));
  NOR2_X1    g00211(.A1(new_n1213_), .A2(new_n1210_), .ZN(new_n1214_));
  INV_X1     g00212(.I(\A[905] ), .ZN(new_n1215_));
  NAND2_X1   g00213(.A1(new_n1215_), .A2(\A[904] ), .ZN(new_n1216_));
  NAND2_X1   g00214(.A1(new_n1212_), .A2(new_n1216_), .ZN(new_n1217_));
  AOI22_X1   g00215(.A1(new_n1217_), .A2(new_n1210_), .B1(new_n1214_), .B2(new_n1212_), .ZN(new_n1218_));
  XOR2_X1    g00216(.A1(new_n1209_), .A2(new_n1218_), .Z(new_n1219_));
  NOR2_X1    g00217(.A1(new_n1215_), .A2(\A[904] ), .ZN(new_n1220_));
  NOR2_X1    g00218(.A1(new_n1220_), .A2(new_n1213_), .ZN(new_n1221_));
  NOR2_X1    g00219(.A1(new_n1211_), .A2(new_n1215_), .ZN(new_n1222_));
  INV_X1     g00220(.I(new_n1222_), .ZN(new_n1223_));
  OAI21_X1   g00221(.A1(new_n1221_), .A2(new_n1210_), .B(new_n1223_), .ZN(new_n1224_));
  NOR2_X1    g00222(.A1(new_n1206_), .A2(\A[901] ), .ZN(new_n1225_));
  NOR2_X1    g00223(.A1(new_n1225_), .A2(new_n1204_), .ZN(new_n1226_));
  NOR2_X1    g00224(.A1(new_n1202_), .A2(new_n1206_), .ZN(new_n1227_));
  INV_X1     g00225(.I(new_n1227_), .ZN(new_n1228_));
  OAI21_X1   g00226(.A1(new_n1226_), .A2(new_n1201_), .B(new_n1228_), .ZN(new_n1229_));
  NOR2_X1    g00227(.A1(new_n1209_), .A2(new_n1218_), .ZN(new_n1230_));
  NAND3_X1   g00228(.A1(new_n1230_), .A2(new_n1224_), .A3(new_n1229_), .ZN(new_n1231_));
  NAND2_X1   g00229(.A1(new_n1219_), .A2(new_n1231_), .ZN(new_n1232_));
  INV_X1     g00230(.I(\A[897] ), .ZN(new_n1233_));
  INV_X1     g00231(.I(\A[895] ), .ZN(new_n1234_));
  NAND2_X1   g00232(.A1(new_n1234_), .A2(\A[896] ), .ZN(new_n1235_));
  NOR2_X1    g00233(.A1(new_n1234_), .A2(\A[896] ), .ZN(new_n1236_));
  NOR2_X1    g00234(.A1(new_n1236_), .A2(new_n1233_), .ZN(new_n1237_));
  INV_X1     g00235(.I(\A[896] ), .ZN(new_n1238_));
  NAND2_X1   g00236(.A1(new_n1238_), .A2(\A[895] ), .ZN(new_n1239_));
  NAND2_X1   g00237(.A1(new_n1235_), .A2(new_n1239_), .ZN(new_n1240_));
  AOI22_X1   g00238(.A1(new_n1240_), .A2(new_n1233_), .B1(new_n1237_), .B2(new_n1235_), .ZN(new_n1241_));
  INV_X1     g00239(.I(\A[900] ), .ZN(new_n1242_));
  INV_X1     g00240(.I(\A[898] ), .ZN(new_n1243_));
  NAND2_X1   g00241(.A1(new_n1243_), .A2(\A[899] ), .ZN(new_n1244_));
  INV_X1     g00242(.I(\A[899] ), .ZN(new_n1245_));
  AOI21_X1   g00243(.A1(\A[898] ), .A2(new_n1245_), .B(new_n1242_), .ZN(new_n1246_));
  NAND2_X1   g00244(.A1(new_n1245_), .A2(\A[898] ), .ZN(new_n1247_));
  NAND2_X1   g00245(.A1(new_n1244_), .A2(new_n1247_), .ZN(new_n1248_));
  AOI22_X1   g00246(.A1(new_n1248_), .A2(new_n1242_), .B1(new_n1244_), .B2(new_n1246_), .ZN(new_n1249_));
  XOR2_X1    g00247(.A1(new_n1241_), .A2(new_n1249_), .Z(new_n1250_));
  XNOR2_X1   g00248(.A1(\A[898] ), .A2(\A[899] ), .ZN(new_n1251_));
  NOR2_X1    g00249(.A1(new_n1243_), .A2(new_n1245_), .ZN(new_n1252_));
  INV_X1     g00250(.I(new_n1252_), .ZN(new_n1253_));
  OAI21_X1   g00251(.A1(new_n1251_), .A2(new_n1242_), .B(new_n1253_), .ZN(new_n1254_));
  NOR2_X1    g00252(.A1(new_n1238_), .A2(\A[895] ), .ZN(new_n1255_));
  NOR2_X1    g00253(.A1(new_n1255_), .A2(new_n1236_), .ZN(new_n1256_));
  NOR2_X1    g00254(.A1(new_n1234_), .A2(new_n1238_), .ZN(new_n1257_));
  INV_X1     g00255(.I(new_n1257_), .ZN(new_n1258_));
  OAI21_X1   g00256(.A1(new_n1256_), .A2(new_n1233_), .B(new_n1258_), .ZN(new_n1259_));
  NOR2_X1    g00257(.A1(new_n1241_), .A2(new_n1249_), .ZN(new_n1260_));
  NAND3_X1   g00258(.A1(new_n1260_), .A2(new_n1254_), .A3(new_n1259_), .ZN(new_n1261_));
  NAND2_X1   g00259(.A1(new_n1250_), .A2(new_n1261_), .ZN(new_n1262_));
  XOR2_X1    g00260(.A1(new_n1232_), .A2(new_n1262_), .Z(new_n1263_));
  XOR2_X1    g00261(.A1(new_n1200_), .A2(new_n1263_), .Z(new_n1264_));
  XNOR2_X1   g00262(.A1(new_n1133_), .A2(new_n1264_), .ZN(new_n1265_));
  INV_X1     g00263(.I(\A[890] ), .ZN(new_n1266_));
  NOR2_X1    g00264(.A1(new_n1266_), .A2(\A[889] ), .ZN(new_n1267_));
  NAND2_X1   g00265(.A1(new_n1266_), .A2(\A[889] ), .ZN(new_n1268_));
  NAND2_X1   g00266(.A1(new_n1268_), .A2(\A[891] ), .ZN(new_n1269_));
  INV_X1     g00267(.I(\A[889] ), .ZN(new_n1270_));
  NOR2_X1    g00268(.A1(new_n1270_), .A2(\A[890] ), .ZN(new_n1271_));
  NOR2_X1    g00269(.A1(new_n1267_), .A2(new_n1271_), .ZN(new_n1272_));
  OAI22_X1   g00270(.A1(new_n1272_), .A2(\A[891] ), .B1(new_n1269_), .B2(new_n1267_), .ZN(new_n1273_));
  INV_X1     g00271(.I(\A[893] ), .ZN(new_n1274_));
  NOR2_X1    g00272(.A1(new_n1274_), .A2(\A[892] ), .ZN(new_n1275_));
  NAND2_X1   g00273(.A1(new_n1274_), .A2(\A[892] ), .ZN(new_n1276_));
  NAND2_X1   g00274(.A1(new_n1276_), .A2(\A[894] ), .ZN(new_n1277_));
  INV_X1     g00275(.I(\A[892] ), .ZN(new_n1278_));
  NOR2_X1    g00276(.A1(new_n1278_), .A2(\A[893] ), .ZN(new_n1279_));
  NOR2_X1    g00277(.A1(new_n1275_), .A2(new_n1279_), .ZN(new_n1280_));
  OAI22_X1   g00278(.A1(new_n1280_), .A2(\A[894] ), .B1(new_n1277_), .B2(new_n1275_), .ZN(new_n1281_));
  XOR2_X1    g00279(.A1(new_n1273_), .A2(new_n1281_), .Z(new_n1282_));
  INV_X1     g00280(.I(\A[894] ), .ZN(new_n1283_));
  NOR2_X1    g00281(.A1(new_n1278_), .A2(new_n1274_), .ZN(new_n1284_));
  INV_X1     g00282(.I(new_n1284_), .ZN(new_n1285_));
  OAI21_X1   g00283(.A1(new_n1280_), .A2(new_n1283_), .B(new_n1285_), .ZN(new_n1286_));
  INV_X1     g00284(.I(\A[891] ), .ZN(new_n1287_));
  NOR2_X1    g00285(.A1(new_n1270_), .A2(new_n1266_), .ZN(new_n1288_));
  INV_X1     g00286(.I(new_n1288_), .ZN(new_n1289_));
  OAI21_X1   g00287(.A1(new_n1272_), .A2(new_n1287_), .B(new_n1289_), .ZN(new_n1290_));
  NAND2_X1   g00288(.A1(new_n1270_), .A2(\A[890] ), .ZN(new_n1291_));
  NOR2_X1    g00289(.A1(new_n1271_), .A2(new_n1287_), .ZN(new_n1292_));
  NAND2_X1   g00290(.A1(new_n1291_), .A2(new_n1268_), .ZN(new_n1293_));
  AOI22_X1   g00291(.A1(new_n1293_), .A2(new_n1287_), .B1(new_n1292_), .B2(new_n1291_), .ZN(new_n1294_));
  NAND2_X1   g00292(.A1(new_n1278_), .A2(\A[893] ), .ZN(new_n1295_));
  NOR2_X1    g00293(.A1(new_n1279_), .A2(new_n1283_), .ZN(new_n1296_));
  NAND2_X1   g00294(.A1(new_n1295_), .A2(new_n1276_), .ZN(new_n1297_));
  AOI22_X1   g00295(.A1(new_n1297_), .A2(new_n1283_), .B1(new_n1296_), .B2(new_n1295_), .ZN(new_n1298_));
  NOR2_X1    g00296(.A1(new_n1294_), .A2(new_n1298_), .ZN(new_n1299_));
  NAND3_X1   g00297(.A1(new_n1299_), .A2(new_n1286_), .A3(new_n1290_), .ZN(new_n1300_));
  NAND2_X1   g00298(.A1(new_n1282_), .A2(new_n1300_), .ZN(new_n1301_));
  INV_X1     g00299(.I(\A[885] ), .ZN(new_n1302_));
  INV_X1     g00300(.I(\A[883] ), .ZN(new_n1303_));
  NAND2_X1   g00301(.A1(new_n1303_), .A2(\A[884] ), .ZN(new_n1304_));
  NOR2_X1    g00302(.A1(new_n1303_), .A2(\A[884] ), .ZN(new_n1305_));
  NOR2_X1    g00303(.A1(new_n1305_), .A2(new_n1302_), .ZN(new_n1306_));
  INV_X1     g00304(.I(\A[884] ), .ZN(new_n1307_));
  NAND2_X1   g00305(.A1(new_n1307_), .A2(\A[883] ), .ZN(new_n1308_));
  NAND2_X1   g00306(.A1(new_n1304_), .A2(new_n1308_), .ZN(new_n1309_));
  AOI22_X1   g00307(.A1(new_n1309_), .A2(new_n1302_), .B1(new_n1306_), .B2(new_n1304_), .ZN(new_n1310_));
  INV_X1     g00308(.I(\A[888] ), .ZN(new_n1311_));
  INV_X1     g00309(.I(\A[886] ), .ZN(new_n1312_));
  NAND2_X1   g00310(.A1(new_n1312_), .A2(\A[887] ), .ZN(new_n1313_));
  INV_X1     g00311(.I(\A[887] ), .ZN(new_n1314_));
  AOI21_X1   g00312(.A1(\A[886] ), .A2(new_n1314_), .B(new_n1311_), .ZN(new_n1315_));
  NAND2_X1   g00313(.A1(new_n1314_), .A2(\A[886] ), .ZN(new_n1316_));
  NAND2_X1   g00314(.A1(new_n1313_), .A2(new_n1316_), .ZN(new_n1317_));
  AOI22_X1   g00315(.A1(new_n1317_), .A2(new_n1311_), .B1(new_n1313_), .B2(new_n1315_), .ZN(new_n1318_));
  XOR2_X1    g00316(.A1(new_n1310_), .A2(new_n1318_), .Z(new_n1319_));
  XNOR2_X1   g00317(.A1(\A[886] ), .A2(\A[887] ), .ZN(new_n1320_));
  NOR2_X1    g00318(.A1(new_n1312_), .A2(new_n1314_), .ZN(new_n1321_));
  INV_X1     g00319(.I(new_n1321_), .ZN(new_n1322_));
  OAI21_X1   g00320(.A1(new_n1320_), .A2(new_n1311_), .B(new_n1322_), .ZN(new_n1323_));
  NOR2_X1    g00321(.A1(new_n1307_), .A2(\A[883] ), .ZN(new_n1324_));
  NOR2_X1    g00322(.A1(new_n1324_), .A2(new_n1305_), .ZN(new_n1325_));
  NOR2_X1    g00323(.A1(new_n1303_), .A2(new_n1307_), .ZN(new_n1326_));
  INV_X1     g00324(.I(new_n1326_), .ZN(new_n1327_));
  OAI21_X1   g00325(.A1(new_n1325_), .A2(new_n1302_), .B(new_n1327_), .ZN(new_n1328_));
  NOR2_X1    g00326(.A1(new_n1310_), .A2(new_n1318_), .ZN(new_n1329_));
  NAND3_X1   g00327(.A1(new_n1329_), .A2(new_n1323_), .A3(new_n1328_), .ZN(new_n1330_));
  NAND2_X1   g00328(.A1(new_n1319_), .A2(new_n1330_), .ZN(new_n1331_));
  XOR2_X1    g00329(.A1(new_n1301_), .A2(new_n1331_), .Z(new_n1332_));
  INV_X1     g00330(.I(\A[879] ), .ZN(new_n1333_));
  INV_X1     g00331(.I(\A[877] ), .ZN(new_n1334_));
  NAND2_X1   g00332(.A1(new_n1334_), .A2(\A[878] ), .ZN(new_n1335_));
  NOR2_X1    g00333(.A1(new_n1334_), .A2(\A[878] ), .ZN(new_n1336_));
  NOR2_X1    g00334(.A1(new_n1336_), .A2(new_n1333_), .ZN(new_n1337_));
  INV_X1     g00335(.I(\A[878] ), .ZN(new_n1338_));
  NAND2_X1   g00336(.A1(new_n1338_), .A2(\A[877] ), .ZN(new_n1339_));
  NAND2_X1   g00337(.A1(new_n1335_), .A2(new_n1339_), .ZN(new_n1340_));
  AOI22_X1   g00338(.A1(new_n1340_), .A2(new_n1333_), .B1(new_n1337_), .B2(new_n1335_), .ZN(new_n1341_));
  INV_X1     g00339(.I(\A[882] ), .ZN(new_n1342_));
  INV_X1     g00340(.I(\A[880] ), .ZN(new_n1343_));
  NAND2_X1   g00341(.A1(new_n1343_), .A2(\A[881] ), .ZN(new_n1344_));
  INV_X1     g00342(.I(\A[881] ), .ZN(new_n1345_));
  AOI21_X1   g00343(.A1(\A[880] ), .A2(new_n1345_), .B(new_n1342_), .ZN(new_n1346_));
  NAND2_X1   g00344(.A1(new_n1345_), .A2(\A[880] ), .ZN(new_n1347_));
  NAND2_X1   g00345(.A1(new_n1344_), .A2(new_n1347_), .ZN(new_n1348_));
  AOI22_X1   g00346(.A1(new_n1348_), .A2(new_n1342_), .B1(new_n1344_), .B2(new_n1346_), .ZN(new_n1349_));
  XOR2_X1    g00347(.A1(new_n1341_), .A2(new_n1349_), .Z(new_n1350_));
  XNOR2_X1   g00348(.A1(\A[880] ), .A2(\A[881] ), .ZN(new_n1351_));
  NOR2_X1    g00349(.A1(new_n1343_), .A2(new_n1345_), .ZN(new_n1352_));
  INV_X1     g00350(.I(new_n1352_), .ZN(new_n1353_));
  OAI21_X1   g00351(.A1(new_n1351_), .A2(new_n1342_), .B(new_n1353_), .ZN(new_n1354_));
  NOR2_X1    g00352(.A1(new_n1338_), .A2(\A[877] ), .ZN(new_n1355_));
  NOR2_X1    g00353(.A1(new_n1355_), .A2(new_n1336_), .ZN(new_n1356_));
  NOR2_X1    g00354(.A1(new_n1334_), .A2(new_n1338_), .ZN(new_n1357_));
  INV_X1     g00355(.I(new_n1357_), .ZN(new_n1358_));
  OAI21_X1   g00356(.A1(new_n1356_), .A2(new_n1333_), .B(new_n1358_), .ZN(new_n1359_));
  NOR2_X1    g00357(.A1(new_n1341_), .A2(new_n1349_), .ZN(new_n1360_));
  NAND3_X1   g00358(.A1(new_n1360_), .A2(new_n1354_), .A3(new_n1359_), .ZN(new_n1361_));
  NAND2_X1   g00359(.A1(new_n1350_), .A2(new_n1361_), .ZN(new_n1362_));
  INV_X1     g00360(.I(\A[873] ), .ZN(new_n1363_));
  INV_X1     g00361(.I(\A[871] ), .ZN(new_n1364_));
  NAND2_X1   g00362(.A1(new_n1364_), .A2(\A[872] ), .ZN(new_n1365_));
  NOR2_X1    g00363(.A1(new_n1364_), .A2(\A[872] ), .ZN(new_n1366_));
  NOR2_X1    g00364(.A1(new_n1366_), .A2(new_n1363_), .ZN(new_n1367_));
  INV_X1     g00365(.I(\A[872] ), .ZN(new_n1368_));
  NAND2_X1   g00366(.A1(new_n1368_), .A2(\A[871] ), .ZN(new_n1369_));
  NAND2_X1   g00367(.A1(new_n1365_), .A2(new_n1369_), .ZN(new_n1370_));
  AOI22_X1   g00368(.A1(new_n1370_), .A2(new_n1363_), .B1(new_n1367_), .B2(new_n1365_), .ZN(new_n1371_));
  INV_X1     g00369(.I(\A[876] ), .ZN(new_n1372_));
  INV_X1     g00370(.I(\A[874] ), .ZN(new_n1373_));
  NAND2_X1   g00371(.A1(new_n1373_), .A2(\A[875] ), .ZN(new_n1374_));
  INV_X1     g00372(.I(\A[875] ), .ZN(new_n1375_));
  AOI21_X1   g00373(.A1(\A[874] ), .A2(new_n1375_), .B(new_n1372_), .ZN(new_n1376_));
  NAND2_X1   g00374(.A1(new_n1375_), .A2(\A[874] ), .ZN(new_n1377_));
  NAND2_X1   g00375(.A1(new_n1374_), .A2(new_n1377_), .ZN(new_n1378_));
  AOI22_X1   g00376(.A1(new_n1378_), .A2(new_n1372_), .B1(new_n1374_), .B2(new_n1376_), .ZN(new_n1379_));
  XOR2_X1    g00377(.A1(new_n1371_), .A2(new_n1379_), .Z(new_n1380_));
  XNOR2_X1   g00378(.A1(\A[874] ), .A2(\A[875] ), .ZN(new_n1381_));
  NOR2_X1    g00379(.A1(new_n1373_), .A2(new_n1375_), .ZN(new_n1382_));
  INV_X1     g00380(.I(new_n1382_), .ZN(new_n1383_));
  OAI21_X1   g00381(.A1(new_n1381_), .A2(new_n1372_), .B(new_n1383_), .ZN(new_n1384_));
  NOR2_X1    g00382(.A1(new_n1368_), .A2(\A[871] ), .ZN(new_n1385_));
  NOR2_X1    g00383(.A1(new_n1385_), .A2(new_n1366_), .ZN(new_n1386_));
  NOR2_X1    g00384(.A1(new_n1364_), .A2(new_n1368_), .ZN(new_n1387_));
  INV_X1     g00385(.I(new_n1387_), .ZN(new_n1388_));
  OAI21_X1   g00386(.A1(new_n1386_), .A2(new_n1363_), .B(new_n1388_), .ZN(new_n1389_));
  NOR2_X1    g00387(.A1(new_n1371_), .A2(new_n1379_), .ZN(new_n1390_));
  NAND3_X1   g00388(.A1(new_n1390_), .A2(new_n1384_), .A3(new_n1389_), .ZN(new_n1391_));
  NAND2_X1   g00389(.A1(new_n1380_), .A2(new_n1391_), .ZN(new_n1392_));
  XOR2_X1    g00390(.A1(new_n1362_), .A2(new_n1392_), .Z(new_n1393_));
  XOR2_X1    g00391(.A1(new_n1332_), .A2(new_n1393_), .Z(new_n1394_));
  INV_X1     g00392(.I(\A[867] ), .ZN(new_n1395_));
  INV_X1     g00393(.I(\A[865] ), .ZN(new_n1396_));
  NAND2_X1   g00394(.A1(new_n1396_), .A2(\A[866] ), .ZN(new_n1397_));
  NOR2_X1    g00395(.A1(new_n1396_), .A2(\A[866] ), .ZN(new_n1398_));
  NOR2_X1    g00396(.A1(new_n1398_), .A2(new_n1395_), .ZN(new_n1399_));
  INV_X1     g00397(.I(\A[866] ), .ZN(new_n1400_));
  NAND2_X1   g00398(.A1(new_n1400_), .A2(\A[865] ), .ZN(new_n1401_));
  NAND2_X1   g00399(.A1(new_n1397_), .A2(new_n1401_), .ZN(new_n1402_));
  AOI22_X1   g00400(.A1(new_n1402_), .A2(new_n1395_), .B1(new_n1399_), .B2(new_n1397_), .ZN(new_n1403_));
  INV_X1     g00401(.I(\A[870] ), .ZN(new_n1404_));
  INV_X1     g00402(.I(\A[868] ), .ZN(new_n1405_));
  NAND2_X1   g00403(.A1(new_n1405_), .A2(\A[869] ), .ZN(new_n1406_));
  NOR2_X1    g00404(.A1(new_n1405_), .A2(\A[869] ), .ZN(new_n1407_));
  NOR2_X1    g00405(.A1(new_n1407_), .A2(new_n1404_), .ZN(new_n1408_));
  INV_X1     g00406(.I(\A[869] ), .ZN(new_n1409_));
  NAND2_X1   g00407(.A1(new_n1409_), .A2(\A[868] ), .ZN(new_n1410_));
  NAND2_X1   g00408(.A1(new_n1406_), .A2(new_n1410_), .ZN(new_n1411_));
  AOI22_X1   g00409(.A1(new_n1411_), .A2(new_n1404_), .B1(new_n1408_), .B2(new_n1406_), .ZN(new_n1412_));
  XOR2_X1    g00410(.A1(new_n1403_), .A2(new_n1412_), .Z(new_n1413_));
  NOR2_X1    g00411(.A1(new_n1409_), .A2(\A[868] ), .ZN(new_n1414_));
  NOR2_X1    g00412(.A1(new_n1414_), .A2(new_n1407_), .ZN(new_n1415_));
  NOR2_X1    g00413(.A1(new_n1405_), .A2(new_n1409_), .ZN(new_n1416_));
  INV_X1     g00414(.I(new_n1416_), .ZN(new_n1417_));
  OAI21_X1   g00415(.A1(new_n1415_), .A2(new_n1404_), .B(new_n1417_), .ZN(new_n1418_));
  NOR2_X1    g00416(.A1(new_n1400_), .A2(\A[865] ), .ZN(new_n1419_));
  NOR2_X1    g00417(.A1(new_n1419_), .A2(new_n1398_), .ZN(new_n1420_));
  NOR2_X1    g00418(.A1(new_n1396_), .A2(new_n1400_), .ZN(new_n1421_));
  INV_X1     g00419(.I(new_n1421_), .ZN(new_n1422_));
  OAI21_X1   g00420(.A1(new_n1420_), .A2(new_n1395_), .B(new_n1422_), .ZN(new_n1423_));
  NOR2_X1    g00421(.A1(new_n1403_), .A2(new_n1412_), .ZN(new_n1424_));
  NAND3_X1   g00422(.A1(new_n1424_), .A2(new_n1418_), .A3(new_n1423_), .ZN(new_n1425_));
  NAND2_X1   g00423(.A1(new_n1413_), .A2(new_n1425_), .ZN(new_n1426_));
  INV_X1     g00424(.I(\A[861] ), .ZN(new_n1427_));
  INV_X1     g00425(.I(\A[859] ), .ZN(new_n1428_));
  NAND2_X1   g00426(.A1(new_n1428_), .A2(\A[860] ), .ZN(new_n1429_));
  NOR2_X1    g00427(.A1(new_n1428_), .A2(\A[860] ), .ZN(new_n1430_));
  NOR2_X1    g00428(.A1(new_n1430_), .A2(new_n1427_), .ZN(new_n1431_));
  INV_X1     g00429(.I(\A[860] ), .ZN(new_n1432_));
  NAND2_X1   g00430(.A1(new_n1432_), .A2(\A[859] ), .ZN(new_n1433_));
  NAND2_X1   g00431(.A1(new_n1429_), .A2(new_n1433_), .ZN(new_n1434_));
  AOI22_X1   g00432(.A1(new_n1434_), .A2(new_n1427_), .B1(new_n1431_), .B2(new_n1429_), .ZN(new_n1435_));
  INV_X1     g00433(.I(\A[864] ), .ZN(new_n1436_));
  INV_X1     g00434(.I(\A[862] ), .ZN(new_n1437_));
  NAND2_X1   g00435(.A1(new_n1437_), .A2(\A[863] ), .ZN(new_n1438_));
  INV_X1     g00436(.I(\A[863] ), .ZN(new_n1439_));
  AOI21_X1   g00437(.A1(\A[862] ), .A2(new_n1439_), .B(new_n1436_), .ZN(new_n1440_));
  NAND2_X1   g00438(.A1(new_n1439_), .A2(\A[862] ), .ZN(new_n1441_));
  NAND2_X1   g00439(.A1(new_n1438_), .A2(new_n1441_), .ZN(new_n1442_));
  AOI22_X1   g00440(.A1(new_n1442_), .A2(new_n1436_), .B1(new_n1438_), .B2(new_n1440_), .ZN(new_n1443_));
  XOR2_X1    g00441(.A1(new_n1435_), .A2(new_n1443_), .Z(new_n1444_));
  XNOR2_X1   g00442(.A1(\A[862] ), .A2(\A[863] ), .ZN(new_n1445_));
  NOR2_X1    g00443(.A1(new_n1437_), .A2(new_n1439_), .ZN(new_n1446_));
  INV_X1     g00444(.I(new_n1446_), .ZN(new_n1447_));
  OAI21_X1   g00445(.A1(new_n1445_), .A2(new_n1436_), .B(new_n1447_), .ZN(new_n1448_));
  NOR2_X1    g00446(.A1(new_n1432_), .A2(\A[859] ), .ZN(new_n1449_));
  NOR2_X1    g00447(.A1(new_n1449_), .A2(new_n1430_), .ZN(new_n1450_));
  NOR2_X1    g00448(.A1(new_n1428_), .A2(new_n1432_), .ZN(new_n1451_));
  INV_X1     g00449(.I(new_n1451_), .ZN(new_n1452_));
  OAI21_X1   g00450(.A1(new_n1450_), .A2(new_n1427_), .B(new_n1452_), .ZN(new_n1453_));
  NOR2_X1    g00451(.A1(new_n1435_), .A2(new_n1443_), .ZN(new_n1454_));
  NAND3_X1   g00452(.A1(new_n1454_), .A2(new_n1448_), .A3(new_n1453_), .ZN(new_n1455_));
  NAND2_X1   g00453(.A1(new_n1444_), .A2(new_n1455_), .ZN(new_n1456_));
  XOR2_X1    g00454(.A1(new_n1426_), .A2(new_n1456_), .Z(new_n1457_));
  INV_X1     g00455(.I(\A[855] ), .ZN(new_n1458_));
  INV_X1     g00456(.I(\A[853] ), .ZN(new_n1459_));
  NAND2_X1   g00457(.A1(new_n1459_), .A2(\A[854] ), .ZN(new_n1460_));
  NOR2_X1    g00458(.A1(new_n1459_), .A2(\A[854] ), .ZN(new_n1461_));
  NOR2_X1    g00459(.A1(new_n1461_), .A2(new_n1458_), .ZN(new_n1462_));
  INV_X1     g00460(.I(\A[854] ), .ZN(new_n1463_));
  NAND2_X1   g00461(.A1(new_n1463_), .A2(\A[853] ), .ZN(new_n1464_));
  NAND2_X1   g00462(.A1(new_n1460_), .A2(new_n1464_), .ZN(new_n1465_));
  AOI22_X1   g00463(.A1(new_n1465_), .A2(new_n1458_), .B1(new_n1462_), .B2(new_n1460_), .ZN(new_n1466_));
  INV_X1     g00464(.I(\A[858] ), .ZN(new_n1467_));
  INV_X1     g00465(.I(\A[856] ), .ZN(new_n1468_));
  NAND2_X1   g00466(.A1(new_n1468_), .A2(\A[857] ), .ZN(new_n1469_));
  NOR2_X1    g00467(.A1(new_n1468_), .A2(\A[857] ), .ZN(new_n1470_));
  NOR2_X1    g00468(.A1(new_n1470_), .A2(new_n1467_), .ZN(new_n1471_));
  INV_X1     g00469(.I(\A[857] ), .ZN(new_n1472_));
  NAND2_X1   g00470(.A1(new_n1472_), .A2(\A[856] ), .ZN(new_n1473_));
  NAND2_X1   g00471(.A1(new_n1469_), .A2(new_n1473_), .ZN(new_n1474_));
  AOI22_X1   g00472(.A1(new_n1474_), .A2(new_n1467_), .B1(new_n1471_), .B2(new_n1469_), .ZN(new_n1475_));
  XOR2_X1    g00473(.A1(new_n1466_), .A2(new_n1475_), .Z(new_n1476_));
  NOR2_X1    g00474(.A1(new_n1472_), .A2(\A[856] ), .ZN(new_n1477_));
  NOR2_X1    g00475(.A1(new_n1477_), .A2(new_n1470_), .ZN(new_n1478_));
  NOR2_X1    g00476(.A1(new_n1468_), .A2(new_n1472_), .ZN(new_n1479_));
  INV_X1     g00477(.I(new_n1479_), .ZN(new_n1480_));
  OAI21_X1   g00478(.A1(new_n1478_), .A2(new_n1467_), .B(new_n1480_), .ZN(new_n1481_));
  NOR2_X1    g00479(.A1(new_n1463_), .A2(\A[853] ), .ZN(new_n1482_));
  NOR2_X1    g00480(.A1(new_n1482_), .A2(new_n1461_), .ZN(new_n1483_));
  NOR2_X1    g00481(.A1(new_n1459_), .A2(new_n1463_), .ZN(new_n1484_));
  INV_X1     g00482(.I(new_n1484_), .ZN(new_n1485_));
  OAI21_X1   g00483(.A1(new_n1483_), .A2(new_n1458_), .B(new_n1485_), .ZN(new_n1486_));
  NOR2_X1    g00484(.A1(new_n1466_), .A2(new_n1475_), .ZN(new_n1487_));
  NAND3_X1   g00485(.A1(new_n1487_), .A2(new_n1481_), .A3(new_n1486_), .ZN(new_n1488_));
  NAND2_X1   g00486(.A1(new_n1476_), .A2(new_n1488_), .ZN(new_n1489_));
  INV_X1     g00487(.I(\A[849] ), .ZN(new_n1490_));
  INV_X1     g00488(.I(\A[847] ), .ZN(new_n1491_));
  NAND2_X1   g00489(.A1(new_n1491_), .A2(\A[848] ), .ZN(new_n1492_));
  NOR2_X1    g00490(.A1(new_n1491_), .A2(\A[848] ), .ZN(new_n1493_));
  NOR2_X1    g00491(.A1(new_n1493_), .A2(new_n1490_), .ZN(new_n1494_));
  INV_X1     g00492(.I(\A[848] ), .ZN(new_n1495_));
  NAND2_X1   g00493(.A1(new_n1495_), .A2(\A[847] ), .ZN(new_n1496_));
  NAND2_X1   g00494(.A1(new_n1492_), .A2(new_n1496_), .ZN(new_n1497_));
  AOI22_X1   g00495(.A1(new_n1497_), .A2(new_n1490_), .B1(new_n1494_), .B2(new_n1492_), .ZN(new_n1498_));
  INV_X1     g00496(.I(\A[852] ), .ZN(new_n1499_));
  INV_X1     g00497(.I(\A[850] ), .ZN(new_n1500_));
  NAND2_X1   g00498(.A1(new_n1500_), .A2(\A[851] ), .ZN(new_n1501_));
  INV_X1     g00499(.I(\A[851] ), .ZN(new_n1502_));
  AOI21_X1   g00500(.A1(\A[850] ), .A2(new_n1502_), .B(new_n1499_), .ZN(new_n1503_));
  NAND2_X1   g00501(.A1(new_n1502_), .A2(\A[850] ), .ZN(new_n1504_));
  NAND2_X1   g00502(.A1(new_n1501_), .A2(new_n1504_), .ZN(new_n1505_));
  AOI22_X1   g00503(.A1(new_n1505_), .A2(new_n1499_), .B1(new_n1501_), .B2(new_n1503_), .ZN(new_n1506_));
  XOR2_X1    g00504(.A1(new_n1498_), .A2(new_n1506_), .Z(new_n1507_));
  NOR2_X1    g00505(.A1(new_n1500_), .A2(new_n1502_), .ZN(new_n1508_));
  INV_X1     g00506(.I(new_n1508_), .ZN(new_n1509_));
  NAND2_X1   g00507(.A1(new_n1505_), .A2(\A[852] ), .ZN(new_n1510_));
  NAND2_X1   g00508(.A1(new_n1510_), .A2(new_n1509_), .ZN(new_n1511_));
  NOR2_X1    g00509(.A1(new_n1495_), .A2(\A[847] ), .ZN(new_n1512_));
  NOR2_X1    g00510(.A1(new_n1512_), .A2(new_n1493_), .ZN(new_n1513_));
  NOR2_X1    g00511(.A1(new_n1491_), .A2(new_n1495_), .ZN(new_n1514_));
  INV_X1     g00512(.I(new_n1514_), .ZN(new_n1515_));
  OAI21_X1   g00513(.A1(new_n1513_), .A2(new_n1490_), .B(new_n1515_), .ZN(new_n1516_));
  NOR2_X1    g00514(.A1(new_n1498_), .A2(new_n1506_), .ZN(new_n1517_));
  NAND3_X1   g00515(.A1(new_n1517_), .A2(new_n1511_), .A3(new_n1516_), .ZN(new_n1518_));
  NAND2_X1   g00516(.A1(new_n1507_), .A2(new_n1518_), .ZN(new_n1519_));
  XOR2_X1    g00517(.A1(new_n1489_), .A2(new_n1519_), .Z(new_n1520_));
  XOR2_X1    g00518(.A1(new_n1457_), .A2(new_n1520_), .Z(new_n1521_));
  XNOR2_X1   g00519(.A1(new_n1394_), .A2(new_n1521_), .ZN(new_n1522_));
  XNOR2_X1   g00520(.A1(new_n1265_), .A2(new_n1522_), .ZN(new_n1523_));
  INV_X1     g00521(.I(\A[988] ), .ZN(new_n1524_));
  INV_X1     g00522(.I(\A[989] ), .ZN(new_n1525_));
  NOR2_X1    g00523(.A1(new_n1524_), .A2(new_n1525_), .ZN(new_n1526_));
  NAND2_X1   g00524(.A1(new_n1525_), .A2(\A[988] ), .ZN(new_n1527_));
  NAND2_X1   g00525(.A1(new_n1524_), .A2(\A[989] ), .ZN(new_n1528_));
  NAND2_X1   g00526(.A1(new_n1527_), .A2(new_n1528_), .ZN(new_n1529_));
  AOI21_X1   g00527(.A1(new_n1529_), .A2(\A[990] ), .B(new_n1526_), .ZN(new_n1530_));
  INV_X1     g00528(.I(new_n1530_), .ZN(new_n1531_));
  INV_X1     g00529(.I(\A[985] ), .ZN(new_n1532_));
  INV_X1     g00530(.I(\A[986] ), .ZN(new_n1533_));
  NOR2_X1    g00531(.A1(new_n1532_), .A2(new_n1533_), .ZN(new_n1534_));
  NAND2_X1   g00532(.A1(new_n1533_), .A2(\A[985] ), .ZN(new_n1535_));
  NAND2_X1   g00533(.A1(new_n1532_), .A2(\A[986] ), .ZN(new_n1536_));
  NAND2_X1   g00534(.A1(new_n1535_), .A2(new_n1536_), .ZN(new_n1537_));
  AOI21_X1   g00535(.A1(new_n1537_), .A2(\A[987] ), .B(new_n1534_), .ZN(new_n1538_));
  INV_X1     g00536(.I(new_n1538_), .ZN(new_n1539_));
  INV_X1     g00537(.I(\A[987] ), .ZN(new_n1540_));
  AOI21_X1   g00538(.A1(\A[985] ), .A2(new_n1533_), .B(new_n1540_), .ZN(new_n1541_));
  AOI22_X1   g00539(.A1(new_n1537_), .A2(new_n1540_), .B1(new_n1536_), .B2(new_n1541_), .ZN(new_n1542_));
  INV_X1     g00540(.I(\A[990] ), .ZN(new_n1543_));
  AOI21_X1   g00541(.A1(\A[988] ), .A2(new_n1525_), .B(new_n1543_), .ZN(new_n1544_));
  AOI22_X1   g00542(.A1(new_n1529_), .A2(new_n1543_), .B1(new_n1528_), .B2(new_n1544_), .ZN(new_n1545_));
  NOR2_X1    g00543(.A1(new_n1542_), .A2(new_n1545_), .ZN(new_n1546_));
  NAND3_X1   g00544(.A1(new_n1546_), .A2(new_n1531_), .A3(new_n1539_), .ZN(new_n1547_));
  XOR2_X1    g00545(.A1(new_n1542_), .A2(new_n1545_), .Z(new_n1548_));
  NAND2_X1   g00546(.A1(new_n1548_), .A2(new_n1547_), .ZN(new_n1549_));
  INV_X1     g00547(.I(\A[981] ), .ZN(new_n1550_));
  INV_X1     g00548(.I(\A[979] ), .ZN(new_n1551_));
  NAND2_X1   g00549(.A1(new_n1551_), .A2(\A[980] ), .ZN(new_n1552_));
  INV_X1     g00550(.I(\A[980] ), .ZN(new_n1553_));
  NAND2_X1   g00551(.A1(new_n1553_), .A2(\A[979] ), .ZN(new_n1554_));
  NAND2_X1   g00552(.A1(new_n1554_), .A2(new_n1552_), .ZN(new_n1555_));
  AOI21_X1   g00553(.A1(\A[979] ), .A2(new_n1553_), .B(new_n1550_), .ZN(new_n1556_));
  AOI22_X1   g00554(.A1(new_n1555_), .A2(new_n1550_), .B1(new_n1552_), .B2(new_n1556_), .ZN(new_n1557_));
  INV_X1     g00555(.I(\A[984] ), .ZN(new_n1558_));
  INV_X1     g00556(.I(\A[982] ), .ZN(new_n1559_));
  NAND2_X1   g00557(.A1(new_n1559_), .A2(\A[983] ), .ZN(new_n1560_));
  INV_X1     g00558(.I(\A[983] ), .ZN(new_n1561_));
  NAND2_X1   g00559(.A1(new_n1561_), .A2(\A[982] ), .ZN(new_n1562_));
  NAND2_X1   g00560(.A1(new_n1562_), .A2(new_n1560_), .ZN(new_n1563_));
  AOI21_X1   g00561(.A1(\A[982] ), .A2(new_n1561_), .B(new_n1558_), .ZN(new_n1564_));
  AOI22_X1   g00562(.A1(new_n1563_), .A2(new_n1558_), .B1(new_n1560_), .B2(new_n1564_), .ZN(new_n1565_));
  XOR2_X1    g00563(.A1(new_n1557_), .A2(new_n1565_), .Z(new_n1566_));
  NOR2_X1    g00564(.A1(new_n1559_), .A2(new_n1561_), .ZN(new_n1567_));
  AOI21_X1   g00565(.A1(new_n1563_), .A2(\A[984] ), .B(new_n1567_), .ZN(new_n1568_));
  NOR2_X1    g00566(.A1(new_n1551_), .A2(new_n1553_), .ZN(new_n1569_));
  AOI21_X1   g00567(.A1(new_n1555_), .A2(\A[981] ), .B(new_n1569_), .ZN(new_n1570_));
  OR4_X2     g00568(.A1(new_n1557_), .A2(new_n1565_), .A3(new_n1568_), .A4(new_n1570_), .Z(new_n1571_));
  NAND2_X1   g00569(.A1(new_n1566_), .A2(new_n1571_), .ZN(new_n1572_));
  XOR2_X1    g00570(.A1(new_n1572_), .A2(new_n1549_), .Z(new_n1573_));
  INV_X1     g00571(.I(\A[976] ), .ZN(new_n1574_));
  INV_X1     g00572(.I(\A[977] ), .ZN(new_n1575_));
  NOR2_X1    g00573(.A1(new_n1574_), .A2(new_n1575_), .ZN(new_n1576_));
  NAND2_X1   g00574(.A1(new_n1575_), .A2(\A[976] ), .ZN(new_n1577_));
  NAND2_X1   g00575(.A1(new_n1574_), .A2(\A[977] ), .ZN(new_n1578_));
  NAND2_X1   g00576(.A1(new_n1577_), .A2(new_n1578_), .ZN(new_n1579_));
  AOI21_X1   g00577(.A1(new_n1579_), .A2(\A[978] ), .B(new_n1576_), .ZN(new_n1580_));
  INV_X1     g00578(.I(new_n1580_), .ZN(new_n1581_));
  INV_X1     g00579(.I(\A[973] ), .ZN(new_n1582_));
  INV_X1     g00580(.I(\A[974] ), .ZN(new_n1583_));
  NOR2_X1    g00581(.A1(new_n1582_), .A2(new_n1583_), .ZN(new_n1584_));
  NAND2_X1   g00582(.A1(new_n1583_), .A2(\A[973] ), .ZN(new_n1585_));
  NAND2_X1   g00583(.A1(new_n1582_), .A2(\A[974] ), .ZN(new_n1586_));
  NAND2_X1   g00584(.A1(new_n1585_), .A2(new_n1586_), .ZN(new_n1587_));
  AOI21_X1   g00585(.A1(new_n1587_), .A2(\A[975] ), .B(new_n1584_), .ZN(new_n1588_));
  INV_X1     g00586(.I(new_n1588_), .ZN(new_n1589_));
  INV_X1     g00587(.I(\A[975] ), .ZN(new_n1590_));
  AOI21_X1   g00588(.A1(\A[973] ), .A2(new_n1583_), .B(new_n1590_), .ZN(new_n1591_));
  AOI22_X1   g00589(.A1(new_n1587_), .A2(new_n1590_), .B1(new_n1586_), .B2(new_n1591_), .ZN(new_n1592_));
  INV_X1     g00590(.I(\A[978] ), .ZN(new_n1593_));
  AOI21_X1   g00591(.A1(\A[976] ), .A2(new_n1575_), .B(new_n1593_), .ZN(new_n1594_));
  AOI22_X1   g00592(.A1(new_n1579_), .A2(new_n1593_), .B1(new_n1578_), .B2(new_n1594_), .ZN(new_n1595_));
  NOR2_X1    g00593(.A1(new_n1592_), .A2(new_n1595_), .ZN(new_n1596_));
  NAND3_X1   g00594(.A1(new_n1596_), .A2(new_n1581_), .A3(new_n1589_), .ZN(new_n1597_));
  XOR2_X1    g00595(.A1(new_n1592_), .A2(new_n1595_), .Z(new_n1598_));
  NAND2_X1   g00596(.A1(new_n1598_), .A2(new_n1597_), .ZN(new_n1599_));
  INV_X1     g00597(.I(\A[969] ), .ZN(new_n1600_));
  INV_X1     g00598(.I(\A[967] ), .ZN(new_n1601_));
  NAND2_X1   g00599(.A1(new_n1601_), .A2(\A[968] ), .ZN(new_n1602_));
  INV_X1     g00600(.I(\A[968] ), .ZN(new_n1603_));
  NAND2_X1   g00601(.A1(new_n1603_), .A2(\A[967] ), .ZN(new_n1604_));
  NAND2_X1   g00602(.A1(new_n1604_), .A2(new_n1602_), .ZN(new_n1605_));
  AOI21_X1   g00603(.A1(\A[967] ), .A2(new_n1603_), .B(new_n1600_), .ZN(new_n1606_));
  AOI22_X1   g00604(.A1(new_n1605_), .A2(new_n1600_), .B1(new_n1602_), .B2(new_n1606_), .ZN(new_n1607_));
  INV_X1     g00605(.I(\A[972] ), .ZN(new_n1608_));
  INV_X1     g00606(.I(\A[970] ), .ZN(new_n1609_));
  NAND2_X1   g00607(.A1(new_n1609_), .A2(\A[971] ), .ZN(new_n1610_));
  INV_X1     g00608(.I(\A[971] ), .ZN(new_n1611_));
  NAND2_X1   g00609(.A1(new_n1611_), .A2(\A[970] ), .ZN(new_n1612_));
  NAND2_X1   g00610(.A1(new_n1612_), .A2(new_n1610_), .ZN(new_n1613_));
  AOI21_X1   g00611(.A1(\A[970] ), .A2(new_n1611_), .B(new_n1608_), .ZN(new_n1614_));
  AOI22_X1   g00612(.A1(new_n1613_), .A2(new_n1608_), .B1(new_n1610_), .B2(new_n1614_), .ZN(new_n1615_));
  XOR2_X1    g00613(.A1(new_n1607_), .A2(new_n1615_), .Z(new_n1616_));
  NOR2_X1    g00614(.A1(new_n1609_), .A2(new_n1611_), .ZN(new_n1617_));
  AOI21_X1   g00615(.A1(new_n1613_), .A2(\A[972] ), .B(new_n1617_), .ZN(new_n1618_));
  NOR2_X1    g00616(.A1(new_n1601_), .A2(new_n1603_), .ZN(new_n1619_));
  AOI21_X1   g00617(.A1(new_n1605_), .A2(\A[969] ), .B(new_n1619_), .ZN(new_n1620_));
  OR4_X2     g00618(.A1(new_n1607_), .A2(new_n1615_), .A3(new_n1618_), .A4(new_n1620_), .Z(new_n1621_));
  NAND2_X1   g00619(.A1(new_n1616_), .A2(new_n1621_), .ZN(new_n1622_));
  XOR2_X1    g00620(.A1(new_n1622_), .A2(new_n1599_), .Z(new_n1623_));
  XNOR2_X1   g00621(.A1(new_n1573_), .A2(new_n1623_), .ZN(new_n1624_));
  INV_X1     g00622(.I(\A[963] ), .ZN(new_n1625_));
  INV_X1     g00623(.I(\A[961] ), .ZN(new_n1626_));
  NAND2_X1   g00624(.A1(new_n1626_), .A2(\A[962] ), .ZN(new_n1627_));
  NOR2_X1    g00625(.A1(new_n1626_), .A2(\A[962] ), .ZN(new_n1628_));
  NOR2_X1    g00626(.A1(new_n1628_), .A2(new_n1625_), .ZN(new_n1629_));
  INV_X1     g00627(.I(\A[962] ), .ZN(new_n1630_));
  NAND2_X1   g00628(.A1(new_n1630_), .A2(\A[961] ), .ZN(new_n1631_));
  NAND2_X1   g00629(.A1(new_n1627_), .A2(new_n1631_), .ZN(new_n1632_));
  AOI22_X1   g00630(.A1(new_n1632_), .A2(new_n1625_), .B1(new_n1629_), .B2(new_n1627_), .ZN(new_n1633_));
  INV_X1     g00631(.I(\A[966] ), .ZN(new_n1634_));
  INV_X1     g00632(.I(\A[964] ), .ZN(new_n1635_));
  NAND2_X1   g00633(.A1(new_n1635_), .A2(\A[965] ), .ZN(new_n1636_));
  NOR2_X1    g00634(.A1(new_n1635_), .A2(\A[965] ), .ZN(new_n1637_));
  NOR2_X1    g00635(.A1(new_n1637_), .A2(new_n1634_), .ZN(new_n1638_));
  INV_X1     g00636(.I(\A[965] ), .ZN(new_n1639_));
  NAND2_X1   g00637(.A1(new_n1639_), .A2(\A[964] ), .ZN(new_n1640_));
  NAND2_X1   g00638(.A1(new_n1636_), .A2(new_n1640_), .ZN(new_n1641_));
  AOI22_X1   g00639(.A1(new_n1641_), .A2(new_n1634_), .B1(new_n1638_), .B2(new_n1636_), .ZN(new_n1642_));
  XOR2_X1    g00640(.A1(new_n1633_), .A2(new_n1642_), .Z(new_n1643_));
  NOR2_X1    g00641(.A1(new_n1635_), .A2(new_n1639_), .ZN(new_n1644_));
  AOI21_X1   g00642(.A1(new_n1641_), .A2(\A[966] ), .B(new_n1644_), .ZN(new_n1645_));
  NOR2_X1    g00643(.A1(new_n1626_), .A2(new_n1630_), .ZN(new_n1646_));
  AOI21_X1   g00644(.A1(new_n1632_), .A2(\A[963] ), .B(new_n1646_), .ZN(new_n1647_));
  OR4_X2     g00645(.A1(new_n1633_), .A2(new_n1642_), .A3(new_n1645_), .A4(new_n1647_), .Z(new_n1648_));
  NAND2_X1   g00646(.A1(new_n1643_), .A2(new_n1648_), .ZN(new_n1649_));
  INV_X1     g00647(.I(\A[957] ), .ZN(new_n1650_));
  INV_X1     g00648(.I(\A[955] ), .ZN(new_n1651_));
  NAND2_X1   g00649(.A1(new_n1651_), .A2(\A[956] ), .ZN(new_n1652_));
  INV_X1     g00650(.I(\A[956] ), .ZN(new_n1653_));
  AOI21_X1   g00651(.A1(\A[955] ), .A2(new_n1653_), .B(new_n1650_), .ZN(new_n1654_));
  NAND2_X1   g00652(.A1(new_n1653_), .A2(\A[955] ), .ZN(new_n1655_));
  NAND2_X1   g00653(.A1(new_n1652_), .A2(new_n1655_), .ZN(new_n1656_));
  AOI22_X1   g00654(.A1(new_n1656_), .A2(new_n1650_), .B1(new_n1654_), .B2(new_n1652_), .ZN(new_n1657_));
  INV_X1     g00655(.I(\A[960] ), .ZN(new_n1658_));
  INV_X1     g00656(.I(\A[958] ), .ZN(new_n1659_));
  NAND2_X1   g00657(.A1(new_n1659_), .A2(\A[959] ), .ZN(new_n1660_));
  NOR2_X1    g00658(.A1(new_n1659_), .A2(\A[959] ), .ZN(new_n1661_));
  NOR2_X1    g00659(.A1(new_n1661_), .A2(new_n1658_), .ZN(new_n1662_));
  INV_X1     g00660(.I(\A[959] ), .ZN(new_n1663_));
  NAND2_X1   g00661(.A1(new_n1663_), .A2(\A[958] ), .ZN(new_n1664_));
  NAND2_X1   g00662(.A1(new_n1660_), .A2(new_n1664_), .ZN(new_n1665_));
  AOI22_X1   g00663(.A1(new_n1665_), .A2(new_n1658_), .B1(new_n1662_), .B2(new_n1660_), .ZN(new_n1666_));
  XOR2_X1    g00664(.A1(new_n1666_), .A2(new_n1657_), .Z(new_n1667_));
  NOR2_X1    g00665(.A1(new_n1659_), .A2(new_n1663_), .ZN(new_n1668_));
  AOI21_X1   g00666(.A1(new_n1665_), .A2(\A[960] ), .B(new_n1668_), .ZN(new_n1669_));
  NOR2_X1    g00667(.A1(new_n1651_), .A2(new_n1653_), .ZN(new_n1670_));
  AOI21_X1   g00668(.A1(new_n1656_), .A2(\A[957] ), .B(new_n1670_), .ZN(new_n1671_));
  OR4_X2     g00669(.A1(new_n1657_), .A2(new_n1666_), .A3(new_n1669_), .A4(new_n1671_), .Z(new_n1672_));
  NAND2_X1   g00670(.A1(new_n1667_), .A2(new_n1672_), .ZN(new_n1673_));
  XOR2_X1    g00671(.A1(new_n1649_), .A2(new_n1673_), .Z(new_n1674_));
  INV_X1     g00672(.I(\A[951] ), .ZN(new_n1675_));
  INV_X1     g00673(.I(\A[949] ), .ZN(new_n1676_));
  NAND2_X1   g00674(.A1(new_n1676_), .A2(\A[950] ), .ZN(new_n1677_));
  INV_X1     g00675(.I(\A[950] ), .ZN(new_n1678_));
  AOI21_X1   g00676(.A1(\A[949] ), .A2(new_n1678_), .B(new_n1675_), .ZN(new_n1679_));
  NAND2_X1   g00677(.A1(new_n1678_), .A2(\A[949] ), .ZN(new_n1680_));
  NAND2_X1   g00678(.A1(new_n1677_), .A2(new_n1680_), .ZN(new_n1681_));
  AOI22_X1   g00679(.A1(new_n1681_), .A2(new_n1675_), .B1(new_n1679_), .B2(new_n1677_), .ZN(new_n1682_));
  INV_X1     g00680(.I(\A[954] ), .ZN(new_n1683_));
  INV_X1     g00681(.I(\A[952] ), .ZN(new_n1684_));
  NAND2_X1   g00682(.A1(new_n1684_), .A2(\A[953] ), .ZN(new_n1685_));
  INV_X1     g00683(.I(\A[953] ), .ZN(new_n1686_));
  AOI21_X1   g00684(.A1(\A[952] ), .A2(new_n1686_), .B(new_n1683_), .ZN(new_n1687_));
  NAND2_X1   g00685(.A1(new_n1686_), .A2(\A[952] ), .ZN(new_n1688_));
  NAND2_X1   g00686(.A1(new_n1685_), .A2(new_n1688_), .ZN(new_n1689_));
  AOI22_X1   g00687(.A1(new_n1689_), .A2(new_n1683_), .B1(new_n1687_), .B2(new_n1685_), .ZN(new_n1690_));
  XOR2_X1    g00688(.A1(new_n1682_), .A2(new_n1690_), .Z(new_n1691_));
  NOR2_X1    g00689(.A1(new_n1684_), .A2(new_n1686_), .ZN(new_n1692_));
  AOI21_X1   g00690(.A1(new_n1689_), .A2(\A[954] ), .B(new_n1692_), .ZN(new_n1693_));
  NOR2_X1    g00691(.A1(new_n1676_), .A2(new_n1678_), .ZN(new_n1694_));
  AOI21_X1   g00692(.A1(new_n1681_), .A2(\A[951] ), .B(new_n1694_), .ZN(new_n1695_));
  OR4_X2     g00693(.A1(new_n1682_), .A2(new_n1690_), .A3(new_n1693_), .A4(new_n1695_), .Z(new_n1696_));
  NAND2_X1   g00694(.A1(new_n1691_), .A2(new_n1696_), .ZN(new_n1697_));
  INV_X1     g00695(.I(\A[945] ), .ZN(new_n1698_));
  INV_X1     g00696(.I(\A[943] ), .ZN(new_n1699_));
  NAND2_X1   g00697(.A1(new_n1699_), .A2(\A[944] ), .ZN(new_n1700_));
  INV_X1     g00698(.I(\A[944] ), .ZN(new_n1701_));
  AOI21_X1   g00699(.A1(\A[943] ), .A2(new_n1701_), .B(new_n1698_), .ZN(new_n1702_));
  NAND2_X1   g00700(.A1(new_n1701_), .A2(\A[943] ), .ZN(new_n1703_));
  NAND2_X1   g00701(.A1(new_n1700_), .A2(new_n1703_), .ZN(new_n1704_));
  AOI22_X1   g00702(.A1(new_n1704_), .A2(new_n1698_), .B1(new_n1702_), .B2(new_n1700_), .ZN(new_n1705_));
  INV_X1     g00703(.I(\A[948] ), .ZN(new_n1706_));
  INV_X1     g00704(.I(\A[946] ), .ZN(new_n1707_));
  NAND2_X1   g00705(.A1(new_n1707_), .A2(\A[947] ), .ZN(new_n1708_));
  INV_X1     g00706(.I(\A[947] ), .ZN(new_n1709_));
  AOI21_X1   g00707(.A1(\A[946] ), .A2(new_n1709_), .B(new_n1706_), .ZN(new_n1710_));
  NAND2_X1   g00708(.A1(new_n1709_), .A2(\A[946] ), .ZN(new_n1711_));
  NAND2_X1   g00709(.A1(new_n1708_), .A2(new_n1711_), .ZN(new_n1712_));
  AOI22_X1   g00710(.A1(new_n1712_), .A2(new_n1706_), .B1(new_n1710_), .B2(new_n1708_), .ZN(new_n1713_));
  XOR2_X1    g00711(.A1(new_n1705_), .A2(new_n1713_), .Z(new_n1714_));
  NOR2_X1    g00712(.A1(new_n1707_), .A2(new_n1709_), .ZN(new_n1715_));
  AOI21_X1   g00713(.A1(new_n1712_), .A2(\A[948] ), .B(new_n1715_), .ZN(new_n1716_));
  NOR2_X1    g00714(.A1(new_n1699_), .A2(new_n1701_), .ZN(new_n1717_));
  AOI21_X1   g00715(.A1(new_n1704_), .A2(\A[945] ), .B(new_n1717_), .ZN(new_n1718_));
  OR4_X2     g00716(.A1(new_n1705_), .A2(new_n1713_), .A3(new_n1716_), .A4(new_n1718_), .Z(new_n1719_));
  NAND2_X1   g00717(.A1(new_n1714_), .A2(new_n1719_), .ZN(new_n1720_));
  XOR2_X1    g00718(.A1(new_n1697_), .A2(new_n1720_), .Z(new_n1721_));
  XNOR2_X1   g00719(.A1(new_n1674_), .A2(new_n1721_), .ZN(new_n1722_));
  XNOR2_X1   g00720(.A1(new_n1624_), .A2(new_n1722_), .ZN(new_n1723_));
  INV_X1     g00721(.I(new_n1723_), .ZN(new_n1724_));
  INV_X1     g00722(.I(\A[76] ), .ZN(new_n1725_));
  INV_X1     g00723(.I(\A[77] ), .ZN(new_n1726_));
  NOR2_X1    g00724(.A1(new_n1725_), .A2(new_n1726_), .ZN(new_n1727_));
  NAND2_X1   g00725(.A1(new_n1726_), .A2(\A[76] ), .ZN(new_n1728_));
  NAND2_X1   g00726(.A1(new_n1725_), .A2(\A[77] ), .ZN(new_n1729_));
  NAND2_X1   g00727(.A1(new_n1728_), .A2(new_n1729_), .ZN(new_n1730_));
  AOI21_X1   g00728(.A1(new_n1730_), .A2(\A[78] ), .B(new_n1727_), .ZN(new_n1731_));
  INV_X1     g00729(.I(\A[73] ), .ZN(new_n1732_));
  INV_X1     g00730(.I(\A[74] ), .ZN(new_n1733_));
  NOR2_X1    g00731(.A1(new_n1732_), .A2(new_n1733_), .ZN(new_n1734_));
  NAND2_X1   g00732(.A1(new_n1733_), .A2(\A[73] ), .ZN(new_n1735_));
  NAND2_X1   g00733(.A1(new_n1732_), .A2(\A[74] ), .ZN(new_n1736_));
  NAND2_X1   g00734(.A1(new_n1735_), .A2(new_n1736_), .ZN(new_n1737_));
  AOI21_X1   g00735(.A1(new_n1737_), .A2(\A[75] ), .B(new_n1734_), .ZN(new_n1738_));
  NOR2_X1    g00736(.A1(new_n1732_), .A2(\A[74] ), .ZN(new_n1739_));
  NOR2_X1    g00737(.A1(new_n1733_), .A2(\A[73] ), .ZN(new_n1740_));
  NOR2_X1    g00738(.A1(new_n1739_), .A2(new_n1740_), .ZN(new_n1741_));
  NOR2_X1    g00739(.A1(new_n1741_), .A2(\A[75] ), .ZN(new_n1742_));
  INV_X1     g00740(.I(\A[75] ), .ZN(new_n1743_));
  NOR3_X1    g00741(.A1(new_n1739_), .A2(new_n1740_), .A3(new_n1743_), .ZN(new_n1744_));
  AOI21_X1   g00742(.A1(new_n1728_), .A2(new_n1729_), .B(\A[78] ), .ZN(new_n1745_));
  INV_X1     g00743(.I(\A[78] ), .ZN(new_n1746_));
  NOR2_X1    g00744(.A1(new_n1725_), .A2(\A[77] ), .ZN(new_n1747_));
  NOR2_X1    g00745(.A1(new_n1726_), .A2(\A[76] ), .ZN(new_n1748_));
  NOR3_X1    g00746(.A1(new_n1747_), .A2(new_n1748_), .A3(new_n1746_), .ZN(new_n1749_));
  OAI22_X1   g00747(.A1(new_n1742_), .A2(new_n1744_), .B1(new_n1749_), .B2(new_n1745_), .ZN(new_n1750_));
  NOR3_X1    g00748(.A1(new_n1750_), .A2(new_n1731_), .A3(new_n1738_), .ZN(new_n1751_));
  AOI21_X1   g00749(.A1(\A[73] ), .A2(new_n1733_), .B(new_n1743_), .ZN(new_n1752_));
  AOI22_X1   g00750(.A1(new_n1737_), .A2(new_n1743_), .B1(new_n1736_), .B2(new_n1752_), .ZN(new_n1753_));
  OAI21_X1   g00751(.A1(new_n1747_), .A2(new_n1748_), .B(new_n1746_), .ZN(new_n1754_));
  NAND3_X1   g00752(.A1(new_n1728_), .A2(new_n1729_), .A3(\A[78] ), .ZN(new_n1755_));
  NAND2_X1   g00753(.A1(new_n1754_), .A2(new_n1755_), .ZN(new_n1756_));
  XOR2_X1    g00754(.A1(new_n1753_), .A2(new_n1756_), .Z(new_n1757_));
  NOR2_X1    g00755(.A1(new_n1757_), .A2(new_n1751_), .ZN(new_n1758_));
  INV_X1     g00756(.I(\A[72] ), .ZN(new_n1759_));
  INV_X1     g00757(.I(\A[70] ), .ZN(new_n1760_));
  INV_X1     g00758(.I(\A[71] ), .ZN(new_n1761_));
  NOR2_X1    g00759(.A1(new_n1760_), .A2(new_n1761_), .ZN(new_n1762_));
  INV_X1     g00760(.I(new_n1762_), .ZN(new_n1763_));
  NOR2_X1    g00761(.A1(new_n1760_), .A2(\A[71] ), .ZN(new_n1764_));
  NOR2_X1    g00762(.A1(new_n1761_), .A2(\A[70] ), .ZN(new_n1765_));
  NOR2_X1    g00763(.A1(new_n1764_), .A2(new_n1765_), .ZN(new_n1766_));
  OAI21_X1   g00764(.A1(new_n1766_), .A2(new_n1759_), .B(new_n1763_), .ZN(new_n1767_));
  INV_X1     g00765(.I(\A[69] ), .ZN(new_n1768_));
  INV_X1     g00766(.I(\A[67] ), .ZN(new_n1769_));
  INV_X1     g00767(.I(\A[68] ), .ZN(new_n1770_));
  NOR2_X1    g00768(.A1(new_n1769_), .A2(new_n1770_), .ZN(new_n1771_));
  INV_X1     g00769(.I(new_n1771_), .ZN(new_n1772_));
  NOR2_X1    g00770(.A1(new_n1769_), .A2(\A[68] ), .ZN(new_n1773_));
  NOR2_X1    g00771(.A1(new_n1770_), .A2(\A[67] ), .ZN(new_n1774_));
  NOR2_X1    g00772(.A1(new_n1773_), .A2(new_n1774_), .ZN(new_n1775_));
  OAI21_X1   g00773(.A1(new_n1775_), .A2(new_n1768_), .B(new_n1772_), .ZN(new_n1776_));
  NAND2_X1   g00774(.A1(new_n1770_), .A2(\A[67] ), .ZN(new_n1777_));
  NAND2_X1   g00775(.A1(new_n1769_), .A2(\A[68] ), .ZN(new_n1778_));
  NAND2_X1   g00776(.A1(new_n1777_), .A2(new_n1778_), .ZN(new_n1779_));
  NAND2_X1   g00777(.A1(new_n1779_), .A2(new_n1768_), .ZN(new_n1780_));
  NOR2_X1    g00778(.A1(new_n1773_), .A2(new_n1768_), .ZN(new_n1781_));
  NAND2_X1   g00779(.A1(new_n1781_), .A2(new_n1778_), .ZN(new_n1782_));
  OAI21_X1   g00780(.A1(new_n1764_), .A2(new_n1765_), .B(new_n1759_), .ZN(new_n1783_));
  NAND2_X1   g00781(.A1(new_n1761_), .A2(\A[70] ), .ZN(new_n1784_));
  NAND2_X1   g00782(.A1(new_n1760_), .A2(\A[71] ), .ZN(new_n1785_));
  NAND3_X1   g00783(.A1(new_n1784_), .A2(new_n1785_), .A3(\A[72] ), .ZN(new_n1786_));
  AOI22_X1   g00784(.A1(new_n1780_), .A2(new_n1782_), .B1(new_n1783_), .B2(new_n1786_), .ZN(new_n1787_));
  NAND3_X1   g00785(.A1(new_n1787_), .A2(new_n1767_), .A3(new_n1776_), .ZN(new_n1788_));
  AOI22_X1   g00786(.A1(new_n1779_), .A2(new_n1768_), .B1(new_n1781_), .B2(new_n1778_), .ZN(new_n1789_));
  NAND2_X1   g00787(.A1(new_n1783_), .A2(new_n1786_), .ZN(new_n1790_));
  NAND2_X1   g00788(.A1(new_n1789_), .A2(new_n1790_), .ZN(new_n1791_));
  NAND2_X1   g00789(.A1(new_n1777_), .A2(\A[69] ), .ZN(new_n1792_));
  OAI22_X1   g00790(.A1(new_n1775_), .A2(\A[69] ), .B1(new_n1792_), .B2(new_n1774_), .ZN(new_n1793_));
  NAND2_X1   g00791(.A1(new_n1784_), .A2(new_n1785_), .ZN(new_n1794_));
  NOR2_X1    g00792(.A1(new_n1764_), .A2(new_n1759_), .ZN(new_n1795_));
  AOI22_X1   g00793(.A1(new_n1794_), .A2(new_n1759_), .B1(new_n1795_), .B2(new_n1785_), .ZN(new_n1796_));
  NAND2_X1   g00794(.A1(new_n1796_), .A2(new_n1793_), .ZN(new_n1797_));
  NAND2_X1   g00795(.A1(new_n1797_), .A2(new_n1791_), .ZN(new_n1798_));
  NAND2_X1   g00796(.A1(new_n1798_), .A2(new_n1788_), .ZN(new_n1799_));
  NAND2_X1   g00797(.A1(new_n1758_), .A2(new_n1799_), .ZN(new_n1800_));
  INV_X1     g00798(.I(new_n1727_), .ZN(new_n1801_));
  NOR2_X1    g00799(.A1(new_n1747_), .A2(new_n1748_), .ZN(new_n1802_));
  OAI21_X1   g00800(.A1(new_n1802_), .A2(new_n1746_), .B(new_n1801_), .ZN(new_n1803_));
  INV_X1     g00801(.I(new_n1734_), .ZN(new_n1804_));
  OAI21_X1   g00802(.A1(new_n1741_), .A2(new_n1743_), .B(new_n1804_), .ZN(new_n1805_));
  NAND2_X1   g00803(.A1(new_n1737_), .A2(new_n1743_), .ZN(new_n1806_));
  NAND2_X1   g00804(.A1(new_n1752_), .A2(new_n1736_), .ZN(new_n1807_));
  AOI22_X1   g00805(.A1(new_n1806_), .A2(new_n1807_), .B1(new_n1754_), .B2(new_n1755_), .ZN(new_n1808_));
  NAND3_X1   g00806(.A1(new_n1808_), .A2(new_n1803_), .A3(new_n1805_), .ZN(new_n1809_));
  OAI21_X1   g00807(.A1(\A[75] ), .A2(new_n1741_), .B(new_n1807_), .ZN(new_n1810_));
  NOR2_X1    g00808(.A1(new_n1745_), .A2(new_n1749_), .ZN(new_n1811_));
  NAND2_X1   g00809(.A1(new_n1810_), .A2(new_n1811_), .ZN(new_n1812_));
  NAND2_X1   g00810(.A1(new_n1753_), .A2(new_n1756_), .ZN(new_n1813_));
  NAND2_X1   g00811(.A1(new_n1812_), .A2(new_n1813_), .ZN(new_n1814_));
  NAND2_X1   g00812(.A1(new_n1814_), .A2(new_n1809_), .ZN(new_n1815_));
  AOI21_X1   g00813(.A1(new_n1794_), .A2(\A[72] ), .B(new_n1762_), .ZN(new_n1816_));
  AOI21_X1   g00814(.A1(new_n1779_), .A2(\A[69] ), .B(new_n1771_), .ZN(new_n1817_));
  NOR4_X1    g00815(.A1(new_n1789_), .A2(new_n1796_), .A3(new_n1816_), .A4(new_n1817_), .ZN(new_n1818_));
  NOR2_X1    g00816(.A1(new_n1796_), .A2(new_n1793_), .ZN(new_n1819_));
  NOR2_X1    g00817(.A1(new_n1789_), .A2(new_n1790_), .ZN(new_n1820_));
  NOR2_X1    g00818(.A1(new_n1819_), .A2(new_n1820_), .ZN(new_n1821_));
  NOR2_X1    g00819(.A1(new_n1821_), .A2(new_n1818_), .ZN(new_n1822_));
  NAND2_X1   g00820(.A1(new_n1822_), .A2(new_n1815_), .ZN(new_n1823_));
  NAND2_X1   g00821(.A1(new_n1800_), .A2(new_n1823_), .ZN(new_n1824_));
  INV_X1     g00822(.I(\A[64] ), .ZN(new_n1825_));
  INV_X1     g00823(.I(\A[65] ), .ZN(new_n1826_));
  NOR2_X1    g00824(.A1(new_n1825_), .A2(new_n1826_), .ZN(new_n1827_));
  NAND2_X1   g00825(.A1(new_n1826_), .A2(\A[64] ), .ZN(new_n1828_));
  NAND2_X1   g00826(.A1(new_n1825_), .A2(\A[65] ), .ZN(new_n1829_));
  NAND2_X1   g00827(.A1(new_n1828_), .A2(new_n1829_), .ZN(new_n1830_));
  AOI21_X1   g00828(.A1(new_n1830_), .A2(\A[66] ), .B(new_n1827_), .ZN(new_n1831_));
  INV_X1     g00829(.I(\A[61] ), .ZN(new_n1832_));
  INV_X1     g00830(.I(\A[62] ), .ZN(new_n1833_));
  NOR2_X1    g00831(.A1(new_n1832_), .A2(new_n1833_), .ZN(new_n1834_));
  NAND2_X1   g00832(.A1(new_n1833_), .A2(\A[61] ), .ZN(new_n1835_));
  NAND2_X1   g00833(.A1(new_n1832_), .A2(\A[62] ), .ZN(new_n1836_));
  NAND2_X1   g00834(.A1(new_n1835_), .A2(new_n1836_), .ZN(new_n1837_));
  AOI21_X1   g00835(.A1(new_n1837_), .A2(\A[63] ), .B(new_n1834_), .ZN(new_n1838_));
  NOR2_X1    g00836(.A1(new_n1833_), .A2(\A[61] ), .ZN(new_n1839_));
  NOR2_X1    g00837(.A1(new_n1832_), .A2(\A[62] ), .ZN(new_n1840_));
  NOR2_X1    g00838(.A1(new_n1840_), .A2(new_n1839_), .ZN(new_n1841_));
  NAND2_X1   g00839(.A1(new_n1835_), .A2(\A[63] ), .ZN(new_n1842_));
  OAI22_X1   g00840(.A1(new_n1841_), .A2(\A[63] ), .B1(new_n1842_), .B2(new_n1839_), .ZN(new_n1843_));
  INV_X1     g00841(.I(\A[66] ), .ZN(new_n1844_));
  NOR2_X1    g00842(.A1(new_n1825_), .A2(\A[65] ), .ZN(new_n1845_));
  NOR2_X1    g00843(.A1(new_n1826_), .A2(\A[64] ), .ZN(new_n1846_));
  OAI21_X1   g00844(.A1(new_n1845_), .A2(new_n1846_), .B(new_n1844_), .ZN(new_n1847_));
  NAND3_X1   g00845(.A1(new_n1828_), .A2(new_n1829_), .A3(\A[66] ), .ZN(new_n1848_));
  NAND2_X1   g00846(.A1(new_n1847_), .A2(new_n1848_), .ZN(new_n1849_));
  NAND2_X1   g00847(.A1(new_n1843_), .A2(new_n1849_), .ZN(new_n1850_));
  NOR3_X1    g00848(.A1(new_n1850_), .A2(new_n1831_), .A3(new_n1838_), .ZN(new_n1851_));
  XNOR2_X1   g00849(.A1(new_n1843_), .A2(new_n1849_), .ZN(new_n1852_));
  NOR2_X1    g00850(.A1(new_n1852_), .A2(new_n1851_), .ZN(new_n1853_));
  INV_X1     g00851(.I(\A[60] ), .ZN(new_n1854_));
  INV_X1     g00852(.I(\A[58] ), .ZN(new_n1855_));
  INV_X1     g00853(.I(\A[59] ), .ZN(new_n1856_));
  NOR2_X1    g00854(.A1(new_n1855_), .A2(new_n1856_), .ZN(new_n1857_));
  INV_X1     g00855(.I(new_n1857_), .ZN(new_n1858_));
  NOR2_X1    g00856(.A1(new_n1855_), .A2(\A[59] ), .ZN(new_n1859_));
  NOR2_X1    g00857(.A1(new_n1856_), .A2(\A[58] ), .ZN(new_n1860_));
  NOR2_X1    g00858(.A1(new_n1859_), .A2(new_n1860_), .ZN(new_n1861_));
  OAI21_X1   g00859(.A1(new_n1861_), .A2(new_n1854_), .B(new_n1858_), .ZN(new_n1862_));
  INV_X1     g00860(.I(\A[57] ), .ZN(new_n1863_));
  INV_X1     g00861(.I(\A[55] ), .ZN(new_n1864_));
  INV_X1     g00862(.I(\A[56] ), .ZN(new_n1865_));
  NOR2_X1    g00863(.A1(new_n1864_), .A2(new_n1865_), .ZN(new_n1866_));
  INV_X1     g00864(.I(new_n1866_), .ZN(new_n1867_));
  NOR2_X1    g00865(.A1(new_n1864_), .A2(\A[56] ), .ZN(new_n1868_));
  NOR2_X1    g00866(.A1(new_n1865_), .A2(\A[55] ), .ZN(new_n1869_));
  NOR2_X1    g00867(.A1(new_n1868_), .A2(new_n1869_), .ZN(new_n1870_));
  OAI21_X1   g00868(.A1(new_n1870_), .A2(new_n1863_), .B(new_n1867_), .ZN(new_n1871_));
  NAND2_X1   g00869(.A1(new_n1864_), .A2(\A[56] ), .ZN(new_n1872_));
  NAND2_X1   g00870(.A1(new_n1865_), .A2(\A[55] ), .ZN(new_n1873_));
  NAND2_X1   g00871(.A1(new_n1873_), .A2(new_n1872_), .ZN(new_n1874_));
  NOR2_X1    g00872(.A1(new_n1868_), .A2(new_n1863_), .ZN(new_n1875_));
  AOI22_X1   g00873(.A1(new_n1874_), .A2(new_n1863_), .B1(new_n1875_), .B2(new_n1872_), .ZN(new_n1876_));
  NAND2_X1   g00874(.A1(new_n1856_), .A2(\A[58] ), .ZN(new_n1877_));
  NAND2_X1   g00875(.A1(new_n1855_), .A2(\A[59] ), .ZN(new_n1878_));
  AOI21_X1   g00876(.A1(new_n1877_), .A2(new_n1878_), .B(\A[60] ), .ZN(new_n1879_));
  NOR3_X1    g00877(.A1(new_n1859_), .A2(new_n1860_), .A3(new_n1854_), .ZN(new_n1880_));
  NOR2_X1    g00878(.A1(new_n1879_), .A2(new_n1880_), .ZN(new_n1881_));
  NOR2_X1    g00879(.A1(new_n1876_), .A2(new_n1881_), .ZN(new_n1882_));
  NAND3_X1   g00880(.A1(new_n1882_), .A2(new_n1862_), .A3(new_n1871_), .ZN(new_n1883_));
  XOR2_X1    g00881(.A1(new_n1876_), .A2(new_n1881_), .Z(new_n1884_));
  NAND2_X1   g00882(.A1(new_n1884_), .A2(new_n1883_), .ZN(new_n1885_));
  NOR2_X1    g00883(.A1(new_n1853_), .A2(new_n1885_), .ZN(new_n1886_));
  INV_X1     g00884(.I(new_n1827_), .ZN(new_n1887_));
  NOR2_X1    g00885(.A1(new_n1845_), .A2(new_n1846_), .ZN(new_n1888_));
  OAI21_X1   g00886(.A1(new_n1888_), .A2(new_n1844_), .B(new_n1887_), .ZN(new_n1889_));
  INV_X1     g00887(.I(\A[63] ), .ZN(new_n1890_));
  INV_X1     g00888(.I(new_n1834_), .ZN(new_n1891_));
  OAI21_X1   g00889(.A1(new_n1841_), .A2(new_n1890_), .B(new_n1891_), .ZN(new_n1892_));
  NAND2_X1   g00890(.A1(new_n1837_), .A2(new_n1890_), .ZN(new_n1893_));
  NAND3_X1   g00891(.A1(new_n1835_), .A2(new_n1836_), .A3(\A[63] ), .ZN(new_n1894_));
  AOI22_X1   g00892(.A1(new_n1893_), .A2(new_n1894_), .B1(new_n1847_), .B2(new_n1848_), .ZN(new_n1895_));
  NAND3_X1   g00893(.A1(new_n1895_), .A2(new_n1889_), .A3(new_n1892_), .ZN(new_n1896_));
  XOR2_X1    g00894(.A1(new_n1843_), .A2(new_n1849_), .Z(new_n1897_));
  NAND2_X1   g00895(.A1(new_n1897_), .A2(new_n1896_), .ZN(new_n1898_));
  NAND2_X1   g00896(.A1(new_n1877_), .A2(new_n1878_), .ZN(new_n1899_));
  AOI21_X1   g00897(.A1(new_n1899_), .A2(\A[60] ), .B(new_n1857_), .ZN(new_n1900_));
  AOI21_X1   g00898(.A1(new_n1874_), .A2(\A[57] ), .B(new_n1866_), .ZN(new_n1901_));
  NOR2_X1    g00899(.A1(new_n1870_), .A2(\A[57] ), .ZN(new_n1902_));
  NAND2_X1   g00900(.A1(new_n1873_), .A2(\A[57] ), .ZN(new_n1903_));
  NOR2_X1    g00901(.A1(new_n1903_), .A2(new_n1869_), .ZN(new_n1904_));
  OAI22_X1   g00902(.A1(new_n1902_), .A2(new_n1904_), .B1(new_n1879_), .B2(new_n1880_), .ZN(new_n1905_));
  NOR3_X1    g00903(.A1(new_n1905_), .A2(new_n1900_), .A3(new_n1901_), .ZN(new_n1906_));
  NOR3_X1    g00904(.A1(new_n1881_), .A2(new_n1902_), .A3(new_n1904_), .ZN(new_n1907_));
  NOR3_X1    g00905(.A1(new_n1876_), .A2(new_n1879_), .A3(new_n1880_), .ZN(new_n1908_));
  NOR2_X1    g00906(.A1(new_n1908_), .A2(new_n1907_), .ZN(new_n1909_));
  NOR2_X1    g00907(.A1(new_n1909_), .A2(new_n1906_), .ZN(new_n1910_));
  NOR2_X1    g00908(.A1(new_n1898_), .A2(new_n1910_), .ZN(new_n1911_));
  NOR2_X1    g00909(.A1(new_n1886_), .A2(new_n1911_), .ZN(new_n1912_));
  NAND2_X1   g00910(.A1(new_n1912_), .A2(new_n1824_), .ZN(new_n1913_));
  NOR2_X1    g00911(.A1(new_n1822_), .A2(new_n1815_), .ZN(new_n1914_));
  NOR2_X1    g00912(.A1(new_n1758_), .A2(new_n1799_), .ZN(new_n1915_));
  NOR2_X1    g00913(.A1(new_n1915_), .A2(new_n1914_), .ZN(new_n1916_));
  NAND2_X1   g00914(.A1(new_n1898_), .A2(new_n1910_), .ZN(new_n1917_));
  NAND2_X1   g00915(.A1(new_n1853_), .A2(new_n1885_), .ZN(new_n1918_));
  NAND2_X1   g00916(.A1(new_n1918_), .A2(new_n1917_), .ZN(new_n1919_));
  NAND2_X1   g00917(.A1(new_n1919_), .A2(new_n1916_), .ZN(new_n1920_));
  NAND2_X1   g00918(.A1(new_n1920_), .A2(new_n1913_), .ZN(new_n1921_));
  INV_X1     g00919(.I(\A[52] ), .ZN(new_n1922_));
  INV_X1     g00920(.I(\A[53] ), .ZN(new_n1923_));
  NOR2_X1    g00921(.A1(new_n1922_), .A2(new_n1923_), .ZN(new_n1924_));
  NAND2_X1   g00922(.A1(new_n1923_), .A2(\A[52] ), .ZN(new_n1925_));
  NAND2_X1   g00923(.A1(new_n1922_), .A2(\A[53] ), .ZN(new_n1926_));
  NAND2_X1   g00924(.A1(new_n1925_), .A2(new_n1926_), .ZN(new_n1927_));
  AOI21_X1   g00925(.A1(new_n1927_), .A2(\A[54] ), .B(new_n1924_), .ZN(new_n1928_));
  INV_X1     g00926(.I(\A[49] ), .ZN(new_n1929_));
  INV_X1     g00927(.I(\A[50] ), .ZN(new_n1930_));
  NOR2_X1    g00928(.A1(new_n1929_), .A2(new_n1930_), .ZN(new_n1931_));
  NAND2_X1   g00929(.A1(new_n1930_), .A2(\A[49] ), .ZN(new_n1932_));
  NAND2_X1   g00930(.A1(new_n1929_), .A2(\A[50] ), .ZN(new_n1933_));
  NAND2_X1   g00931(.A1(new_n1932_), .A2(new_n1933_), .ZN(new_n1934_));
  AOI21_X1   g00932(.A1(new_n1934_), .A2(\A[51] ), .B(new_n1931_), .ZN(new_n1935_));
  NOR2_X1    g00933(.A1(new_n1929_), .A2(\A[50] ), .ZN(new_n1936_));
  NOR2_X1    g00934(.A1(new_n1930_), .A2(\A[49] ), .ZN(new_n1937_));
  NOR2_X1    g00935(.A1(new_n1936_), .A2(new_n1937_), .ZN(new_n1938_));
  NAND3_X1   g00936(.A1(new_n1932_), .A2(new_n1933_), .A3(\A[51] ), .ZN(new_n1939_));
  OAI21_X1   g00937(.A1(\A[51] ), .A2(new_n1938_), .B(new_n1939_), .ZN(new_n1940_));
  INV_X1     g00938(.I(\A[54] ), .ZN(new_n1941_));
  NOR2_X1    g00939(.A1(new_n1922_), .A2(\A[53] ), .ZN(new_n1942_));
  NOR2_X1    g00940(.A1(new_n1923_), .A2(\A[52] ), .ZN(new_n1943_));
  OAI21_X1   g00941(.A1(new_n1942_), .A2(new_n1943_), .B(new_n1941_), .ZN(new_n1944_));
  NAND3_X1   g00942(.A1(new_n1925_), .A2(new_n1926_), .A3(\A[54] ), .ZN(new_n1945_));
  NAND2_X1   g00943(.A1(new_n1944_), .A2(new_n1945_), .ZN(new_n1946_));
  NAND2_X1   g00944(.A1(new_n1940_), .A2(new_n1946_), .ZN(new_n1947_));
  NOR3_X1    g00945(.A1(new_n1947_), .A2(new_n1928_), .A3(new_n1935_), .ZN(new_n1948_));
  INV_X1     g00946(.I(\A[51] ), .ZN(new_n1949_));
  NAND2_X1   g00947(.A1(new_n1934_), .A2(new_n1949_), .ZN(new_n1950_));
  AOI21_X1   g00948(.A1(new_n1950_), .A2(new_n1939_), .B(new_n1946_), .ZN(new_n1951_));
  AOI21_X1   g00949(.A1(new_n1944_), .A2(new_n1945_), .B(new_n1940_), .ZN(new_n1952_));
  NOR2_X1    g00950(.A1(new_n1952_), .A2(new_n1951_), .ZN(new_n1953_));
  NOR2_X1    g00951(.A1(new_n1953_), .A2(new_n1948_), .ZN(new_n1954_));
  INV_X1     g00952(.I(\A[48] ), .ZN(new_n1955_));
  INV_X1     g00953(.I(\A[46] ), .ZN(new_n1956_));
  INV_X1     g00954(.I(\A[47] ), .ZN(new_n1957_));
  NOR2_X1    g00955(.A1(new_n1956_), .A2(new_n1957_), .ZN(new_n1958_));
  INV_X1     g00956(.I(new_n1958_), .ZN(new_n1959_));
  NOR2_X1    g00957(.A1(new_n1956_), .A2(\A[47] ), .ZN(new_n1960_));
  NOR2_X1    g00958(.A1(new_n1957_), .A2(\A[46] ), .ZN(new_n1961_));
  NOR2_X1    g00959(.A1(new_n1960_), .A2(new_n1961_), .ZN(new_n1962_));
  OAI21_X1   g00960(.A1(new_n1962_), .A2(new_n1955_), .B(new_n1959_), .ZN(new_n1963_));
  INV_X1     g00961(.I(\A[45] ), .ZN(new_n1964_));
  INV_X1     g00962(.I(\A[43] ), .ZN(new_n1965_));
  INV_X1     g00963(.I(\A[44] ), .ZN(new_n1966_));
  NOR2_X1    g00964(.A1(new_n1965_), .A2(new_n1966_), .ZN(new_n1967_));
  INV_X1     g00965(.I(new_n1967_), .ZN(new_n1968_));
  NOR2_X1    g00966(.A1(new_n1965_), .A2(\A[44] ), .ZN(new_n1969_));
  NOR2_X1    g00967(.A1(new_n1966_), .A2(\A[43] ), .ZN(new_n1970_));
  NOR2_X1    g00968(.A1(new_n1969_), .A2(new_n1970_), .ZN(new_n1971_));
  OAI21_X1   g00969(.A1(new_n1971_), .A2(new_n1964_), .B(new_n1968_), .ZN(new_n1972_));
  NAND2_X1   g00970(.A1(new_n1966_), .A2(\A[43] ), .ZN(new_n1973_));
  NAND2_X1   g00971(.A1(new_n1973_), .A2(\A[45] ), .ZN(new_n1974_));
  OAI22_X1   g00972(.A1(new_n1971_), .A2(\A[45] ), .B1(new_n1974_), .B2(new_n1970_), .ZN(new_n1975_));
  OAI21_X1   g00973(.A1(new_n1960_), .A2(new_n1961_), .B(new_n1955_), .ZN(new_n1976_));
  NAND2_X1   g00974(.A1(new_n1957_), .A2(\A[46] ), .ZN(new_n1977_));
  NAND2_X1   g00975(.A1(new_n1956_), .A2(\A[47] ), .ZN(new_n1978_));
  NAND3_X1   g00976(.A1(new_n1977_), .A2(new_n1978_), .A3(\A[48] ), .ZN(new_n1979_));
  NAND2_X1   g00977(.A1(new_n1976_), .A2(new_n1979_), .ZN(new_n1980_));
  NAND4_X1   g00978(.A1(new_n1975_), .A2(new_n1980_), .A3(new_n1963_), .A4(new_n1972_), .ZN(new_n1981_));
  XOR2_X1    g00979(.A1(new_n1975_), .A2(new_n1980_), .Z(new_n1982_));
  NAND2_X1   g00980(.A1(new_n1982_), .A2(new_n1981_), .ZN(new_n1983_));
  NAND2_X1   g00981(.A1(new_n1954_), .A2(new_n1983_), .ZN(new_n1984_));
  INV_X1     g00982(.I(new_n1924_), .ZN(new_n1985_));
  NOR2_X1    g00983(.A1(new_n1942_), .A2(new_n1943_), .ZN(new_n1986_));
  OAI21_X1   g00984(.A1(new_n1986_), .A2(new_n1941_), .B(new_n1985_), .ZN(new_n1987_));
  INV_X1     g00985(.I(new_n1931_), .ZN(new_n1988_));
  OAI21_X1   g00986(.A1(new_n1938_), .A2(new_n1949_), .B(new_n1988_), .ZN(new_n1989_));
  AOI22_X1   g00987(.A1(new_n1950_), .A2(new_n1939_), .B1(new_n1944_), .B2(new_n1945_), .ZN(new_n1990_));
  NAND3_X1   g00988(.A1(new_n1990_), .A2(new_n1987_), .A3(new_n1989_), .ZN(new_n1991_));
  XOR2_X1    g00989(.A1(new_n1940_), .A2(new_n1946_), .Z(new_n1992_));
  NAND2_X1   g00990(.A1(new_n1992_), .A2(new_n1991_), .ZN(new_n1993_));
  INV_X1     g00991(.I(new_n1981_), .ZN(new_n1994_));
  XNOR2_X1   g00992(.A1(new_n1975_), .A2(new_n1980_), .ZN(new_n1995_));
  NOR2_X1    g00993(.A1(new_n1995_), .A2(new_n1994_), .ZN(new_n1996_));
  NAND2_X1   g00994(.A1(new_n1996_), .A2(new_n1993_), .ZN(new_n1997_));
  NAND2_X1   g00995(.A1(new_n1997_), .A2(new_n1984_), .ZN(new_n1998_));
  INV_X1     g00996(.I(\A[42] ), .ZN(new_n1999_));
  INV_X1     g00997(.I(\A[40] ), .ZN(new_n2000_));
  INV_X1     g00998(.I(\A[41] ), .ZN(new_n2001_));
  NOR2_X1    g00999(.A1(new_n2000_), .A2(new_n2001_), .ZN(new_n2002_));
  INV_X1     g01000(.I(new_n2002_), .ZN(new_n2003_));
  NOR2_X1    g01001(.A1(new_n2000_), .A2(\A[41] ), .ZN(new_n2004_));
  NOR2_X1    g01002(.A1(new_n2001_), .A2(\A[40] ), .ZN(new_n2005_));
  NOR2_X1    g01003(.A1(new_n2004_), .A2(new_n2005_), .ZN(new_n2006_));
  OAI21_X1   g01004(.A1(new_n2006_), .A2(new_n1999_), .B(new_n2003_), .ZN(new_n2007_));
  INV_X1     g01005(.I(\A[39] ), .ZN(new_n2008_));
  INV_X1     g01006(.I(\A[37] ), .ZN(new_n2009_));
  INV_X1     g01007(.I(\A[38] ), .ZN(new_n2010_));
  NOR2_X1    g01008(.A1(new_n2009_), .A2(new_n2010_), .ZN(new_n2011_));
  INV_X1     g01009(.I(new_n2011_), .ZN(new_n2012_));
  NOR2_X1    g01010(.A1(new_n2009_), .A2(\A[38] ), .ZN(new_n2013_));
  NOR2_X1    g01011(.A1(new_n2010_), .A2(\A[37] ), .ZN(new_n2014_));
  NOR2_X1    g01012(.A1(new_n2013_), .A2(new_n2014_), .ZN(new_n2015_));
  OAI21_X1   g01013(.A1(new_n2015_), .A2(new_n2008_), .B(new_n2012_), .ZN(new_n2016_));
  NAND2_X1   g01014(.A1(new_n2009_), .A2(\A[38] ), .ZN(new_n2017_));
  NAND2_X1   g01015(.A1(new_n2010_), .A2(\A[37] ), .ZN(new_n2018_));
  NAND2_X1   g01016(.A1(new_n2018_), .A2(new_n2017_), .ZN(new_n2019_));
  NOR2_X1    g01017(.A1(new_n2013_), .A2(new_n2008_), .ZN(new_n2020_));
  AOI22_X1   g01018(.A1(new_n2019_), .A2(new_n2008_), .B1(new_n2020_), .B2(new_n2017_), .ZN(new_n2021_));
  NAND2_X1   g01019(.A1(new_n2000_), .A2(\A[41] ), .ZN(new_n2022_));
  NAND2_X1   g01020(.A1(new_n2001_), .A2(\A[40] ), .ZN(new_n2023_));
  NAND2_X1   g01021(.A1(new_n2023_), .A2(new_n2022_), .ZN(new_n2024_));
  AOI21_X1   g01022(.A1(\A[40] ), .A2(new_n2001_), .B(new_n1999_), .ZN(new_n2025_));
  AOI22_X1   g01023(.A1(new_n2024_), .A2(new_n1999_), .B1(new_n2022_), .B2(new_n2025_), .ZN(new_n2026_));
  NOR2_X1    g01024(.A1(new_n2021_), .A2(new_n2026_), .ZN(new_n2027_));
  NAND3_X1   g01025(.A1(new_n2027_), .A2(new_n2007_), .A3(new_n2016_), .ZN(new_n2028_));
  XOR2_X1    g01026(.A1(new_n2021_), .A2(new_n2026_), .Z(new_n2029_));
  NAND2_X1   g01027(.A1(new_n2029_), .A2(new_n2028_), .ZN(new_n2030_));
  INV_X1     g01028(.I(\A[34] ), .ZN(new_n2031_));
  INV_X1     g01029(.I(\A[35] ), .ZN(new_n2032_));
  NOR2_X1    g01030(.A1(new_n2031_), .A2(new_n2032_), .ZN(new_n2033_));
  NAND2_X1   g01031(.A1(new_n2032_), .A2(\A[34] ), .ZN(new_n2034_));
  NAND2_X1   g01032(.A1(new_n2031_), .A2(\A[35] ), .ZN(new_n2035_));
  NAND2_X1   g01033(.A1(new_n2034_), .A2(new_n2035_), .ZN(new_n2036_));
  AOI21_X1   g01034(.A1(new_n2036_), .A2(\A[36] ), .B(new_n2033_), .ZN(new_n2037_));
  INV_X1     g01035(.I(\A[31] ), .ZN(new_n2038_));
  INV_X1     g01036(.I(\A[32] ), .ZN(new_n2039_));
  NOR2_X1    g01037(.A1(new_n2038_), .A2(new_n2039_), .ZN(new_n2040_));
  NAND2_X1   g01038(.A1(new_n2039_), .A2(\A[31] ), .ZN(new_n2041_));
  NAND2_X1   g01039(.A1(new_n2038_), .A2(\A[32] ), .ZN(new_n2042_));
  NAND2_X1   g01040(.A1(new_n2041_), .A2(new_n2042_), .ZN(new_n2043_));
  AOI21_X1   g01041(.A1(new_n2043_), .A2(\A[33] ), .B(new_n2040_), .ZN(new_n2044_));
  INV_X1     g01042(.I(\A[33] ), .ZN(new_n2045_));
  NOR2_X1    g01043(.A1(new_n2038_), .A2(\A[32] ), .ZN(new_n2046_));
  NOR2_X1    g01044(.A1(new_n2046_), .A2(new_n2045_), .ZN(new_n2047_));
  AOI22_X1   g01045(.A1(new_n2043_), .A2(new_n2045_), .B1(new_n2047_), .B2(new_n2042_), .ZN(new_n2048_));
  INV_X1     g01046(.I(\A[36] ), .ZN(new_n2049_));
  AOI21_X1   g01047(.A1(\A[34] ), .A2(new_n2032_), .B(new_n2049_), .ZN(new_n2050_));
  AOI22_X1   g01048(.A1(new_n2036_), .A2(new_n2049_), .B1(new_n2035_), .B2(new_n2050_), .ZN(new_n2051_));
  NOR4_X1    g01049(.A1(new_n2048_), .A2(new_n2051_), .A3(new_n2037_), .A4(new_n2044_), .ZN(new_n2052_));
  XNOR2_X1   g01050(.A1(new_n2048_), .A2(new_n2051_), .ZN(new_n2053_));
  NOR2_X1    g01051(.A1(new_n2053_), .A2(new_n2052_), .ZN(new_n2054_));
  NAND2_X1   g01052(.A1(new_n2054_), .A2(new_n2030_), .ZN(new_n2055_));
  INV_X1     g01053(.I(new_n2052_), .ZN(new_n2056_));
  XOR2_X1    g01054(.A1(new_n2048_), .A2(new_n2051_), .Z(new_n2057_));
  NAND2_X1   g01055(.A1(new_n2057_), .A2(new_n2056_), .ZN(new_n2058_));
  NAND3_X1   g01056(.A1(new_n2058_), .A2(new_n2028_), .A3(new_n2029_), .ZN(new_n2059_));
  NAND3_X1   g01057(.A1(new_n1998_), .A2(new_n2055_), .A3(new_n2059_), .ZN(new_n2060_));
  NAND2_X1   g01058(.A1(new_n2055_), .A2(new_n2059_), .ZN(new_n2061_));
  NAND3_X1   g01059(.A1(new_n2061_), .A2(new_n1984_), .A3(new_n1997_), .ZN(new_n2062_));
  NAND2_X1   g01060(.A1(new_n2062_), .A2(new_n2060_), .ZN(new_n2063_));
  XNOR2_X1   g01061(.A1(new_n2063_), .A2(new_n1921_), .ZN(new_n2064_));
  INV_X1     g01062(.I(\A[993] ), .ZN(new_n2065_));
  INV_X1     g01063(.I(\A[991] ), .ZN(new_n2066_));
  NAND2_X1   g01064(.A1(new_n2066_), .A2(\A[992] ), .ZN(new_n2067_));
  INV_X1     g01065(.I(\A[992] ), .ZN(new_n2068_));
  AOI21_X1   g01066(.A1(\A[991] ), .A2(new_n2068_), .B(new_n2065_), .ZN(new_n2069_));
  NAND2_X1   g01067(.A1(new_n2068_), .A2(\A[991] ), .ZN(new_n2070_));
  NAND2_X1   g01068(.A1(new_n2067_), .A2(new_n2070_), .ZN(new_n2071_));
  AOI22_X1   g01069(.A1(new_n2071_), .A2(new_n2065_), .B1(new_n2069_), .B2(new_n2067_), .ZN(new_n2072_));
  INV_X1     g01070(.I(\A[996] ), .ZN(new_n2073_));
  INV_X1     g01071(.I(\A[994] ), .ZN(new_n2074_));
  NAND2_X1   g01072(.A1(new_n2074_), .A2(\A[995] ), .ZN(new_n2075_));
  NOR2_X1    g01073(.A1(new_n2074_), .A2(\A[995] ), .ZN(new_n2076_));
  NOR2_X1    g01074(.A1(new_n2076_), .A2(new_n2073_), .ZN(new_n2077_));
  INV_X1     g01075(.I(\A[995] ), .ZN(new_n2078_));
  NAND2_X1   g01076(.A1(new_n2078_), .A2(\A[994] ), .ZN(new_n2079_));
  NAND2_X1   g01077(.A1(new_n2075_), .A2(new_n2079_), .ZN(new_n2080_));
  AOI22_X1   g01078(.A1(new_n2080_), .A2(new_n2073_), .B1(new_n2077_), .B2(new_n2075_), .ZN(new_n2081_));
  NOR2_X1    g01079(.A1(new_n2074_), .A2(new_n2078_), .ZN(new_n2082_));
  AOI21_X1   g01080(.A1(new_n2080_), .A2(\A[996] ), .B(new_n2082_), .ZN(new_n2083_));
  NOR2_X1    g01081(.A1(new_n2066_), .A2(new_n2068_), .ZN(new_n2084_));
  AOI21_X1   g01082(.A1(new_n2071_), .A2(\A[993] ), .B(new_n2084_), .ZN(new_n2085_));
  XOR2_X1    g01083(.A1(new_n2081_), .A2(new_n2072_), .Z(new_n2086_));
  INV_X1     g01084(.I(new_n2086_), .ZN(new_n2087_));
  INV_X1     g01085(.I(\A[5] ), .ZN(new_n2088_));
  XOR2_X1    g01086(.A1(\A[3] ), .A2(\A[4] ), .Z(new_n2089_));
  INV_X1     g01087(.I(\A[4] ), .ZN(new_n2090_));
  NOR2_X1    g01088(.A1(new_n2090_), .A2(\A[3] ), .ZN(new_n2091_));
  INV_X1     g01089(.I(\A[3] ), .ZN(new_n2092_));
  OAI21_X1   g01090(.A1(new_n2092_), .A2(\A[4] ), .B(\A[5] ), .ZN(new_n2093_));
  NOR2_X1    g01091(.A1(new_n2093_), .A2(new_n2091_), .ZN(new_n2094_));
  AOI21_X1   g01092(.A1(new_n2088_), .A2(new_n2089_), .B(new_n2094_), .ZN(new_n2095_));
  INV_X1     g01093(.I(\A[0] ), .ZN(new_n2096_));
  NAND2_X1   g01094(.A1(new_n2096_), .A2(\A[1] ), .ZN(new_n2097_));
  INV_X1     g01095(.I(\A[1] ), .ZN(new_n2098_));
  NAND2_X1   g01096(.A1(new_n2098_), .A2(\A[0] ), .ZN(new_n2099_));
  NAND3_X1   g01097(.A1(new_n2097_), .A2(new_n2099_), .A3(\A[2] ), .ZN(new_n2100_));
  INV_X1     g01098(.I(\A[2] ), .ZN(new_n2101_));
  NOR2_X1    g01099(.A1(new_n2098_), .A2(\A[0] ), .ZN(new_n2102_));
  NOR2_X1    g01100(.A1(new_n2096_), .A2(\A[1] ), .ZN(new_n2103_));
  OAI21_X1   g01101(.A1(new_n2102_), .A2(new_n2103_), .B(new_n2101_), .ZN(new_n2104_));
  AOI21_X1   g01102(.A1(new_n2104_), .A2(new_n2100_), .B(\A[6] ), .ZN(new_n2105_));
  INV_X1     g01103(.I(\A[6] ), .ZN(new_n2106_));
  NOR3_X1    g01104(.A1(new_n2102_), .A2(new_n2103_), .A3(new_n2101_), .ZN(new_n2107_));
  AOI21_X1   g01105(.A1(new_n2097_), .A2(new_n2099_), .B(\A[2] ), .ZN(new_n2108_));
  NOR3_X1    g01106(.A1(new_n2108_), .A2(new_n2107_), .A3(new_n2106_), .ZN(new_n2109_));
  OAI21_X1   g01107(.A1(new_n2109_), .A2(new_n2105_), .B(new_n2095_), .ZN(new_n2110_));
  NOR2_X1    g01108(.A1(new_n2092_), .A2(\A[4] ), .ZN(new_n2111_));
  NOR2_X1    g01109(.A1(new_n2111_), .A2(new_n2091_), .ZN(new_n2112_));
  OAI22_X1   g01110(.A1(new_n2112_), .A2(\A[5] ), .B1(new_n2091_), .B2(new_n2093_), .ZN(new_n2113_));
  OAI21_X1   g01111(.A1(new_n2108_), .A2(new_n2107_), .B(new_n2106_), .ZN(new_n2114_));
  NAND3_X1   g01112(.A1(new_n2104_), .A2(new_n2100_), .A3(\A[6] ), .ZN(new_n2115_));
  NAND3_X1   g01113(.A1(new_n2113_), .A2(new_n2114_), .A3(new_n2115_), .ZN(new_n2116_));
  INV_X1     g01114(.I(\A[998] ), .ZN(new_n2117_));
  NOR2_X1    g01115(.A1(new_n2117_), .A2(\A[997] ), .ZN(new_n2118_));
  INV_X1     g01116(.I(new_n2118_), .ZN(new_n2119_));
  INV_X1     g01117(.I(\A[999] ), .ZN(new_n2120_));
  INV_X1     g01118(.I(\A[997] ), .ZN(new_n2121_));
  NOR2_X1    g01119(.A1(new_n2121_), .A2(\A[998] ), .ZN(new_n2122_));
  NOR2_X1    g01120(.A1(new_n2122_), .A2(new_n2120_), .ZN(new_n2123_));
  NAND2_X1   g01121(.A1(new_n2123_), .A2(new_n2119_), .ZN(new_n2124_));
  NOR2_X1    g01122(.A1(new_n2118_), .A2(new_n2122_), .ZN(new_n2125_));
  OAI21_X1   g01123(.A1(\A[999] ), .A2(new_n2125_), .B(new_n2124_), .ZN(new_n2126_));
  NAND3_X1   g01124(.A1(new_n2110_), .A2(new_n2116_), .A3(new_n2126_), .ZN(new_n2127_));
  AOI21_X1   g01125(.A1(new_n2114_), .A2(new_n2115_), .B(new_n2113_), .ZN(new_n2128_));
  NOR3_X1    g01126(.A1(new_n2095_), .A2(new_n2109_), .A3(new_n2105_), .ZN(new_n2129_));
  INV_X1     g01127(.I(new_n2125_), .ZN(new_n2130_));
  AOI22_X1   g01128(.A1(new_n2130_), .A2(new_n2120_), .B1(new_n2123_), .B2(new_n2119_), .ZN(new_n2131_));
  OAI21_X1   g01129(.A1(new_n2129_), .A2(new_n2128_), .B(new_n2131_), .ZN(new_n2132_));
  NAND2_X1   g01130(.A1(new_n2132_), .A2(new_n2127_), .ZN(new_n2133_));
  XOR2_X1    g01131(.A1(new_n2133_), .A2(new_n2087_), .Z(new_n2134_));
  INV_X1     g01132(.I(new_n2134_), .ZN(new_n2135_));
  INV_X1     g01133(.I(\A[28] ), .ZN(new_n2136_));
  INV_X1     g01134(.I(\A[29] ), .ZN(new_n2137_));
  NOR2_X1    g01135(.A1(new_n2136_), .A2(new_n2137_), .ZN(new_n2138_));
  NAND2_X1   g01136(.A1(new_n2137_), .A2(\A[28] ), .ZN(new_n2139_));
  NAND2_X1   g01137(.A1(new_n2136_), .A2(\A[29] ), .ZN(new_n2140_));
  NAND2_X1   g01138(.A1(new_n2139_), .A2(new_n2140_), .ZN(new_n2141_));
  AOI21_X1   g01139(.A1(new_n2141_), .A2(\A[30] ), .B(new_n2138_), .ZN(new_n2142_));
  INV_X1     g01140(.I(\A[25] ), .ZN(new_n2143_));
  INV_X1     g01141(.I(\A[26] ), .ZN(new_n2144_));
  NOR2_X1    g01142(.A1(new_n2143_), .A2(new_n2144_), .ZN(new_n2145_));
  NAND2_X1   g01143(.A1(new_n2144_), .A2(\A[25] ), .ZN(new_n2146_));
  NAND2_X1   g01144(.A1(new_n2143_), .A2(\A[26] ), .ZN(new_n2147_));
  NAND2_X1   g01145(.A1(new_n2146_), .A2(new_n2147_), .ZN(new_n2148_));
  AOI21_X1   g01146(.A1(new_n2148_), .A2(\A[27] ), .B(new_n2145_), .ZN(new_n2149_));
  NOR2_X1    g01147(.A1(new_n2143_), .A2(\A[26] ), .ZN(new_n2150_));
  NOR2_X1    g01148(.A1(new_n2144_), .A2(\A[25] ), .ZN(new_n2151_));
  NOR2_X1    g01149(.A1(new_n2150_), .A2(new_n2151_), .ZN(new_n2152_));
  NOR2_X1    g01150(.A1(new_n2152_), .A2(\A[27] ), .ZN(new_n2153_));
  INV_X1     g01151(.I(\A[27] ), .ZN(new_n2154_));
  NOR3_X1    g01152(.A1(new_n2150_), .A2(new_n2151_), .A3(new_n2154_), .ZN(new_n2155_));
  AOI21_X1   g01153(.A1(new_n2139_), .A2(new_n2140_), .B(\A[30] ), .ZN(new_n2156_));
  INV_X1     g01154(.I(\A[30] ), .ZN(new_n2157_));
  NOR2_X1    g01155(.A1(new_n2136_), .A2(\A[29] ), .ZN(new_n2158_));
  NOR2_X1    g01156(.A1(new_n2137_), .A2(\A[28] ), .ZN(new_n2159_));
  NOR3_X1    g01157(.A1(new_n2158_), .A2(new_n2159_), .A3(new_n2157_), .ZN(new_n2160_));
  OAI22_X1   g01158(.A1(new_n2153_), .A2(new_n2155_), .B1(new_n2160_), .B2(new_n2156_), .ZN(new_n2161_));
  NOR3_X1    g01159(.A1(new_n2161_), .A2(new_n2142_), .A3(new_n2149_), .ZN(new_n2162_));
  AOI21_X1   g01160(.A1(\A[25] ), .A2(new_n2144_), .B(new_n2154_), .ZN(new_n2163_));
  AOI22_X1   g01161(.A1(new_n2148_), .A2(new_n2154_), .B1(new_n2147_), .B2(new_n2163_), .ZN(new_n2164_));
  OAI21_X1   g01162(.A1(new_n2158_), .A2(new_n2159_), .B(new_n2157_), .ZN(new_n2165_));
  AOI21_X1   g01163(.A1(\A[28] ), .A2(new_n2137_), .B(new_n2157_), .ZN(new_n2166_));
  NAND2_X1   g01164(.A1(new_n2166_), .A2(new_n2140_), .ZN(new_n2167_));
  NAND2_X1   g01165(.A1(new_n2167_), .A2(new_n2165_), .ZN(new_n2168_));
  NOR2_X1    g01166(.A1(new_n2164_), .A2(new_n2168_), .ZN(new_n2169_));
  NAND2_X1   g01167(.A1(new_n2163_), .A2(new_n2147_), .ZN(new_n2170_));
  OAI21_X1   g01168(.A1(\A[27] ), .A2(new_n2152_), .B(new_n2170_), .ZN(new_n2171_));
  NOR2_X1    g01169(.A1(new_n2156_), .A2(new_n2160_), .ZN(new_n2172_));
  NOR2_X1    g01170(.A1(new_n2171_), .A2(new_n2172_), .ZN(new_n2173_));
  NOR2_X1    g01171(.A1(new_n2173_), .A2(new_n2169_), .ZN(new_n2174_));
  NOR2_X1    g01172(.A1(new_n2174_), .A2(new_n2162_), .ZN(new_n2175_));
  INV_X1     g01173(.I(\A[24] ), .ZN(new_n2176_));
  INV_X1     g01174(.I(\A[22] ), .ZN(new_n2177_));
  INV_X1     g01175(.I(\A[23] ), .ZN(new_n2178_));
  NOR2_X1    g01176(.A1(new_n2177_), .A2(new_n2178_), .ZN(new_n2179_));
  INV_X1     g01177(.I(new_n2179_), .ZN(new_n2180_));
  NOR2_X1    g01178(.A1(new_n2177_), .A2(\A[23] ), .ZN(new_n2181_));
  NOR2_X1    g01179(.A1(new_n2178_), .A2(\A[22] ), .ZN(new_n2182_));
  NOR2_X1    g01180(.A1(new_n2181_), .A2(new_n2182_), .ZN(new_n2183_));
  OAI21_X1   g01181(.A1(new_n2183_), .A2(new_n2176_), .B(new_n2180_), .ZN(new_n2184_));
  INV_X1     g01182(.I(\A[21] ), .ZN(new_n2185_));
  INV_X1     g01183(.I(\A[19] ), .ZN(new_n2186_));
  INV_X1     g01184(.I(\A[20] ), .ZN(new_n2187_));
  NOR2_X1    g01185(.A1(new_n2186_), .A2(new_n2187_), .ZN(new_n2188_));
  INV_X1     g01186(.I(new_n2188_), .ZN(new_n2189_));
  NOR2_X1    g01187(.A1(new_n2186_), .A2(\A[20] ), .ZN(new_n2190_));
  NOR2_X1    g01188(.A1(new_n2187_), .A2(\A[19] ), .ZN(new_n2191_));
  NOR2_X1    g01189(.A1(new_n2190_), .A2(new_n2191_), .ZN(new_n2192_));
  OAI21_X1   g01190(.A1(new_n2192_), .A2(new_n2185_), .B(new_n2189_), .ZN(new_n2193_));
  NAND2_X1   g01191(.A1(new_n2187_), .A2(\A[19] ), .ZN(new_n2194_));
  NAND2_X1   g01192(.A1(new_n2186_), .A2(\A[20] ), .ZN(new_n2195_));
  NAND2_X1   g01193(.A1(new_n2194_), .A2(new_n2195_), .ZN(new_n2196_));
  NAND2_X1   g01194(.A1(new_n2196_), .A2(new_n2185_), .ZN(new_n2197_));
  NAND3_X1   g01195(.A1(new_n2194_), .A2(new_n2195_), .A3(\A[21] ), .ZN(new_n2198_));
  OAI21_X1   g01196(.A1(new_n2181_), .A2(new_n2182_), .B(new_n2176_), .ZN(new_n2199_));
  NAND2_X1   g01197(.A1(new_n2177_), .A2(\A[23] ), .ZN(new_n2200_));
  AOI21_X1   g01198(.A1(\A[22] ), .A2(new_n2178_), .B(new_n2176_), .ZN(new_n2201_));
  NAND2_X1   g01199(.A1(new_n2201_), .A2(new_n2200_), .ZN(new_n2202_));
  AOI22_X1   g01200(.A1(new_n2197_), .A2(new_n2198_), .B1(new_n2199_), .B2(new_n2202_), .ZN(new_n2203_));
  NAND3_X1   g01201(.A1(new_n2203_), .A2(new_n2184_), .A3(new_n2193_), .ZN(new_n2204_));
  NOR2_X1    g01202(.A1(new_n2190_), .A2(new_n2185_), .ZN(new_n2205_));
  AOI22_X1   g01203(.A1(new_n2196_), .A2(new_n2185_), .B1(new_n2205_), .B2(new_n2195_), .ZN(new_n2206_));
  NAND2_X1   g01204(.A1(new_n2202_), .A2(new_n2199_), .ZN(new_n2207_));
  NAND2_X1   g01205(.A1(new_n2206_), .A2(new_n2207_), .ZN(new_n2208_));
  OAI21_X1   g01206(.A1(\A[21] ), .A2(new_n2192_), .B(new_n2198_), .ZN(new_n2209_));
  NAND2_X1   g01207(.A1(new_n2178_), .A2(\A[22] ), .ZN(new_n2210_));
  NAND2_X1   g01208(.A1(new_n2210_), .A2(new_n2200_), .ZN(new_n2211_));
  AOI22_X1   g01209(.A1(new_n2211_), .A2(new_n2176_), .B1(new_n2200_), .B2(new_n2201_), .ZN(new_n2212_));
  NAND2_X1   g01210(.A1(new_n2209_), .A2(new_n2212_), .ZN(new_n2213_));
  NAND2_X1   g01211(.A1(new_n2213_), .A2(new_n2208_), .ZN(new_n2214_));
  NAND2_X1   g01212(.A1(new_n2214_), .A2(new_n2204_), .ZN(new_n2215_));
  NAND2_X1   g01213(.A1(new_n2175_), .A2(new_n2215_), .ZN(new_n2216_));
  INV_X1     g01214(.I(new_n2138_), .ZN(new_n2217_));
  NOR2_X1    g01215(.A1(new_n2158_), .A2(new_n2159_), .ZN(new_n2218_));
  OAI21_X1   g01216(.A1(new_n2218_), .A2(new_n2157_), .B(new_n2217_), .ZN(new_n2219_));
  INV_X1     g01217(.I(new_n2145_), .ZN(new_n2220_));
  OAI21_X1   g01218(.A1(new_n2152_), .A2(new_n2154_), .B(new_n2220_), .ZN(new_n2221_));
  NAND2_X1   g01219(.A1(new_n2148_), .A2(new_n2154_), .ZN(new_n2222_));
  AOI22_X1   g01220(.A1(new_n2222_), .A2(new_n2170_), .B1(new_n2165_), .B2(new_n2167_), .ZN(new_n2223_));
  NAND3_X1   g01221(.A1(new_n2223_), .A2(new_n2219_), .A3(new_n2221_), .ZN(new_n2224_));
  NAND2_X1   g01222(.A1(new_n2171_), .A2(new_n2172_), .ZN(new_n2225_));
  NAND2_X1   g01223(.A1(new_n2164_), .A2(new_n2168_), .ZN(new_n2226_));
  NAND2_X1   g01224(.A1(new_n2225_), .A2(new_n2226_), .ZN(new_n2227_));
  NAND2_X1   g01225(.A1(new_n2227_), .A2(new_n2224_), .ZN(new_n2228_));
  AOI21_X1   g01226(.A1(new_n2211_), .A2(\A[24] ), .B(new_n2179_), .ZN(new_n2229_));
  AOI21_X1   g01227(.A1(new_n2196_), .A2(\A[21] ), .B(new_n2188_), .ZN(new_n2230_));
  NOR4_X1    g01228(.A1(new_n2206_), .A2(new_n2212_), .A3(new_n2229_), .A4(new_n2230_), .ZN(new_n2231_));
  NOR2_X1    g01229(.A1(new_n2209_), .A2(new_n2212_), .ZN(new_n2232_));
  NOR2_X1    g01230(.A1(new_n2206_), .A2(new_n2207_), .ZN(new_n2233_));
  NOR2_X1    g01231(.A1(new_n2232_), .A2(new_n2233_), .ZN(new_n2234_));
  NOR2_X1    g01232(.A1(new_n2234_), .A2(new_n2231_), .ZN(new_n2235_));
  NAND2_X1   g01233(.A1(new_n2235_), .A2(new_n2228_), .ZN(new_n2236_));
  NAND2_X1   g01234(.A1(new_n2216_), .A2(new_n2236_), .ZN(new_n2237_));
  INV_X1     g01235(.I(\A[18] ), .ZN(new_n2238_));
  INV_X1     g01236(.I(\A[16] ), .ZN(new_n2239_));
  INV_X1     g01237(.I(\A[17] ), .ZN(new_n2240_));
  NOR2_X1    g01238(.A1(new_n2239_), .A2(new_n2240_), .ZN(new_n2241_));
  INV_X1     g01239(.I(new_n2241_), .ZN(new_n2242_));
  NOR2_X1    g01240(.A1(new_n2239_), .A2(\A[17] ), .ZN(new_n2243_));
  NOR2_X1    g01241(.A1(new_n2240_), .A2(\A[16] ), .ZN(new_n2244_));
  NOR2_X1    g01242(.A1(new_n2243_), .A2(new_n2244_), .ZN(new_n2245_));
  OAI21_X1   g01243(.A1(new_n2245_), .A2(new_n2238_), .B(new_n2242_), .ZN(new_n2246_));
  INV_X1     g01244(.I(\A[15] ), .ZN(new_n2247_));
  INV_X1     g01245(.I(\A[13] ), .ZN(new_n2248_));
  INV_X1     g01246(.I(\A[14] ), .ZN(new_n2249_));
  NOR2_X1    g01247(.A1(new_n2248_), .A2(new_n2249_), .ZN(new_n2250_));
  INV_X1     g01248(.I(new_n2250_), .ZN(new_n2251_));
  NOR2_X1    g01249(.A1(new_n2248_), .A2(\A[14] ), .ZN(new_n2252_));
  NOR2_X1    g01250(.A1(new_n2249_), .A2(\A[13] ), .ZN(new_n2253_));
  NOR2_X1    g01251(.A1(new_n2252_), .A2(new_n2253_), .ZN(new_n2254_));
  OAI21_X1   g01252(.A1(new_n2254_), .A2(new_n2247_), .B(new_n2251_), .ZN(new_n2255_));
  NAND2_X1   g01253(.A1(new_n2249_), .A2(\A[13] ), .ZN(new_n2256_));
  NAND2_X1   g01254(.A1(new_n2248_), .A2(\A[14] ), .ZN(new_n2257_));
  NAND2_X1   g01255(.A1(new_n2256_), .A2(new_n2257_), .ZN(new_n2258_));
  NAND2_X1   g01256(.A1(new_n2258_), .A2(new_n2247_), .ZN(new_n2259_));
  NAND3_X1   g01257(.A1(new_n2256_), .A2(new_n2257_), .A3(\A[15] ), .ZN(new_n2260_));
  OAI21_X1   g01258(.A1(new_n2243_), .A2(new_n2244_), .B(new_n2238_), .ZN(new_n2261_));
  NAND2_X1   g01259(.A1(new_n2240_), .A2(\A[16] ), .ZN(new_n2262_));
  NAND2_X1   g01260(.A1(new_n2239_), .A2(\A[17] ), .ZN(new_n2263_));
  NAND3_X1   g01261(.A1(new_n2262_), .A2(new_n2263_), .A3(\A[18] ), .ZN(new_n2264_));
  AOI22_X1   g01262(.A1(new_n2259_), .A2(new_n2260_), .B1(new_n2261_), .B2(new_n2264_), .ZN(new_n2265_));
  NAND3_X1   g01263(.A1(new_n2265_), .A2(new_n2246_), .A3(new_n2255_), .ZN(new_n2266_));
  NAND2_X1   g01264(.A1(new_n2259_), .A2(new_n2260_), .ZN(new_n2267_));
  NAND2_X1   g01265(.A1(new_n2261_), .A2(new_n2264_), .ZN(new_n2268_));
  INV_X1     g01266(.I(new_n2268_), .ZN(new_n2269_));
  NAND2_X1   g01267(.A1(new_n2269_), .A2(new_n2267_), .ZN(new_n2270_));
  NOR2_X1    g01268(.A1(new_n2252_), .A2(new_n2247_), .ZN(new_n2271_));
  AOI22_X1   g01269(.A1(new_n2258_), .A2(new_n2247_), .B1(new_n2271_), .B2(new_n2257_), .ZN(new_n2272_));
  NAND2_X1   g01270(.A1(new_n2272_), .A2(new_n2268_), .ZN(new_n2273_));
  NAND2_X1   g01271(.A1(new_n2270_), .A2(new_n2273_), .ZN(new_n2274_));
  NAND2_X1   g01272(.A1(new_n2274_), .A2(new_n2266_), .ZN(new_n2275_));
  INV_X1     g01273(.I(\A[12] ), .ZN(new_n2276_));
  INV_X1     g01274(.I(\A[10] ), .ZN(new_n2277_));
  INV_X1     g01275(.I(\A[11] ), .ZN(new_n2278_));
  NOR2_X1    g01276(.A1(new_n2277_), .A2(new_n2278_), .ZN(new_n2279_));
  INV_X1     g01277(.I(new_n2279_), .ZN(new_n2280_));
  NOR2_X1    g01278(.A1(new_n2277_), .A2(\A[11] ), .ZN(new_n2281_));
  NOR2_X1    g01279(.A1(new_n2278_), .A2(\A[10] ), .ZN(new_n2282_));
  NOR2_X1    g01280(.A1(new_n2281_), .A2(new_n2282_), .ZN(new_n2283_));
  OAI21_X1   g01281(.A1(new_n2283_), .A2(new_n2276_), .B(new_n2280_), .ZN(new_n2284_));
  INV_X1     g01282(.I(\A[9] ), .ZN(new_n2285_));
  INV_X1     g01283(.I(\A[7] ), .ZN(new_n2286_));
  INV_X1     g01284(.I(\A[8] ), .ZN(new_n2287_));
  NOR2_X1    g01285(.A1(new_n2286_), .A2(new_n2287_), .ZN(new_n2288_));
  INV_X1     g01286(.I(new_n2288_), .ZN(new_n2289_));
  NOR2_X1    g01287(.A1(new_n2286_), .A2(\A[8] ), .ZN(new_n2290_));
  NOR2_X1    g01288(.A1(new_n2287_), .A2(\A[7] ), .ZN(new_n2291_));
  NOR2_X1    g01289(.A1(new_n2290_), .A2(new_n2291_), .ZN(new_n2292_));
  OAI21_X1   g01290(.A1(new_n2292_), .A2(new_n2285_), .B(new_n2289_), .ZN(new_n2293_));
  NAND2_X1   g01291(.A1(new_n2287_), .A2(\A[7] ), .ZN(new_n2294_));
  NAND2_X1   g01292(.A1(new_n2294_), .A2(\A[9] ), .ZN(new_n2295_));
  OAI22_X1   g01293(.A1(new_n2292_), .A2(\A[9] ), .B1(new_n2295_), .B2(new_n2291_), .ZN(new_n2296_));
  OAI21_X1   g01294(.A1(new_n2277_), .A2(\A[11] ), .B(\A[12] ), .ZN(new_n2297_));
  OAI22_X1   g01295(.A1(new_n2283_), .A2(\A[12] ), .B1(new_n2282_), .B2(new_n2297_), .ZN(new_n2298_));
  NAND4_X1   g01296(.A1(new_n2296_), .A2(new_n2298_), .A3(new_n2284_), .A4(new_n2293_), .ZN(new_n2299_));
  INV_X1     g01297(.I(new_n2299_), .ZN(new_n2300_));
  NAND2_X1   g01298(.A1(new_n2277_), .A2(\A[11] ), .ZN(new_n2301_));
  NAND2_X1   g01299(.A1(new_n2278_), .A2(\A[10] ), .ZN(new_n2302_));
  NAND2_X1   g01300(.A1(new_n2302_), .A2(new_n2301_), .ZN(new_n2303_));
  NOR2_X1    g01301(.A1(new_n2281_), .A2(new_n2276_), .ZN(new_n2304_));
  AOI22_X1   g01302(.A1(new_n2303_), .A2(new_n2276_), .B1(new_n2304_), .B2(new_n2301_), .ZN(new_n2305_));
  NOR2_X1    g01303(.A1(new_n2305_), .A2(new_n2296_), .ZN(new_n2306_));
  NAND2_X1   g01304(.A1(new_n2286_), .A2(\A[8] ), .ZN(new_n2307_));
  NAND2_X1   g01305(.A1(new_n2294_), .A2(new_n2307_), .ZN(new_n2308_));
  NOR2_X1    g01306(.A1(new_n2290_), .A2(new_n2285_), .ZN(new_n2309_));
  AOI22_X1   g01307(.A1(new_n2308_), .A2(new_n2285_), .B1(new_n2309_), .B2(new_n2307_), .ZN(new_n2310_));
  NOR2_X1    g01308(.A1(new_n2310_), .A2(new_n2298_), .ZN(new_n2311_));
  NOR2_X1    g01309(.A1(new_n2306_), .A2(new_n2311_), .ZN(new_n2312_));
  NOR2_X1    g01310(.A1(new_n2300_), .A2(new_n2312_), .ZN(new_n2313_));
  NAND2_X1   g01311(.A1(new_n2275_), .A2(new_n2313_), .ZN(new_n2314_));
  NAND2_X1   g01312(.A1(new_n2262_), .A2(new_n2263_), .ZN(new_n2315_));
  AOI21_X1   g01313(.A1(new_n2315_), .A2(\A[18] ), .B(new_n2241_), .ZN(new_n2316_));
  AOI21_X1   g01314(.A1(new_n2258_), .A2(\A[15] ), .B(new_n2250_), .ZN(new_n2317_));
  NOR4_X1    g01315(.A1(new_n2269_), .A2(new_n2316_), .A3(new_n2317_), .A4(new_n2272_), .ZN(new_n2318_));
  XOR2_X1    g01316(.A1(new_n2272_), .A2(new_n2268_), .Z(new_n2319_));
  NOR2_X1    g01317(.A1(new_n2319_), .A2(new_n2318_), .ZN(new_n2320_));
  NAND2_X1   g01318(.A1(new_n2310_), .A2(new_n2298_), .ZN(new_n2321_));
  NAND2_X1   g01319(.A1(new_n2305_), .A2(new_n2296_), .ZN(new_n2322_));
  NAND2_X1   g01320(.A1(new_n2322_), .A2(new_n2321_), .ZN(new_n2323_));
  NAND2_X1   g01321(.A1(new_n2323_), .A2(new_n2299_), .ZN(new_n2324_));
  NAND2_X1   g01322(.A1(new_n2320_), .A2(new_n2324_), .ZN(new_n2325_));
  NAND3_X1   g01323(.A1(new_n2237_), .A2(new_n2314_), .A3(new_n2325_), .ZN(new_n2326_));
  INV_X1     g01324(.I(new_n2326_), .ZN(new_n2327_));
  NOR2_X1    g01325(.A1(new_n2235_), .A2(new_n2228_), .ZN(new_n2328_));
  NOR2_X1    g01326(.A1(new_n2175_), .A2(new_n2215_), .ZN(new_n2329_));
  NOR2_X1    g01327(.A1(new_n2328_), .A2(new_n2329_), .ZN(new_n2330_));
  NAND2_X1   g01328(.A1(new_n2314_), .A2(new_n2325_), .ZN(new_n2331_));
  NAND2_X1   g01329(.A1(new_n2331_), .A2(new_n2330_), .ZN(new_n2332_));
  NAND2_X1   g01330(.A1(new_n2332_), .A2(new_n2326_), .ZN(new_n2333_));
  INV_X1     g01331(.I(new_n2333_), .ZN(new_n2334_));
  NAND2_X1   g01332(.A1(new_n2135_), .A2(new_n2332_), .ZN(new_n2335_));
  OAI22_X1   g01333(.A1(new_n2334_), .A2(new_n2135_), .B1(new_n2335_), .B2(new_n2327_), .ZN(new_n2336_));
  NOR2_X1    g01334(.A1(new_n2064_), .A2(new_n2336_), .ZN(new_n2337_));
  INV_X1     g01335(.I(new_n2064_), .ZN(new_n2338_));
  INV_X1     g01336(.I(new_n2336_), .ZN(new_n2339_));
  NOR2_X1    g01337(.A1(new_n2338_), .A2(new_n2339_), .ZN(new_n2340_));
  NOR2_X1    g01338(.A1(new_n2340_), .A2(new_n2337_), .ZN(new_n2341_));
  NOR2_X1    g01339(.A1(new_n2341_), .A2(new_n1724_), .ZN(new_n2342_));
  NOR3_X1    g01340(.A1(new_n2340_), .A2(new_n1723_), .A3(new_n2337_), .ZN(new_n2343_));
  NOR2_X1    g01341(.A1(new_n2342_), .A2(new_n2343_), .ZN(new_n2344_));
  NOR2_X1    g01342(.A1(new_n2344_), .A2(new_n1523_), .ZN(new_n2345_));
  INV_X1     g01343(.I(new_n2345_), .ZN(new_n2346_));
  XOR2_X1    g01344(.A1(new_n1716_), .A2(new_n1718_), .Z(new_n2347_));
  NOR2_X1    g01345(.A1(new_n1705_), .A2(new_n1713_), .ZN(new_n2348_));
  INV_X1     g01346(.I(new_n2348_), .ZN(new_n2349_));
  XOR2_X1    g01347(.A1(new_n2347_), .A2(new_n2349_), .Z(new_n2350_));
  XNOR2_X1   g01348(.A1(new_n1705_), .A2(new_n1713_), .ZN(new_n2351_));
  NOR2_X1    g01349(.A1(new_n1716_), .A2(new_n1718_), .ZN(new_n2352_));
  AOI21_X1   g01350(.A1(new_n2347_), .A2(new_n2348_), .B(new_n2352_), .ZN(new_n2353_));
  NOR2_X1    g01351(.A1(new_n2353_), .A2(new_n2351_), .ZN(new_n2354_));
  NOR2_X1    g01352(.A1(new_n2350_), .A2(new_n2354_), .ZN(new_n2355_));
  XOR2_X1    g01353(.A1(new_n1693_), .A2(new_n1695_), .Z(new_n2356_));
  NOR2_X1    g01354(.A1(new_n1682_), .A2(new_n1690_), .ZN(new_n2357_));
  NOR2_X1    g01355(.A1(new_n1693_), .A2(new_n1695_), .ZN(new_n2358_));
  AOI21_X1   g01356(.A1(new_n2356_), .A2(new_n2357_), .B(new_n2358_), .ZN(new_n2359_));
  XOR2_X1    g01357(.A1(new_n2356_), .A2(new_n2357_), .Z(new_n2360_));
  INV_X1     g01358(.I(new_n1691_), .ZN(new_n2361_));
  NOR2_X1    g01359(.A1(new_n2361_), .A2(new_n2351_), .ZN(new_n2362_));
  INV_X1     g01360(.I(new_n1719_), .ZN(new_n2363_));
  NOR2_X1    g01361(.A1(new_n2359_), .A2(new_n2361_), .ZN(new_n2364_));
  NOR2_X1    g01362(.A1(new_n2364_), .A2(new_n2363_), .ZN(new_n2365_));
  NAND4_X1   g01363(.A1(new_n2365_), .A2(new_n2359_), .A3(new_n2360_), .A4(new_n2362_), .ZN(new_n2366_));
  INV_X1     g01364(.I(new_n2366_), .ZN(new_n2367_));
  AND3_X2    g01365(.A1(new_n2362_), .A2(new_n1696_), .A3(new_n1719_), .Z(new_n2368_));
  XNOR2_X1   g01366(.A1(new_n2356_), .A2(new_n2357_), .ZN(new_n2369_));
  NOR2_X1    g01367(.A1(new_n2369_), .A2(new_n2364_), .ZN(new_n2370_));
  NOR2_X1    g01368(.A1(new_n2368_), .A2(new_n2370_), .ZN(new_n2371_));
  OAI21_X1   g01369(.A1(new_n2367_), .A2(new_n2371_), .B(new_n2355_), .ZN(new_n2372_));
  XOR2_X1    g01370(.A1(new_n2347_), .A2(new_n2348_), .Z(new_n2373_));
  OAI21_X1   g01371(.A1(new_n2351_), .A2(new_n2353_), .B(new_n2373_), .ZN(new_n2374_));
  OAI21_X1   g01372(.A1(new_n2361_), .A2(new_n2359_), .B(new_n2360_), .ZN(new_n2375_));
  NOR2_X1    g01373(.A1(new_n2375_), .A2(new_n2368_), .ZN(new_n2376_));
  NAND3_X1   g01374(.A1(new_n2362_), .A2(new_n1696_), .A3(new_n1719_), .ZN(new_n2377_));
  NOR2_X1    g01375(.A1(new_n2370_), .A2(new_n2377_), .ZN(new_n2378_));
  OAI21_X1   g01376(.A1(new_n2376_), .A2(new_n2378_), .B(new_n2374_), .ZN(new_n2379_));
  NAND2_X1   g01377(.A1(new_n2372_), .A2(new_n2379_), .ZN(new_n2380_));
  XOR2_X1    g01378(.A1(new_n1669_), .A2(new_n1671_), .Z(new_n2381_));
  NOR2_X1    g01379(.A1(new_n1666_), .A2(new_n1657_), .ZN(new_n2382_));
  INV_X1     g01380(.I(new_n2382_), .ZN(new_n2383_));
  XOR2_X1    g01381(.A1(new_n2381_), .A2(new_n2383_), .Z(new_n2384_));
  INV_X1     g01382(.I(new_n1667_), .ZN(new_n2385_));
  NOR2_X1    g01383(.A1(new_n1669_), .A2(new_n1671_), .ZN(new_n2386_));
  AOI21_X1   g01384(.A1(new_n2381_), .A2(new_n2382_), .B(new_n2386_), .ZN(new_n2387_));
  NOR2_X1    g01385(.A1(new_n2387_), .A2(new_n2385_), .ZN(new_n2388_));
  NOR2_X1    g01386(.A1(new_n2384_), .A2(new_n2388_), .ZN(new_n2389_));
  INV_X1     g01387(.I(new_n1648_), .ZN(new_n2390_));
  INV_X1     g01388(.I(new_n1672_), .ZN(new_n2391_));
  XOR2_X1    g01389(.A1(new_n1645_), .A2(new_n1647_), .Z(new_n2392_));
  NOR2_X1    g01390(.A1(new_n1633_), .A2(new_n1642_), .ZN(new_n2393_));
  XOR2_X1    g01391(.A1(new_n2392_), .A2(new_n2393_), .Z(new_n2394_));
  INV_X1     g01392(.I(new_n1643_), .ZN(new_n2395_));
  NOR2_X1    g01393(.A1(new_n2395_), .A2(new_n2385_), .ZN(new_n2396_));
  NAND2_X1   g01394(.A1(new_n2394_), .A2(new_n2396_), .ZN(new_n2397_));
  NOR2_X1    g01395(.A1(new_n1645_), .A2(new_n1647_), .ZN(new_n2398_));
  AOI21_X1   g01396(.A1(new_n2392_), .A2(new_n2393_), .B(new_n2398_), .ZN(new_n2399_));
  NOR2_X1    g01397(.A1(new_n2399_), .A2(new_n2395_), .ZN(new_n2400_));
  NOR4_X1    g01398(.A1(new_n2397_), .A2(new_n2390_), .A3(new_n2391_), .A4(new_n2400_), .ZN(new_n2401_));
  NOR4_X1    g01399(.A1(new_n2395_), .A2(new_n2385_), .A3(new_n2390_), .A4(new_n2391_), .ZN(new_n2402_));
  INV_X1     g01400(.I(new_n2393_), .ZN(new_n2403_));
  XOR2_X1    g01401(.A1(new_n2392_), .A2(new_n2403_), .Z(new_n2404_));
  NOR2_X1    g01402(.A1(new_n2404_), .A2(new_n2400_), .ZN(new_n2405_));
  NOR2_X1    g01403(.A1(new_n2405_), .A2(new_n2402_), .ZN(new_n2406_));
  OAI21_X1   g01404(.A1(new_n2401_), .A2(new_n2406_), .B(new_n2389_), .ZN(new_n2407_));
  XOR2_X1    g01405(.A1(new_n2381_), .A2(new_n2382_), .Z(new_n2408_));
  OAI21_X1   g01406(.A1(new_n2385_), .A2(new_n2387_), .B(new_n2408_), .ZN(new_n2409_));
  INV_X1     g01407(.I(new_n2402_), .ZN(new_n2410_));
  NOR2_X1    g01408(.A1(new_n2405_), .A2(new_n2410_), .ZN(new_n2411_));
  NOR3_X1    g01409(.A1(new_n2402_), .A2(new_n2404_), .A3(new_n2400_), .ZN(new_n2412_));
  OAI21_X1   g01410(.A1(new_n2411_), .A2(new_n2412_), .B(new_n2409_), .ZN(new_n2413_));
  NAND2_X1   g01411(.A1(new_n1674_), .A2(new_n1721_), .ZN(new_n2414_));
  INV_X1     g01412(.I(new_n2414_), .ZN(new_n2415_));
  NAND3_X1   g01413(.A1(new_n2407_), .A2(new_n2415_), .A3(new_n2413_), .ZN(new_n2416_));
  NAND2_X1   g01414(.A1(new_n2407_), .A2(new_n2413_), .ZN(new_n2417_));
  NAND2_X1   g01415(.A1(new_n2417_), .A2(new_n2414_), .ZN(new_n2418_));
  AOI21_X1   g01416(.A1(new_n2418_), .A2(new_n2416_), .B(new_n2380_), .ZN(new_n2419_));
  NAND2_X1   g01417(.A1(new_n2375_), .A2(new_n2377_), .ZN(new_n2420_));
  AOI21_X1   g01418(.A1(new_n2420_), .A2(new_n2366_), .B(new_n2374_), .ZN(new_n2421_));
  XNOR2_X1   g01419(.A1(new_n2370_), .A2(new_n2377_), .ZN(new_n2422_));
  AOI21_X1   g01420(.A1(new_n2422_), .A2(new_n2374_), .B(new_n2421_), .ZN(new_n2423_));
  NAND3_X1   g01421(.A1(new_n2407_), .A2(new_n2413_), .A3(new_n2414_), .ZN(new_n2424_));
  NOR2_X1    g01422(.A1(new_n2400_), .A2(new_n2391_), .ZN(new_n2425_));
  NAND4_X1   g01423(.A1(new_n2425_), .A2(new_n2399_), .A3(new_n2394_), .A4(new_n2396_), .ZN(new_n2426_));
  INV_X1     g01424(.I(new_n2406_), .ZN(new_n2427_));
  AOI21_X1   g01425(.A1(new_n2427_), .A2(new_n2426_), .B(new_n2409_), .ZN(new_n2428_));
  OAI21_X1   g01426(.A1(new_n2395_), .A2(new_n2399_), .B(new_n2394_), .ZN(new_n2429_));
  NAND2_X1   g01427(.A1(new_n2429_), .A2(new_n2402_), .ZN(new_n2430_));
  INV_X1     g01428(.I(new_n2412_), .ZN(new_n2431_));
  AOI21_X1   g01429(.A1(new_n2430_), .A2(new_n2431_), .B(new_n2389_), .ZN(new_n2432_));
  OAI21_X1   g01430(.A1(new_n2428_), .A2(new_n2432_), .B(new_n2415_), .ZN(new_n2433_));
  AOI21_X1   g01431(.A1(new_n2424_), .A2(new_n2433_), .B(new_n2423_), .ZN(new_n2434_));
  NOR2_X1    g01432(.A1(new_n2419_), .A2(new_n2434_), .ZN(new_n2435_));
  NOR2_X1    g01433(.A1(new_n1722_), .A2(new_n1624_), .ZN(new_n2436_));
  INV_X1     g01434(.I(new_n1616_), .ZN(new_n2437_));
  XOR2_X1    g01435(.A1(new_n1618_), .A2(new_n1620_), .Z(new_n2438_));
  NOR2_X1    g01436(.A1(new_n1607_), .A2(new_n1615_), .ZN(new_n2439_));
  NOR2_X1    g01437(.A1(new_n1618_), .A2(new_n1620_), .ZN(new_n2440_));
  AOI21_X1   g01438(.A1(new_n2438_), .A2(new_n2439_), .B(new_n2440_), .ZN(new_n2441_));
  XOR2_X1    g01439(.A1(new_n2438_), .A2(new_n2439_), .Z(new_n2442_));
  OAI21_X1   g01440(.A1(new_n2437_), .A2(new_n2441_), .B(new_n2442_), .ZN(new_n2443_));
  INV_X1     g01441(.I(new_n1597_), .ZN(new_n2444_));
  INV_X1     g01442(.I(new_n1621_), .ZN(new_n2445_));
  NAND2_X1   g01443(.A1(new_n1616_), .A2(new_n1598_), .ZN(new_n2446_));
  NOR3_X1    g01444(.A1(new_n2446_), .A2(new_n2444_), .A3(new_n2445_), .ZN(new_n2447_));
  INV_X1     g01445(.I(new_n2447_), .ZN(new_n2448_));
  INV_X1     g01446(.I(new_n1596_), .ZN(new_n2449_));
  XOR2_X1    g01447(.A1(new_n1580_), .A2(new_n1588_), .Z(new_n2450_));
  XOR2_X1    g01448(.A1(new_n2450_), .A2(new_n2449_), .Z(new_n2451_));
  NOR2_X1    g01449(.A1(new_n1580_), .A2(new_n1588_), .ZN(new_n2452_));
  AOI21_X1   g01450(.A1(new_n2450_), .A2(new_n1596_), .B(new_n2452_), .ZN(new_n2453_));
  INV_X1     g01451(.I(new_n1598_), .ZN(new_n2454_));
  NOR2_X1    g01452(.A1(new_n2453_), .A2(new_n2454_), .ZN(new_n2455_));
  NOR2_X1    g01453(.A1(new_n2451_), .A2(new_n2455_), .ZN(new_n2456_));
  NAND2_X1   g01454(.A1(new_n2456_), .A2(new_n2448_), .ZN(new_n2457_));
  INV_X1     g01455(.I(new_n2457_), .ZN(new_n2458_));
  NOR2_X1    g01456(.A1(new_n2456_), .A2(new_n2448_), .ZN(new_n2459_));
  OAI21_X1   g01457(.A1(new_n2458_), .A2(new_n2459_), .B(new_n2443_), .ZN(new_n2460_));
  INV_X1     g01458(.I(new_n2439_), .ZN(new_n2461_));
  XOR2_X1    g01459(.A1(new_n2438_), .A2(new_n2461_), .Z(new_n2462_));
  NOR2_X1    g01460(.A1(new_n2441_), .A2(new_n2437_), .ZN(new_n2463_));
  NOR2_X1    g01461(.A1(new_n2462_), .A2(new_n2463_), .ZN(new_n2464_));
  XOR2_X1    g01462(.A1(new_n2450_), .A2(new_n1596_), .Z(new_n2465_));
  INV_X1     g01463(.I(new_n2446_), .ZN(new_n2466_));
  NAND2_X1   g01464(.A1(new_n2465_), .A2(new_n2466_), .ZN(new_n2467_));
  NOR4_X1    g01465(.A1(new_n2467_), .A2(new_n2444_), .A3(new_n2445_), .A4(new_n2455_), .ZN(new_n2468_));
  NOR2_X1    g01466(.A1(new_n2456_), .A2(new_n2447_), .ZN(new_n2469_));
  OAI21_X1   g01467(.A1(new_n2468_), .A2(new_n2469_), .B(new_n2464_), .ZN(new_n2470_));
  NAND2_X1   g01468(.A1(new_n2460_), .A2(new_n2470_), .ZN(new_n2471_));
  XOR2_X1    g01469(.A1(new_n1568_), .A2(new_n1570_), .Z(new_n2472_));
  NOR2_X1    g01470(.A1(new_n1557_), .A2(new_n1565_), .ZN(new_n2473_));
  INV_X1     g01471(.I(new_n2473_), .ZN(new_n2474_));
  XOR2_X1    g01472(.A1(new_n2472_), .A2(new_n2474_), .Z(new_n2475_));
  INV_X1     g01473(.I(new_n1566_), .ZN(new_n2476_));
  NOR2_X1    g01474(.A1(new_n1568_), .A2(new_n1570_), .ZN(new_n2477_));
  AOI21_X1   g01475(.A1(new_n2472_), .A2(new_n2473_), .B(new_n2477_), .ZN(new_n2478_));
  NOR2_X1    g01476(.A1(new_n2478_), .A2(new_n2476_), .ZN(new_n2479_));
  NOR2_X1    g01477(.A1(new_n2475_), .A2(new_n2479_), .ZN(new_n2480_));
  INV_X1     g01478(.I(new_n1571_), .ZN(new_n2481_));
  XOR2_X1    g01479(.A1(new_n1530_), .A2(new_n1538_), .Z(new_n2482_));
  XOR2_X1    g01480(.A1(new_n2482_), .A2(new_n1546_), .Z(new_n2483_));
  INV_X1     g01481(.I(new_n1548_), .ZN(new_n2484_));
  NOR2_X1    g01482(.A1(new_n2484_), .A2(new_n2476_), .ZN(new_n2485_));
  NAND3_X1   g01483(.A1(new_n2483_), .A2(new_n2485_), .A3(new_n1547_), .ZN(new_n2486_));
  NOR2_X1    g01484(.A1(new_n1530_), .A2(new_n1538_), .ZN(new_n2487_));
  AOI21_X1   g01485(.A1(new_n2482_), .A2(new_n1546_), .B(new_n2487_), .ZN(new_n2488_));
  NOR2_X1    g01486(.A1(new_n2488_), .A2(new_n2484_), .ZN(new_n2489_));
  NOR3_X1    g01487(.A1(new_n2486_), .A2(new_n2481_), .A3(new_n2489_), .ZN(new_n2490_));
  AND4_X2    g01488(.A1(new_n1547_), .A2(new_n1548_), .A3(new_n1566_), .A4(new_n1571_), .Z(new_n2491_));
  INV_X1     g01489(.I(new_n1546_), .ZN(new_n2492_));
  XOR2_X1    g01490(.A1(new_n2482_), .A2(new_n2492_), .Z(new_n2493_));
  NOR2_X1    g01491(.A1(new_n2493_), .A2(new_n2489_), .ZN(new_n2494_));
  NOR2_X1    g01492(.A1(new_n2494_), .A2(new_n2491_), .ZN(new_n2495_));
  OAI21_X1   g01493(.A1(new_n2490_), .A2(new_n2495_), .B(new_n2480_), .ZN(new_n2496_));
  XOR2_X1    g01494(.A1(new_n2472_), .A2(new_n2473_), .Z(new_n2497_));
  XNOR2_X1   g01495(.A1(new_n1568_), .A2(new_n1570_), .ZN(new_n2498_));
  INV_X1     g01496(.I(new_n2477_), .ZN(new_n2499_));
  OAI21_X1   g01497(.A1(new_n2498_), .A2(new_n2474_), .B(new_n2499_), .ZN(new_n2500_));
  NAND2_X1   g01498(.A1(new_n2500_), .A2(new_n1566_), .ZN(new_n2501_));
  NAND2_X1   g01499(.A1(new_n2497_), .A2(new_n2501_), .ZN(new_n2502_));
  INV_X1     g01500(.I(new_n2487_), .ZN(new_n2503_));
  XNOR2_X1   g01501(.A1(new_n1530_), .A2(new_n1538_), .ZN(new_n2504_));
  OAI21_X1   g01502(.A1(new_n2504_), .A2(new_n2492_), .B(new_n2503_), .ZN(new_n2505_));
  NAND2_X1   g01503(.A1(new_n2505_), .A2(new_n1548_), .ZN(new_n2506_));
  NAND2_X1   g01504(.A1(new_n2483_), .A2(new_n2506_), .ZN(new_n2507_));
  NOR2_X1    g01505(.A1(new_n2507_), .A2(new_n2491_), .ZN(new_n2508_));
  INV_X1     g01506(.I(new_n2491_), .ZN(new_n2509_));
  NOR2_X1    g01507(.A1(new_n2494_), .A2(new_n2509_), .ZN(new_n2510_));
  OAI21_X1   g01508(.A1(new_n2510_), .A2(new_n2508_), .B(new_n2502_), .ZN(new_n2511_));
  NAND2_X1   g01509(.A1(new_n1573_), .A2(new_n1623_), .ZN(new_n2512_));
  INV_X1     g01510(.I(new_n2512_), .ZN(new_n2513_));
  NAND3_X1   g01511(.A1(new_n2496_), .A2(new_n2511_), .A3(new_n2513_), .ZN(new_n2514_));
  NOR2_X1    g01512(.A1(new_n2489_), .A2(new_n2481_), .ZN(new_n2515_));
  NAND4_X1   g01513(.A1(new_n2515_), .A2(new_n2488_), .A3(new_n2483_), .A4(new_n2485_), .ZN(new_n2516_));
  NAND2_X1   g01514(.A1(new_n2507_), .A2(new_n2509_), .ZN(new_n2517_));
  AOI21_X1   g01515(.A1(new_n2516_), .A2(new_n2517_), .B(new_n2502_), .ZN(new_n2518_));
  NAND2_X1   g01516(.A1(new_n2494_), .A2(new_n2509_), .ZN(new_n2519_));
  NAND2_X1   g01517(.A1(new_n2507_), .A2(new_n2491_), .ZN(new_n2520_));
  AOI21_X1   g01518(.A1(new_n2519_), .A2(new_n2520_), .B(new_n2480_), .ZN(new_n2521_));
  OAI21_X1   g01519(.A1(new_n2518_), .A2(new_n2521_), .B(new_n2512_), .ZN(new_n2522_));
  AOI21_X1   g01520(.A1(new_n2522_), .A2(new_n2514_), .B(new_n2471_), .ZN(new_n2523_));
  INV_X1     g01521(.I(new_n2456_), .ZN(new_n2524_));
  NAND2_X1   g01522(.A1(new_n2524_), .A2(new_n2447_), .ZN(new_n2525_));
  AOI21_X1   g01523(.A1(new_n2525_), .A2(new_n2457_), .B(new_n2464_), .ZN(new_n2526_));
  NOR2_X1    g01524(.A1(new_n2455_), .A2(new_n2445_), .ZN(new_n2527_));
  NAND4_X1   g01525(.A1(new_n2527_), .A2(new_n2453_), .A3(new_n2465_), .A4(new_n2466_), .ZN(new_n2528_));
  INV_X1     g01526(.I(new_n2469_), .ZN(new_n2529_));
  AOI21_X1   g01527(.A1(new_n2529_), .A2(new_n2528_), .B(new_n2443_), .ZN(new_n2530_));
  NOR2_X1    g01528(.A1(new_n2530_), .A2(new_n2526_), .ZN(new_n2531_));
  NAND3_X1   g01529(.A1(new_n2496_), .A2(new_n2511_), .A3(new_n2512_), .ZN(new_n2532_));
  OAI21_X1   g01530(.A1(new_n2518_), .A2(new_n2521_), .B(new_n2513_), .ZN(new_n2533_));
  AOI21_X1   g01531(.A1(new_n2532_), .A2(new_n2533_), .B(new_n2531_), .ZN(new_n2534_));
  NOR2_X1    g01532(.A1(new_n2534_), .A2(new_n2523_), .ZN(new_n2535_));
  NOR2_X1    g01533(.A1(new_n2535_), .A2(new_n2436_), .ZN(new_n2536_));
  INV_X1     g01534(.I(new_n2436_), .ZN(new_n2537_));
  NOR3_X1    g01535(.A1(new_n2534_), .A2(new_n2523_), .A3(new_n2537_), .ZN(new_n2538_));
  OAI21_X1   g01536(.A1(new_n2536_), .A2(new_n2538_), .B(new_n2435_), .ZN(new_n2539_));
  NOR2_X1    g01537(.A1(new_n2535_), .A2(new_n2537_), .ZN(new_n2540_));
  NOR3_X1    g01538(.A1(new_n2534_), .A2(new_n2523_), .A3(new_n2436_), .ZN(new_n2541_));
  OAI22_X1   g01539(.A1(new_n2540_), .A2(new_n2541_), .B1(new_n2419_), .B2(new_n2434_), .ZN(new_n2542_));
  NAND2_X1   g01540(.A1(new_n2542_), .A2(new_n2539_), .ZN(new_n2543_));
  INV_X1     g01541(.I(new_n2543_), .ZN(new_n2544_));
  XNOR2_X1   g01542(.A1(new_n2081_), .A2(new_n2072_), .ZN(new_n2545_));
  INV_X1     g01543(.I(new_n2545_), .ZN(new_n2546_));
  XOR2_X1    g01544(.A1(new_n2083_), .A2(new_n2085_), .Z(new_n2547_));
  NOR2_X1    g01545(.A1(new_n2081_), .A2(new_n2072_), .ZN(new_n2548_));
  NOR2_X1    g01546(.A1(new_n2083_), .A2(new_n2085_), .ZN(new_n2549_));
  AOI21_X1   g01547(.A1(new_n2547_), .A2(new_n2548_), .B(new_n2549_), .ZN(new_n2550_));
  INV_X1     g01548(.I(new_n2550_), .ZN(new_n2551_));
  XNOR2_X1   g01549(.A1(new_n2547_), .A2(new_n2548_), .ZN(new_n2552_));
  AOI21_X1   g01550(.A1(new_n2546_), .A2(new_n2551_), .B(new_n2552_), .ZN(new_n2553_));
  NAND2_X1   g01551(.A1(new_n2133_), .A2(new_n2086_), .ZN(new_n2554_));
  NOR2_X1    g01552(.A1(new_n2121_), .A2(new_n2117_), .ZN(new_n2555_));
  AOI21_X1   g01553(.A1(new_n2130_), .A2(\A[999] ), .B(new_n2555_), .ZN(new_n2556_));
  AOI21_X1   g01554(.A1(new_n2110_), .A2(new_n2116_), .B(new_n2131_), .ZN(new_n2557_));
  NOR2_X1    g01555(.A1(new_n2092_), .A2(new_n2090_), .ZN(new_n2558_));
  AOI21_X1   g01556(.A1(new_n2089_), .A2(\A[5] ), .B(new_n2558_), .ZN(new_n2559_));
  INV_X1     g01557(.I(new_n2559_), .ZN(new_n2560_));
  NAND2_X1   g01558(.A1(new_n2097_), .A2(new_n2099_), .ZN(new_n2561_));
  NOR2_X1    g01559(.A1(new_n2096_), .A2(new_n2098_), .ZN(new_n2562_));
  AOI21_X1   g01560(.A1(new_n2561_), .A2(\A[2] ), .B(new_n2562_), .ZN(new_n2563_));
  NOR2_X1    g01561(.A1(new_n2560_), .A2(new_n2563_), .ZN(new_n2564_));
  NOR2_X1    g01562(.A1(new_n2102_), .A2(new_n2103_), .ZN(new_n2565_));
  INV_X1     g01563(.I(new_n2562_), .ZN(new_n2566_));
  OAI21_X1   g01564(.A1(new_n2565_), .A2(new_n2101_), .B(new_n2566_), .ZN(new_n2567_));
  NOR2_X1    g01565(.A1(new_n2567_), .A2(new_n2559_), .ZN(new_n2568_));
  AOI21_X1   g01566(.A1(new_n2114_), .A2(new_n2115_), .B(new_n2095_), .ZN(new_n2569_));
  AOI21_X1   g01567(.A1(new_n2104_), .A2(new_n2100_), .B(new_n2106_), .ZN(new_n2570_));
  OAI22_X1   g01568(.A1(new_n2569_), .A2(new_n2570_), .B1(new_n2564_), .B2(new_n2568_), .ZN(new_n2571_));
  NAND2_X1   g01569(.A1(new_n2567_), .A2(new_n2559_), .ZN(new_n2572_));
  NAND2_X1   g01570(.A1(new_n2560_), .A2(new_n2563_), .ZN(new_n2573_));
  OAI21_X1   g01571(.A1(new_n2109_), .A2(new_n2105_), .B(new_n2113_), .ZN(new_n2574_));
  INV_X1     g01572(.I(new_n2570_), .ZN(new_n2575_));
  NAND4_X1   g01573(.A1(new_n2574_), .A2(new_n2573_), .A3(new_n2572_), .A4(new_n2575_), .ZN(new_n2576_));
  NAND3_X1   g01574(.A1(new_n2571_), .A2(new_n2557_), .A3(new_n2576_), .ZN(new_n2577_));
  OAI21_X1   g01575(.A1(new_n2129_), .A2(new_n2128_), .B(new_n2126_), .ZN(new_n2578_));
  AOI22_X1   g01576(.A1(new_n2574_), .A2(new_n2575_), .B1(new_n2573_), .B2(new_n2572_), .ZN(new_n2579_));
  NOR4_X1    g01577(.A1(new_n2569_), .A2(new_n2564_), .A3(new_n2568_), .A4(new_n2570_), .ZN(new_n2580_));
  OAI21_X1   g01578(.A1(new_n2580_), .A2(new_n2579_), .B(new_n2578_), .ZN(new_n2581_));
  AOI21_X1   g01579(.A1(new_n2581_), .A2(new_n2577_), .B(new_n2556_), .ZN(new_n2582_));
  INV_X1     g01580(.I(new_n2556_), .ZN(new_n2583_));
  NOR3_X1    g01581(.A1(new_n2579_), .A2(new_n2580_), .A3(new_n2578_), .ZN(new_n2584_));
  AOI21_X1   g01582(.A1(new_n2571_), .A2(new_n2576_), .B(new_n2557_), .ZN(new_n2585_));
  NOR3_X1    g01583(.A1(new_n2584_), .A2(new_n2585_), .A3(new_n2583_), .ZN(new_n2586_));
  OAI21_X1   g01584(.A1(new_n2586_), .A2(new_n2582_), .B(new_n2554_), .ZN(new_n2587_));
  INV_X1     g01585(.I(new_n2554_), .ZN(new_n2588_));
  OAI21_X1   g01586(.A1(new_n2584_), .A2(new_n2585_), .B(new_n2583_), .ZN(new_n2589_));
  NAND3_X1   g01587(.A1(new_n2581_), .A2(new_n2577_), .A3(new_n2556_), .ZN(new_n2590_));
  NAND3_X1   g01588(.A1(new_n2588_), .A2(new_n2589_), .A3(new_n2590_), .ZN(new_n2591_));
  AOI21_X1   g01589(.A1(new_n2591_), .A2(new_n2587_), .B(new_n2553_), .ZN(new_n2592_));
  XOR2_X1    g01590(.A1(new_n2547_), .A2(new_n2548_), .Z(new_n2593_));
  OAI21_X1   g01591(.A1(new_n2545_), .A2(new_n2550_), .B(new_n2593_), .ZN(new_n2594_));
  OAI21_X1   g01592(.A1(new_n2586_), .A2(new_n2582_), .B(new_n2588_), .ZN(new_n2595_));
  NAND3_X1   g01593(.A1(new_n2589_), .A2(new_n2590_), .A3(new_n2554_), .ZN(new_n2596_));
  AOI21_X1   g01594(.A1(new_n2595_), .A2(new_n2596_), .B(new_n2594_), .ZN(new_n2597_));
  NOR2_X1    g01595(.A1(new_n2592_), .A2(new_n2597_), .ZN(new_n2598_));
  INV_X1     g01596(.I(new_n2598_), .ZN(new_n2599_));
  NAND2_X1   g01597(.A1(new_n2333_), .A2(new_n2135_), .ZN(new_n2600_));
  AOI21_X1   g01598(.A1(new_n2308_), .A2(\A[9] ), .B(new_n2288_), .ZN(new_n2601_));
  NAND2_X1   g01599(.A1(new_n2284_), .A2(new_n2601_), .ZN(new_n2602_));
  AOI21_X1   g01600(.A1(new_n2303_), .A2(\A[12] ), .B(new_n2279_), .ZN(new_n2603_));
  NAND2_X1   g01601(.A1(new_n2293_), .A2(new_n2603_), .ZN(new_n2604_));
  NAND2_X1   g01602(.A1(new_n2296_), .A2(new_n2298_), .ZN(new_n2605_));
  AOI21_X1   g01603(.A1(new_n2602_), .A2(new_n2604_), .B(new_n2605_), .ZN(new_n2606_));
  NOR2_X1    g01604(.A1(new_n2603_), .A2(new_n2601_), .ZN(new_n2607_));
  NOR2_X1    g01605(.A1(new_n2606_), .A2(new_n2607_), .ZN(new_n2608_));
  NAND4_X1   g01606(.A1(new_n2602_), .A2(new_n2604_), .A3(new_n2296_), .A4(new_n2298_), .ZN(new_n2609_));
  NOR2_X1    g01607(.A1(new_n2293_), .A2(new_n2603_), .ZN(new_n2610_));
  NOR2_X1    g01608(.A1(new_n2284_), .A2(new_n2601_), .ZN(new_n2611_));
  OAI21_X1   g01609(.A1(new_n2610_), .A2(new_n2611_), .B(new_n2605_), .ZN(new_n2612_));
  NAND2_X1   g01610(.A1(new_n2612_), .A2(new_n2609_), .ZN(new_n2613_));
  OAI21_X1   g01611(.A1(new_n2608_), .A2(new_n2312_), .B(new_n2613_), .ZN(new_n2614_));
  NOR2_X1    g01612(.A1(new_n2246_), .A2(new_n2317_), .ZN(new_n2615_));
  NOR2_X1    g01613(.A1(new_n2255_), .A2(new_n2316_), .ZN(new_n2616_));
  NOR4_X1    g01614(.A1(new_n2615_), .A2(new_n2616_), .A3(new_n2272_), .A4(new_n2269_), .ZN(new_n2617_));
  NAND2_X1   g01615(.A1(new_n2255_), .A2(new_n2316_), .ZN(new_n2618_));
  NAND2_X1   g01616(.A1(new_n2246_), .A2(new_n2317_), .ZN(new_n2619_));
  AOI21_X1   g01617(.A1(new_n2618_), .A2(new_n2619_), .B(new_n2265_), .ZN(new_n2620_));
  NOR2_X1    g01618(.A1(new_n2617_), .A2(new_n2620_), .ZN(new_n2621_));
  NOR4_X1    g01619(.A1(new_n2319_), .A2(new_n2300_), .A3(new_n2312_), .A4(new_n2318_), .ZN(new_n2622_));
  NOR2_X1    g01620(.A1(new_n2316_), .A2(new_n2317_), .ZN(new_n2623_));
  NAND2_X1   g01621(.A1(new_n2618_), .A2(new_n2619_), .ZN(new_n2624_));
  AOI21_X1   g01622(.A1(new_n2624_), .A2(new_n2265_), .B(new_n2623_), .ZN(new_n2625_));
  NOR2_X1    g01623(.A1(new_n2625_), .A2(new_n2319_), .ZN(new_n2626_));
  NOR3_X1    g01624(.A1(new_n2626_), .A2(new_n2622_), .A3(new_n2621_), .ZN(new_n2627_));
  AOI22_X1   g01625(.A1(new_n2270_), .A2(new_n2273_), .B1(new_n2321_), .B2(new_n2322_), .ZN(new_n2628_));
  NAND3_X1   g01626(.A1(new_n2628_), .A2(new_n2266_), .A3(new_n2299_), .ZN(new_n2629_));
  INV_X1     g01627(.I(new_n2623_), .ZN(new_n2630_));
  OAI21_X1   g01628(.A1(new_n2615_), .A2(new_n2616_), .B(new_n2265_), .ZN(new_n2631_));
  NAND2_X1   g01629(.A1(new_n2631_), .A2(new_n2630_), .ZN(new_n2632_));
  NAND3_X1   g01630(.A1(new_n2618_), .A2(new_n2265_), .A3(new_n2619_), .ZN(new_n2633_));
  OAI22_X1   g01631(.A1(new_n2615_), .A2(new_n2616_), .B1(new_n2272_), .B2(new_n2269_), .ZN(new_n2634_));
  AOI22_X1   g01632(.A1(new_n2632_), .A2(new_n2274_), .B1(new_n2633_), .B2(new_n2634_), .ZN(new_n2635_));
  NOR2_X1    g01633(.A1(new_n2635_), .A2(new_n2629_), .ZN(new_n2636_));
  OAI21_X1   g01634(.A1(new_n2636_), .A2(new_n2627_), .B(new_n2614_), .ZN(new_n2637_));
  NOR2_X1    g01635(.A1(new_n2610_), .A2(new_n2611_), .ZN(new_n2638_));
  INV_X1     g01636(.I(new_n2607_), .ZN(new_n2639_));
  OAI21_X1   g01637(.A1(new_n2638_), .A2(new_n2605_), .B(new_n2639_), .ZN(new_n2640_));
  AOI22_X1   g01638(.A1(new_n2640_), .A2(new_n2323_), .B1(new_n2609_), .B2(new_n2612_), .ZN(new_n2641_));
  NAND2_X1   g01639(.A1(new_n2634_), .A2(new_n2633_), .ZN(new_n2642_));
  NAND3_X1   g01640(.A1(new_n2642_), .A2(new_n2266_), .A3(new_n2628_), .ZN(new_n2643_));
  OAI21_X1   g01641(.A1(new_n2625_), .A2(new_n2319_), .B(new_n2299_), .ZN(new_n2644_));
  NOR2_X1    g01642(.A1(new_n2643_), .A2(new_n2644_), .ZN(new_n2645_));
  NOR2_X1    g01643(.A1(new_n2635_), .A2(new_n2622_), .ZN(new_n2646_));
  OAI21_X1   g01644(.A1(new_n2646_), .A2(new_n2645_), .B(new_n2641_), .ZN(new_n2647_));
  NAND2_X1   g01645(.A1(new_n2647_), .A2(new_n2637_), .ZN(new_n2648_));
  NOR2_X1    g01646(.A1(new_n2193_), .A2(new_n2229_), .ZN(new_n2649_));
  NOR2_X1    g01647(.A1(new_n2184_), .A2(new_n2230_), .ZN(new_n2650_));
  OAI21_X1   g01648(.A1(new_n2649_), .A2(new_n2650_), .B(new_n2203_), .ZN(new_n2651_));
  NOR2_X1    g01649(.A1(new_n2229_), .A2(new_n2230_), .ZN(new_n2652_));
  INV_X1     g01650(.I(new_n2652_), .ZN(new_n2653_));
  NAND2_X1   g01651(.A1(new_n2651_), .A2(new_n2653_), .ZN(new_n2654_));
  NAND2_X1   g01652(.A1(new_n2184_), .A2(new_n2230_), .ZN(new_n2655_));
  NAND2_X1   g01653(.A1(new_n2193_), .A2(new_n2229_), .ZN(new_n2656_));
  NAND3_X1   g01654(.A1(new_n2655_), .A2(new_n2203_), .A3(new_n2656_), .ZN(new_n2657_));
  OAI22_X1   g01655(.A1(new_n2649_), .A2(new_n2650_), .B1(new_n2206_), .B2(new_n2212_), .ZN(new_n2658_));
  AOI22_X1   g01656(.A1(new_n2654_), .A2(new_n2214_), .B1(new_n2657_), .B2(new_n2658_), .ZN(new_n2659_));
  NAND2_X1   g01657(.A1(new_n2221_), .A2(new_n2142_), .ZN(new_n2660_));
  NAND2_X1   g01658(.A1(new_n2219_), .A2(new_n2149_), .ZN(new_n2661_));
  NAND3_X1   g01659(.A1(new_n2660_), .A2(new_n2223_), .A3(new_n2661_), .ZN(new_n2662_));
  NOR2_X1    g01660(.A1(new_n2219_), .A2(new_n2149_), .ZN(new_n2663_));
  NOR2_X1    g01661(.A1(new_n2221_), .A2(new_n2142_), .ZN(new_n2664_));
  OAI21_X1   g01662(.A1(new_n2663_), .A2(new_n2664_), .B(new_n2161_), .ZN(new_n2665_));
  NAND2_X1   g01663(.A1(new_n2665_), .A2(new_n2662_), .ZN(new_n2666_));
  NAND4_X1   g01664(.A1(new_n2666_), .A2(new_n2224_), .A3(new_n2227_), .A4(new_n2214_), .ZN(new_n2667_));
  NOR2_X1    g01665(.A1(new_n2142_), .A2(new_n2149_), .ZN(new_n2668_));
  AOI21_X1   g01666(.A1(new_n2660_), .A2(new_n2661_), .B(new_n2161_), .ZN(new_n2669_));
  OAI21_X1   g01667(.A1(new_n2669_), .A2(new_n2668_), .B(new_n2227_), .ZN(new_n2670_));
  NAND2_X1   g01668(.A1(new_n2670_), .A2(new_n2204_), .ZN(new_n2671_));
  NOR2_X1    g01669(.A1(new_n2667_), .A2(new_n2671_), .ZN(new_n2672_));
  OAI22_X1   g01670(.A1(new_n2169_), .A2(new_n2173_), .B1(new_n2232_), .B2(new_n2233_), .ZN(new_n2673_));
  NOR3_X1    g01671(.A1(new_n2673_), .A2(new_n2162_), .A3(new_n2231_), .ZN(new_n2674_));
  AOI21_X1   g01672(.A1(new_n2666_), .A2(new_n2670_), .B(new_n2674_), .ZN(new_n2675_));
  OAI21_X1   g01673(.A1(new_n2672_), .A2(new_n2675_), .B(new_n2659_), .ZN(new_n2676_));
  NAND2_X1   g01674(.A1(new_n2655_), .A2(new_n2656_), .ZN(new_n2677_));
  AOI21_X1   g01675(.A1(new_n2677_), .A2(new_n2203_), .B(new_n2652_), .ZN(new_n2678_));
  NOR4_X1    g01676(.A1(new_n2649_), .A2(new_n2650_), .A3(new_n2206_), .A4(new_n2212_), .ZN(new_n2679_));
  AOI21_X1   g01677(.A1(new_n2655_), .A2(new_n2656_), .B(new_n2203_), .ZN(new_n2680_));
  OAI22_X1   g01678(.A1(new_n2678_), .A2(new_n2234_), .B1(new_n2679_), .B2(new_n2680_), .ZN(new_n2681_));
  NOR3_X1    g01679(.A1(new_n2663_), .A2(new_n2161_), .A3(new_n2664_), .ZN(new_n2682_));
  AOI21_X1   g01680(.A1(new_n2660_), .A2(new_n2661_), .B(new_n2223_), .ZN(new_n2683_));
  NOR2_X1    g01681(.A1(new_n2683_), .A2(new_n2682_), .ZN(new_n2684_));
  INV_X1     g01682(.I(new_n2668_), .ZN(new_n2685_));
  OAI21_X1   g01683(.A1(new_n2663_), .A2(new_n2664_), .B(new_n2223_), .ZN(new_n2686_));
  AOI21_X1   g01684(.A1(new_n2685_), .A2(new_n2686_), .B(new_n2174_), .ZN(new_n2687_));
  NOR3_X1    g01685(.A1(new_n2674_), .A2(new_n2687_), .A3(new_n2684_), .ZN(new_n2688_));
  NAND4_X1   g01686(.A1(new_n2227_), .A2(new_n2214_), .A3(new_n2224_), .A4(new_n2204_), .ZN(new_n2689_));
  AOI21_X1   g01687(.A1(new_n2666_), .A2(new_n2670_), .B(new_n2689_), .ZN(new_n2690_));
  OAI21_X1   g01688(.A1(new_n2688_), .A2(new_n2690_), .B(new_n2681_), .ZN(new_n2691_));
  AOI22_X1   g01689(.A1(new_n2314_), .A2(new_n2325_), .B1(new_n2216_), .B2(new_n2236_), .ZN(new_n2692_));
  NAND3_X1   g01690(.A1(new_n2676_), .A2(new_n2691_), .A3(new_n2692_), .ZN(new_n2693_));
  NOR3_X1    g01691(.A1(new_n2684_), .A2(new_n2162_), .A3(new_n2673_), .ZN(new_n2694_));
  NAND2_X1   g01692(.A1(new_n2686_), .A2(new_n2685_), .ZN(new_n2695_));
  AOI21_X1   g01693(.A1(new_n2695_), .A2(new_n2227_), .B(new_n2231_), .ZN(new_n2696_));
  NAND2_X1   g01694(.A1(new_n2694_), .A2(new_n2696_), .ZN(new_n2697_));
  NAND2_X1   g01695(.A1(new_n2670_), .A2(new_n2666_), .ZN(new_n2698_));
  NAND2_X1   g01696(.A1(new_n2698_), .A2(new_n2689_), .ZN(new_n2699_));
  AOI21_X1   g01697(.A1(new_n2697_), .A2(new_n2699_), .B(new_n2681_), .ZN(new_n2700_));
  NAND3_X1   g01698(.A1(new_n2689_), .A2(new_n2670_), .A3(new_n2666_), .ZN(new_n2701_));
  NAND2_X1   g01699(.A1(new_n2698_), .A2(new_n2674_), .ZN(new_n2702_));
  AOI21_X1   g01700(.A1(new_n2702_), .A2(new_n2701_), .B(new_n2659_), .ZN(new_n2703_));
  NOR2_X1    g01701(.A1(new_n2320_), .A2(new_n2324_), .ZN(new_n2704_));
  NOR2_X1    g01702(.A1(new_n2275_), .A2(new_n2313_), .ZN(new_n2705_));
  OAI22_X1   g01703(.A1(new_n2705_), .A2(new_n2704_), .B1(new_n2328_), .B2(new_n2329_), .ZN(new_n2706_));
  OAI21_X1   g01704(.A1(new_n2700_), .A2(new_n2703_), .B(new_n2706_), .ZN(new_n2707_));
  AOI21_X1   g01705(.A1(new_n2707_), .A2(new_n2693_), .B(new_n2648_), .ZN(new_n2708_));
  NAND2_X1   g01706(.A1(new_n2635_), .A2(new_n2629_), .ZN(new_n2709_));
  OAI21_X1   g01707(.A1(new_n2625_), .A2(new_n2319_), .B(new_n2642_), .ZN(new_n2710_));
  NAND2_X1   g01708(.A1(new_n2710_), .A2(new_n2622_), .ZN(new_n2711_));
  AOI21_X1   g01709(.A1(new_n2711_), .A2(new_n2709_), .B(new_n2641_), .ZN(new_n2712_));
  AOI21_X1   g01710(.A1(new_n2632_), .A2(new_n2274_), .B(new_n2300_), .ZN(new_n2713_));
  NAND4_X1   g01711(.A1(new_n2713_), .A2(new_n2625_), .A3(new_n2642_), .A4(new_n2628_), .ZN(new_n2714_));
  OAI21_X1   g01712(.A1(new_n2626_), .A2(new_n2621_), .B(new_n2629_), .ZN(new_n2715_));
  AOI21_X1   g01713(.A1(new_n2714_), .A2(new_n2715_), .B(new_n2614_), .ZN(new_n2716_));
  NOR2_X1    g01714(.A1(new_n2712_), .A2(new_n2716_), .ZN(new_n2717_));
  NAND3_X1   g01715(.A1(new_n2676_), .A2(new_n2691_), .A3(new_n2706_), .ZN(new_n2718_));
  OAI21_X1   g01716(.A1(new_n2700_), .A2(new_n2703_), .B(new_n2692_), .ZN(new_n2719_));
  AOI21_X1   g01717(.A1(new_n2718_), .A2(new_n2719_), .B(new_n2717_), .ZN(new_n2720_));
  OAI21_X1   g01718(.A1(new_n2720_), .A2(new_n2708_), .B(new_n2600_), .ZN(new_n2721_));
  INV_X1     g01719(.I(new_n2600_), .ZN(new_n2722_));
  NOR3_X1    g01720(.A1(new_n2700_), .A2(new_n2703_), .A3(new_n2706_), .ZN(new_n2723_));
  AOI21_X1   g01721(.A1(new_n2676_), .A2(new_n2691_), .B(new_n2692_), .ZN(new_n2724_));
  OAI21_X1   g01722(.A1(new_n2723_), .A2(new_n2724_), .B(new_n2717_), .ZN(new_n2725_));
  NOR3_X1    g01723(.A1(new_n2700_), .A2(new_n2703_), .A3(new_n2692_), .ZN(new_n2726_));
  AOI21_X1   g01724(.A1(new_n2676_), .A2(new_n2691_), .B(new_n2706_), .ZN(new_n2727_));
  OAI21_X1   g01725(.A1(new_n2727_), .A2(new_n2726_), .B(new_n2648_), .ZN(new_n2728_));
  NAND3_X1   g01726(.A1(new_n2722_), .A2(new_n2725_), .A3(new_n2728_), .ZN(new_n2729_));
  AOI21_X1   g01727(.A1(new_n2729_), .A2(new_n2721_), .B(new_n2599_), .ZN(new_n2730_));
  OAI21_X1   g01728(.A1(new_n2720_), .A2(new_n2708_), .B(new_n2722_), .ZN(new_n2731_));
  NAND3_X1   g01729(.A1(new_n2725_), .A2(new_n2728_), .A3(new_n2600_), .ZN(new_n2732_));
  AOI21_X1   g01730(.A1(new_n2731_), .A2(new_n2732_), .B(new_n2598_), .ZN(new_n2733_));
  NOR2_X1    g01731(.A1(new_n2730_), .A2(new_n2733_), .ZN(new_n2734_));
  INV_X1     g01732(.I(new_n2040_), .ZN(new_n2735_));
  NOR2_X1    g01733(.A1(new_n2039_), .A2(\A[31] ), .ZN(new_n2736_));
  NOR2_X1    g01734(.A1(new_n2046_), .A2(new_n2736_), .ZN(new_n2737_));
  OAI21_X1   g01735(.A1(new_n2737_), .A2(new_n2045_), .B(new_n2735_), .ZN(new_n2738_));
  NOR2_X1    g01736(.A1(new_n2738_), .A2(new_n2037_), .ZN(new_n2739_));
  INV_X1     g01737(.I(new_n2033_), .ZN(new_n2740_));
  XNOR2_X1   g01738(.A1(\A[34] ), .A2(\A[35] ), .ZN(new_n2741_));
  OAI21_X1   g01739(.A1(new_n2741_), .A2(new_n2049_), .B(new_n2740_), .ZN(new_n2742_));
  NOR2_X1    g01740(.A1(new_n2742_), .A2(new_n2044_), .ZN(new_n2743_));
  NOR2_X1    g01741(.A1(new_n2048_), .A2(new_n2051_), .ZN(new_n2744_));
  OAI21_X1   g01742(.A1(new_n2739_), .A2(new_n2743_), .B(new_n2744_), .ZN(new_n2745_));
  NOR2_X1    g01743(.A1(new_n2037_), .A2(new_n2044_), .ZN(new_n2746_));
  INV_X1     g01744(.I(new_n2746_), .ZN(new_n2747_));
  NAND2_X1   g01745(.A1(new_n2745_), .A2(new_n2747_), .ZN(new_n2748_));
  NOR4_X1    g01746(.A1(new_n2739_), .A2(new_n2743_), .A3(new_n2048_), .A4(new_n2051_), .ZN(new_n2749_));
  NAND2_X1   g01747(.A1(new_n2742_), .A2(new_n2044_), .ZN(new_n2750_));
  NAND2_X1   g01748(.A1(new_n2738_), .A2(new_n2037_), .ZN(new_n2751_));
  AOI21_X1   g01749(.A1(new_n2750_), .A2(new_n2751_), .B(new_n2744_), .ZN(new_n2752_));
  NOR2_X1    g01750(.A1(new_n2752_), .A2(new_n2749_), .ZN(new_n2753_));
  AOI21_X1   g01751(.A1(new_n2748_), .A2(new_n2057_), .B(new_n2753_), .ZN(new_n2754_));
  AOI21_X1   g01752(.A1(new_n2019_), .A2(\A[39] ), .B(new_n2011_), .ZN(new_n2755_));
  NAND2_X1   g01753(.A1(new_n2007_), .A2(new_n2755_), .ZN(new_n2756_));
  AOI21_X1   g01754(.A1(new_n2024_), .A2(\A[42] ), .B(new_n2002_), .ZN(new_n2757_));
  NAND2_X1   g01755(.A1(new_n2016_), .A2(new_n2757_), .ZN(new_n2758_));
  NAND3_X1   g01756(.A1(new_n2027_), .A2(new_n2756_), .A3(new_n2758_), .ZN(new_n2759_));
  NOR2_X1    g01757(.A1(new_n2016_), .A2(new_n2757_), .ZN(new_n2760_));
  NOR2_X1    g01758(.A1(new_n2007_), .A2(new_n2755_), .ZN(new_n2761_));
  NAND2_X1   g01759(.A1(new_n2018_), .A2(\A[39] ), .ZN(new_n2762_));
  OAI22_X1   g01760(.A1(new_n2015_), .A2(\A[39] ), .B1(new_n2762_), .B2(new_n2014_), .ZN(new_n2763_));
  NAND2_X1   g01761(.A1(new_n2023_), .A2(\A[42] ), .ZN(new_n2764_));
  OAI22_X1   g01762(.A1(new_n2006_), .A2(\A[42] ), .B1(new_n2764_), .B2(new_n2005_), .ZN(new_n2765_));
  NAND2_X1   g01763(.A1(new_n2763_), .A2(new_n2765_), .ZN(new_n2766_));
  OAI21_X1   g01764(.A1(new_n2760_), .A2(new_n2761_), .B(new_n2766_), .ZN(new_n2767_));
  NAND2_X1   g01765(.A1(new_n2767_), .A2(new_n2759_), .ZN(new_n2768_));
  NAND4_X1   g01766(.A1(new_n2029_), .A2(new_n2057_), .A3(new_n2028_), .A4(new_n2056_), .ZN(new_n2769_));
  AOI21_X1   g01767(.A1(new_n2756_), .A2(new_n2758_), .B(new_n2766_), .ZN(new_n2770_));
  NOR2_X1    g01768(.A1(new_n2757_), .A2(new_n2755_), .ZN(new_n2771_));
  OAI21_X1   g01769(.A1(new_n2770_), .A2(new_n2771_), .B(new_n2029_), .ZN(new_n2772_));
  NAND3_X1   g01770(.A1(new_n2769_), .A2(new_n2772_), .A3(new_n2768_), .ZN(new_n2773_));
  NOR3_X1    g01771(.A1(new_n2766_), .A2(new_n2757_), .A3(new_n2755_), .ZN(new_n2774_));
  XOR2_X1    g01772(.A1(new_n2763_), .A2(new_n2026_), .Z(new_n2775_));
  NOR4_X1    g01773(.A1(new_n2053_), .A2(new_n2775_), .A3(new_n2774_), .A4(new_n2052_), .ZN(new_n2776_));
  NAND2_X1   g01774(.A1(new_n2772_), .A2(new_n2768_), .ZN(new_n2777_));
  NAND2_X1   g01775(.A1(new_n2777_), .A2(new_n2776_), .ZN(new_n2778_));
  AOI21_X1   g01776(.A1(new_n2778_), .A2(new_n2773_), .B(new_n2754_), .ZN(new_n2779_));
  NAND2_X1   g01777(.A1(new_n2750_), .A2(new_n2751_), .ZN(new_n2780_));
  AOI21_X1   g01778(.A1(new_n2780_), .A2(new_n2744_), .B(new_n2746_), .ZN(new_n2781_));
  NAND3_X1   g01779(.A1(new_n2744_), .A2(new_n2750_), .A3(new_n2751_), .ZN(new_n2782_));
  OAI22_X1   g01780(.A1(new_n2739_), .A2(new_n2743_), .B1(new_n2048_), .B2(new_n2051_), .ZN(new_n2783_));
  NAND2_X1   g01781(.A1(new_n2783_), .A2(new_n2782_), .ZN(new_n2784_));
  OAI21_X1   g01782(.A1(new_n2781_), .A2(new_n2053_), .B(new_n2784_), .ZN(new_n2785_));
  NAND2_X1   g01783(.A1(new_n2777_), .A2(new_n2769_), .ZN(new_n2786_));
  NOR3_X1    g01784(.A1(new_n2766_), .A2(new_n2760_), .A3(new_n2761_), .ZN(new_n2787_));
  AOI21_X1   g01785(.A1(new_n2756_), .A2(new_n2758_), .B(new_n2027_), .ZN(new_n2788_));
  NOR2_X1    g01786(.A1(new_n2788_), .A2(new_n2787_), .ZN(new_n2789_));
  NOR4_X1    g01787(.A1(new_n2789_), .A2(new_n2774_), .A3(new_n2775_), .A4(new_n2053_), .ZN(new_n2790_));
  NOR2_X1    g01788(.A1(new_n2760_), .A2(new_n2761_), .ZN(new_n2791_));
  INV_X1     g01789(.I(new_n2771_), .ZN(new_n2792_));
  OAI21_X1   g01790(.A1(new_n2791_), .A2(new_n2766_), .B(new_n2792_), .ZN(new_n2793_));
  AOI21_X1   g01791(.A1(new_n2793_), .A2(new_n2029_), .B(new_n2052_), .ZN(new_n2794_));
  NAND2_X1   g01792(.A1(new_n2790_), .A2(new_n2794_), .ZN(new_n2795_));
  AOI21_X1   g01793(.A1(new_n2786_), .A2(new_n2795_), .B(new_n2785_), .ZN(new_n2796_));
  NOR2_X1    g01794(.A1(new_n2796_), .A2(new_n2779_), .ZN(new_n2797_));
  NAND2_X1   g01795(.A1(new_n1965_), .A2(\A[44] ), .ZN(new_n2798_));
  NAND2_X1   g01796(.A1(new_n1973_), .A2(new_n2798_), .ZN(new_n2799_));
  AOI21_X1   g01797(.A1(new_n2799_), .A2(\A[45] ), .B(new_n1967_), .ZN(new_n2800_));
  NAND2_X1   g01798(.A1(new_n1963_), .A2(new_n2800_), .ZN(new_n2801_));
  NAND2_X1   g01799(.A1(new_n1977_), .A2(new_n1978_), .ZN(new_n2802_));
  AOI21_X1   g01800(.A1(new_n2802_), .A2(\A[48] ), .B(new_n1958_), .ZN(new_n2803_));
  NAND2_X1   g01801(.A1(new_n1972_), .A2(new_n2803_), .ZN(new_n2804_));
  NAND2_X1   g01802(.A1(new_n1975_), .A2(new_n1980_), .ZN(new_n2805_));
  AOI21_X1   g01803(.A1(new_n2801_), .A2(new_n2804_), .B(new_n2805_), .ZN(new_n2806_));
  NOR2_X1    g01804(.A1(new_n2803_), .A2(new_n2800_), .ZN(new_n2807_));
  NOR2_X1    g01805(.A1(new_n2806_), .A2(new_n2807_), .ZN(new_n2808_));
  NAND4_X1   g01806(.A1(new_n2801_), .A2(new_n2804_), .A3(new_n1975_), .A4(new_n1980_), .ZN(new_n2809_));
  NOR2_X1    g01807(.A1(new_n1972_), .A2(new_n2803_), .ZN(new_n2810_));
  NOR2_X1    g01808(.A1(new_n1963_), .A2(new_n2800_), .ZN(new_n2811_));
  OAI21_X1   g01809(.A1(new_n2810_), .A2(new_n2811_), .B(new_n2805_), .ZN(new_n2812_));
  NAND2_X1   g01810(.A1(new_n2812_), .A2(new_n2809_), .ZN(new_n2813_));
  OAI21_X1   g01811(.A1(new_n2808_), .A2(new_n1995_), .B(new_n2813_), .ZN(new_n2814_));
  NOR2_X1    g01812(.A1(new_n1987_), .A2(new_n1935_), .ZN(new_n2815_));
  NOR2_X1    g01813(.A1(new_n1989_), .A2(new_n1928_), .ZN(new_n2816_));
  NOR3_X1    g01814(.A1(new_n1947_), .A2(new_n2815_), .A3(new_n2816_), .ZN(new_n2817_));
  NAND2_X1   g01815(.A1(new_n1989_), .A2(new_n1928_), .ZN(new_n2818_));
  NAND2_X1   g01816(.A1(new_n1987_), .A2(new_n1935_), .ZN(new_n2819_));
  AOI21_X1   g01817(.A1(new_n2818_), .A2(new_n2819_), .B(new_n1990_), .ZN(new_n2820_));
  NOR2_X1    g01818(.A1(new_n2820_), .A2(new_n2817_), .ZN(new_n2821_));
  NAND4_X1   g01819(.A1(new_n1992_), .A2(new_n1982_), .A3(new_n1991_), .A4(new_n1981_), .ZN(new_n2822_));
  NOR2_X1    g01820(.A1(new_n1928_), .A2(new_n1935_), .ZN(new_n2823_));
  NAND2_X1   g01821(.A1(new_n2818_), .A2(new_n2819_), .ZN(new_n2824_));
  AOI21_X1   g01822(.A1(new_n2824_), .A2(new_n1990_), .B(new_n2823_), .ZN(new_n2825_));
  NOR2_X1    g01823(.A1(new_n2825_), .A2(new_n1953_), .ZN(new_n2826_));
  OAI21_X1   g01824(.A1(new_n2826_), .A2(new_n2821_), .B(new_n2822_), .ZN(new_n2827_));
  NAND3_X1   g01825(.A1(new_n2818_), .A2(new_n1990_), .A3(new_n2819_), .ZN(new_n2828_));
  OAI21_X1   g01826(.A1(new_n2815_), .A2(new_n2816_), .B(new_n1947_), .ZN(new_n2829_));
  NAND2_X1   g01827(.A1(new_n2829_), .A2(new_n2828_), .ZN(new_n2830_));
  NOR2_X1    g01828(.A1(new_n1995_), .A2(new_n1953_), .ZN(new_n2831_));
  INV_X1     g01829(.I(new_n2823_), .ZN(new_n2832_));
  NOR2_X1    g01830(.A1(new_n2815_), .A2(new_n2816_), .ZN(new_n2833_));
  OAI21_X1   g01831(.A1(new_n2833_), .A2(new_n1947_), .B(new_n2832_), .ZN(new_n2834_));
  AOI21_X1   g01832(.A1(new_n2834_), .A2(new_n1992_), .B(new_n1994_), .ZN(new_n2835_));
  NAND4_X1   g01833(.A1(new_n2835_), .A2(new_n2825_), .A3(new_n2830_), .A4(new_n2831_), .ZN(new_n2836_));
  AOI21_X1   g01834(.A1(new_n2836_), .A2(new_n2827_), .B(new_n2814_), .ZN(new_n2837_));
  NOR2_X1    g01835(.A1(new_n2810_), .A2(new_n2811_), .ZN(new_n2838_));
  INV_X1     g01836(.I(new_n2807_), .ZN(new_n2839_));
  OAI21_X1   g01837(.A1(new_n2838_), .A2(new_n2805_), .B(new_n2839_), .ZN(new_n2840_));
  NOR3_X1    g01838(.A1(new_n2810_), .A2(new_n2805_), .A3(new_n2811_), .ZN(new_n2841_));
  AOI22_X1   g01839(.A1(new_n2801_), .A2(new_n2804_), .B1(new_n1975_), .B2(new_n1980_), .ZN(new_n2842_));
  NOR2_X1    g01840(.A1(new_n2842_), .A2(new_n2841_), .ZN(new_n2843_));
  AOI21_X1   g01841(.A1(new_n2840_), .A2(new_n1982_), .B(new_n2843_), .ZN(new_n2844_));
  AOI22_X1   g01842(.A1(new_n2834_), .A2(new_n1992_), .B1(new_n2828_), .B2(new_n2829_), .ZN(new_n2845_));
  NAND2_X1   g01843(.A1(new_n2845_), .A2(new_n2822_), .ZN(new_n2846_));
  NOR4_X1    g01844(.A1(new_n1995_), .A2(new_n1953_), .A3(new_n1994_), .A4(new_n1948_), .ZN(new_n2847_));
  OAI21_X1   g01845(.A1(new_n2826_), .A2(new_n2821_), .B(new_n2847_), .ZN(new_n2848_));
  AOI21_X1   g01846(.A1(new_n2846_), .A2(new_n2848_), .B(new_n2844_), .ZN(new_n2849_));
  NAND2_X1   g01847(.A1(new_n2061_), .A2(new_n1998_), .ZN(new_n2850_));
  NOR3_X1    g01848(.A1(new_n2837_), .A2(new_n2850_), .A3(new_n2849_), .ZN(new_n2851_));
  NOR2_X1    g01849(.A1(new_n2845_), .A2(new_n2847_), .ZN(new_n2852_));
  NAND3_X1   g01850(.A1(new_n2831_), .A2(new_n2830_), .A3(new_n1991_), .ZN(new_n2853_));
  OAI21_X1   g01851(.A1(new_n2825_), .A2(new_n1953_), .B(new_n1981_), .ZN(new_n2854_));
  NOR2_X1    g01852(.A1(new_n2853_), .A2(new_n2854_), .ZN(new_n2855_));
  OAI21_X1   g01853(.A1(new_n2855_), .A2(new_n2852_), .B(new_n2844_), .ZN(new_n2856_));
  NOR3_X1    g01854(.A1(new_n2826_), .A2(new_n2847_), .A3(new_n2821_), .ZN(new_n2857_));
  NOR2_X1    g01855(.A1(new_n2845_), .A2(new_n2822_), .ZN(new_n2858_));
  OAI21_X1   g01856(.A1(new_n2858_), .A2(new_n2857_), .B(new_n2814_), .ZN(new_n2859_));
  AOI22_X1   g01857(.A1(new_n2055_), .A2(new_n2059_), .B1(new_n1997_), .B2(new_n1984_), .ZN(new_n2860_));
  AOI21_X1   g01858(.A1(new_n2856_), .A2(new_n2859_), .B(new_n2860_), .ZN(new_n2861_));
  OAI21_X1   g01859(.A1(new_n2851_), .A2(new_n2861_), .B(new_n2797_), .ZN(new_n2862_));
  NOR2_X1    g01860(.A1(new_n2770_), .A2(new_n2771_), .ZN(new_n2863_));
  NOR2_X1    g01861(.A1(new_n2863_), .A2(new_n2775_), .ZN(new_n2864_));
  NOR3_X1    g01862(.A1(new_n2864_), .A2(new_n2789_), .A3(new_n2776_), .ZN(new_n2865_));
  AOI21_X1   g01863(.A1(new_n2768_), .A2(new_n2772_), .B(new_n2769_), .ZN(new_n2866_));
  OAI21_X1   g01864(.A1(new_n2865_), .A2(new_n2866_), .B(new_n2785_), .ZN(new_n2867_));
  AOI21_X1   g01865(.A1(new_n2768_), .A2(new_n2772_), .B(new_n2776_), .ZN(new_n2868_));
  NAND4_X1   g01866(.A1(new_n2768_), .A2(new_n2028_), .A3(new_n2029_), .A4(new_n2057_), .ZN(new_n2869_));
  OAI21_X1   g01867(.A1(new_n2863_), .A2(new_n2775_), .B(new_n2056_), .ZN(new_n2870_));
  NOR2_X1    g01868(.A1(new_n2869_), .A2(new_n2870_), .ZN(new_n2871_));
  OAI21_X1   g01869(.A1(new_n2871_), .A2(new_n2868_), .B(new_n2754_), .ZN(new_n2872_));
  NAND2_X1   g01870(.A1(new_n2872_), .A2(new_n2867_), .ZN(new_n2873_));
  NOR3_X1    g01871(.A1(new_n2837_), .A2(new_n2849_), .A3(new_n2860_), .ZN(new_n2874_));
  AOI21_X1   g01872(.A1(new_n2856_), .A2(new_n2859_), .B(new_n2850_), .ZN(new_n2875_));
  OAI21_X1   g01873(.A1(new_n2875_), .A2(new_n2874_), .B(new_n2873_), .ZN(new_n2876_));
  NAND2_X1   g01874(.A1(new_n2862_), .A2(new_n2876_), .ZN(new_n2877_));
  NOR2_X1    g01875(.A1(new_n1871_), .A2(new_n1900_), .ZN(new_n2878_));
  NOR2_X1    g01876(.A1(new_n1862_), .A2(new_n1901_), .ZN(new_n2879_));
  NOR2_X1    g01877(.A1(new_n2878_), .A2(new_n2879_), .ZN(new_n2880_));
  NOR2_X1    g01878(.A1(new_n1900_), .A2(new_n1901_), .ZN(new_n2881_));
  INV_X1     g01879(.I(new_n2881_), .ZN(new_n2882_));
  OAI21_X1   g01880(.A1(new_n2880_), .A2(new_n1905_), .B(new_n2882_), .ZN(new_n2883_));
  NOR3_X1    g01881(.A1(new_n2878_), .A2(new_n1905_), .A3(new_n2879_), .ZN(new_n2884_));
  NAND2_X1   g01882(.A1(new_n1862_), .A2(new_n1901_), .ZN(new_n2885_));
  NAND2_X1   g01883(.A1(new_n1871_), .A2(new_n1900_), .ZN(new_n2886_));
  AOI21_X1   g01884(.A1(new_n2885_), .A2(new_n2886_), .B(new_n1882_), .ZN(new_n2887_));
  NOR2_X1    g01885(.A1(new_n2887_), .A2(new_n2884_), .ZN(new_n2888_));
  AOI21_X1   g01886(.A1(new_n2883_), .A2(new_n1884_), .B(new_n2888_), .ZN(new_n2889_));
  NAND2_X1   g01887(.A1(new_n1892_), .A2(new_n1831_), .ZN(new_n2890_));
  NAND2_X1   g01888(.A1(new_n1889_), .A2(new_n1838_), .ZN(new_n2891_));
  NAND3_X1   g01889(.A1(new_n2890_), .A2(new_n1895_), .A3(new_n2891_), .ZN(new_n2892_));
  NOR2_X1    g01890(.A1(new_n1889_), .A2(new_n1838_), .ZN(new_n2893_));
  NOR2_X1    g01891(.A1(new_n1892_), .A2(new_n1831_), .ZN(new_n2894_));
  OAI21_X1   g01892(.A1(new_n2893_), .A2(new_n2894_), .B(new_n1850_), .ZN(new_n2895_));
  NAND2_X1   g01893(.A1(new_n2895_), .A2(new_n2892_), .ZN(new_n2896_));
  NAND4_X1   g01894(.A1(new_n1884_), .A2(new_n1897_), .A3(new_n1883_), .A4(new_n1896_), .ZN(new_n2897_));
  NOR2_X1    g01895(.A1(new_n1831_), .A2(new_n1838_), .ZN(new_n2898_));
  INV_X1     g01896(.I(new_n2898_), .ZN(new_n2899_));
  OAI21_X1   g01897(.A1(new_n2893_), .A2(new_n2894_), .B(new_n1895_), .ZN(new_n2900_));
  NAND2_X1   g01898(.A1(new_n2900_), .A2(new_n2899_), .ZN(new_n2901_));
  NAND2_X1   g01899(.A1(new_n2901_), .A2(new_n1897_), .ZN(new_n2902_));
  NAND3_X1   g01900(.A1(new_n2902_), .A2(new_n2896_), .A3(new_n2897_), .ZN(new_n2903_));
  NOR3_X1    g01901(.A1(new_n2893_), .A2(new_n1850_), .A3(new_n2894_), .ZN(new_n2904_));
  AOI21_X1   g01902(.A1(new_n2890_), .A2(new_n2891_), .B(new_n1895_), .ZN(new_n2905_));
  NOR2_X1    g01903(.A1(new_n2905_), .A2(new_n2904_), .ZN(new_n2906_));
  NOR4_X1    g01904(.A1(new_n1852_), .A2(new_n1909_), .A3(new_n1851_), .A4(new_n1906_), .ZN(new_n2907_));
  NAND2_X1   g01905(.A1(new_n2890_), .A2(new_n2891_), .ZN(new_n2908_));
  AOI21_X1   g01906(.A1(new_n2908_), .A2(new_n1895_), .B(new_n2898_), .ZN(new_n2909_));
  NOR2_X1    g01907(.A1(new_n2909_), .A2(new_n1852_), .ZN(new_n2910_));
  OAI21_X1   g01908(.A1(new_n2910_), .A2(new_n2906_), .B(new_n2907_), .ZN(new_n2911_));
  AOI21_X1   g01909(.A1(new_n2911_), .A2(new_n2903_), .B(new_n2889_), .ZN(new_n2912_));
  NAND2_X1   g01910(.A1(new_n2885_), .A2(new_n2886_), .ZN(new_n2913_));
  AOI21_X1   g01911(.A1(new_n2913_), .A2(new_n1882_), .B(new_n2881_), .ZN(new_n2914_));
  OAI22_X1   g01912(.A1(new_n2914_), .A2(new_n1909_), .B1(new_n2884_), .B2(new_n2887_), .ZN(new_n2915_));
  NOR2_X1    g01913(.A1(new_n1852_), .A2(new_n1909_), .ZN(new_n2916_));
  AOI21_X1   g01914(.A1(new_n2901_), .A2(new_n1897_), .B(new_n1906_), .ZN(new_n2917_));
  NAND4_X1   g01915(.A1(new_n2917_), .A2(new_n2909_), .A3(new_n2896_), .A4(new_n2916_), .ZN(new_n2918_));
  OAI21_X1   g01916(.A1(new_n2910_), .A2(new_n2906_), .B(new_n2897_), .ZN(new_n2919_));
  AOI21_X1   g01917(.A1(new_n2918_), .A2(new_n2919_), .B(new_n2915_), .ZN(new_n2920_));
  NOR2_X1    g01918(.A1(new_n2920_), .A2(new_n2912_), .ZN(new_n2921_));
  NOR2_X1    g01919(.A1(new_n1776_), .A2(new_n1816_), .ZN(new_n2922_));
  NOR2_X1    g01920(.A1(new_n1767_), .A2(new_n1817_), .ZN(new_n2923_));
  OAI21_X1   g01921(.A1(new_n2922_), .A2(new_n2923_), .B(new_n1787_), .ZN(new_n2924_));
  NOR2_X1    g01922(.A1(new_n1816_), .A2(new_n1817_), .ZN(new_n2925_));
  INV_X1     g01923(.I(new_n2925_), .ZN(new_n2926_));
  NAND2_X1   g01924(.A1(new_n2924_), .A2(new_n2926_), .ZN(new_n2927_));
  NAND2_X1   g01925(.A1(new_n1767_), .A2(new_n1817_), .ZN(new_n2928_));
  NAND2_X1   g01926(.A1(new_n1776_), .A2(new_n1816_), .ZN(new_n2929_));
  NAND3_X1   g01927(.A1(new_n2928_), .A2(new_n1787_), .A3(new_n2929_), .ZN(new_n2930_));
  OAI22_X1   g01928(.A1(new_n2922_), .A2(new_n2923_), .B1(new_n1789_), .B2(new_n1796_), .ZN(new_n2931_));
  AOI22_X1   g01929(.A1(new_n2927_), .A2(new_n1798_), .B1(new_n2930_), .B2(new_n2931_), .ZN(new_n2932_));
  NAND2_X1   g01930(.A1(new_n1805_), .A2(new_n1731_), .ZN(new_n2933_));
  NAND2_X1   g01931(.A1(new_n1803_), .A2(new_n1738_), .ZN(new_n2934_));
  NAND3_X1   g01932(.A1(new_n2933_), .A2(new_n1808_), .A3(new_n2934_), .ZN(new_n2935_));
  NOR2_X1    g01933(.A1(new_n1803_), .A2(new_n1738_), .ZN(new_n2936_));
  NOR2_X1    g01934(.A1(new_n1805_), .A2(new_n1731_), .ZN(new_n2937_));
  OAI21_X1   g01935(.A1(new_n2936_), .A2(new_n2937_), .B(new_n1750_), .ZN(new_n2938_));
  NAND2_X1   g01936(.A1(new_n2938_), .A2(new_n2935_), .ZN(new_n2939_));
  AOI22_X1   g01937(.A1(new_n1812_), .A2(new_n1813_), .B1(new_n1797_), .B2(new_n1791_), .ZN(new_n2940_));
  NAND3_X1   g01938(.A1(new_n2939_), .A2(new_n1809_), .A3(new_n2940_), .ZN(new_n2941_));
  NOR2_X1    g01939(.A1(new_n1731_), .A2(new_n1738_), .ZN(new_n2942_));
  AOI21_X1   g01940(.A1(new_n2933_), .A2(new_n2934_), .B(new_n1750_), .ZN(new_n2943_));
  OAI21_X1   g01941(.A1(new_n2943_), .A2(new_n2942_), .B(new_n1814_), .ZN(new_n2944_));
  NAND2_X1   g01942(.A1(new_n2944_), .A2(new_n1788_), .ZN(new_n2945_));
  NOR2_X1    g01943(.A1(new_n2945_), .A2(new_n2941_), .ZN(new_n2946_));
  NOR4_X1    g01944(.A1(new_n1757_), .A2(new_n1821_), .A3(new_n1751_), .A4(new_n1818_), .ZN(new_n2947_));
  INV_X1     g01945(.I(new_n2942_), .ZN(new_n2948_));
  NOR2_X1    g01946(.A1(new_n2936_), .A2(new_n2937_), .ZN(new_n2949_));
  OAI21_X1   g01947(.A1(new_n2949_), .A2(new_n1750_), .B(new_n2948_), .ZN(new_n2950_));
  AOI22_X1   g01948(.A1(new_n2950_), .A2(new_n1814_), .B1(new_n2935_), .B2(new_n2938_), .ZN(new_n2951_));
  NOR2_X1    g01949(.A1(new_n2951_), .A2(new_n2947_), .ZN(new_n2952_));
  OAI21_X1   g01950(.A1(new_n2946_), .A2(new_n2952_), .B(new_n2932_), .ZN(new_n2953_));
  NAND2_X1   g01951(.A1(new_n2928_), .A2(new_n2929_), .ZN(new_n2954_));
  AOI21_X1   g01952(.A1(new_n2954_), .A2(new_n1787_), .B(new_n2925_), .ZN(new_n2955_));
  NOR4_X1    g01953(.A1(new_n2922_), .A2(new_n2923_), .A3(new_n1789_), .A4(new_n1796_), .ZN(new_n2956_));
  AOI21_X1   g01954(.A1(new_n2928_), .A2(new_n2929_), .B(new_n1787_), .ZN(new_n2957_));
  OAI22_X1   g01955(.A1(new_n2955_), .A2(new_n1821_), .B1(new_n2956_), .B2(new_n2957_), .ZN(new_n2958_));
  NAND2_X1   g01956(.A1(new_n2944_), .A2(new_n2939_), .ZN(new_n2959_));
  NOR2_X1    g01957(.A1(new_n2959_), .A2(new_n2947_), .ZN(new_n2960_));
  NAND3_X1   g01958(.A1(new_n2940_), .A2(new_n1809_), .A3(new_n1788_), .ZN(new_n2961_));
  AOI21_X1   g01959(.A1(new_n2939_), .A2(new_n2944_), .B(new_n2961_), .ZN(new_n2962_));
  OAI21_X1   g01960(.A1(new_n2960_), .A2(new_n2962_), .B(new_n2958_), .ZN(new_n2963_));
  NAND2_X1   g01961(.A1(new_n1919_), .A2(new_n1824_), .ZN(new_n2964_));
  NAND3_X1   g01962(.A1(new_n2953_), .A2(new_n2963_), .A3(new_n2964_), .ZN(new_n2965_));
  NAND2_X1   g01963(.A1(new_n2933_), .A2(new_n2934_), .ZN(new_n2966_));
  AOI21_X1   g01964(.A1(new_n2966_), .A2(new_n1808_), .B(new_n2942_), .ZN(new_n2967_));
  AOI21_X1   g01965(.A1(new_n2950_), .A2(new_n1814_), .B(new_n1818_), .ZN(new_n2968_));
  NAND4_X1   g01966(.A1(new_n2968_), .A2(new_n2967_), .A3(new_n2939_), .A4(new_n2940_), .ZN(new_n2969_));
  NAND2_X1   g01967(.A1(new_n2959_), .A2(new_n2961_), .ZN(new_n2970_));
  AOI21_X1   g01968(.A1(new_n2969_), .A2(new_n2970_), .B(new_n2958_), .ZN(new_n2971_));
  NAND2_X1   g01969(.A1(new_n2951_), .A2(new_n2961_), .ZN(new_n2972_));
  NAND2_X1   g01970(.A1(new_n2959_), .A2(new_n2947_), .ZN(new_n2973_));
  AOI21_X1   g01971(.A1(new_n2972_), .A2(new_n2973_), .B(new_n2932_), .ZN(new_n2974_));
  NOR2_X1    g01972(.A1(new_n1912_), .A2(new_n1916_), .ZN(new_n2975_));
  OAI21_X1   g01973(.A1(new_n2971_), .A2(new_n2974_), .B(new_n2975_), .ZN(new_n2976_));
  AOI21_X1   g01974(.A1(new_n2976_), .A2(new_n2965_), .B(new_n2921_), .ZN(new_n2977_));
  NOR3_X1    g01975(.A1(new_n2910_), .A2(new_n2907_), .A3(new_n2906_), .ZN(new_n2978_));
  AOI22_X1   g01976(.A1(new_n2901_), .A2(new_n1897_), .B1(new_n2892_), .B2(new_n2895_), .ZN(new_n2979_));
  NOR2_X1    g01977(.A1(new_n2979_), .A2(new_n2897_), .ZN(new_n2980_));
  OAI21_X1   g01978(.A1(new_n2980_), .A2(new_n2978_), .B(new_n2915_), .ZN(new_n2981_));
  NAND4_X1   g01979(.A1(new_n2896_), .A2(new_n1896_), .A3(new_n1897_), .A4(new_n1884_), .ZN(new_n2982_));
  OAI21_X1   g01980(.A1(new_n2909_), .A2(new_n1852_), .B(new_n1883_), .ZN(new_n2983_));
  NOR2_X1    g01981(.A1(new_n2982_), .A2(new_n2983_), .ZN(new_n2984_));
  NOR2_X1    g01982(.A1(new_n2979_), .A2(new_n2907_), .ZN(new_n2985_));
  OAI21_X1   g01983(.A1(new_n2984_), .A2(new_n2985_), .B(new_n2889_), .ZN(new_n2986_));
  NAND2_X1   g01984(.A1(new_n2986_), .A2(new_n2981_), .ZN(new_n2987_));
  NAND3_X1   g01985(.A1(new_n2953_), .A2(new_n2963_), .A3(new_n2975_), .ZN(new_n2988_));
  OAI21_X1   g01986(.A1(new_n2971_), .A2(new_n2974_), .B(new_n2964_), .ZN(new_n2989_));
  AOI21_X1   g01987(.A1(new_n2989_), .A2(new_n2988_), .B(new_n2987_), .ZN(new_n2990_));
  AOI22_X1   g01988(.A1(new_n2062_), .A2(new_n2060_), .B1(new_n1920_), .B2(new_n1913_), .ZN(new_n2991_));
  NOR3_X1    g01989(.A1(new_n2990_), .A2(new_n2977_), .A3(new_n2991_), .ZN(new_n2992_));
  NOR3_X1    g01990(.A1(new_n2971_), .A2(new_n2974_), .A3(new_n2975_), .ZN(new_n2993_));
  AOI21_X1   g01991(.A1(new_n2953_), .A2(new_n2963_), .B(new_n2964_), .ZN(new_n2994_));
  OAI21_X1   g01992(.A1(new_n2993_), .A2(new_n2994_), .B(new_n2987_), .ZN(new_n2995_));
  NOR3_X1    g01993(.A1(new_n2971_), .A2(new_n2974_), .A3(new_n2964_), .ZN(new_n2996_));
  AOI21_X1   g01994(.A1(new_n2953_), .A2(new_n2963_), .B(new_n2975_), .ZN(new_n2997_));
  OAI21_X1   g01995(.A1(new_n2996_), .A2(new_n2997_), .B(new_n2921_), .ZN(new_n2998_));
  INV_X1     g01996(.I(new_n2991_), .ZN(new_n2999_));
  AOI21_X1   g01997(.A1(new_n2998_), .A2(new_n2995_), .B(new_n2999_), .ZN(new_n3000_));
  OAI21_X1   g01998(.A1(new_n3000_), .A2(new_n2992_), .B(new_n2877_), .ZN(new_n3001_));
  NAND3_X1   g01999(.A1(new_n2856_), .A2(new_n2859_), .A3(new_n2860_), .ZN(new_n3002_));
  OAI21_X1   g02000(.A1(new_n2837_), .A2(new_n2849_), .B(new_n2850_), .ZN(new_n3003_));
  AOI21_X1   g02001(.A1(new_n3003_), .A2(new_n3002_), .B(new_n2873_), .ZN(new_n3004_));
  NAND3_X1   g02002(.A1(new_n2856_), .A2(new_n2850_), .A3(new_n2859_), .ZN(new_n3005_));
  OAI21_X1   g02003(.A1(new_n2837_), .A2(new_n2849_), .B(new_n2860_), .ZN(new_n3006_));
  AOI21_X1   g02004(.A1(new_n3005_), .A2(new_n3006_), .B(new_n2797_), .ZN(new_n3007_));
  NOR2_X1    g02005(.A1(new_n3007_), .A2(new_n3004_), .ZN(new_n3008_));
  NOR3_X1    g02006(.A1(new_n2990_), .A2(new_n2977_), .A3(new_n2999_), .ZN(new_n3009_));
  AOI21_X1   g02007(.A1(new_n2998_), .A2(new_n2995_), .B(new_n2991_), .ZN(new_n3010_));
  OAI21_X1   g02008(.A1(new_n3010_), .A2(new_n3009_), .B(new_n3008_), .ZN(new_n3011_));
  NOR2_X1    g02009(.A1(new_n2339_), .A2(new_n2064_), .ZN(new_n3012_));
  INV_X1     g02010(.I(new_n3012_), .ZN(new_n3013_));
  NAND3_X1   g02011(.A1(new_n3013_), .A2(new_n3001_), .A3(new_n3011_), .ZN(new_n3014_));
  NAND2_X1   g02012(.A1(new_n3011_), .A2(new_n3001_), .ZN(new_n3015_));
  NAND2_X1   g02013(.A1(new_n3015_), .A2(new_n3012_), .ZN(new_n3016_));
  AOI21_X1   g02014(.A1(new_n3016_), .A2(new_n3014_), .B(new_n2734_), .ZN(new_n3017_));
  INV_X1     g02015(.I(new_n2734_), .ZN(new_n3018_));
  NAND3_X1   g02016(.A1(new_n3011_), .A2(new_n3001_), .A3(new_n3012_), .ZN(new_n3019_));
  NAND2_X1   g02017(.A1(new_n3015_), .A2(new_n3013_), .ZN(new_n3020_));
  AOI21_X1   g02018(.A1(new_n3020_), .A2(new_n3019_), .B(new_n3018_), .ZN(new_n3021_));
  NOR2_X1    g02019(.A1(new_n2341_), .A2(new_n1723_), .ZN(new_n3022_));
  INV_X1     g02020(.I(new_n3022_), .ZN(new_n3023_));
  NOR3_X1    g02021(.A1(new_n3021_), .A2(new_n3017_), .A3(new_n3023_), .ZN(new_n3024_));
  OAI21_X1   g02022(.A1(new_n3021_), .A2(new_n3017_), .B(new_n3023_), .ZN(new_n3025_));
  INV_X1     g02023(.I(new_n3025_), .ZN(new_n3026_));
  OAI21_X1   g02024(.A1(new_n3026_), .A2(new_n3024_), .B(new_n2544_), .ZN(new_n3027_));
  NOR3_X1    g02025(.A1(new_n3021_), .A2(new_n3017_), .A3(new_n3022_), .ZN(new_n3028_));
  OAI21_X1   g02026(.A1(new_n3021_), .A2(new_n3017_), .B(new_n3022_), .ZN(new_n3029_));
  INV_X1     g02027(.I(new_n3029_), .ZN(new_n3030_));
  OAI21_X1   g02028(.A1(new_n3030_), .A2(new_n3028_), .B(new_n2543_), .ZN(new_n3031_));
  AOI21_X1   g02029(.A1(new_n3027_), .A2(new_n3031_), .B(new_n2346_), .ZN(new_n3032_));
  AOI21_X1   g02030(.A1(new_n1505_), .A2(\A[852] ), .B(new_n1508_), .ZN(new_n3033_));
  XOR2_X1    g02031(.A1(new_n1516_), .A2(new_n3033_), .Z(new_n3034_));
  INV_X1     g02032(.I(new_n1517_), .ZN(new_n3035_));
  AOI21_X1   g02033(.A1(new_n1497_), .A2(\A[849] ), .B(new_n1514_), .ZN(new_n3036_));
  NOR2_X1    g02034(.A1(new_n3033_), .A2(new_n3036_), .ZN(new_n3037_));
  INV_X1     g02035(.I(new_n3037_), .ZN(new_n3038_));
  OAI21_X1   g02036(.A1(new_n3034_), .A2(new_n3035_), .B(new_n3038_), .ZN(new_n3039_));
  NAND2_X1   g02037(.A1(new_n1511_), .A2(new_n3036_), .ZN(new_n3040_));
  NAND2_X1   g02038(.A1(new_n1516_), .A2(new_n3033_), .ZN(new_n3041_));
  NAND3_X1   g02039(.A1(new_n3040_), .A2(new_n1517_), .A3(new_n3041_), .ZN(new_n3042_));
  NAND2_X1   g02040(.A1(new_n3040_), .A2(new_n3041_), .ZN(new_n3043_));
  NAND2_X1   g02041(.A1(new_n3043_), .A2(new_n3035_), .ZN(new_n3044_));
  AOI22_X1   g02042(.A1(new_n3039_), .A2(new_n1507_), .B1(new_n3044_), .B2(new_n3042_), .ZN(new_n3045_));
  INV_X1     g02043(.I(new_n3045_), .ZN(new_n3046_));
  AOI21_X1   g02044(.A1(new_n1465_), .A2(\A[855] ), .B(new_n1484_), .ZN(new_n3047_));
  NAND2_X1   g02045(.A1(new_n1481_), .A2(new_n3047_), .ZN(new_n3048_));
  AOI21_X1   g02046(.A1(new_n1474_), .A2(\A[858] ), .B(new_n1479_), .ZN(new_n3049_));
  NAND2_X1   g02047(.A1(new_n1486_), .A2(new_n3049_), .ZN(new_n3050_));
  NAND2_X1   g02048(.A1(new_n3048_), .A2(new_n3050_), .ZN(new_n3051_));
  XOR2_X1    g02049(.A1(new_n3051_), .A2(new_n1487_), .Z(new_n3052_));
  NOR2_X1    g02050(.A1(new_n3049_), .A2(new_n3047_), .ZN(new_n3053_));
  AOI21_X1   g02051(.A1(new_n3051_), .A2(new_n1487_), .B(new_n3053_), .ZN(new_n3054_));
  XNOR2_X1   g02052(.A1(new_n1466_), .A2(new_n1475_), .ZN(new_n3055_));
  XNOR2_X1   g02053(.A1(new_n1498_), .A2(new_n1506_), .ZN(new_n3056_));
  NOR2_X1    g02054(.A1(new_n3055_), .A2(new_n3056_), .ZN(new_n3057_));
  INV_X1     g02055(.I(new_n1518_), .ZN(new_n3058_));
  NOR2_X1    g02056(.A1(new_n3054_), .A2(new_n3055_), .ZN(new_n3059_));
  NOR2_X1    g02057(.A1(new_n3059_), .A2(new_n3058_), .ZN(new_n3060_));
  NAND4_X1   g02058(.A1(new_n3060_), .A2(new_n3052_), .A3(new_n3054_), .A4(new_n3057_), .ZN(new_n3061_));
  AND4_X2    g02059(.A1(new_n1476_), .A2(new_n1507_), .A3(new_n1488_), .A4(new_n1518_), .Z(new_n3062_));
  INV_X1     g02060(.I(new_n3062_), .ZN(new_n3063_));
  XOR2_X1    g02061(.A1(new_n1481_), .A2(new_n3047_), .Z(new_n3064_));
  INV_X1     g02062(.I(new_n1487_), .ZN(new_n3065_));
  INV_X1     g02063(.I(new_n3053_), .ZN(new_n3066_));
  OAI21_X1   g02064(.A1(new_n3064_), .A2(new_n3065_), .B(new_n3066_), .ZN(new_n3067_));
  NAND2_X1   g02065(.A1(new_n3067_), .A2(new_n1476_), .ZN(new_n3068_));
  NAND2_X1   g02066(.A1(new_n3068_), .A2(new_n3052_), .ZN(new_n3069_));
  NAND2_X1   g02067(.A1(new_n3069_), .A2(new_n3063_), .ZN(new_n3070_));
  AOI21_X1   g02068(.A1(new_n3070_), .A2(new_n3061_), .B(new_n3046_), .ZN(new_n3071_));
  XNOR2_X1   g02069(.A1(new_n3051_), .A2(new_n1487_), .ZN(new_n3072_));
  NOR2_X1    g02070(.A1(new_n3072_), .A2(new_n3059_), .ZN(new_n3073_));
  XOR2_X1    g02071(.A1(new_n3073_), .A2(new_n3062_), .Z(new_n3074_));
  AOI21_X1   g02072(.A1(new_n3074_), .A2(new_n3046_), .B(new_n3071_), .ZN(new_n3075_));
  NAND2_X1   g02073(.A1(new_n1433_), .A2(\A[861] ), .ZN(new_n3076_));
  OAI22_X1   g02074(.A1(new_n1450_), .A2(\A[861] ), .B1(new_n3076_), .B2(new_n1449_), .ZN(new_n3077_));
  XOR2_X1    g02075(.A1(new_n3077_), .A2(new_n1443_), .Z(new_n3078_));
  AOI21_X1   g02076(.A1(new_n1434_), .A2(\A[861] ), .B(new_n1451_), .ZN(new_n3079_));
  NAND2_X1   g02077(.A1(new_n1448_), .A2(new_n3079_), .ZN(new_n3080_));
  AOI21_X1   g02078(.A1(new_n1442_), .A2(\A[864] ), .B(new_n1446_), .ZN(new_n3081_));
  NAND2_X1   g02079(.A1(new_n1453_), .A2(new_n3081_), .ZN(new_n3082_));
  NAND2_X1   g02080(.A1(new_n3080_), .A2(new_n3082_), .ZN(new_n3083_));
  NOR2_X1    g02081(.A1(new_n3081_), .A2(new_n3079_), .ZN(new_n3084_));
  AOI21_X1   g02082(.A1(new_n3083_), .A2(new_n1454_), .B(new_n3084_), .ZN(new_n3085_));
  NAND2_X1   g02083(.A1(new_n1440_), .A2(new_n1438_), .ZN(new_n3086_));
  OAI21_X1   g02084(.A1(\A[864] ), .A2(new_n1445_), .B(new_n3086_), .ZN(new_n3087_));
  NAND2_X1   g02085(.A1(new_n3087_), .A2(new_n3077_), .ZN(new_n3088_));
  NOR2_X1    g02086(.A1(new_n3083_), .A2(new_n3088_), .ZN(new_n3089_));
  AOI21_X1   g02087(.A1(new_n3080_), .A2(new_n3082_), .B(new_n1454_), .ZN(new_n3090_));
  OAI22_X1   g02088(.A1(new_n3085_), .A2(new_n3078_), .B1(new_n3089_), .B2(new_n3090_), .ZN(new_n3091_));
  AOI21_X1   g02089(.A1(new_n1402_), .A2(\A[867] ), .B(new_n1421_), .ZN(new_n3092_));
  NAND2_X1   g02090(.A1(new_n1418_), .A2(new_n3092_), .ZN(new_n3093_));
  AOI21_X1   g02091(.A1(new_n1411_), .A2(\A[870] ), .B(new_n1416_), .ZN(new_n3094_));
  NAND2_X1   g02092(.A1(new_n1423_), .A2(new_n3094_), .ZN(new_n3095_));
  NAND3_X1   g02093(.A1(new_n1424_), .A2(new_n3093_), .A3(new_n3095_), .ZN(new_n3096_));
  NAND2_X1   g02094(.A1(new_n3093_), .A2(new_n3095_), .ZN(new_n3097_));
  INV_X1     g02095(.I(new_n1424_), .ZN(new_n3098_));
  NAND2_X1   g02096(.A1(new_n3097_), .A2(new_n3098_), .ZN(new_n3099_));
  NAND2_X1   g02097(.A1(new_n3099_), .A2(new_n3096_), .ZN(new_n3100_));
  NOR2_X1    g02098(.A1(new_n3094_), .A2(new_n3092_), .ZN(new_n3101_));
  AOI21_X1   g02099(.A1(new_n3097_), .A2(new_n1424_), .B(new_n3101_), .ZN(new_n3102_));
  XNOR2_X1   g02100(.A1(new_n1403_), .A2(new_n1412_), .ZN(new_n3103_));
  NOR2_X1    g02101(.A1(new_n3103_), .A2(new_n3078_), .ZN(new_n3104_));
  INV_X1     g02102(.I(new_n1455_), .ZN(new_n3105_));
  NOR2_X1    g02103(.A1(new_n3102_), .A2(new_n3103_), .ZN(new_n3106_));
  NOR2_X1    g02104(.A1(new_n3106_), .A2(new_n3105_), .ZN(new_n3107_));
  NAND4_X1   g02105(.A1(new_n3107_), .A2(new_n3100_), .A3(new_n3102_), .A4(new_n3104_), .ZN(new_n3108_));
  NAND3_X1   g02106(.A1(new_n3104_), .A2(new_n1425_), .A3(new_n1455_), .ZN(new_n3109_));
  OAI21_X1   g02107(.A1(new_n3103_), .A2(new_n3102_), .B(new_n3100_), .ZN(new_n3110_));
  NAND2_X1   g02108(.A1(new_n3110_), .A2(new_n3109_), .ZN(new_n3111_));
  AOI21_X1   g02109(.A1(new_n3111_), .A2(new_n3108_), .B(new_n3091_), .ZN(new_n3112_));
  INV_X1     g02110(.I(new_n3091_), .ZN(new_n3113_));
  INV_X1     g02111(.I(new_n1425_), .ZN(new_n3114_));
  NOR4_X1    g02112(.A1(new_n3114_), .A2(new_n3105_), .A3(new_n3103_), .A4(new_n3078_), .ZN(new_n3115_));
  NAND2_X1   g02113(.A1(new_n3110_), .A2(new_n3115_), .ZN(new_n3116_));
  INV_X1     g02114(.I(new_n3096_), .ZN(new_n3117_));
  AOI21_X1   g02115(.A1(new_n3093_), .A2(new_n3095_), .B(new_n1424_), .ZN(new_n3118_));
  NOR2_X1    g02116(.A1(new_n3117_), .A2(new_n3118_), .ZN(new_n3119_));
  NOR2_X1    g02117(.A1(new_n3106_), .A2(new_n3119_), .ZN(new_n3120_));
  NAND2_X1   g02118(.A1(new_n3120_), .A2(new_n3109_), .ZN(new_n3121_));
  AOI21_X1   g02119(.A1(new_n3116_), .A2(new_n3121_), .B(new_n3113_), .ZN(new_n3122_));
  NAND2_X1   g02120(.A1(new_n1457_), .A2(new_n1520_), .ZN(new_n3123_));
  NOR3_X1    g02121(.A1(new_n3112_), .A2(new_n3122_), .A3(new_n3123_), .ZN(new_n3124_));
  XNOR2_X1   g02122(.A1(new_n1426_), .A2(new_n1456_), .ZN(new_n3125_));
  XNOR2_X1   g02123(.A1(new_n1489_), .A2(new_n1519_), .ZN(new_n3126_));
  NOR2_X1    g02124(.A1(new_n3126_), .A2(new_n3125_), .ZN(new_n3127_));
  NOR2_X1    g02125(.A1(new_n3112_), .A2(new_n3122_), .ZN(new_n3128_));
  NOR2_X1    g02126(.A1(new_n3128_), .A2(new_n3127_), .ZN(new_n3129_));
  OAI21_X1   g02127(.A1(new_n3129_), .A2(new_n3124_), .B(new_n3075_), .ZN(new_n3130_));
  NAND3_X1   g02128(.A1(new_n3052_), .A2(new_n1488_), .A3(new_n3057_), .ZN(new_n3131_));
  NAND2_X1   g02129(.A1(new_n3068_), .A2(new_n1518_), .ZN(new_n3132_));
  NOR2_X1    g02130(.A1(new_n3131_), .A2(new_n3132_), .ZN(new_n3133_));
  NOR2_X1    g02131(.A1(new_n3073_), .A2(new_n3062_), .ZN(new_n3134_));
  OAI21_X1   g02132(.A1(new_n3133_), .A2(new_n3134_), .B(new_n3045_), .ZN(new_n3135_));
  NOR2_X1    g02133(.A1(new_n3069_), .A2(new_n3062_), .ZN(new_n3136_));
  NOR2_X1    g02134(.A1(new_n3073_), .A2(new_n3063_), .ZN(new_n3137_));
  OAI21_X1   g02135(.A1(new_n3137_), .A2(new_n3136_), .B(new_n3046_), .ZN(new_n3138_));
  NAND2_X1   g02136(.A1(new_n3138_), .A2(new_n3135_), .ZN(new_n3139_));
  NOR3_X1    g02137(.A1(new_n3112_), .A2(new_n3122_), .A3(new_n3127_), .ZN(new_n3140_));
  NAND2_X1   g02138(.A1(new_n3100_), .A2(new_n3104_), .ZN(new_n3141_));
  NOR4_X1    g02139(.A1(new_n3141_), .A2(new_n3114_), .A3(new_n3105_), .A4(new_n3106_), .ZN(new_n3142_));
  NOR2_X1    g02140(.A1(new_n3120_), .A2(new_n3115_), .ZN(new_n3143_));
  OAI21_X1   g02141(.A1(new_n3142_), .A2(new_n3143_), .B(new_n3113_), .ZN(new_n3144_));
  NOR2_X1    g02142(.A1(new_n3120_), .A2(new_n3109_), .ZN(new_n3145_));
  NOR3_X1    g02143(.A1(new_n3115_), .A2(new_n3106_), .A3(new_n3119_), .ZN(new_n3146_));
  OAI21_X1   g02144(.A1(new_n3145_), .A2(new_n3146_), .B(new_n3091_), .ZN(new_n3147_));
  AOI21_X1   g02145(.A1(new_n3144_), .A2(new_n3147_), .B(new_n3123_), .ZN(new_n3148_));
  OAI21_X1   g02146(.A1(new_n3140_), .A2(new_n3148_), .B(new_n3139_), .ZN(new_n3149_));
  NAND2_X1   g02147(.A1(new_n3130_), .A2(new_n3149_), .ZN(new_n3150_));
  AOI21_X1   g02148(.A1(new_n1370_), .A2(\A[873] ), .B(new_n1387_), .ZN(new_n3151_));
  NAND2_X1   g02149(.A1(new_n1384_), .A2(new_n3151_), .ZN(new_n3152_));
  AOI21_X1   g02150(.A1(new_n1378_), .A2(\A[876] ), .B(new_n1382_), .ZN(new_n3153_));
  NAND2_X1   g02151(.A1(new_n1389_), .A2(new_n3153_), .ZN(new_n3154_));
  NAND2_X1   g02152(.A1(new_n3152_), .A2(new_n3154_), .ZN(new_n3155_));
  NOR2_X1    g02153(.A1(new_n3153_), .A2(new_n3151_), .ZN(new_n3156_));
  AOI21_X1   g02154(.A1(new_n3155_), .A2(new_n1390_), .B(new_n3156_), .ZN(new_n3157_));
  INV_X1     g02155(.I(new_n3157_), .ZN(new_n3158_));
  NAND3_X1   g02156(.A1(new_n1390_), .A2(new_n3152_), .A3(new_n3154_), .ZN(new_n3159_));
  NAND2_X1   g02157(.A1(new_n1369_), .A2(\A[873] ), .ZN(new_n3160_));
  OAI22_X1   g02158(.A1(new_n1386_), .A2(\A[873] ), .B1(new_n3160_), .B2(new_n1385_), .ZN(new_n3161_));
  NAND2_X1   g02159(.A1(new_n1376_), .A2(new_n1374_), .ZN(new_n3162_));
  OAI21_X1   g02160(.A1(\A[876] ), .A2(new_n1381_), .B(new_n3162_), .ZN(new_n3163_));
  NAND2_X1   g02161(.A1(new_n3163_), .A2(new_n3161_), .ZN(new_n3164_));
  NAND2_X1   g02162(.A1(new_n3155_), .A2(new_n3164_), .ZN(new_n3165_));
  AOI22_X1   g02163(.A1(new_n3158_), .A2(new_n1380_), .B1(new_n3165_), .B2(new_n3159_), .ZN(new_n3166_));
  AOI21_X1   g02164(.A1(new_n1348_), .A2(\A[882] ), .B(new_n1352_), .ZN(new_n3167_));
  AOI21_X1   g02165(.A1(new_n1340_), .A2(\A[879] ), .B(new_n1357_), .ZN(new_n3168_));
  NAND2_X1   g02166(.A1(new_n1339_), .A2(\A[879] ), .ZN(new_n3169_));
  OAI22_X1   g02167(.A1(new_n1356_), .A2(\A[879] ), .B1(new_n3169_), .B2(new_n1355_), .ZN(new_n3170_));
  NAND2_X1   g02168(.A1(new_n1346_), .A2(new_n1344_), .ZN(new_n3171_));
  OAI21_X1   g02169(.A1(\A[882] ), .A2(new_n1351_), .B(new_n3171_), .ZN(new_n3172_));
  NAND2_X1   g02170(.A1(new_n3172_), .A2(new_n3170_), .ZN(new_n3173_));
  NOR3_X1    g02171(.A1(new_n3173_), .A2(new_n3167_), .A3(new_n3168_), .ZN(new_n3174_));
  NOR3_X1    g02172(.A1(new_n3164_), .A2(new_n3153_), .A3(new_n3151_), .ZN(new_n3175_));
  NAND2_X1   g02173(.A1(new_n1354_), .A2(new_n3168_), .ZN(new_n3176_));
  NAND2_X1   g02174(.A1(new_n1359_), .A2(new_n3167_), .ZN(new_n3177_));
  NAND3_X1   g02175(.A1(new_n1360_), .A2(new_n3176_), .A3(new_n3177_), .ZN(new_n3178_));
  NAND2_X1   g02176(.A1(new_n3176_), .A2(new_n3177_), .ZN(new_n3179_));
  NAND2_X1   g02177(.A1(new_n3179_), .A2(new_n3173_), .ZN(new_n3180_));
  NAND2_X1   g02178(.A1(new_n3180_), .A2(new_n3178_), .ZN(new_n3181_));
  XOR2_X1    g02179(.A1(new_n3170_), .A2(new_n1349_), .Z(new_n3182_));
  XOR2_X1    g02180(.A1(new_n3161_), .A2(new_n1379_), .Z(new_n3183_));
  NOR2_X1    g02181(.A1(new_n3182_), .A2(new_n3183_), .ZN(new_n3184_));
  NAND2_X1   g02182(.A1(new_n3181_), .A2(new_n3184_), .ZN(new_n3185_));
  NOR2_X1    g02183(.A1(new_n3167_), .A2(new_n3168_), .ZN(new_n3186_));
  AOI21_X1   g02184(.A1(new_n3179_), .A2(new_n1360_), .B(new_n3186_), .ZN(new_n3187_));
  NOR2_X1    g02185(.A1(new_n3187_), .A2(new_n3182_), .ZN(new_n3188_));
  NOR4_X1    g02186(.A1(new_n3185_), .A2(new_n3174_), .A3(new_n3175_), .A4(new_n3188_), .ZN(new_n3189_));
  XOR2_X1    g02187(.A1(new_n1354_), .A2(new_n3168_), .Z(new_n3190_));
  INV_X1     g02188(.I(new_n3186_), .ZN(new_n3191_));
  OAI21_X1   g02189(.A1(new_n3190_), .A2(new_n3173_), .B(new_n3191_), .ZN(new_n3192_));
  NAND2_X1   g02190(.A1(new_n3192_), .A2(new_n1350_), .ZN(new_n3193_));
  NOR4_X1    g02191(.A1(new_n3182_), .A2(new_n3183_), .A3(new_n3174_), .A4(new_n3175_), .ZN(new_n3194_));
  AOI21_X1   g02192(.A1(new_n3193_), .A2(new_n3181_), .B(new_n3194_), .ZN(new_n3195_));
  OAI21_X1   g02193(.A1(new_n3189_), .A2(new_n3195_), .B(new_n3166_), .ZN(new_n3196_));
  NAND2_X1   g02194(.A1(new_n3165_), .A2(new_n3159_), .ZN(new_n3197_));
  OAI21_X1   g02195(.A1(new_n3183_), .A2(new_n3157_), .B(new_n3197_), .ZN(new_n3198_));
  NAND2_X1   g02196(.A1(new_n3193_), .A2(new_n3181_), .ZN(new_n3199_));
  NOR2_X1    g02197(.A1(new_n3199_), .A2(new_n3194_), .ZN(new_n3200_));
  INV_X1     g02198(.I(new_n3194_), .ZN(new_n3201_));
  INV_X1     g02199(.I(new_n3178_), .ZN(new_n3202_));
  AOI21_X1   g02200(.A1(new_n3176_), .A2(new_n3177_), .B(new_n1360_), .ZN(new_n3203_));
  NOR2_X1    g02201(.A1(new_n3202_), .A2(new_n3203_), .ZN(new_n3204_));
  NOR2_X1    g02202(.A1(new_n3188_), .A2(new_n3204_), .ZN(new_n3205_));
  NOR2_X1    g02203(.A1(new_n3205_), .A2(new_n3201_), .ZN(new_n3206_));
  OAI21_X1   g02204(.A1(new_n3200_), .A2(new_n3206_), .B(new_n3198_), .ZN(new_n3207_));
  NAND2_X1   g02205(.A1(new_n3207_), .A2(new_n3196_), .ZN(new_n3208_));
  NAND2_X1   g02206(.A1(new_n1332_), .A2(new_n1393_), .ZN(new_n3209_));
  NAND2_X1   g02207(.A1(new_n1308_), .A2(\A[885] ), .ZN(new_n3210_));
  OAI22_X1   g02208(.A1(new_n1325_), .A2(\A[885] ), .B1(new_n3210_), .B2(new_n1324_), .ZN(new_n3211_));
  XOR2_X1    g02209(.A1(new_n3211_), .A2(new_n1318_), .Z(new_n3212_));
  AOI21_X1   g02210(.A1(new_n1309_), .A2(\A[885] ), .B(new_n1326_), .ZN(new_n3213_));
  NAND2_X1   g02211(.A1(new_n1323_), .A2(new_n3213_), .ZN(new_n3214_));
  AOI21_X1   g02212(.A1(new_n1317_), .A2(\A[888] ), .B(new_n1321_), .ZN(new_n3215_));
  NAND2_X1   g02213(.A1(new_n1328_), .A2(new_n3215_), .ZN(new_n3216_));
  NAND2_X1   g02214(.A1(new_n3214_), .A2(new_n3216_), .ZN(new_n3217_));
  NOR2_X1    g02215(.A1(new_n3215_), .A2(new_n3213_), .ZN(new_n3218_));
  AOI21_X1   g02216(.A1(new_n3217_), .A2(new_n1329_), .B(new_n3218_), .ZN(new_n3219_));
  NAND3_X1   g02217(.A1(new_n1329_), .A2(new_n3214_), .A3(new_n3216_), .ZN(new_n3220_));
  NAND2_X1   g02218(.A1(new_n1315_), .A2(new_n1313_), .ZN(new_n3221_));
  OAI21_X1   g02219(.A1(\A[888] ), .A2(new_n1320_), .B(new_n3221_), .ZN(new_n3222_));
  NAND2_X1   g02220(.A1(new_n3222_), .A2(new_n3211_), .ZN(new_n3223_));
  NAND2_X1   g02221(.A1(new_n3217_), .A2(new_n3223_), .ZN(new_n3224_));
  NAND2_X1   g02222(.A1(new_n3224_), .A2(new_n3220_), .ZN(new_n3225_));
  OAI21_X1   g02223(.A1(new_n3212_), .A2(new_n3219_), .B(new_n3225_), .ZN(new_n3226_));
  AOI21_X1   g02224(.A1(new_n1293_), .A2(\A[891] ), .B(new_n1288_), .ZN(new_n3227_));
  NAND2_X1   g02225(.A1(new_n1286_), .A2(new_n3227_), .ZN(new_n3228_));
  AOI21_X1   g02226(.A1(new_n1297_), .A2(\A[894] ), .B(new_n1284_), .ZN(new_n3229_));
  NAND2_X1   g02227(.A1(new_n1290_), .A2(new_n3229_), .ZN(new_n3230_));
  NAND3_X1   g02228(.A1(new_n1299_), .A2(new_n3228_), .A3(new_n3230_), .ZN(new_n3231_));
  NOR2_X1    g02229(.A1(new_n1290_), .A2(new_n3229_), .ZN(new_n3232_));
  NOR2_X1    g02230(.A1(new_n1286_), .A2(new_n3227_), .ZN(new_n3233_));
  NAND2_X1   g02231(.A1(new_n1273_), .A2(new_n1281_), .ZN(new_n3234_));
  OAI21_X1   g02232(.A1(new_n3232_), .A2(new_n3233_), .B(new_n3234_), .ZN(new_n3235_));
  NAND2_X1   g02233(.A1(new_n3235_), .A2(new_n3231_), .ZN(new_n3236_));
  NAND2_X1   g02234(.A1(new_n3228_), .A2(new_n3230_), .ZN(new_n3237_));
  NOR2_X1    g02235(.A1(new_n3229_), .A2(new_n3227_), .ZN(new_n3238_));
  AOI21_X1   g02236(.A1(new_n3237_), .A2(new_n1299_), .B(new_n3238_), .ZN(new_n3239_));
  XOR2_X1    g02237(.A1(new_n1294_), .A2(new_n1281_), .Z(new_n3240_));
  NOR2_X1    g02238(.A1(new_n3240_), .A2(new_n3212_), .ZN(new_n3241_));
  NOR2_X1    g02239(.A1(new_n3232_), .A2(new_n3233_), .ZN(new_n3242_));
  INV_X1     g02240(.I(new_n3238_), .ZN(new_n3243_));
  OAI21_X1   g02241(.A1(new_n3242_), .A2(new_n3234_), .B(new_n3243_), .ZN(new_n3244_));
  NOR3_X1    g02242(.A1(new_n3223_), .A2(new_n3215_), .A3(new_n3213_), .ZN(new_n3245_));
  AOI21_X1   g02243(.A1(new_n3244_), .A2(new_n1282_), .B(new_n3245_), .ZN(new_n3246_));
  NAND4_X1   g02244(.A1(new_n3246_), .A2(new_n3236_), .A3(new_n3239_), .A4(new_n3241_), .ZN(new_n3247_));
  NAND4_X1   g02245(.A1(new_n1282_), .A2(new_n1319_), .A3(new_n1300_), .A4(new_n1330_), .ZN(new_n3248_));
  OAI21_X1   g02246(.A1(new_n3240_), .A2(new_n3239_), .B(new_n3236_), .ZN(new_n3249_));
  NAND2_X1   g02247(.A1(new_n3249_), .A2(new_n3248_), .ZN(new_n3250_));
  AOI21_X1   g02248(.A1(new_n3250_), .A2(new_n3247_), .B(new_n3226_), .ZN(new_n3251_));
  INV_X1     g02249(.I(new_n3219_), .ZN(new_n3252_));
  INV_X1     g02250(.I(new_n3220_), .ZN(new_n3253_));
  AOI21_X1   g02251(.A1(new_n3214_), .A2(new_n3216_), .B(new_n1329_), .ZN(new_n3254_));
  NOR2_X1    g02252(.A1(new_n3253_), .A2(new_n3254_), .ZN(new_n3255_));
  AOI21_X1   g02253(.A1(new_n1319_), .A2(new_n3252_), .B(new_n3255_), .ZN(new_n3256_));
  NOR3_X1    g02254(.A1(new_n3234_), .A2(new_n3229_), .A3(new_n3227_), .ZN(new_n3257_));
  NOR4_X1    g02255(.A1(new_n3240_), .A2(new_n3212_), .A3(new_n3245_), .A4(new_n3257_), .ZN(new_n3258_));
  NAND2_X1   g02256(.A1(new_n3249_), .A2(new_n3258_), .ZN(new_n3259_));
  NAND2_X1   g02257(.A1(new_n3244_), .A2(new_n1282_), .ZN(new_n3260_));
  NAND3_X1   g02258(.A1(new_n3260_), .A2(new_n3248_), .A3(new_n3236_), .ZN(new_n3261_));
  AOI21_X1   g02259(.A1(new_n3259_), .A2(new_n3261_), .B(new_n3256_), .ZN(new_n3262_));
  NOR2_X1    g02260(.A1(new_n3251_), .A2(new_n3262_), .ZN(new_n3263_));
  NOR2_X1    g02261(.A1(new_n3263_), .A2(new_n3209_), .ZN(new_n3264_));
  XNOR2_X1   g02262(.A1(new_n1301_), .A2(new_n1331_), .ZN(new_n3265_));
  XNOR2_X1   g02263(.A1(new_n1362_), .A2(new_n1392_), .ZN(new_n3266_));
  NOR2_X1    g02264(.A1(new_n3265_), .A2(new_n3266_), .ZN(new_n3267_));
  NOR3_X1    g02265(.A1(new_n3267_), .A2(new_n3251_), .A3(new_n3262_), .ZN(new_n3268_));
  OAI21_X1   g02266(.A1(new_n3264_), .A2(new_n3268_), .B(new_n3208_), .ZN(new_n3269_));
  NOR2_X1    g02267(.A1(new_n3188_), .A2(new_n3175_), .ZN(new_n3270_));
  NAND4_X1   g02268(.A1(new_n3270_), .A2(new_n3181_), .A3(new_n3187_), .A4(new_n3184_), .ZN(new_n3271_));
  INV_X1     g02269(.I(new_n3195_), .ZN(new_n3272_));
  AOI21_X1   g02270(.A1(new_n3271_), .A2(new_n3272_), .B(new_n3198_), .ZN(new_n3273_));
  NAND2_X1   g02271(.A1(new_n3205_), .A2(new_n3201_), .ZN(new_n3274_));
  NAND2_X1   g02272(.A1(new_n3199_), .A2(new_n3194_), .ZN(new_n3275_));
  AOI21_X1   g02273(.A1(new_n3275_), .A2(new_n3274_), .B(new_n3166_), .ZN(new_n3276_));
  NOR2_X1    g02274(.A1(new_n3273_), .A2(new_n3276_), .ZN(new_n3277_));
  NOR2_X1    g02275(.A1(new_n3263_), .A2(new_n3267_), .ZN(new_n3278_));
  NOR3_X1    g02276(.A1(new_n3209_), .A2(new_n3251_), .A3(new_n3262_), .ZN(new_n3279_));
  OAI21_X1   g02277(.A1(new_n3278_), .A2(new_n3279_), .B(new_n3277_), .ZN(new_n3280_));
  NAND2_X1   g02278(.A1(new_n1394_), .A2(new_n1521_), .ZN(new_n3281_));
  INV_X1     g02279(.I(new_n3281_), .ZN(new_n3282_));
  NAND3_X1   g02280(.A1(new_n3282_), .A2(new_n3269_), .A3(new_n3280_), .ZN(new_n3283_));
  NAND2_X1   g02281(.A1(new_n3269_), .A2(new_n3280_), .ZN(new_n3284_));
  NAND2_X1   g02282(.A1(new_n3284_), .A2(new_n3281_), .ZN(new_n3285_));
  AOI21_X1   g02283(.A1(new_n3285_), .A2(new_n3283_), .B(new_n3150_), .ZN(new_n3286_));
  NAND3_X1   g02284(.A1(new_n3269_), .A2(new_n3280_), .A3(new_n3281_), .ZN(new_n3287_));
  NAND2_X1   g02285(.A1(new_n3284_), .A2(new_n3282_), .ZN(new_n3288_));
  AOI22_X1   g02286(.A1(new_n3288_), .A2(new_n3287_), .B1(new_n3130_), .B2(new_n3149_), .ZN(new_n3289_));
  NOR2_X1    g02287(.A1(new_n3289_), .A2(new_n3286_), .ZN(new_n3290_));
  AOI21_X1   g02288(.A1(new_n1240_), .A2(\A[897] ), .B(new_n1257_), .ZN(new_n3291_));
  NAND2_X1   g02289(.A1(new_n1254_), .A2(new_n3291_), .ZN(new_n3292_));
  AOI21_X1   g02290(.A1(new_n1248_), .A2(\A[900] ), .B(new_n1252_), .ZN(new_n3293_));
  NAND2_X1   g02291(.A1(new_n1259_), .A2(new_n3293_), .ZN(new_n3294_));
  NAND2_X1   g02292(.A1(new_n3292_), .A2(new_n3294_), .ZN(new_n3295_));
  NOR2_X1    g02293(.A1(new_n3293_), .A2(new_n3291_), .ZN(new_n3296_));
  AOI21_X1   g02294(.A1(new_n3295_), .A2(new_n1260_), .B(new_n3296_), .ZN(new_n3297_));
  INV_X1     g02295(.I(new_n3297_), .ZN(new_n3298_));
  NAND3_X1   g02296(.A1(new_n1260_), .A2(new_n3292_), .A3(new_n3294_), .ZN(new_n3299_));
  INV_X1     g02297(.I(new_n1260_), .ZN(new_n3300_));
  NAND2_X1   g02298(.A1(new_n3295_), .A2(new_n3300_), .ZN(new_n3301_));
  AOI22_X1   g02299(.A1(new_n3298_), .A2(new_n1250_), .B1(new_n3301_), .B2(new_n3299_), .ZN(new_n3302_));
  INV_X1     g02300(.I(new_n1231_), .ZN(new_n3303_));
  INV_X1     g02301(.I(new_n1261_), .ZN(new_n3304_));
  AOI21_X1   g02302(.A1(new_n1208_), .A2(\A[903] ), .B(new_n1227_), .ZN(new_n3305_));
  NAND2_X1   g02303(.A1(new_n1224_), .A2(new_n3305_), .ZN(new_n3306_));
  AOI21_X1   g02304(.A1(new_n1217_), .A2(\A[906] ), .B(new_n1222_), .ZN(new_n3307_));
  NAND2_X1   g02305(.A1(new_n1229_), .A2(new_n3307_), .ZN(new_n3308_));
  NAND3_X1   g02306(.A1(new_n1230_), .A2(new_n3306_), .A3(new_n3308_), .ZN(new_n3309_));
  NAND2_X1   g02307(.A1(new_n3306_), .A2(new_n3308_), .ZN(new_n3310_));
  INV_X1     g02308(.I(new_n1230_), .ZN(new_n3311_));
  NAND2_X1   g02309(.A1(new_n3310_), .A2(new_n3311_), .ZN(new_n3312_));
  NAND2_X1   g02310(.A1(new_n3312_), .A2(new_n3309_), .ZN(new_n3313_));
  NAND2_X1   g02311(.A1(new_n1207_), .A2(\A[903] ), .ZN(new_n3314_));
  OAI22_X1   g02312(.A1(new_n1226_), .A2(\A[903] ), .B1(new_n3314_), .B2(new_n1225_), .ZN(new_n3315_));
  XOR2_X1    g02313(.A1(new_n1218_), .A2(new_n3315_), .Z(new_n3316_));
  NAND2_X1   g02314(.A1(new_n1239_), .A2(\A[897] ), .ZN(new_n3317_));
  OAI22_X1   g02315(.A1(new_n1256_), .A2(\A[897] ), .B1(new_n3317_), .B2(new_n1255_), .ZN(new_n3318_));
  XOR2_X1    g02316(.A1(new_n3318_), .A2(new_n1249_), .Z(new_n3319_));
  NOR2_X1    g02317(.A1(new_n3316_), .A2(new_n3319_), .ZN(new_n3320_));
  NAND2_X1   g02318(.A1(new_n3313_), .A2(new_n3320_), .ZN(new_n3321_));
  NOR2_X1    g02319(.A1(new_n3307_), .A2(new_n3305_), .ZN(new_n3322_));
  AOI21_X1   g02320(.A1(new_n3310_), .A2(new_n1230_), .B(new_n3322_), .ZN(new_n3323_));
  NOR2_X1    g02321(.A1(new_n3323_), .A2(new_n3316_), .ZN(new_n3324_));
  NOR4_X1    g02322(.A1(new_n3321_), .A2(new_n3303_), .A3(new_n3304_), .A4(new_n3324_), .ZN(new_n3325_));
  NOR4_X1    g02323(.A1(new_n3303_), .A2(new_n3304_), .A3(new_n3316_), .A4(new_n3319_), .ZN(new_n3326_));
  INV_X1     g02324(.I(new_n3309_), .ZN(new_n3327_));
  AOI21_X1   g02325(.A1(new_n3306_), .A2(new_n3308_), .B(new_n1230_), .ZN(new_n3328_));
  NOR2_X1    g02326(.A1(new_n3327_), .A2(new_n3328_), .ZN(new_n3329_));
  NOR2_X1    g02327(.A1(new_n3324_), .A2(new_n3329_), .ZN(new_n3330_));
  NOR2_X1    g02328(.A1(new_n3330_), .A2(new_n3326_), .ZN(new_n3331_));
  OAI21_X1   g02329(.A1(new_n3325_), .A2(new_n3331_), .B(new_n3302_), .ZN(new_n3332_));
  INV_X1     g02330(.I(new_n3302_), .ZN(new_n3333_));
  NOR3_X1    g02331(.A1(new_n3326_), .A2(new_n3324_), .A3(new_n3329_), .ZN(new_n3334_));
  INV_X1     g02332(.I(new_n3326_), .ZN(new_n3335_));
  NOR2_X1    g02333(.A1(new_n3335_), .A2(new_n3330_), .ZN(new_n3336_));
  OAI21_X1   g02334(.A1(new_n3336_), .A2(new_n3334_), .B(new_n3333_), .ZN(new_n3337_));
  AND2_X2    g02335(.A1(new_n3337_), .A2(new_n3332_), .Z(new_n3338_));
  NAND2_X1   g02336(.A1(new_n1176_), .A2(\A[909] ), .ZN(new_n3339_));
  OAI22_X1   g02337(.A1(new_n1193_), .A2(\A[909] ), .B1(new_n3339_), .B2(new_n1192_), .ZN(new_n3340_));
  XOR2_X1    g02338(.A1(new_n3340_), .A2(new_n1186_), .Z(new_n3341_));
  AOI21_X1   g02339(.A1(new_n1177_), .A2(\A[909] ), .B(new_n1194_), .ZN(new_n3342_));
  NAND2_X1   g02340(.A1(new_n1191_), .A2(new_n3342_), .ZN(new_n3343_));
  AOI21_X1   g02341(.A1(new_n1185_), .A2(\A[912] ), .B(new_n1189_), .ZN(new_n3344_));
  NAND2_X1   g02342(.A1(new_n1196_), .A2(new_n3344_), .ZN(new_n3345_));
  NAND2_X1   g02343(.A1(new_n3343_), .A2(new_n3345_), .ZN(new_n3346_));
  NOR2_X1    g02344(.A1(new_n3344_), .A2(new_n3342_), .ZN(new_n3347_));
  AOI21_X1   g02345(.A1(new_n3346_), .A2(new_n1197_), .B(new_n3347_), .ZN(new_n3348_));
  NAND3_X1   g02346(.A1(new_n3343_), .A2(new_n1197_), .A3(new_n3345_), .ZN(new_n3349_));
  INV_X1     g02347(.I(new_n1186_), .ZN(new_n3350_));
  NAND2_X1   g02348(.A1(new_n3350_), .A2(new_n3340_), .ZN(new_n3351_));
  NAND2_X1   g02349(.A1(new_n3346_), .A2(new_n3351_), .ZN(new_n3352_));
  NAND2_X1   g02350(.A1(new_n3352_), .A2(new_n3349_), .ZN(new_n3353_));
  OAI21_X1   g02351(.A1(new_n3341_), .A2(new_n3348_), .B(new_n3353_), .ZN(new_n3354_));
  AOI21_X1   g02352(.A1(new_n1161_), .A2(\A[915] ), .B(new_n1156_), .ZN(new_n3355_));
  NAND2_X1   g02353(.A1(new_n1154_), .A2(new_n3355_), .ZN(new_n3356_));
  AOI21_X1   g02354(.A1(new_n1165_), .A2(\A[918] ), .B(new_n1152_), .ZN(new_n3357_));
  NAND2_X1   g02355(.A1(new_n1158_), .A2(new_n3357_), .ZN(new_n3358_));
  NAND2_X1   g02356(.A1(new_n3356_), .A2(new_n3358_), .ZN(new_n3359_));
  NAND2_X1   g02357(.A1(new_n1141_), .A2(new_n1149_), .ZN(new_n3360_));
  NOR2_X1    g02358(.A1(new_n3359_), .A2(new_n3360_), .ZN(new_n3361_));
  NOR2_X1    g02359(.A1(new_n1158_), .A2(new_n3357_), .ZN(new_n3362_));
  NOR2_X1    g02360(.A1(new_n1154_), .A2(new_n3355_), .ZN(new_n3363_));
  NOR2_X1    g02361(.A1(new_n3362_), .A2(new_n3363_), .ZN(new_n3364_));
  NOR2_X1    g02362(.A1(new_n3364_), .A2(new_n1167_), .ZN(new_n3365_));
  NOR2_X1    g02363(.A1(new_n3365_), .A2(new_n3361_), .ZN(new_n3366_));
  NAND2_X1   g02364(.A1(new_n1150_), .A2(new_n1187_), .ZN(new_n3367_));
  NOR2_X1    g02365(.A1(new_n3366_), .A2(new_n3367_), .ZN(new_n3368_));
  NOR2_X1    g02366(.A1(new_n3357_), .A2(new_n3355_), .ZN(new_n3369_));
  INV_X1     g02367(.I(new_n3369_), .ZN(new_n3370_));
  OAI21_X1   g02368(.A1(new_n3364_), .A2(new_n3360_), .B(new_n3370_), .ZN(new_n3371_));
  NAND2_X1   g02369(.A1(new_n3371_), .A2(new_n1150_), .ZN(new_n3372_));
  NAND4_X1   g02370(.A1(new_n3368_), .A2(new_n1168_), .A3(new_n1198_), .A4(new_n3372_), .ZN(new_n3373_));
  NAND4_X1   g02371(.A1(new_n1150_), .A2(new_n1187_), .A3(new_n1168_), .A4(new_n1198_), .ZN(new_n3374_));
  NAND3_X1   g02372(.A1(new_n1167_), .A2(new_n3356_), .A3(new_n3358_), .ZN(new_n3375_));
  OAI21_X1   g02373(.A1(new_n3362_), .A2(new_n3363_), .B(new_n3360_), .ZN(new_n3376_));
  NAND2_X1   g02374(.A1(new_n3376_), .A2(new_n3375_), .ZN(new_n3377_));
  NAND2_X1   g02375(.A1(new_n3372_), .A2(new_n3377_), .ZN(new_n3378_));
  NAND2_X1   g02376(.A1(new_n3378_), .A2(new_n3374_), .ZN(new_n3379_));
  AOI21_X1   g02377(.A1(new_n3373_), .A2(new_n3379_), .B(new_n3354_), .ZN(new_n3380_));
  INV_X1     g02378(.I(new_n3348_), .ZN(new_n3381_));
  INV_X1     g02379(.I(new_n3349_), .ZN(new_n3382_));
  AOI21_X1   g02380(.A1(new_n3343_), .A2(new_n3345_), .B(new_n1197_), .ZN(new_n3383_));
  NOR2_X1    g02381(.A1(new_n3382_), .A2(new_n3383_), .ZN(new_n3384_));
  AOI21_X1   g02382(.A1(new_n1187_), .A2(new_n3381_), .B(new_n3384_), .ZN(new_n3385_));
  XOR2_X1    g02383(.A1(new_n1162_), .A2(new_n1149_), .Z(new_n3386_));
  NOR3_X1    g02384(.A1(new_n3360_), .A2(new_n3357_), .A3(new_n3355_), .ZN(new_n3387_));
  NOR3_X1    g02385(.A1(new_n3351_), .A2(new_n3344_), .A3(new_n3342_), .ZN(new_n3388_));
  NOR4_X1    g02386(.A1(new_n3388_), .A2(new_n3386_), .A3(new_n3341_), .A4(new_n3387_), .ZN(new_n3389_));
  NAND2_X1   g02387(.A1(new_n3378_), .A2(new_n3389_), .ZN(new_n3390_));
  NAND3_X1   g02388(.A1(new_n3372_), .A2(new_n3374_), .A3(new_n3377_), .ZN(new_n3391_));
  AOI21_X1   g02389(.A1(new_n3390_), .A2(new_n3391_), .B(new_n3385_), .ZN(new_n3392_));
  NAND2_X1   g02390(.A1(new_n1200_), .A2(new_n1263_), .ZN(new_n3393_));
  NOR3_X1    g02391(.A1(new_n3380_), .A2(new_n3392_), .A3(new_n3393_), .ZN(new_n3394_));
  AOI21_X1   g02392(.A1(new_n3359_), .A2(new_n1167_), .B(new_n3369_), .ZN(new_n3395_));
  NAND4_X1   g02393(.A1(new_n3377_), .A2(new_n1150_), .A3(new_n3395_), .A4(new_n1187_), .ZN(new_n3396_));
  NOR2_X1    g02394(.A1(new_n3395_), .A2(new_n3386_), .ZN(new_n3397_));
  NOR3_X1    g02395(.A1(new_n3396_), .A2(new_n3388_), .A3(new_n3397_), .ZN(new_n3398_));
  AOI21_X1   g02396(.A1(new_n3377_), .A2(new_n3372_), .B(new_n3389_), .ZN(new_n3399_));
  OAI21_X1   g02397(.A1(new_n3398_), .A2(new_n3399_), .B(new_n3385_), .ZN(new_n3400_));
  NOR2_X1    g02398(.A1(new_n3397_), .A2(new_n3366_), .ZN(new_n3401_));
  NOR2_X1    g02399(.A1(new_n3401_), .A2(new_n3374_), .ZN(new_n3402_));
  INV_X1     g02400(.I(new_n3391_), .ZN(new_n3403_));
  OAI21_X1   g02401(.A1(new_n3402_), .A2(new_n3403_), .B(new_n3354_), .ZN(new_n3404_));
  XNOR2_X1   g02402(.A1(new_n1169_), .A2(new_n1199_), .ZN(new_n3405_));
  XNOR2_X1   g02403(.A1(new_n1232_), .A2(new_n1262_), .ZN(new_n3406_));
  NOR2_X1    g02404(.A1(new_n3406_), .A2(new_n3405_), .ZN(new_n3407_));
  AOI21_X1   g02405(.A1(new_n3400_), .A2(new_n3404_), .B(new_n3407_), .ZN(new_n3408_));
  OAI21_X1   g02406(.A1(new_n3408_), .A2(new_n3394_), .B(new_n3338_), .ZN(new_n3409_));
  NAND2_X1   g02407(.A1(new_n3337_), .A2(new_n3332_), .ZN(new_n3410_));
  NAND3_X1   g02408(.A1(new_n3404_), .A2(new_n3393_), .A3(new_n3400_), .ZN(new_n3411_));
  OAI21_X1   g02409(.A1(new_n3380_), .A2(new_n3392_), .B(new_n3407_), .ZN(new_n3412_));
  NAND2_X1   g02410(.A1(new_n3412_), .A2(new_n3411_), .ZN(new_n3413_));
  NAND2_X1   g02411(.A1(new_n3413_), .A2(new_n3410_), .ZN(new_n3414_));
  NAND2_X1   g02412(.A1(new_n3409_), .A2(new_n3414_), .ZN(new_n3415_));
  INV_X1     g02413(.I(new_n3415_), .ZN(new_n3416_));
  AOI21_X1   g02414(.A1(new_n1109_), .A2(\A[921] ), .B(new_n1126_), .ZN(new_n3417_));
  NAND2_X1   g02415(.A1(new_n1123_), .A2(new_n3417_), .ZN(new_n3418_));
  AOI21_X1   g02416(.A1(new_n1117_), .A2(\A[924] ), .B(new_n1121_), .ZN(new_n3419_));
  NAND2_X1   g02417(.A1(new_n1128_), .A2(new_n3419_), .ZN(new_n3420_));
  NAND2_X1   g02418(.A1(new_n3418_), .A2(new_n3420_), .ZN(new_n3421_));
  NAND2_X1   g02419(.A1(new_n3421_), .A2(new_n1129_), .ZN(new_n3422_));
  NOR2_X1    g02420(.A1(new_n3419_), .A2(new_n3417_), .ZN(new_n3423_));
  INV_X1     g02421(.I(new_n3423_), .ZN(new_n3424_));
  NAND2_X1   g02422(.A1(new_n3422_), .A2(new_n3424_), .ZN(new_n3425_));
  OR2_X2     g02423(.A1(new_n1110_), .A2(new_n1118_), .Z(new_n3426_));
  NOR2_X1    g02424(.A1(new_n3421_), .A2(new_n3426_), .ZN(new_n3427_));
  AOI21_X1   g02425(.A1(new_n3418_), .A2(new_n3420_), .B(new_n1129_), .ZN(new_n3428_));
  NOR2_X1    g02426(.A1(new_n3427_), .A2(new_n3428_), .ZN(new_n3429_));
  AOI21_X1   g02427(.A1(new_n1119_), .A2(new_n3425_), .B(new_n3429_), .ZN(new_n3430_));
  AOI21_X1   g02428(.A1(new_n1079_), .A2(\A[927] ), .B(new_n1096_), .ZN(new_n3431_));
  NAND2_X1   g02429(.A1(new_n1093_), .A2(new_n3431_), .ZN(new_n3432_));
  AOI21_X1   g02430(.A1(new_n1087_), .A2(\A[930] ), .B(new_n1091_), .ZN(new_n3433_));
  NAND2_X1   g02431(.A1(new_n1098_), .A2(new_n3433_), .ZN(new_n3434_));
  NAND3_X1   g02432(.A1(new_n3432_), .A2(new_n1099_), .A3(new_n3434_), .ZN(new_n3435_));
  INV_X1     g02433(.I(new_n3435_), .ZN(new_n3436_));
  AOI21_X1   g02434(.A1(new_n3432_), .A2(new_n3434_), .B(new_n1099_), .ZN(new_n3437_));
  NOR2_X1    g02435(.A1(new_n3436_), .A2(new_n3437_), .ZN(new_n3438_));
  XOR2_X1    g02436(.A1(new_n1098_), .A2(new_n3433_), .Z(new_n3439_));
  INV_X1     g02437(.I(new_n1099_), .ZN(new_n3440_));
  NOR2_X1    g02438(.A1(new_n3433_), .A2(new_n3431_), .ZN(new_n3441_));
  INV_X1     g02439(.I(new_n3441_), .ZN(new_n3442_));
  OAI21_X1   g02440(.A1(new_n3439_), .A2(new_n3440_), .B(new_n3442_), .ZN(new_n3443_));
  NAND2_X1   g02441(.A1(new_n1089_), .A2(new_n1119_), .ZN(new_n3444_));
  INV_X1     g02442(.I(new_n1089_), .ZN(new_n3445_));
  NAND2_X1   g02443(.A1(new_n3432_), .A2(new_n3434_), .ZN(new_n3446_));
  AOI21_X1   g02444(.A1(new_n3446_), .A2(new_n1099_), .B(new_n3441_), .ZN(new_n3447_));
  OAI21_X1   g02445(.A1(new_n3447_), .A2(new_n3445_), .B(new_n1130_), .ZN(new_n3448_));
  NOR4_X1    g02446(.A1(new_n3448_), .A2(new_n3438_), .A3(new_n3443_), .A4(new_n3444_), .ZN(new_n3449_));
  NAND2_X1   g02447(.A1(new_n3446_), .A2(new_n3440_), .ZN(new_n3450_));
  NAND2_X1   g02448(.A1(new_n3450_), .A2(new_n3435_), .ZN(new_n3451_));
  NAND2_X1   g02449(.A1(new_n3443_), .A2(new_n1089_), .ZN(new_n3452_));
  NAND4_X1   g02450(.A1(new_n1089_), .A2(new_n1119_), .A3(new_n1100_), .A4(new_n1130_), .ZN(new_n3453_));
  INV_X1     g02451(.I(new_n3453_), .ZN(new_n3454_));
  AOI21_X1   g02452(.A1(new_n3451_), .A2(new_n3452_), .B(new_n3454_), .ZN(new_n3455_));
  OAI21_X1   g02453(.A1(new_n3455_), .A2(new_n3449_), .B(new_n3430_), .ZN(new_n3456_));
  XOR2_X1    g02454(.A1(new_n3421_), .A2(new_n1129_), .Z(new_n3457_));
  AOI21_X1   g02455(.A1(new_n3418_), .A2(new_n3420_), .B(new_n3426_), .ZN(new_n3458_));
  OAI21_X1   g02456(.A1(new_n3458_), .A2(new_n3423_), .B(new_n1119_), .ZN(new_n3459_));
  NAND2_X1   g02457(.A1(new_n3457_), .A2(new_n3459_), .ZN(new_n3460_));
  NOR2_X1    g02458(.A1(new_n3447_), .A2(new_n3445_), .ZN(new_n3461_));
  NOR3_X1    g02459(.A1(new_n3454_), .A2(new_n3461_), .A3(new_n3438_), .ZN(new_n3462_));
  AOI21_X1   g02460(.A1(new_n3452_), .A2(new_n3451_), .B(new_n3453_), .ZN(new_n3463_));
  OAI21_X1   g02461(.A1(new_n3462_), .A2(new_n3463_), .B(new_n3460_), .ZN(new_n3464_));
  NAND2_X1   g02462(.A1(new_n3456_), .A2(new_n3464_), .ZN(new_n3465_));
  XNOR2_X1   g02463(.A1(new_n1038_), .A2(new_n1070_), .ZN(new_n3466_));
  XNOR2_X1   g02464(.A1(new_n1101_), .A2(new_n1131_), .ZN(new_n3467_));
  NOR2_X1    g02465(.A1(new_n3466_), .A2(new_n3467_), .ZN(new_n3468_));
  NAND2_X1   g02466(.A1(new_n1045_), .A2(\A[933] ), .ZN(new_n3469_));
  OAI22_X1   g02467(.A1(new_n1064_), .A2(\A[933] ), .B1(new_n3469_), .B2(new_n1063_), .ZN(new_n3470_));
  XOR2_X1    g02468(.A1(new_n3470_), .A2(new_n1055_), .Z(new_n3471_));
  AOI21_X1   g02469(.A1(new_n1046_), .A2(\A[933] ), .B(new_n1065_), .ZN(new_n3472_));
  NAND2_X1   g02470(.A1(new_n1062_), .A2(new_n3472_), .ZN(new_n3473_));
  AOI21_X1   g02471(.A1(new_n1054_), .A2(\A[936] ), .B(new_n1060_), .ZN(new_n3474_));
  NAND2_X1   g02472(.A1(new_n1067_), .A2(new_n3474_), .ZN(new_n3475_));
  NAND2_X1   g02473(.A1(new_n3473_), .A2(new_n3475_), .ZN(new_n3476_));
  NOR2_X1    g02474(.A1(new_n3474_), .A2(new_n3472_), .ZN(new_n3477_));
  AOI21_X1   g02475(.A1(new_n3476_), .A2(new_n1068_), .B(new_n3477_), .ZN(new_n3478_));
  NAND3_X1   g02476(.A1(new_n1068_), .A2(new_n3473_), .A3(new_n3475_), .ZN(new_n3479_));
  NOR2_X1    g02477(.A1(new_n1067_), .A2(new_n3474_), .ZN(new_n3480_));
  NOR2_X1    g02478(.A1(new_n1062_), .A2(new_n3472_), .ZN(new_n3481_));
  NAND2_X1   g02479(.A1(new_n1053_), .A2(\A[936] ), .ZN(new_n3482_));
  OAI22_X1   g02480(.A1(new_n1059_), .A2(\A[936] ), .B1(new_n3482_), .B2(new_n1057_), .ZN(new_n3483_));
  NAND2_X1   g02481(.A1(new_n3470_), .A2(new_n3483_), .ZN(new_n3484_));
  OAI21_X1   g02482(.A1(new_n3480_), .A2(new_n3481_), .B(new_n3484_), .ZN(new_n3485_));
  NAND2_X1   g02483(.A1(new_n3485_), .A2(new_n3479_), .ZN(new_n3486_));
  OAI21_X1   g02484(.A1(new_n3471_), .A2(new_n3478_), .B(new_n3486_), .ZN(new_n3487_));
  AOI21_X1   g02485(.A1(new_n1030_), .A2(\A[939] ), .B(new_n1025_), .ZN(new_n3488_));
  NAND2_X1   g02486(.A1(new_n1023_), .A2(new_n3488_), .ZN(new_n3489_));
  AOI21_X1   g02487(.A1(new_n1034_), .A2(\A[942] ), .B(new_n1021_), .ZN(new_n3490_));
  NAND2_X1   g02488(.A1(new_n1027_), .A2(new_n3490_), .ZN(new_n3491_));
  NAND3_X1   g02489(.A1(new_n1036_), .A2(new_n3489_), .A3(new_n3491_), .ZN(new_n3492_));
  NOR2_X1    g02490(.A1(new_n1027_), .A2(new_n3490_), .ZN(new_n3493_));
  NOR2_X1    g02491(.A1(new_n1023_), .A2(new_n3488_), .ZN(new_n3494_));
  NAND2_X1   g02492(.A1(new_n1010_), .A2(new_n1018_), .ZN(new_n3495_));
  OAI21_X1   g02493(.A1(new_n3493_), .A2(new_n3494_), .B(new_n3495_), .ZN(new_n3496_));
  NAND2_X1   g02494(.A1(new_n3496_), .A2(new_n3492_), .ZN(new_n3497_));
  NAND2_X1   g02495(.A1(new_n3489_), .A2(new_n3491_), .ZN(new_n3498_));
  NOR2_X1    g02496(.A1(new_n3490_), .A2(new_n3488_), .ZN(new_n3499_));
  AOI21_X1   g02497(.A1(new_n3498_), .A2(new_n1036_), .B(new_n3499_), .ZN(new_n3500_));
  XOR2_X1    g02498(.A1(new_n1031_), .A2(new_n1018_), .Z(new_n3501_));
  NOR2_X1    g02499(.A1(new_n3501_), .A2(new_n3471_), .ZN(new_n3502_));
  NOR2_X1    g02500(.A1(new_n3493_), .A2(new_n3494_), .ZN(new_n3503_));
  INV_X1     g02501(.I(new_n3499_), .ZN(new_n3504_));
  OAI21_X1   g02502(.A1(new_n3503_), .A2(new_n3495_), .B(new_n3504_), .ZN(new_n3505_));
  NOR3_X1    g02503(.A1(new_n3484_), .A2(new_n3474_), .A3(new_n3472_), .ZN(new_n3506_));
  AOI21_X1   g02504(.A1(new_n3505_), .A2(new_n1019_), .B(new_n3506_), .ZN(new_n3507_));
  NAND4_X1   g02505(.A1(new_n3507_), .A2(new_n3497_), .A3(new_n3500_), .A4(new_n3502_), .ZN(new_n3508_));
  NAND2_X1   g02506(.A1(new_n3505_), .A2(new_n1019_), .ZN(new_n3509_));
  NOR3_X1    g02507(.A1(new_n3495_), .A2(new_n3490_), .A3(new_n3488_), .ZN(new_n3510_));
  NOR4_X1    g02508(.A1(new_n3501_), .A2(new_n3471_), .A3(new_n3510_), .A4(new_n3506_), .ZN(new_n3511_));
  AOI21_X1   g02509(.A1(new_n3497_), .A2(new_n3509_), .B(new_n3511_), .ZN(new_n3512_));
  INV_X1     g02510(.I(new_n3512_), .ZN(new_n3513_));
  AOI21_X1   g02511(.A1(new_n3513_), .A2(new_n3508_), .B(new_n3487_), .ZN(new_n3514_));
  INV_X1     g02512(.I(new_n3478_), .ZN(new_n3515_));
  AOI22_X1   g02513(.A1(new_n3515_), .A2(new_n1056_), .B1(new_n3479_), .B2(new_n3485_), .ZN(new_n3516_));
  NAND4_X1   g02514(.A1(new_n1019_), .A2(new_n1056_), .A3(new_n1037_), .A4(new_n1069_), .ZN(new_n3517_));
  AOI21_X1   g02515(.A1(new_n3509_), .A2(new_n3497_), .B(new_n3517_), .ZN(new_n3518_));
  INV_X1     g02516(.I(new_n3518_), .ZN(new_n3519_));
  NAND3_X1   g02517(.A1(new_n3509_), .A2(new_n3517_), .A3(new_n3497_), .ZN(new_n3520_));
  AOI21_X1   g02518(.A1(new_n3519_), .A2(new_n3520_), .B(new_n3516_), .ZN(new_n3521_));
  OAI21_X1   g02519(.A1(new_n3514_), .A2(new_n3521_), .B(new_n3468_), .ZN(new_n3522_));
  NAND2_X1   g02520(.A1(new_n1071_), .A2(new_n1132_), .ZN(new_n3523_));
  NAND2_X1   g02521(.A1(new_n3502_), .A2(new_n3497_), .ZN(new_n3524_));
  NOR2_X1    g02522(.A1(new_n3500_), .A2(new_n3501_), .ZN(new_n3525_));
  NOR4_X1    g02523(.A1(new_n3524_), .A2(new_n3510_), .A3(new_n3506_), .A4(new_n3525_), .ZN(new_n3526_));
  OAI21_X1   g02524(.A1(new_n3526_), .A2(new_n3512_), .B(new_n3516_), .ZN(new_n3527_));
  INV_X1     g02525(.I(new_n3520_), .ZN(new_n3528_));
  OAI21_X1   g02526(.A1(new_n3528_), .A2(new_n3518_), .B(new_n3487_), .ZN(new_n3529_));
  NAND3_X1   g02527(.A1(new_n3523_), .A2(new_n3529_), .A3(new_n3527_), .ZN(new_n3530_));
  NAND2_X1   g02528(.A1(new_n3522_), .A2(new_n3530_), .ZN(new_n3531_));
  NAND2_X1   g02529(.A1(new_n3531_), .A2(new_n3465_), .ZN(new_n3532_));
  INV_X1     g02530(.I(new_n3465_), .ZN(new_n3533_));
  AOI21_X1   g02531(.A1(new_n3527_), .A2(new_n3529_), .B(new_n3468_), .ZN(new_n3534_));
  NOR3_X1    g02532(.A1(new_n3514_), .A2(new_n3521_), .A3(new_n3523_), .ZN(new_n3535_));
  OAI21_X1   g02533(.A1(new_n3534_), .A2(new_n3535_), .B(new_n3533_), .ZN(new_n3536_));
  NAND2_X1   g02534(.A1(new_n1133_), .A2(new_n1264_), .ZN(new_n3537_));
  NAND3_X1   g02535(.A1(new_n3532_), .A2(new_n3536_), .A3(new_n3537_), .ZN(new_n3538_));
  AOI21_X1   g02536(.A1(new_n3522_), .A2(new_n3530_), .B(new_n3533_), .ZN(new_n3539_));
  NOR2_X1    g02537(.A1(new_n3534_), .A2(new_n3535_), .ZN(new_n3540_));
  NOR2_X1    g02538(.A1(new_n3540_), .A2(new_n3465_), .ZN(new_n3541_));
  AND2_X2    g02539(.A1(new_n1133_), .A2(new_n1264_), .Z(new_n3542_));
  OAI21_X1   g02540(.A1(new_n3541_), .A2(new_n3539_), .B(new_n3542_), .ZN(new_n3543_));
  AOI21_X1   g02541(.A1(new_n3538_), .A2(new_n3543_), .B(new_n3416_), .ZN(new_n3544_));
  NOR3_X1    g02542(.A1(new_n3541_), .A2(new_n3539_), .A3(new_n3537_), .ZN(new_n3545_));
  AOI21_X1   g02543(.A1(new_n3532_), .A2(new_n3536_), .B(new_n3542_), .ZN(new_n3546_));
  NOR2_X1    g02544(.A1(new_n3545_), .A2(new_n3546_), .ZN(new_n3547_));
  NOR2_X1    g02545(.A1(new_n3547_), .A2(new_n3415_), .ZN(new_n3548_));
  NOR2_X1    g02546(.A1(new_n1265_), .A2(new_n1522_), .ZN(new_n3549_));
  INV_X1     g02547(.I(new_n3549_), .ZN(new_n3550_));
  NOR3_X1    g02548(.A1(new_n3548_), .A2(new_n3544_), .A3(new_n3550_), .ZN(new_n3551_));
  NAND2_X1   g02549(.A1(new_n3543_), .A2(new_n3538_), .ZN(new_n3552_));
  NAND2_X1   g02550(.A1(new_n3552_), .A2(new_n3415_), .ZN(new_n3553_));
  OAI21_X1   g02551(.A1(new_n3545_), .A2(new_n3546_), .B(new_n3416_), .ZN(new_n3554_));
  AOI21_X1   g02552(.A1(new_n3554_), .A2(new_n3553_), .B(new_n3549_), .ZN(new_n3555_));
  OAI21_X1   g02553(.A1(new_n3551_), .A2(new_n3555_), .B(new_n3290_), .ZN(new_n3556_));
  NOR3_X1    g02554(.A1(new_n3548_), .A2(new_n3544_), .A3(new_n3549_), .ZN(new_n3557_));
  AOI21_X1   g02555(.A1(new_n3554_), .A2(new_n3553_), .B(new_n3550_), .ZN(new_n3558_));
  OAI22_X1   g02556(.A1(new_n3557_), .A2(new_n3558_), .B1(new_n3286_), .B2(new_n3289_), .ZN(new_n3559_));
  NAND2_X1   g02557(.A1(new_n3559_), .A2(new_n3556_), .ZN(new_n3560_));
  NAND3_X1   g02558(.A1(new_n3027_), .A2(new_n3031_), .A3(new_n2346_), .ZN(new_n3561_));
  AOI21_X1   g02559(.A1(new_n3560_), .A2(new_n3561_), .B(new_n3032_), .ZN(new_n3562_));
  OAI22_X1   g02560(.A1(new_n2541_), .A2(new_n2435_), .B1(new_n2535_), .B2(new_n2537_), .ZN(new_n3563_));
  INV_X1     g02561(.I(new_n3563_), .ZN(new_n3564_));
  NOR3_X1    g02562(.A1(new_n2428_), .A2(new_n2432_), .A3(new_n2415_), .ZN(new_n3565_));
  OAI21_X1   g02563(.A1(new_n2423_), .A2(new_n3565_), .B(new_n2433_), .ZN(new_n3566_));
  AND2_X2    g02564(.A1(new_n2356_), .A2(new_n2357_), .Z(new_n3567_));
  OAI22_X1   g02565(.A1(new_n2369_), .A2(new_n2361_), .B1(new_n3567_), .B2(new_n2358_), .ZN(new_n3568_));
  AOI21_X1   g02566(.A1(new_n2373_), .A2(new_n1714_), .B(new_n2353_), .ZN(new_n3569_));
  NAND2_X1   g02567(.A1(new_n3568_), .A2(new_n3569_), .ZN(new_n3570_));
  AOI21_X1   g02568(.A1(new_n2360_), .A2(new_n1691_), .B(new_n2359_), .ZN(new_n3571_));
  AND2_X2    g02569(.A1(new_n2347_), .A2(new_n2348_), .Z(new_n3572_));
  OAI22_X1   g02570(.A1(new_n2350_), .A2(new_n2351_), .B1(new_n3572_), .B2(new_n2352_), .ZN(new_n3573_));
  NAND2_X1   g02571(.A1(new_n3573_), .A2(new_n3571_), .ZN(new_n3574_));
  NAND2_X1   g02572(.A1(new_n3570_), .A2(new_n3574_), .ZN(new_n3575_));
  OAI21_X1   g02573(.A1(new_n2368_), .A2(new_n2370_), .B(new_n2355_), .ZN(new_n3576_));
  NAND2_X1   g02574(.A1(new_n3576_), .A2(new_n2366_), .ZN(new_n3577_));
  NOR2_X1    g02575(.A1(new_n3573_), .A2(new_n3571_), .ZN(new_n3578_));
  NOR2_X1    g02576(.A1(new_n3568_), .A2(new_n3569_), .ZN(new_n3579_));
  NOR3_X1    g02577(.A1(new_n2367_), .A2(new_n3579_), .A3(new_n3578_), .ZN(new_n3580_));
  AOI22_X1   g02578(.A1(new_n3580_), .A2(new_n3576_), .B1(new_n3575_), .B2(new_n3577_), .ZN(new_n3581_));
  AOI21_X1   g02579(.A1(new_n2394_), .A2(new_n1643_), .B(new_n2399_), .ZN(new_n3582_));
  XNOR2_X1   g02580(.A1(new_n1669_), .A2(new_n1671_), .ZN(new_n3583_));
  NOR2_X1    g02581(.A1(new_n3583_), .A2(new_n2383_), .ZN(new_n3584_));
  OAI22_X1   g02582(.A1(new_n2384_), .A2(new_n2385_), .B1(new_n3584_), .B2(new_n2386_), .ZN(new_n3585_));
  NOR2_X1    g02583(.A1(new_n3585_), .A2(new_n3582_), .ZN(new_n3586_));
  AND2_X2    g02584(.A1(new_n2392_), .A2(new_n2393_), .Z(new_n3587_));
  OAI22_X1   g02585(.A1(new_n2404_), .A2(new_n2395_), .B1(new_n3587_), .B2(new_n2398_), .ZN(new_n3588_));
  AOI21_X1   g02586(.A1(new_n2408_), .A2(new_n1667_), .B(new_n2387_), .ZN(new_n3589_));
  NOR2_X1    g02587(.A1(new_n3588_), .A2(new_n3589_), .ZN(new_n3590_));
  NOR2_X1    g02588(.A1(new_n2406_), .A2(new_n2409_), .ZN(new_n3591_));
  OAI22_X1   g02589(.A1(new_n3591_), .A2(new_n2401_), .B1(new_n3586_), .B2(new_n3590_), .ZN(new_n3592_));
  NAND2_X1   g02590(.A1(new_n3588_), .A2(new_n3589_), .ZN(new_n3593_));
  NAND2_X1   g02591(.A1(new_n3585_), .A2(new_n3582_), .ZN(new_n3594_));
  OAI21_X1   g02592(.A1(new_n2402_), .A2(new_n2405_), .B(new_n2389_), .ZN(new_n3595_));
  NAND4_X1   g02593(.A1(new_n3593_), .A2(new_n3595_), .A3(new_n3594_), .A4(new_n2426_), .ZN(new_n3596_));
  NAND2_X1   g02594(.A1(new_n3592_), .A2(new_n3596_), .ZN(new_n3597_));
  NOR2_X1    g02595(.A1(new_n3581_), .A2(new_n3597_), .ZN(new_n3598_));
  AOI21_X1   g02596(.A1(new_n2377_), .A2(new_n2375_), .B(new_n2374_), .ZN(new_n3599_));
  OAI22_X1   g02597(.A1(new_n3599_), .A2(new_n2367_), .B1(new_n3578_), .B2(new_n3579_), .ZN(new_n3600_));
  NAND4_X1   g02598(.A1(new_n3576_), .A2(new_n3570_), .A3(new_n3574_), .A4(new_n2366_), .ZN(new_n3601_));
  NAND2_X1   g02599(.A1(new_n3600_), .A2(new_n3601_), .ZN(new_n3602_));
  NAND2_X1   g02600(.A1(new_n3593_), .A2(new_n3594_), .ZN(new_n3603_));
  NAND2_X1   g02601(.A1(new_n3595_), .A2(new_n2426_), .ZN(new_n3604_));
  NOR3_X1    g02602(.A1(new_n3586_), .A2(new_n3590_), .A3(new_n2401_), .ZN(new_n3605_));
  AOI22_X1   g02603(.A1(new_n3605_), .A2(new_n3595_), .B1(new_n3603_), .B2(new_n3604_), .ZN(new_n3606_));
  NOR2_X1    g02604(.A1(new_n3602_), .A2(new_n3606_), .ZN(new_n3607_));
  OAI21_X1   g02605(.A1(new_n3598_), .A2(new_n3607_), .B(new_n3566_), .ZN(new_n3608_));
  AOI22_X1   g02606(.A1(new_n2380_), .A2(new_n2424_), .B1(new_n2415_), .B2(new_n2417_), .ZN(new_n3609_));
  NAND2_X1   g02607(.A1(new_n3602_), .A2(new_n3606_), .ZN(new_n3610_));
  NAND2_X1   g02608(.A1(new_n3581_), .A2(new_n3597_), .ZN(new_n3611_));
  NAND3_X1   g02609(.A1(new_n3610_), .A2(new_n3611_), .A3(new_n3609_), .ZN(new_n3612_));
  NAND2_X1   g02610(.A1(new_n3608_), .A2(new_n3612_), .ZN(new_n3613_));
  AOI21_X1   g02611(.A1(new_n2496_), .A2(new_n2511_), .B(new_n2512_), .ZN(new_n3614_));
  AOI21_X1   g02612(.A1(new_n2471_), .A2(new_n2532_), .B(new_n3614_), .ZN(new_n3615_));
  AOI21_X1   g02613(.A1(new_n2465_), .A2(new_n1598_), .B(new_n2453_), .ZN(new_n3616_));
  XNOR2_X1   g02614(.A1(new_n1618_), .A2(new_n1620_), .ZN(new_n3617_));
  INV_X1     g02615(.I(new_n2440_), .ZN(new_n3618_));
  OAI21_X1   g02616(.A1(new_n3617_), .A2(new_n2461_), .B(new_n3618_), .ZN(new_n3619_));
  OAI21_X1   g02617(.A1(new_n2462_), .A2(new_n2437_), .B(new_n3619_), .ZN(new_n3620_));
  NOR2_X1    g02618(.A1(new_n3616_), .A2(new_n3620_), .ZN(new_n3621_));
  AND2_X2    g02619(.A1(new_n2450_), .A2(new_n1596_), .Z(new_n3622_));
  OAI22_X1   g02620(.A1(new_n2451_), .A2(new_n2454_), .B1(new_n2452_), .B2(new_n3622_), .ZN(new_n3623_));
  AOI21_X1   g02621(.A1(new_n2442_), .A2(new_n1616_), .B(new_n2441_), .ZN(new_n3624_));
  NOR2_X1    g02622(.A1(new_n3623_), .A2(new_n3624_), .ZN(new_n3625_));
  NOR2_X1    g02623(.A1(new_n2469_), .A2(new_n2443_), .ZN(new_n3626_));
  OAI22_X1   g02624(.A1(new_n3626_), .A2(new_n2468_), .B1(new_n3625_), .B2(new_n3621_), .ZN(new_n3627_));
  NAND2_X1   g02625(.A1(new_n3623_), .A2(new_n3624_), .ZN(new_n3628_));
  NAND2_X1   g02626(.A1(new_n3616_), .A2(new_n3620_), .ZN(new_n3629_));
  OAI21_X1   g02627(.A1(new_n2447_), .A2(new_n2456_), .B(new_n2464_), .ZN(new_n3630_));
  NAND4_X1   g02628(.A1(new_n3628_), .A2(new_n3630_), .A3(new_n3629_), .A4(new_n2528_), .ZN(new_n3631_));
  NAND2_X1   g02629(.A1(new_n3627_), .A2(new_n3631_), .ZN(new_n3632_));
  OAI21_X1   g02630(.A1(new_n2493_), .A2(new_n2484_), .B(new_n2505_), .ZN(new_n3633_));
  AOI21_X1   g02631(.A1(new_n2497_), .A2(new_n1566_), .B(new_n2478_), .ZN(new_n3634_));
  NAND2_X1   g02632(.A1(new_n3634_), .A2(new_n3633_), .ZN(new_n3635_));
  AOI21_X1   g02633(.A1(new_n2483_), .A2(new_n1548_), .B(new_n2488_), .ZN(new_n3636_));
  OAI21_X1   g02634(.A1(new_n2475_), .A2(new_n2476_), .B(new_n2500_), .ZN(new_n3637_));
  NAND2_X1   g02635(.A1(new_n3636_), .A2(new_n3637_), .ZN(new_n3638_));
  OAI21_X1   g02636(.A1(new_n2491_), .A2(new_n2494_), .B(new_n2480_), .ZN(new_n3639_));
  AOI22_X1   g02637(.A1(new_n3635_), .A2(new_n3638_), .B1(new_n3639_), .B2(new_n2516_), .ZN(new_n3640_));
  NOR2_X1    g02638(.A1(new_n3636_), .A2(new_n3637_), .ZN(new_n3641_));
  NOR2_X1    g02639(.A1(new_n3634_), .A2(new_n3633_), .ZN(new_n3642_));
  AOI21_X1   g02640(.A1(new_n2509_), .A2(new_n2507_), .B(new_n2502_), .ZN(new_n3643_));
  NOR4_X1    g02641(.A1(new_n3641_), .A2(new_n3643_), .A3(new_n3642_), .A4(new_n2490_), .ZN(new_n3644_));
  NOR2_X1    g02642(.A1(new_n3644_), .A2(new_n3640_), .ZN(new_n3645_));
  NAND2_X1   g02643(.A1(new_n3632_), .A2(new_n3645_), .ZN(new_n3646_));
  NAND2_X1   g02644(.A1(new_n3628_), .A2(new_n3629_), .ZN(new_n3647_));
  NAND2_X1   g02645(.A1(new_n3630_), .A2(new_n2528_), .ZN(new_n3648_));
  NOR3_X1    g02646(.A1(new_n2468_), .A2(new_n3625_), .A3(new_n3621_), .ZN(new_n3649_));
  AOI22_X1   g02647(.A1(new_n3649_), .A2(new_n3630_), .B1(new_n3647_), .B2(new_n3648_), .ZN(new_n3650_));
  OAI22_X1   g02648(.A1(new_n3641_), .A2(new_n3642_), .B1(new_n3643_), .B2(new_n2490_), .ZN(new_n3651_));
  NAND4_X1   g02649(.A1(new_n3635_), .A2(new_n3639_), .A3(new_n3638_), .A4(new_n2516_), .ZN(new_n3652_));
  NAND2_X1   g02650(.A1(new_n3651_), .A2(new_n3652_), .ZN(new_n3653_));
  NAND2_X1   g02651(.A1(new_n3650_), .A2(new_n3653_), .ZN(new_n3654_));
  AOI21_X1   g02652(.A1(new_n3646_), .A2(new_n3654_), .B(new_n3615_), .ZN(new_n3655_));
  NOR3_X1    g02653(.A1(new_n2518_), .A2(new_n2513_), .A3(new_n2521_), .ZN(new_n3656_));
  OAI21_X1   g02654(.A1(new_n2531_), .A2(new_n3656_), .B(new_n2533_), .ZN(new_n3657_));
  NOR2_X1    g02655(.A1(new_n3650_), .A2(new_n3653_), .ZN(new_n3658_));
  NOR2_X1    g02656(.A1(new_n3632_), .A2(new_n3645_), .ZN(new_n3659_));
  NOR3_X1    g02657(.A1(new_n3659_), .A2(new_n3657_), .A3(new_n3658_), .ZN(new_n3660_));
  NOR2_X1    g02658(.A1(new_n3660_), .A2(new_n3655_), .ZN(new_n3661_));
  NAND2_X1   g02659(.A1(new_n3613_), .A2(new_n3661_), .ZN(new_n3662_));
  AOI21_X1   g02660(.A1(new_n3611_), .A2(new_n3610_), .B(new_n3609_), .ZN(new_n3663_));
  NOR3_X1    g02661(.A1(new_n3566_), .A2(new_n3598_), .A3(new_n3607_), .ZN(new_n3664_));
  NOR2_X1    g02662(.A1(new_n3664_), .A2(new_n3663_), .ZN(new_n3665_));
  OAI21_X1   g02663(.A1(new_n3659_), .A2(new_n3658_), .B(new_n3657_), .ZN(new_n3666_));
  NAND3_X1   g02664(.A1(new_n3646_), .A2(new_n3654_), .A3(new_n3615_), .ZN(new_n3667_));
  NAND2_X1   g02665(.A1(new_n3666_), .A2(new_n3667_), .ZN(new_n3668_));
  NAND2_X1   g02666(.A1(new_n3665_), .A2(new_n3668_), .ZN(new_n3669_));
  AOI21_X1   g02667(.A1(new_n3669_), .A2(new_n3662_), .B(new_n3564_), .ZN(new_n3670_));
  NOR2_X1    g02668(.A1(new_n3665_), .A2(new_n3668_), .ZN(new_n3671_));
  NOR2_X1    g02669(.A1(new_n3613_), .A2(new_n3661_), .ZN(new_n3672_));
  NOR3_X1    g02670(.A1(new_n3671_), .A2(new_n3672_), .A3(new_n3563_), .ZN(new_n3673_));
  NOR2_X1    g02671(.A1(new_n3670_), .A2(new_n3673_), .ZN(new_n3674_));
  AOI22_X1   g02672(.A1(new_n3018_), .A2(new_n3014_), .B1(new_n3012_), .B2(new_n3015_), .ZN(new_n3675_));
  NAND3_X1   g02673(.A1(new_n2998_), .A2(new_n2995_), .A3(new_n2999_), .ZN(new_n3676_));
  AOI21_X1   g02674(.A1(new_n2877_), .A2(new_n3676_), .B(new_n3000_), .ZN(new_n3677_));
  AOI21_X1   g02675(.A1(new_n2768_), .A2(new_n2029_), .B(new_n2863_), .ZN(new_n3678_));
  OAI21_X1   g02676(.A1(new_n2753_), .A2(new_n2053_), .B(new_n2748_), .ZN(new_n3679_));
  NOR2_X1    g02677(.A1(new_n3678_), .A2(new_n3679_), .ZN(new_n3680_));
  OAI21_X1   g02678(.A1(new_n2789_), .A2(new_n2775_), .B(new_n2793_), .ZN(new_n3681_));
  AOI21_X1   g02679(.A1(new_n2784_), .A2(new_n2057_), .B(new_n2781_), .ZN(new_n3682_));
  NOR2_X1    g02680(.A1(new_n3681_), .A2(new_n3682_), .ZN(new_n3683_));
  AOI21_X1   g02681(.A1(new_n2777_), .A2(new_n2769_), .B(new_n2785_), .ZN(new_n3684_));
  OAI22_X1   g02682(.A1(new_n3684_), .A2(new_n2871_), .B1(new_n3680_), .B2(new_n3683_), .ZN(new_n3685_));
  NAND2_X1   g02683(.A1(new_n3681_), .A2(new_n3682_), .ZN(new_n3686_));
  NAND2_X1   g02684(.A1(new_n3678_), .A2(new_n3679_), .ZN(new_n3687_));
  AOI21_X1   g02685(.A1(new_n2793_), .A2(new_n2029_), .B(new_n2789_), .ZN(new_n3688_));
  OAI21_X1   g02686(.A1(new_n3688_), .A2(new_n2776_), .B(new_n2754_), .ZN(new_n3689_));
  NAND4_X1   g02687(.A1(new_n3689_), .A2(new_n3686_), .A3(new_n3687_), .A4(new_n2795_), .ZN(new_n3690_));
  NAND2_X1   g02688(.A1(new_n3690_), .A2(new_n3685_), .ZN(new_n3691_));
  OAI21_X1   g02689(.A1(new_n2821_), .A2(new_n1953_), .B(new_n2834_), .ZN(new_n3692_));
  AOI21_X1   g02690(.A1(new_n2813_), .A2(new_n1982_), .B(new_n2808_), .ZN(new_n3693_));
  NAND2_X1   g02691(.A1(new_n3693_), .A2(new_n3692_), .ZN(new_n3694_));
  AOI21_X1   g02692(.A1(new_n2830_), .A2(new_n1992_), .B(new_n2825_), .ZN(new_n3695_));
  OAI21_X1   g02693(.A1(new_n2843_), .A2(new_n1995_), .B(new_n2840_), .ZN(new_n3696_));
  NAND2_X1   g02694(.A1(new_n3696_), .A2(new_n3695_), .ZN(new_n3697_));
  NAND2_X1   g02695(.A1(new_n2827_), .A2(new_n2844_), .ZN(new_n3698_));
  AOI22_X1   g02696(.A1(new_n3698_), .A2(new_n2836_), .B1(new_n3694_), .B2(new_n3697_), .ZN(new_n3699_));
  NOR2_X1    g02697(.A1(new_n3696_), .A2(new_n3695_), .ZN(new_n3700_));
  NOR2_X1    g02698(.A1(new_n3693_), .A2(new_n3692_), .ZN(new_n3701_));
  OAI21_X1   g02699(.A1(new_n2825_), .A2(new_n1953_), .B(new_n2830_), .ZN(new_n3702_));
  AOI21_X1   g02700(.A1(new_n3702_), .A2(new_n2822_), .B(new_n2814_), .ZN(new_n3703_));
  NOR4_X1    g02701(.A1(new_n3703_), .A2(new_n3701_), .A3(new_n2855_), .A4(new_n3700_), .ZN(new_n3704_));
  NOR2_X1    g02702(.A1(new_n3704_), .A2(new_n3699_), .ZN(new_n3705_));
  NAND2_X1   g02703(.A1(new_n3691_), .A2(new_n3705_), .ZN(new_n3706_));
  AOI22_X1   g02704(.A1(new_n3689_), .A2(new_n2795_), .B1(new_n3686_), .B2(new_n3687_), .ZN(new_n3707_));
  NOR4_X1    g02705(.A1(new_n3684_), .A2(new_n3680_), .A3(new_n3683_), .A4(new_n2871_), .ZN(new_n3708_));
  NOR2_X1    g02706(.A1(new_n3707_), .A2(new_n3708_), .ZN(new_n3709_));
  OAI22_X1   g02707(.A1(new_n3703_), .A2(new_n2855_), .B1(new_n3701_), .B2(new_n3700_), .ZN(new_n3710_));
  NAND4_X1   g02708(.A1(new_n3698_), .A2(new_n3694_), .A3(new_n3697_), .A4(new_n2836_), .ZN(new_n3711_));
  NAND2_X1   g02709(.A1(new_n3710_), .A2(new_n3711_), .ZN(new_n3712_));
  NAND2_X1   g02710(.A1(new_n3709_), .A2(new_n3712_), .ZN(new_n3713_));
  AOI21_X1   g02711(.A1(new_n2873_), .A2(new_n3005_), .B(new_n2875_), .ZN(new_n3714_));
  NAND3_X1   g02712(.A1(new_n3706_), .A2(new_n3713_), .A3(new_n3714_), .ZN(new_n3715_));
  NOR2_X1    g02713(.A1(new_n3709_), .A2(new_n3712_), .ZN(new_n3716_));
  NOR2_X1    g02714(.A1(new_n3691_), .A2(new_n3705_), .ZN(new_n3717_));
  OAI21_X1   g02715(.A1(new_n2797_), .A2(new_n2874_), .B(new_n3006_), .ZN(new_n3718_));
  OAI21_X1   g02716(.A1(new_n3717_), .A2(new_n3716_), .B(new_n3718_), .ZN(new_n3719_));
  NAND2_X1   g02717(.A1(new_n3719_), .A2(new_n3715_), .ZN(new_n3720_));
  AOI21_X1   g02718(.A1(new_n2987_), .A2(new_n2965_), .B(new_n2994_), .ZN(new_n3721_));
  AOI21_X1   g02719(.A1(new_n2896_), .A2(new_n1897_), .B(new_n2909_), .ZN(new_n3722_));
  OAI21_X1   g02720(.A1(new_n2888_), .A2(new_n1909_), .B(new_n2883_), .ZN(new_n3723_));
  NOR2_X1    g02721(.A1(new_n3723_), .A2(new_n3722_), .ZN(new_n3724_));
  OAI21_X1   g02722(.A1(new_n2906_), .A2(new_n1852_), .B(new_n2901_), .ZN(new_n3725_));
  NAND3_X1   g02723(.A1(new_n1882_), .A2(new_n2885_), .A3(new_n2886_), .ZN(new_n3726_));
  OAI21_X1   g02724(.A1(new_n2878_), .A2(new_n2879_), .B(new_n1905_), .ZN(new_n3727_));
  NAND2_X1   g02725(.A1(new_n3727_), .A2(new_n3726_), .ZN(new_n3728_));
  AOI21_X1   g02726(.A1(new_n3728_), .A2(new_n1884_), .B(new_n2914_), .ZN(new_n3729_));
  NOR2_X1    g02727(.A1(new_n3725_), .A2(new_n3729_), .ZN(new_n3730_));
  OAI21_X1   g02728(.A1(new_n2909_), .A2(new_n1852_), .B(new_n2896_), .ZN(new_n3731_));
  AOI21_X1   g02729(.A1(new_n3731_), .A2(new_n2897_), .B(new_n2915_), .ZN(new_n3732_));
  OAI22_X1   g02730(.A1(new_n3732_), .A2(new_n2984_), .B1(new_n3730_), .B2(new_n3724_), .ZN(new_n3733_));
  NAND2_X1   g02731(.A1(new_n3725_), .A2(new_n3729_), .ZN(new_n3734_));
  NAND2_X1   g02732(.A1(new_n3723_), .A2(new_n3722_), .ZN(new_n3735_));
  NAND2_X1   g02733(.A1(new_n2919_), .A2(new_n2889_), .ZN(new_n3736_));
  NAND4_X1   g02734(.A1(new_n3736_), .A2(new_n3734_), .A3(new_n3735_), .A4(new_n2918_), .ZN(new_n3737_));
  NAND2_X1   g02735(.A1(new_n3737_), .A2(new_n3733_), .ZN(new_n3738_));
  NOR3_X1    g02736(.A1(new_n2936_), .A2(new_n1750_), .A3(new_n2937_), .ZN(new_n3739_));
  AOI21_X1   g02737(.A1(new_n2933_), .A2(new_n2934_), .B(new_n1808_), .ZN(new_n3740_));
  NOR2_X1    g02738(.A1(new_n3740_), .A2(new_n3739_), .ZN(new_n3741_));
  OAI21_X1   g02739(.A1(new_n3741_), .A2(new_n1757_), .B(new_n2950_), .ZN(new_n3742_));
  NAND2_X1   g02740(.A1(new_n2931_), .A2(new_n2930_), .ZN(new_n3743_));
  AOI21_X1   g02741(.A1(new_n3743_), .A2(new_n1798_), .B(new_n2955_), .ZN(new_n3744_));
  NAND2_X1   g02742(.A1(new_n3742_), .A2(new_n3744_), .ZN(new_n3745_));
  AOI21_X1   g02743(.A1(new_n2939_), .A2(new_n1814_), .B(new_n2967_), .ZN(new_n3746_));
  NOR2_X1    g02744(.A1(new_n2956_), .A2(new_n2957_), .ZN(new_n3747_));
  OAI21_X1   g02745(.A1(new_n3747_), .A2(new_n1821_), .B(new_n2927_), .ZN(new_n3748_));
  NAND2_X1   g02746(.A1(new_n3748_), .A2(new_n3746_), .ZN(new_n3749_));
  OAI21_X1   g02747(.A1(new_n2947_), .A2(new_n2951_), .B(new_n2932_), .ZN(new_n3750_));
  AOI22_X1   g02748(.A1(new_n3750_), .A2(new_n2969_), .B1(new_n3745_), .B2(new_n3749_), .ZN(new_n3751_));
  NOR2_X1    g02749(.A1(new_n3748_), .A2(new_n3746_), .ZN(new_n3752_));
  NOR2_X1    g02750(.A1(new_n3742_), .A2(new_n3744_), .ZN(new_n3753_));
  AOI21_X1   g02751(.A1(new_n2961_), .A2(new_n2959_), .B(new_n2958_), .ZN(new_n3754_));
  NOR4_X1    g02752(.A1(new_n3754_), .A2(new_n3752_), .A3(new_n3753_), .A4(new_n2946_), .ZN(new_n3755_));
  NOR2_X1    g02753(.A1(new_n3751_), .A2(new_n3755_), .ZN(new_n3756_));
  NAND2_X1   g02754(.A1(new_n3738_), .A2(new_n3756_), .ZN(new_n3757_));
  AOI22_X1   g02755(.A1(new_n3736_), .A2(new_n2918_), .B1(new_n3735_), .B2(new_n3734_), .ZN(new_n3758_));
  NOR4_X1    g02756(.A1(new_n3732_), .A2(new_n3724_), .A3(new_n3730_), .A4(new_n2984_), .ZN(new_n3759_));
  NOR2_X1    g02757(.A1(new_n3758_), .A2(new_n3759_), .ZN(new_n3760_));
  OAI22_X1   g02758(.A1(new_n2946_), .A2(new_n3754_), .B1(new_n3752_), .B2(new_n3753_), .ZN(new_n3761_));
  NAND4_X1   g02759(.A1(new_n3750_), .A2(new_n3745_), .A3(new_n3749_), .A4(new_n2969_), .ZN(new_n3762_));
  NAND2_X1   g02760(.A1(new_n3761_), .A2(new_n3762_), .ZN(new_n3763_));
  NAND2_X1   g02761(.A1(new_n3760_), .A2(new_n3763_), .ZN(new_n3764_));
  AOI21_X1   g02762(.A1(new_n3757_), .A2(new_n3764_), .B(new_n3721_), .ZN(new_n3765_));
  OAI21_X1   g02763(.A1(new_n2921_), .A2(new_n2993_), .B(new_n2976_), .ZN(new_n3766_));
  NOR2_X1    g02764(.A1(new_n3760_), .A2(new_n3763_), .ZN(new_n3767_));
  NOR2_X1    g02765(.A1(new_n3738_), .A2(new_n3756_), .ZN(new_n3768_));
  NOR3_X1    g02766(.A1(new_n3768_), .A2(new_n3767_), .A3(new_n3766_), .ZN(new_n3769_));
  NOR2_X1    g02767(.A1(new_n3769_), .A2(new_n3765_), .ZN(new_n3770_));
  NAND2_X1   g02768(.A1(new_n3720_), .A2(new_n3770_), .ZN(new_n3771_));
  OAI21_X1   g02769(.A1(new_n3768_), .A2(new_n3767_), .B(new_n3766_), .ZN(new_n3772_));
  NAND3_X1   g02770(.A1(new_n3757_), .A2(new_n3764_), .A3(new_n3721_), .ZN(new_n3773_));
  NAND2_X1   g02771(.A1(new_n3772_), .A2(new_n3773_), .ZN(new_n3774_));
  NAND3_X1   g02772(.A1(new_n3774_), .A2(new_n3715_), .A3(new_n3719_), .ZN(new_n3775_));
  AOI21_X1   g02773(.A1(new_n3771_), .A2(new_n3775_), .B(new_n3677_), .ZN(new_n3776_));
  NOR2_X1    g02774(.A1(new_n2990_), .A2(new_n2977_), .ZN(new_n3777_));
  OAI22_X1   g02775(.A1(new_n2992_), .A2(new_n3008_), .B1(new_n3777_), .B2(new_n2999_), .ZN(new_n3778_));
  NOR3_X1    g02776(.A1(new_n3717_), .A2(new_n3716_), .A3(new_n3718_), .ZN(new_n3779_));
  AOI21_X1   g02777(.A1(new_n3706_), .A2(new_n3713_), .B(new_n3714_), .ZN(new_n3780_));
  NOR2_X1    g02778(.A1(new_n3780_), .A2(new_n3779_), .ZN(new_n3781_));
  NOR2_X1    g02779(.A1(new_n3781_), .A2(new_n3774_), .ZN(new_n3782_));
  NOR2_X1    g02780(.A1(new_n3720_), .A2(new_n3770_), .ZN(new_n3783_));
  NOR3_X1    g02781(.A1(new_n3783_), .A2(new_n3782_), .A3(new_n3778_), .ZN(new_n3784_));
  NAND2_X1   g02782(.A1(new_n2725_), .A2(new_n2728_), .ZN(new_n3785_));
  AOI22_X1   g02783(.A1(new_n2732_), .A2(new_n2599_), .B1(new_n3785_), .B2(new_n2722_), .ZN(new_n3786_));
  NOR2_X1    g02784(.A1(new_n2588_), .A2(new_n2582_), .ZN(new_n3787_));
  AOI21_X1   g02785(.A1(new_n3787_), .A2(new_n2590_), .B(new_n2594_), .ZN(new_n3788_));
  OAI21_X1   g02786(.A1(new_n2552_), .A2(new_n2545_), .B(new_n2551_), .ZN(new_n3789_));
  OAI21_X1   g02787(.A1(new_n2559_), .A2(new_n2563_), .B(new_n2571_), .ZN(new_n3790_));
  NAND2_X1   g02788(.A1(new_n2581_), .A2(new_n2583_), .ZN(new_n3791_));
  AOI21_X1   g02789(.A1(new_n3791_), .A2(new_n2577_), .B(new_n3790_), .ZN(new_n3792_));
  AOI21_X1   g02790(.A1(new_n2560_), .A2(new_n2567_), .B(new_n2579_), .ZN(new_n3793_));
  NOR2_X1    g02791(.A1(new_n2585_), .A2(new_n2556_), .ZN(new_n3794_));
  NOR3_X1    g02792(.A1(new_n3794_), .A2(new_n2584_), .A3(new_n3793_), .ZN(new_n3795_));
  OAI21_X1   g02793(.A1(new_n3795_), .A2(new_n3792_), .B(new_n3789_), .ZN(new_n3796_));
  AOI21_X1   g02794(.A1(new_n2593_), .A2(new_n2546_), .B(new_n2550_), .ZN(new_n3797_));
  OAI21_X1   g02795(.A1(new_n3794_), .A2(new_n2584_), .B(new_n3793_), .ZN(new_n3798_));
  NAND3_X1   g02796(.A1(new_n3791_), .A2(new_n2577_), .A3(new_n3790_), .ZN(new_n3799_));
  NAND3_X1   g02797(.A1(new_n3798_), .A2(new_n3799_), .A3(new_n3797_), .ZN(new_n3800_));
  NAND3_X1   g02798(.A1(new_n3796_), .A2(new_n3800_), .A3(new_n2595_), .ZN(new_n3801_));
  AOI21_X1   g02799(.A1(new_n2589_), .A2(new_n2590_), .B(new_n2554_), .ZN(new_n3802_));
  NOR2_X1    g02800(.A1(new_n3788_), .A2(new_n3802_), .ZN(new_n3803_));
  NAND2_X1   g02801(.A1(new_n3798_), .A2(new_n3799_), .ZN(new_n3804_));
  NOR2_X1    g02802(.A1(new_n3795_), .A2(new_n3789_), .ZN(new_n3805_));
  AOI22_X1   g02803(.A1(new_n3804_), .A2(new_n3789_), .B1(new_n3805_), .B2(new_n3798_), .ZN(new_n3806_));
  OAI22_X1   g02804(.A1(new_n3806_), .A2(new_n3803_), .B1(new_n3801_), .B2(new_n3788_), .ZN(new_n3807_));
  AOI21_X1   g02805(.A1(new_n2642_), .A2(new_n2274_), .B(new_n2625_), .ZN(new_n3808_));
  NOR3_X1    g02806(.A1(new_n2605_), .A2(new_n2610_), .A3(new_n2611_), .ZN(new_n3809_));
  AOI22_X1   g02807(.A1(new_n2602_), .A2(new_n2604_), .B1(new_n2296_), .B2(new_n2298_), .ZN(new_n3810_));
  NOR2_X1    g02808(.A1(new_n3810_), .A2(new_n3809_), .ZN(new_n3811_));
  OAI21_X1   g02809(.A1(new_n3811_), .A2(new_n2312_), .B(new_n2640_), .ZN(new_n3812_));
  NOR2_X1    g02810(.A1(new_n3812_), .A2(new_n3808_), .ZN(new_n3813_));
  OAI21_X1   g02811(.A1(new_n2621_), .A2(new_n2319_), .B(new_n2632_), .ZN(new_n3814_));
  AOI21_X1   g02812(.A1(new_n2613_), .A2(new_n2323_), .B(new_n2608_), .ZN(new_n3815_));
  NOR2_X1    g02813(.A1(new_n3815_), .A2(new_n3814_), .ZN(new_n3816_));
  AOI21_X1   g02814(.A1(new_n2710_), .A2(new_n2629_), .B(new_n2614_), .ZN(new_n3817_));
  OAI22_X1   g02815(.A1(new_n3817_), .A2(new_n2645_), .B1(new_n3816_), .B2(new_n3813_), .ZN(new_n3818_));
  NAND2_X1   g02816(.A1(new_n3815_), .A2(new_n3814_), .ZN(new_n3819_));
  NAND2_X1   g02817(.A1(new_n3812_), .A2(new_n3808_), .ZN(new_n3820_));
  OAI21_X1   g02818(.A1(new_n2622_), .A2(new_n2635_), .B(new_n2641_), .ZN(new_n3821_));
  NAND4_X1   g02819(.A1(new_n3821_), .A2(new_n3819_), .A3(new_n3820_), .A4(new_n2714_), .ZN(new_n3822_));
  NAND2_X1   g02820(.A1(new_n3818_), .A2(new_n3822_), .ZN(new_n3823_));
  OAI21_X1   g02821(.A1(new_n2684_), .A2(new_n2174_), .B(new_n2695_), .ZN(new_n3824_));
  NAND2_X1   g02822(.A1(new_n2658_), .A2(new_n2657_), .ZN(new_n3825_));
  AOI21_X1   g02823(.A1(new_n3825_), .A2(new_n2214_), .B(new_n2678_), .ZN(new_n3826_));
  NAND2_X1   g02824(.A1(new_n3824_), .A2(new_n3826_), .ZN(new_n3827_));
  NAND2_X1   g02825(.A1(new_n2660_), .A2(new_n2661_), .ZN(new_n3828_));
  AOI21_X1   g02826(.A1(new_n3828_), .A2(new_n2223_), .B(new_n2668_), .ZN(new_n3829_));
  AOI21_X1   g02827(.A1(new_n2666_), .A2(new_n2227_), .B(new_n3829_), .ZN(new_n3830_));
  NOR2_X1    g02828(.A1(new_n2679_), .A2(new_n2680_), .ZN(new_n3831_));
  OAI21_X1   g02829(.A1(new_n3831_), .A2(new_n2234_), .B(new_n2654_), .ZN(new_n3832_));
  NAND2_X1   g02830(.A1(new_n3832_), .A2(new_n3830_), .ZN(new_n3833_));
  NOR2_X1    g02831(.A1(new_n2687_), .A2(new_n2684_), .ZN(new_n3834_));
  OAI21_X1   g02832(.A1(new_n2674_), .A2(new_n3834_), .B(new_n2659_), .ZN(new_n3835_));
  AOI22_X1   g02833(.A1(new_n3835_), .A2(new_n2697_), .B1(new_n3827_), .B2(new_n3833_), .ZN(new_n3836_));
  NOR2_X1    g02834(.A1(new_n3832_), .A2(new_n3830_), .ZN(new_n3837_));
  NOR2_X1    g02835(.A1(new_n3824_), .A2(new_n3826_), .ZN(new_n3838_));
  AOI21_X1   g02836(.A1(new_n2689_), .A2(new_n2698_), .B(new_n2681_), .ZN(new_n3839_));
  NOR4_X1    g02837(.A1(new_n3839_), .A2(new_n3837_), .A3(new_n3838_), .A4(new_n2672_), .ZN(new_n3840_));
  NOR2_X1    g02838(.A1(new_n3836_), .A2(new_n3840_), .ZN(new_n3841_));
  NOR2_X1    g02839(.A1(new_n3823_), .A2(new_n3841_), .ZN(new_n3842_));
  AOI22_X1   g02840(.A1(new_n3821_), .A2(new_n2714_), .B1(new_n3819_), .B2(new_n3820_), .ZN(new_n3843_));
  NOR4_X1    g02841(.A1(new_n3817_), .A2(new_n2645_), .A3(new_n3813_), .A4(new_n3816_), .ZN(new_n3844_));
  NOR2_X1    g02842(.A1(new_n3844_), .A2(new_n3843_), .ZN(new_n3845_));
  OAI22_X1   g02843(.A1(new_n2672_), .A2(new_n3839_), .B1(new_n3837_), .B2(new_n3838_), .ZN(new_n3846_));
  NAND4_X1   g02844(.A1(new_n3835_), .A2(new_n3827_), .A3(new_n3833_), .A4(new_n2697_), .ZN(new_n3847_));
  NAND2_X1   g02845(.A1(new_n3846_), .A2(new_n3847_), .ZN(new_n3848_));
  NOR2_X1    g02846(.A1(new_n3845_), .A2(new_n3848_), .ZN(new_n3849_));
  OAI21_X1   g02847(.A1(new_n2717_), .A2(new_n2726_), .B(new_n2719_), .ZN(new_n3850_));
  OAI21_X1   g02848(.A1(new_n3842_), .A2(new_n3849_), .B(new_n3850_), .ZN(new_n3851_));
  NAND2_X1   g02849(.A1(new_n3845_), .A2(new_n3848_), .ZN(new_n3852_));
  NAND2_X1   g02850(.A1(new_n3823_), .A2(new_n3841_), .ZN(new_n3853_));
  AOI21_X1   g02851(.A1(new_n2648_), .A2(new_n2718_), .B(new_n2727_), .ZN(new_n3854_));
  NAND3_X1   g02852(.A1(new_n3853_), .A2(new_n3852_), .A3(new_n3854_), .ZN(new_n3855_));
  NAND3_X1   g02853(.A1(new_n3851_), .A2(new_n3855_), .A3(new_n3807_), .ZN(new_n3856_));
  NOR2_X1    g02854(.A1(new_n3801_), .A2(new_n3788_), .ZN(new_n3857_));
  NOR2_X1    g02855(.A1(new_n3806_), .A2(new_n3803_), .ZN(new_n3858_));
  NOR2_X1    g02856(.A1(new_n3858_), .A2(new_n3857_), .ZN(new_n3859_));
  AOI21_X1   g02857(.A1(new_n3853_), .A2(new_n3852_), .B(new_n3854_), .ZN(new_n3860_));
  NOR3_X1    g02858(.A1(new_n3842_), .A2(new_n3849_), .A3(new_n3850_), .ZN(new_n3861_));
  OAI21_X1   g02859(.A1(new_n3860_), .A2(new_n3861_), .B(new_n3859_), .ZN(new_n3862_));
  AOI21_X1   g02860(.A1(new_n3862_), .A2(new_n3856_), .B(new_n3786_), .ZN(new_n3863_));
  NOR3_X1    g02861(.A1(new_n2722_), .A2(new_n2720_), .A3(new_n2708_), .ZN(new_n3864_));
  OAI21_X1   g02862(.A1(new_n2598_), .A2(new_n3864_), .B(new_n2731_), .ZN(new_n3865_));
  NOR3_X1    g02863(.A1(new_n3860_), .A2(new_n3861_), .A3(new_n3859_), .ZN(new_n3866_));
  AOI21_X1   g02864(.A1(new_n3851_), .A2(new_n3855_), .B(new_n3807_), .ZN(new_n3867_));
  NOR3_X1    g02865(.A1(new_n3866_), .A2(new_n3867_), .A3(new_n3865_), .ZN(new_n3868_));
  NOR2_X1    g02866(.A1(new_n3868_), .A2(new_n3863_), .ZN(new_n3869_));
  OAI21_X1   g02867(.A1(new_n3776_), .A2(new_n3784_), .B(new_n3869_), .ZN(new_n3870_));
  OAI21_X1   g02868(.A1(new_n3783_), .A2(new_n3782_), .B(new_n3778_), .ZN(new_n3871_));
  NAND3_X1   g02869(.A1(new_n3771_), .A2(new_n3775_), .A3(new_n3677_), .ZN(new_n3872_));
  OAI21_X1   g02870(.A1(new_n3866_), .A2(new_n3867_), .B(new_n3865_), .ZN(new_n3873_));
  NAND3_X1   g02871(.A1(new_n3862_), .A2(new_n3856_), .A3(new_n3786_), .ZN(new_n3874_));
  NAND2_X1   g02872(.A1(new_n3873_), .A2(new_n3874_), .ZN(new_n3875_));
  NAND3_X1   g02873(.A1(new_n3875_), .A2(new_n3871_), .A3(new_n3872_), .ZN(new_n3876_));
  AOI21_X1   g02874(.A1(new_n3870_), .A2(new_n3876_), .B(new_n3675_), .ZN(new_n3877_));
  INV_X1     g02875(.I(new_n3001_), .ZN(new_n3878_));
  INV_X1     g02876(.I(new_n3011_), .ZN(new_n3879_));
  NOR3_X1    g02877(.A1(new_n3879_), .A2(new_n3878_), .A3(new_n3012_), .ZN(new_n3880_));
  OAI21_X1   g02878(.A1(new_n2734_), .A2(new_n3880_), .B(new_n3016_), .ZN(new_n3881_));
  AOI21_X1   g02879(.A1(new_n3871_), .A2(new_n3872_), .B(new_n3875_), .ZN(new_n3882_));
  NOR3_X1    g02880(.A1(new_n3869_), .A2(new_n3784_), .A3(new_n3776_), .ZN(new_n3883_));
  NOR3_X1    g02881(.A1(new_n3882_), .A2(new_n3883_), .A3(new_n3881_), .ZN(new_n3884_));
  OAI21_X1   g02882(.A1(new_n3877_), .A2(new_n3884_), .B(new_n3674_), .ZN(new_n3885_));
  OAI21_X1   g02883(.A1(new_n3671_), .A2(new_n3672_), .B(new_n3563_), .ZN(new_n3886_));
  NAND3_X1   g02884(.A1(new_n3564_), .A2(new_n3669_), .A3(new_n3662_), .ZN(new_n3887_));
  NAND2_X1   g02885(.A1(new_n3887_), .A2(new_n3886_), .ZN(new_n3888_));
  OAI21_X1   g02886(.A1(new_n3882_), .A2(new_n3883_), .B(new_n3881_), .ZN(new_n3889_));
  NAND3_X1   g02887(.A1(new_n3870_), .A2(new_n3876_), .A3(new_n3675_), .ZN(new_n3890_));
  NAND3_X1   g02888(.A1(new_n3889_), .A2(new_n3890_), .A3(new_n3888_), .ZN(new_n3891_));
  OAI21_X1   g02889(.A1(new_n2544_), .A2(new_n3028_), .B(new_n3029_), .ZN(new_n3892_));
  INV_X1     g02890(.I(new_n3892_), .ZN(new_n3893_));
  NAND3_X1   g02891(.A1(new_n3893_), .A2(new_n3885_), .A3(new_n3891_), .ZN(new_n3894_));
  AOI21_X1   g02892(.A1(new_n3889_), .A2(new_n3890_), .B(new_n3888_), .ZN(new_n3895_));
  NOR3_X1    g02893(.A1(new_n3877_), .A2(new_n3884_), .A3(new_n3674_), .ZN(new_n3896_));
  OAI21_X1   g02894(.A1(new_n3896_), .A2(new_n3895_), .B(new_n3892_), .ZN(new_n3897_));
  INV_X1     g02895(.I(new_n3558_), .ZN(new_n3898_));
  OAI21_X1   g02896(.A1(new_n3290_), .A2(new_n3557_), .B(new_n3898_), .ZN(new_n3899_));
  AOI22_X1   g02897(.A1(new_n3150_), .A2(new_n3287_), .B1(new_n3284_), .B2(new_n3282_), .ZN(new_n3900_));
  OAI22_X1   g02898(.A1(new_n3075_), .A2(new_n3140_), .B1(new_n3123_), .B2(new_n3128_), .ZN(new_n3901_));
  OAI21_X1   g02899(.A1(new_n3072_), .A2(new_n3055_), .B(new_n3067_), .ZN(new_n3902_));
  NAND2_X1   g02900(.A1(new_n3043_), .A2(new_n1517_), .ZN(new_n3903_));
  NAND2_X1   g02901(.A1(new_n3044_), .A2(new_n3042_), .ZN(new_n3904_));
  AOI22_X1   g02902(.A1(new_n3904_), .A2(new_n1507_), .B1(new_n3903_), .B2(new_n3038_), .ZN(new_n3905_));
  NAND2_X1   g02903(.A1(new_n3902_), .A2(new_n3905_), .ZN(new_n3906_));
  AOI21_X1   g02904(.A1(new_n3052_), .A2(new_n1476_), .B(new_n3054_), .ZN(new_n3907_));
  XOR2_X1    g02905(.A1(new_n3034_), .A2(new_n1517_), .Z(new_n3908_));
  OAI21_X1   g02906(.A1(new_n3908_), .A2(new_n3056_), .B(new_n3039_), .ZN(new_n3909_));
  NAND2_X1   g02907(.A1(new_n3909_), .A2(new_n3907_), .ZN(new_n3910_));
  OAI21_X1   g02908(.A1(new_n3073_), .A2(new_n3062_), .B(new_n3045_), .ZN(new_n3911_));
  AOI22_X1   g02909(.A1(new_n3910_), .A2(new_n3906_), .B1(new_n3911_), .B2(new_n3061_), .ZN(new_n3912_));
  NOR2_X1    g02910(.A1(new_n3909_), .A2(new_n3907_), .ZN(new_n3913_));
  NOR2_X1    g02911(.A1(new_n3902_), .A2(new_n3905_), .ZN(new_n3914_));
  AOI21_X1   g02912(.A1(new_n3063_), .A2(new_n3069_), .B(new_n3046_), .ZN(new_n3915_));
  NOR4_X1    g02913(.A1(new_n3915_), .A2(new_n3913_), .A3(new_n3914_), .A4(new_n3133_), .ZN(new_n3916_));
  NOR2_X1    g02914(.A1(new_n3916_), .A2(new_n3912_), .ZN(new_n3917_));
  AOI21_X1   g02915(.A1(new_n3100_), .A2(new_n1413_), .B(new_n3102_), .ZN(new_n3918_));
  INV_X1     g02916(.I(new_n3085_), .ZN(new_n3919_));
  NOR2_X1    g02917(.A1(new_n3089_), .A2(new_n3090_), .ZN(new_n3920_));
  OAI21_X1   g02918(.A1(new_n3920_), .A2(new_n3078_), .B(new_n3919_), .ZN(new_n3921_));
  NOR2_X1    g02919(.A1(new_n3921_), .A2(new_n3918_), .ZN(new_n3922_));
  INV_X1     g02920(.I(new_n3102_), .ZN(new_n3923_));
  OAI21_X1   g02921(.A1(new_n3119_), .A2(new_n3103_), .B(new_n3923_), .ZN(new_n3924_));
  XOR2_X1    g02922(.A1(new_n3083_), .A2(new_n1454_), .Z(new_n3925_));
  AOI21_X1   g02923(.A1(new_n3925_), .A2(new_n1444_), .B(new_n3085_), .ZN(new_n3926_));
  NOR2_X1    g02924(.A1(new_n3926_), .A2(new_n3924_), .ZN(new_n3927_));
  AOI21_X1   g02925(.A1(new_n3110_), .A2(new_n3109_), .B(new_n3091_), .ZN(new_n3928_));
  OAI22_X1   g02926(.A1(new_n3142_), .A2(new_n3928_), .B1(new_n3927_), .B2(new_n3922_), .ZN(new_n3929_));
  NAND2_X1   g02927(.A1(new_n3926_), .A2(new_n3924_), .ZN(new_n3930_));
  NAND2_X1   g02928(.A1(new_n3921_), .A2(new_n3918_), .ZN(new_n3931_));
  OAI21_X1   g02929(.A1(new_n3115_), .A2(new_n3120_), .B(new_n3113_), .ZN(new_n3932_));
  NAND4_X1   g02930(.A1(new_n3932_), .A2(new_n3108_), .A3(new_n3930_), .A4(new_n3931_), .ZN(new_n3933_));
  NAND2_X1   g02931(.A1(new_n3929_), .A2(new_n3933_), .ZN(new_n3934_));
  NOR2_X1    g02932(.A1(new_n3917_), .A2(new_n3934_), .ZN(new_n3935_));
  OAI22_X1   g02933(.A1(new_n3915_), .A2(new_n3133_), .B1(new_n3913_), .B2(new_n3914_), .ZN(new_n3936_));
  NAND4_X1   g02934(.A1(new_n3910_), .A2(new_n3906_), .A3(new_n3911_), .A4(new_n3061_), .ZN(new_n3937_));
  NAND2_X1   g02935(.A1(new_n3936_), .A2(new_n3937_), .ZN(new_n3938_));
  AOI22_X1   g02936(.A1(new_n3932_), .A2(new_n3108_), .B1(new_n3930_), .B2(new_n3931_), .ZN(new_n3939_));
  NOR4_X1    g02937(.A1(new_n3928_), .A2(new_n3927_), .A3(new_n3142_), .A4(new_n3922_), .ZN(new_n3940_));
  NOR2_X1    g02938(.A1(new_n3939_), .A2(new_n3940_), .ZN(new_n3941_));
  NOR2_X1    g02939(.A1(new_n3938_), .A2(new_n3941_), .ZN(new_n3942_));
  OAI21_X1   g02940(.A1(new_n3935_), .A2(new_n3942_), .B(new_n3901_), .ZN(new_n3943_));
  NAND3_X1   g02941(.A1(new_n3144_), .A2(new_n3147_), .A3(new_n3123_), .ZN(new_n3944_));
  AOI21_X1   g02942(.A1(new_n3139_), .A2(new_n3944_), .B(new_n3148_), .ZN(new_n3945_));
  NAND2_X1   g02943(.A1(new_n3938_), .A2(new_n3941_), .ZN(new_n3946_));
  NAND2_X1   g02944(.A1(new_n3917_), .A2(new_n3934_), .ZN(new_n3947_));
  NAND3_X1   g02945(.A1(new_n3947_), .A2(new_n3946_), .A3(new_n3945_), .ZN(new_n3948_));
  NAND2_X1   g02946(.A1(new_n3943_), .A2(new_n3948_), .ZN(new_n3949_));
  NAND2_X1   g02947(.A1(new_n3241_), .A2(new_n3236_), .ZN(new_n3950_));
  NOR2_X1    g02948(.A1(new_n3239_), .A2(new_n3240_), .ZN(new_n3951_));
  NOR4_X1    g02949(.A1(new_n3950_), .A2(new_n3257_), .A3(new_n3245_), .A4(new_n3951_), .ZN(new_n3952_));
  AOI21_X1   g02950(.A1(new_n3236_), .A2(new_n3260_), .B(new_n3258_), .ZN(new_n3953_));
  OAI21_X1   g02951(.A1(new_n3952_), .A2(new_n3953_), .B(new_n3256_), .ZN(new_n3954_));
  AOI21_X1   g02952(.A1(new_n3260_), .A2(new_n3236_), .B(new_n3248_), .ZN(new_n3955_));
  INV_X1     g02953(.I(new_n3261_), .ZN(new_n3956_));
  OAI21_X1   g02954(.A1(new_n3956_), .A2(new_n3955_), .B(new_n3226_), .ZN(new_n3957_));
  NAND2_X1   g02955(.A1(new_n3957_), .A2(new_n3954_), .ZN(new_n3958_));
  NAND3_X1   g02956(.A1(new_n3209_), .A2(new_n3957_), .A3(new_n3954_), .ZN(new_n3959_));
  AOI22_X1   g02957(.A1(new_n3959_), .A2(new_n3208_), .B1(new_n3958_), .B2(new_n3267_), .ZN(new_n3960_));
  AOI21_X1   g02958(.A1(new_n3181_), .A2(new_n1350_), .B(new_n3187_), .ZN(new_n3961_));
  AOI21_X1   g02959(.A1(new_n3197_), .A2(new_n1380_), .B(new_n3157_), .ZN(new_n3962_));
  INV_X1     g02960(.I(new_n3962_), .ZN(new_n3963_));
  NOR2_X1    g02961(.A1(new_n3963_), .A2(new_n3961_), .ZN(new_n3964_));
  OAI21_X1   g02962(.A1(new_n3204_), .A2(new_n3182_), .B(new_n3192_), .ZN(new_n3965_));
  NOR2_X1    g02963(.A1(new_n3965_), .A2(new_n3962_), .ZN(new_n3966_));
  NOR2_X1    g02964(.A1(new_n3195_), .A2(new_n3198_), .ZN(new_n3967_));
  OAI22_X1   g02965(.A1(new_n3964_), .A2(new_n3966_), .B1(new_n3967_), .B2(new_n3189_), .ZN(new_n3968_));
  NAND2_X1   g02966(.A1(new_n3965_), .A2(new_n3962_), .ZN(new_n3969_));
  NAND2_X1   g02967(.A1(new_n3963_), .A2(new_n3961_), .ZN(new_n3970_));
  OAI21_X1   g02968(.A1(new_n3205_), .A2(new_n3194_), .B(new_n3166_), .ZN(new_n3971_));
  NAND4_X1   g02969(.A1(new_n3970_), .A2(new_n3971_), .A3(new_n3271_), .A4(new_n3969_), .ZN(new_n3972_));
  NAND2_X1   g02970(.A1(new_n3968_), .A2(new_n3972_), .ZN(new_n3973_));
  NAND2_X1   g02971(.A1(new_n3236_), .A2(new_n1282_), .ZN(new_n3974_));
  NAND2_X1   g02972(.A1(new_n3974_), .A2(new_n3244_), .ZN(new_n3975_));
  AOI21_X1   g02973(.A1(new_n3225_), .A2(new_n1319_), .B(new_n3219_), .ZN(new_n3976_));
  NAND2_X1   g02974(.A1(new_n3975_), .A2(new_n3976_), .ZN(new_n3977_));
  AOI21_X1   g02975(.A1(new_n3236_), .A2(new_n1282_), .B(new_n3239_), .ZN(new_n3978_));
  OAI21_X1   g02976(.A1(new_n3255_), .A2(new_n3212_), .B(new_n3252_), .ZN(new_n3979_));
  NAND2_X1   g02977(.A1(new_n3979_), .A2(new_n3978_), .ZN(new_n3980_));
  NAND2_X1   g02978(.A1(new_n3250_), .A2(new_n3256_), .ZN(new_n3981_));
  AOI22_X1   g02979(.A1(new_n3981_), .A2(new_n3247_), .B1(new_n3977_), .B2(new_n3980_), .ZN(new_n3982_));
  NOR2_X1    g02980(.A1(new_n3979_), .A2(new_n3978_), .ZN(new_n3983_));
  NOR2_X1    g02981(.A1(new_n3975_), .A2(new_n3976_), .ZN(new_n3984_));
  NOR2_X1    g02982(.A1(new_n3953_), .A2(new_n3226_), .ZN(new_n3985_));
  NOR4_X1    g02983(.A1(new_n3985_), .A2(new_n3984_), .A3(new_n3983_), .A4(new_n3952_), .ZN(new_n3986_));
  NOR2_X1    g02984(.A1(new_n3982_), .A2(new_n3986_), .ZN(new_n3987_));
  NAND2_X1   g02985(.A1(new_n3973_), .A2(new_n3987_), .ZN(new_n3988_));
  NAND2_X1   g02986(.A1(new_n3970_), .A2(new_n3969_), .ZN(new_n3989_));
  NAND2_X1   g02987(.A1(new_n3971_), .A2(new_n3271_), .ZN(new_n3990_));
  NOR3_X1    g02988(.A1(new_n3964_), .A2(new_n3189_), .A3(new_n3966_), .ZN(new_n3991_));
  AOI22_X1   g02989(.A1(new_n3991_), .A2(new_n3971_), .B1(new_n3989_), .B2(new_n3990_), .ZN(new_n3992_));
  OAI22_X1   g02990(.A1(new_n3952_), .A2(new_n3985_), .B1(new_n3984_), .B2(new_n3983_), .ZN(new_n3993_));
  NAND4_X1   g02991(.A1(new_n3981_), .A2(new_n3247_), .A3(new_n3977_), .A4(new_n3980_), .ZN(new_n3994_));
  NAND2_X1   g02992(.A1(new_n3994_), .A2(new_n3993_), .ZN(new_n3995_));
  NAND2_X1   g02993(.A1(new_n3992_), .A2(new_n3995_), .ZN(new_n3996_));
  AOI21_X1   g02994(.A1(new_n3996_), .A2(new_n3988_), .B(new_n3960_), .ZN(new_n3997_));
  OAI22_X1   g02995(.A1(new_n3277_), .A2(new_n3268_), .B1(new_n3209_), .B2(new_n3263_), .ZN(new_n3998_));
  NOR2_X1    g02996(.A1(new_n3992_), .A2(new_n3995_), .ZN(new_n3999_));
  NOR2_X1    g02997(.A1(new_n3973_), .A2(new_n3987_), .ZN(new_n4000_));
  NOR3_X1    g02998(.A1(new_n3999_), .A2(new_n4000_), .A3(new_n3998_), .ZN(new_n4001_));
  NOR2_X1    g02999(.A1(new_n3997_), .A2(new_n4001_), .ZN(new_n4002_));
  NAND2_X1   g03000(.A1(new_n3949_), .A2(new_n4002_), .ZN(new_n4003_));
  AOI21_X1   g03001(.A1(new_n3947_), .A2(new_n3946_), .B(new_n3945_), .ZN(new_n4004_));
  NOR3_X1    g03002(.A1(new_n3901_), .A2(new_n3935_), .A3(new_n3942_), .ZN(new_n4005_));
  NOR2_X1    g03003(.A1(new_n4005_), .A2(new_n4004_), .ZN(new_n4006_));
  OAI21_X1   g03004(.A1(new_n3999_), .A2(new_n4000_), .B(new_n3998_), .ZN(new_n4007_));
  NAND3_X1   g03005(.A1(new_n3996_), .A2(new_n3988_), .A3(new_n3960_), .ZN(new_n4008_));
  NAND2_X1   g03006(.A1(new_n4007_), .A2(new_n4008_), .ZN(new_n4009_));
  NAND2_X1   g03007(.A1(new_n4006_), .A2(new_n4009_), .ZN(new_n4010_));
  AOI21_X1   g03008(.A1(new_n4003_), .A2(new_n4010_), .B(new_n3900_), .ZN(new_n4011_));
  NAND2_X1   g03009(.A1(new_n3150_), .A2(new_n3287_), .ZN(new_n4012_));
  NAND2_X1   g03010(.A1(new_n4012_), .A2(new_n3288_), .ZN(new_n4013_));
  NOR2_X1    g03011(.A1(new_n4006_), .A2(new_n4009_), .ZN(new_n4014_));
  NOR2_X1    g03012(.A1(new_n3949_), .A2(new_n4002_), .ZN(new_n4015_));
  NOR3_X1    g03013(.A1(new_n4015_), .A2(new_n4014_), .A3(new_n4013_), .ZN(new_n4016_));
  NOR2_X1    g03014(.A1(new_n4011_), .A2(new_n4016_), .ZN(new_n4017_));
  NOR3_X1    g03015(.A1(new_n3541_), .A2(new_n3539_), .A3(new_n3542_), .ZN(new_n4018_));
  OAI21_X1   g03016(.A1(new_n3416_), .A2(new_n4018_), .B(new_n3543_), .ZN(new_n4019_));
  NOR3_X1    g03017(.A1(new_n3380_), .A2(new_n3407_), .A3(new_n3392_), .ZN(new_n4020_));
  OAI21_X1   g03018(.A1(new_n3338_), .A2(new_n4020_), .B(new_n3412_), .ZN(new_n4021_));
  INV_X1     g03019(.I(new_n3323_), .ZN(new_n4022_));
  OAI21_X1   g03020(.A1(new_n3329_), .A2(new_n3316_), .B(new_n4022_), .ZN(new_n4023_));
  NAND2_X1   g03021(.A1(new_n3301_), .A2(new_n3299_), .ZN(new_n4024_));
  AOI21_X1   g03022(.A1(new_n4024_), .A2(new_n1250_), .B(new_n3297_), .ZN(new_n4025_));
  NAND2_X1   g03023(.A1(new_n4023_), .A2(new_n4025_), .ZN(new_n4026_));
  AOI21_X1   g03024(.A1(new_n3313_), .A2(new_n1219_), .B(new_n3323_), .ZN(new_n4027_));
  INV_X1     g03025(.I(new_n4025_), .ZN(new_n4028_));
  NAND2_X1   g03026(.A1(new_n4028_), .A2(new_n4027_), .ZN(new_n4029_));
  NAND2_X1   g03027(.A1(new_n4029_), .A2(new_n4026_), .ZN(new_n4030_));
  OAI21_X1   g03028(.A1(new_n3330_), .A2(new_n3326_), .B(new_n3302_), .ZN(new_n4031_));
  NOR2_X1    g03029(.A1(new_n3324_), .A2(new_n3304_), .ZN(new_n4032_));
  NAND4_X1   g03030(.A1(new_n4032_), .A2(new_n3313_), .A3(new_n3323_), .A4(new_n3320_), .ZN(new_n4033_));
  NAND2_X1   g03031(.A1(new_n4031_), .A2(new_n4033_), .ZN(new_n4034_));
  NOR2_X1    g03032(.A1(new_n4028_), .A2(new_n4027_), .ZN(new_n4035_));
  NOR2_X1    g03033(.A1(new_n4023_), .A2(new_n4025_), .ZN(new_n4036_));
  NOR3_X1    g03034(.A1(new_n4035_), .A2(new_n3325_), .A3(new_n4036_), .ZN(new_n4037_));
  AOI22_X1   g03035(.A1(new_n4037_), .A2(new_n4031_), .B1(new_n4030_), .B2(new_n4034_), .ZN(new_n4038_));
  AOI21_X1   g03036(.A1(new_n3377_), .A2(new_n1150_), .B(new_n3395_), .ZN(new_n4039_));
  OAI21_X1   g03037(.A1(new_n3384_), .A2(new_n3341_), .B(new_n3381_), .ZN(new_n4040_));
  NOR2_X1    g03038(.A1(new_n4040_), .A2(new_n4039_), .ZN(new_n4041_));
  INV_X1     g03039(.I(new_n4039_), .ZN(new_n4042_));
  AOI21_X1   g03040(.A1(new_n3353_), .A2(new_n1187_), .B(new_n3348_), .ZN(new_n4043_));
  NOR2_X1    g03041(.A1(new_n4042_), .A2(new_n4043_), .ZN(new_n4044_));
  NOR2_X1    g03042(.A1(new_n3399_), .A2(new_n3354_), .ZN(new_n4045_));
  OAI22_X1   g03043(.A1(new_n4045_), .A2(new_n3398_), .B1(new_n4041_), .B2(new_n4044_), .ZN(new_n4046_));
  NAND2_X1   g03044(.A1(new_n4042_), .A2(new_n4043_), .ZN(new_n4047_));
  NAND2_X1   g03045(.A1(new_n4040_), .A2(new_n4039_), .ZN(new_n4048_));
  NAND2_X1   g03046(.A1(new_n3379_), .A2(new_n3385_), .ZN(new_n4049_));
  NAND4_X1   g03047(.A1(new_n4049_), .A2(new_n3373_), .A3(new_n4047_), .A4(new_n4048_), .ZN(new_n4050_));
  NAND2_X1   g03048(.A1(new_n4050_), .A2(new_n4046_), .ZN(new_n4051_));
  NOR2_X1    g03049(.A1(new_n4038_), .A2(new_n4051_), .ZN(new_n4052_));
  NOR2_X1    g03050(.A1(new_n3331_), .A2(new_n3333_), .ZN(new_n4053_));
  OAI22_X1   g03051(.A1(new_n4053_), .A2(new_n3325_), .B1(new_n4035_), .B2(new_n4036_), .ZN(new_n4054_));
  NAND4_X1   g03052(.A1(new_n4029_), .A2(new_n4031_), .A3(new_n4033_), .A4(new_n4026_), .ZN(new_n4055_));
  NAND2_X1   g03053(.A1(new_n4054_), .A2(new_n4055_), .ZN(new_n4056_));
  NAND2_X1   g03054(.A1(new_n4048_), .A2(new_n4047_), .ZN(new_n4057_));
  NAND2_X1   g03055(.A1(new_n4049_), .A2(new_n3373_), .ZN(new_n4058_));
  NOR3_X1    g03056(.A1(new_n4041_), .A2(new_n4044_), .A3(new_n3398_), .ZN(new_n4059_));
  AOI22_X1   g03057(.A1(new_n4058_), .A2(new_n4057_), .B1(new_n4059_), .B2(new_n4049_), .ZN(new_n4060_));
  NOR2_X1    g03058(.A1(new_n4056_), .A2(new_n4060_), .ZN(new_n4061_));
  OAI21_X1   g03059(.A1(new_n4061_), .A2(new_n4052_), .B(new_n4021_), .ZN(new_n4062_));
  NAND2_X1   g03060(.A1(new_n3404_), .A2(new_n3400_), .ZN(new_n4063_));
  AOI22_X1   g03061(.A1(new_n3410_), .A2(new_n3411_), .B1(new_n3407_), .B2(new_n4063_), .ZN(new_n4064_));
  NAND2_X1   g03062(.A1(new_n4056_), .A2(new_n4060_), .ZN(new_n4065_));
  NAND2_X1   g03063(.A1(new_n4038_), .A2(new_n4051_), .ZN(new_n4066_));
  NAND3_X1   g03064(.A1(new_n4065_), .A2(new_n4066_), .A3(new_n4064_), .ZN(new_n4067_));
  NOR3_X1    g03065(.A1(new_n3468_), .A2(new_n3514_), .A3(new_n3521_), .ZN(new_n4068_));
  OAI21_X1   g03066(.A1(new_n3533_), .A2(new_n4068_), .B(new_n3522_), .ZN(new_n4069_));
  NOR2_X1    g03067(.A1(new_n3438_), .A2(new_n3444_), .ZN(new_n4070_));
  NAND4_X1   g03068(.A1(new_n4070_), .A2(new_n1100_), .A3(new_n1130_), .A4(new_n3452_), .ZN(new_n4071_));
  OAI21_X1   g03069(.A1(new_n3438_), .A2(new_n3445_), .B(new_n3443_), .ZN(new_n4072_));
  NOR2_X1    g03070(.A1(new_n3458_), .A2(new_n3423_), .ZN(new_n4073_));
  AOI21_X1   g03071(.A1(new_n3457_), .A2(new_n1119_), .B(new_n4073_), .ZN(new_n4074_));
  NAND2_X1   g03072(.A1(new_n4074_), .A2(new_n4072_), .ZN(new_n4075_));
  AOI21_X1   g03073(.A1(new_n3451_), .A2(new_n1089_), .B(new_n3447_), .ZN(new_n4076_));
  INV_X1     g03074(.I(new_n1119_), .ZN(new_n4077_));
  OAI21_X1   g03075(.A1(new_n3429_), .A2(new_n4077_), .B(new_n3425_), .ZN(new_n4078_));
  NAND2_X1   g03076(.A1(new_n4078_), .A2(new_n4076_), .ZN(new_n4079_));
  NOR2_X1    g03077(.A1(new_n3461_), .A2(new_n3438_), .ZN(new_n4080_));
  OAI21_X1   g03078(.A1(new_n3454_), .A2(new_n4080_), .B(new_n3430_), .ZN(new_n4081_));
  AOI22_X1   g03079(.A1(new_n4081_), .A2(new_n4071_), .B1(new_n4075_), .B2(new_n4079_), .ZN(new_n4082_));
  NOR2_X1    g03080(.A1(new_n4078_), .A2(new_n4076_), .ZN(new_n4083_));
  NOR2_X1    g03081(.A1(new_n4074_), .A2(new_n4072_), .ZN(new_n4084_));
  NAND2_X1   g03082(.A1(new_n3452_), .A2(new_n3451_), .ZN(new_n4085_));
  AOI21_X1   g03083(.A1(new_n3453_), .A2(new_n4085_), .B(new_n3460_), .ZN(new_n4086_));
  NOR4_X1    g03084(.A1(new_n4086_), .A2(new_n4083_), .A3(new_n4084_), .A4(new_n3449_), .ZN(new_n4087_));
  NOR2_X1    g03085(.A1(new_n4087_), .A2(new_n4082_), .ZN(new_n4088_));
  AOI21_X1   g03086(.A1(new_n3497_), .A2(new_n1019_), .B(new_n3500_), .ZN(new_n4089_));
  AOI21_X1   g03087(.A1(new_n3486_), .A2(new_n1056_), .B(new_n3478_), .ZN(new_n4090_));
  INV_X1     g03088(.I(new_n4090_), .ZN(new_n4091_));
  NOR2_X1    g03089(.A1(new_n4091_), .A2(new_n4089_), .ZN(new_n4092_));
  NOR2_X1    g03090(.A1(new_n3498_), .A2(new_n3495_), .ZN(new_n4093_));
  NOR2_X1    g03091(.A1(new_n3503_), .A2(new_n1036_), .ZN(new_n4094_));
  NOR2_X1    g03092(.A1(new_n4094_), .A2(new_n4093_), .ZN(new_n4095_));
  OAI21_X1   g03093(.A1(new_n4095_), .A2(new_n3501_), .B(new_n3505_), .ZN(new_n4096_));
  NOR2_X1    g03094(.A1(new_n4096_), .A2(new_n4090_), .ZN(new_n4097_));
  NOR2_X1    g03095(.A1(new_n3512_), .A2(new_n3487_), .ZN(new_n4098_));
  OAI22_X1   g03096(.A1(new_n4098_), .A2(new_n3526_), .B1(new_n4092_), .B2(new_n4097_), .ZN(new_n4099_));
  NAND2_X1   g03097(.A1(new_n4096_), .A2(new_n4090_), .ZN(new_n4100_));
  NAND2_X1   g03098(.A1(new_n4091_), .A2(new_n4089_), .ZN(new_n4101_));
  NOR2_X1    g03099(.A1(new_n3525_), .A2(new_n4095_), .ZN(new_n4102_));
  OAI21_X1   g03100(.A1(new_n4102_), .A2(new_n3511_), .B(new_n3516_), .ZN(new_n4103_));
  NAND4_X1   g03101(.A1(new_n4103_), .A2(new_n3508_), .A3(new_n4101_), .A4(new_n4100_), .ZN(new_n4104_));
  NAND2_X1   g03102(.A1(new_n4099_), .A2(new_n4104_), .ZN(new_n4105_));
  NOR2_X1    g03103(.A1(new_n4088_), .A2(new_n4105_), .ZN(new_n4106_));
  OAI22_X1   g03104(.A1(new_n4086_), .A2(new_n3449_), .B1(new_n4084_), .B2(new_n4083_), .ZN(new_n4107_));
  NAND4_X1   g03105(.A1(new_n4081_), .A2(new_n4075_), .A3(new_n4079_), .A4(new_n4071_), .ZN(new_n4108_));
  NAND2_X1   g03106(.A1(new_n4107_), .A2(new_n4108_), .ZN(new_n4109_));
  AOI22_X1   g03107(.A1(new_n4103_), .A2(new_n3508_), .B1(new_n4101_), .B2(new_n4100_), .ZN(new_n4110_));
  NOR4_X1    g03108(.A1(new_n4098_), .A2(new_n4092_), .A3(new_n4097_), .A4(new_n3526_), .ZN(new_n4111_));
  NOR2_X1    g03109(.A1(new_n4110_), .A2(new_n4111_), .ZN(new_n4112_));
  NOR2_X1    g03110(.A1(new_n4109_), .A2(new_n4112_), .ZN(new_n4113_));
  OAI21_X1   g03111(.A1(new_n4106_), .A2(new_n4113_), .B(new_n4069_), .ZN(new_n4114_));
  NAND2_X1   g03112(.A1(new_n3529_), .A2(new_n3527_), .ZN(new_n4115_));
  AOI22_X1   g03113(.A1(new_n3530_), .A2(new_n3465_), .B1(new_n4115_), .B2(new_n3468_), .ZN(new_n4116_));
  NAND2_X1   g03114(.A1(new_n4109_), .A2(new_n4112_), .ZN(new_n4117_));
  NAND2_X1   g03115(.A1(new_n4088_), .A2(new_n4105_), .ZN(new_n4118_));
  NAND3_X1   g03116(.A1(new_n4118_), .A2(new_n4117_), .A3(new_n4116_), .ZN(new_n4119_));
  NAND2_X1   g03117(.A1(new_n4114_), .A2(new_n4119_), .ZN(new_n4120_));
  AOI21_X1   g03118(.A1(new_n4062_), .A2(new_n4067_), .B(new_n4120_), .ZN(new_n4121_));
  NAND2_X1   g03119(.A1(new_n4062_), .A2(new_n4067_), .ZN(new_n4122_));
  AOI21_X1   g03120(.A1(new_n4118_), .A2(new_n4117_), .B(new_n4116_), .ZN(new_n4123_));
  NOR3_X1    g03121(.A1(new_n4106_), .A2(new_n4113_), .A3(new_n4069_), .ZN(new_n4124_));
  NOR2_X1    g03122(.A1(new_n4124_), .A2(new_n4123_), .ZN(new_n4125_));
  NOR2_X1    g03123(.A1(new_n4122_), .A2(new_n4125_), .ZN(new_n4126_));
  OAI21_X1   g03124(.A1(new_n4121_), .A2(new_n4126_), .B(new_n4019_), .ZN(new_n4127_));
  NAND2_X1   g03125(.A1(new_n3532_), .A2(new_n3536_), .ZN(new_n4128_));
  AOI22_X1   g03126(.A1(new_n3415_), .A2(new_n3538_), .B1(new_n4128_), .B2(new_n3542_), .ZN(new_n4129_));
  NAND2_X1   g03127(.A1(new_n4122_), .A2(new_n4125_), .ZN(new_n4130_));
  NAND3_X1   g03128(.A1(new_n4120_), .A2(new_n4062_), .A3(new_n4067_), .ZN(new_n4131_));
  NAND3_X1   g03129(.A1(new_n4130_), .A2(new_n4131_), .A3(new_n4129_), .ZN(new_n4132_));
  NAND2_X1   g03130(.A1(new_n4127_), .A2(new_n4132_), .ZN(new_n4133_));
  NOR2_X1    g03131(.A1(new_n4017_), .A2(new_n4133_), .ZN(new_n4134_));
  OAI21_X1   g03132(.A1(new_n4015_), .A2(new_n4014_), .B(new_n4013_), .ZN(new_n4135_));
  NAND3_X1   g03133(.A1(new_n4003_), .A2(new_n4010_), .A3(new_n3900_), .ZN(new_n4136_));
  NAND2_X1   g03134(.A1(new_n4135_), .A2(new_n4136_), .ZN(new_n4137_));
  AOI21_X1   g03135(.A1(new_n4130_), .A2(new_n4131_), .B(new_n4129_), .ZN(new_n4138_));
  NOR3_X1    g03136(.A1(new_n4121_), .A2(new_n4126_), .A3(new_n4019_), .ZN(new_n4139_));
  NOR2_X1    g03137(.A1(new_n4139_), .A2(new_n4138_), .ZN(new_n4140_));
  NOR2_X1    g03138(.A1(new_n4137_), .A2(new_n4140_), .ZN(new_n4141_));
  OAI21_X1   g03139(.A1(new_n4141_), .A2(new_n4134_), .B(new_n3899_), .ZN(new_n4142_));
  NOR2_X1    g03140(.A1(new_n3557_), .A2(new_n3290_), .ZN(new_n4143_));
  NOR2_X1    g03141(.A1(new_n4143_), .A2(new_n3558_), .ZN(new_n4144_));
  NAND2_X1   g03142(.A1(new_n4137_), .A2(new_n4140_), .ZN(new_n4145_));
  NAND2_X1   g03143(.A1(new_n4017_), .A2(new_n4133_), .ZN(new_n4146_));
  NAND3_X1   g03144(.A1(new_n4145_), .A2(new_n4146_), .A3(new_n4144_), .ZN(new_n4147_));
  NAND2_X1   g03145(.A1(new_n4142_), .A2(new_n4147_), .ZN(new_n4148_));
  NAND3_X1   g03146(.A1(new_n3894_), .A2(new_n3897_), .A3(new_n4148_), .ZN(new_n4149_));
  NOR3_X1    g03147(.A1(new_n3896_), .A2(new_n3895_), .A3(new_n3892_), .ZN(new_n4150_));
  AOI21_X1   g03148(.A1(new_n3885_), .A2(new_n3891_), .B(new_n3893_), .ZN(new_n4151_));
  AOI21_X1   g03149(.A1(new_n4145_), .A2(new_n4146_), .B(new_n4144_), .ZN(new_n4152_));
  NOR3_X1    g03150(.A1(new_n3899_), .A2(new_n4141_), .A3(new_n4134_), .ZN(new_n4153_));
  NOR2_X1    g03151(.A1(new_n4153_), .A2(new_n4152_), .ZN(new_n4154_));
  OAI21_X1   g03152(.A1(new_n4151_), .A2(new_n4150_), .B(new_n4154_), .ZN(new_n4155_));
  AOI21_X1   g03153(.A1(new_n4155_), .A2(new_n4149_), .B(new_n3562_), .ZN(new_n4156_));
  INV_X1     g03154(.I(new_n3024_), .ZN(new_n4157_));
  AOI21_X1   g03155(.A1(new_n4157_), .A2(new_n3025_), .B(new_n2543_), .ZN(new_n4158_));
  INV_X1     g03156(.I(new_n3017_), .ZN(new_n4159_));
  NAND2_X1   g03157(.A1(new_n3020_), .A2(new_n3019_), .ZN(new_n4160_));
  NAND2_X1   g03158(.A1(new_n4160_), .A2(new_n2734_), .ZN(new_n4161_));
  NAND3_X1   g03159(.A1(new_n4159_), .A2(new_n4161_), .A3(new_n3023_), .ZN(new_n4162_));
  AOI21_X1   g03160(.A1(new_n4162_), .A2(new_n3029_), .B(new_n2544_), .ZN(new_n4163_));
  NOR2_X1    g03161(.A1(new_n4158_), .A2(new_n4163_), .ZN(new_n4164_));
  INV_X1     g03162(.I(new_n3560_), .ZN(new_n4165_));
  NOR3_X1    g03163(.A1(new_n4158_), .A2(new_n4163_), .A3(new_n2345_), .ZN(new_n4166_));
  OAI22_X1   g03164(.A1(new_n4166_), .A2(new_n4165_), .B1(new_n4164_), .B2(new_n2346_), .ZN(new_n4167_));
  NOR3_X1    g03165(.A1(new_n4151_), .A2(new_n4150_), .A3(new_n4154_), .ZN(new_n4168_));
  AOI21_X1   g03166(.A1(new_n3894_), .A2(new_n3897_), .B(new_n4148_), .ZN(new_n4169_));
  NOR3_X1    g03167(.A1(new_n4168_), .A2(new_n4169_), .A3(new_n4167_), .ZN(new_n4170_));
  NOR2_X1    g03168(.A1(new_n4156_), .A2(new_n4170_), .ZN(new_n4171_));
  INV_X1     g03169(.I(\A[414] ), .ZN(new_n4172_));
  NAND2_X1   g03170(.A1(\A[412] ), .A2(\A[413] ), .ZN(new_n4173_));
  XNOR2_X1   g03171(.A1(\A[412] ), .A2(\A[413] ), .ZN(new_n4174_));
  OAI21_X1   g03172(.A1(new_n4174_), .A2(new_n4172_), .B(new_n4173_), .ZN(new_n4175_));
  INV_X1     g03173(.I(\A[411] ), .ZN(new_n4176_));
  NAND2_X1   g03174(.A1(\A[409] ), .A2(\A[410] ), .ZN(new_n4177_));
  XNOR2_X1   g03175(.A1(\A[409] ), .A2(\A[410] ), .ZN(new_n4178_));
  OAI21_X1   g03176(.A1(new_n4178_), .A2(new_n4176_), .B(new_n4177_), .ZN(new_n4179_));
  INV_X1     g03177(.I(\A[409] ), .ZN(new_n4180_));
  NOR2_X1    g03178(.A1(new_n4180_), .A2(\A[410] ), .ZN(new_n4181_));
  INV_X1     g03179(.I(\A[410] ), .ZN(new_n4182_));
  NOR2_X1    g03180(.A1(new_n4182_), .A2(\A[409] ), .ZN(new_n4183_));
  OAI21_X1   g03181(.A1(new_n4181_), .A2(new_n4183_), .B(new_n4176_), .ZN(new_n4184_));
  NAND2_X1   g03182(.A1(new_n4182_), .A2(\A[409] ), .ZN(new_n4185_));
  NAND2_X1   g03183(.A1(new_n4180_), .A2(\A[410] ), .ZN(new_n4186_));
  NAND3_X1   g03184(.A1(new_n4185_), .A2(new_n4186_), .A3(\A[411] ), .ZN(new_n4187_));
  INV_X1     g03185(.I(\A[412] ), .ZN(new_n4188_));
  NOR2_X1    g03186(.A1(new_n4188_), .A2(\A[413] ), .ZN(new_n4189_));
  INV_X1     g03187(.I(\A[413] ), .ZN(new_n4190_));
  NOR2_X1    g03188(.A1(new_n4190_), .A2(\A[412] ), .ZN(new_n4191_));
  OAI21_X1   g03189(.A1(new_n4189_), .A2(new_n4191_), .B(new_n4172_), .ZN(new_n4192_));
  NAND2_X1   g03190(.A1(new_n4190_), .A2(\A[412] ), .ZN(new_n4193_));
  NAND2_X1   g03191(.A1(new_n4188_), .A2(\A[413] ), .ZN(new_n4194_));
  NAND3_X1   g03192(.A1(new_n4193_), .A2(new_n4194_), .A3(\A[414] ), .ZN(new_n4195_));
  AOI22_X1   g03193(.A1(new_n4184_), .A2(new_n4187_), .B1(new_n4192_), .B2(new_n4195_), .ZN(new_n4196_));
  NAND3_X1   g03194(.A1(new_n4196_), .A2(new_n4175_), .A3(new_n4179_), .ZN(new_n4197_));
  AOI21_X1   g03195(.A1(new_n4185_), .A2(new_n4186_), .B(\A[411] ), .ZN(new_n4198_));
  NOR3_X1    g03196(.A1(new_n4181_), .A2(new_n4183_), .A3(new_n4176_), .ZN(new_n4199_));
  NOR2_X1    g03197(.A1(new_n4198_), .A2(new_n4199_), .ZN(new_n4200_));
  NAND2_X1   g03198(.A1(new_n4192_), .A2(new_n4195_), .ZN(new_n4201_));
  NAND2_X1   g03199(.A1(new_n4200_), .A2(new_n4201_), .ZN(new_n4202_));
  NAND2_X1   g03200(.A1(new_n4184_), .A2(new_n4187_), .ZN(new_n4203_));
  AOI21_X1   g03201(.A1(new_n4193_), .A2(new_n4194_), .B(\A[414] ), .ZN(new_n4204_));
  OAI21_X1   g03202(.A1(new_n4188_), .A2(\A[413] ), .B(\A[414] ), .ZN(new_n4205_));
  NOR2_X1    g03203(.A1(new_n4205_), .A2(new_n4191_), .ZN(new_n4206_));
  NOR2_X1    g03204(.A1(new_n4204_), .A2(new_n4206_), .ZN(new_n4207_));
  NAND2_X1   g03205(.A1(new_n4203_), .A2(new_n4207_), .ZN(new_n4208_));
  NAND2_X1   g03206(.A1(new_n4202_), .A2(new_n4208_), .ZN(new_n4209_));
  NAND2_X1   g03207(.A1(new_n4209_), .A2(new_n4197_), .ZN(new_n4210_));
  INV_X1     g03208(.I(\A[404] ), .ZN(new_n4211_));
  NOR2_X1    g03209(.A1(new_n4211_), .A2(\A[403] ), .ZN(new_n4212_));
  XNOR2_X1   g03210(.A1(\A[403] ), .A2(\A[404] ), .ZN(new_n4213_));
  INV_X1     g03211(.I(\A[403] ), .ZN(new_n4214_));
  OAI21_X1   g03212(.A1(new_n4214_), .A2(\A[404] ), .B(\A[405] ), .ZN(new_n4215_));
  OAI22_X1   g03213(.A1(new_n4213_), .A2(\A[405] ), .B1(new_n4212_), .B2(new_n4215_), .ZN(new_n4216_));
  INV_X1     g03214(.I(\A[408] ), .ZN(new_n4217_));
  INV_X1     g03215(.I(\A[406] ), .ZN(new_n4218_));
  NAND2_X1   g03216(.A1(new_n4218_), .A2(\A[407] ), .ZN(new_n4219_));
  XOR2_X1    g03217(.A1(\A[406] ), .A2(\A[407] ), .Z(new_n4220_));
  INV_X1     g03218(.I(\A[407] ), .ZN(new_n4221_));
  AOI21_X1   g03219(.A1(\A[406] ), .A2(new_n4221_), .B(new_n4217_), .ZN(new_n4222_));
  AOI22_X1   g03220(.A1(new_n4220_), .A2(new_n4217_), .B1(new_n4219_), .B2(new_n4222_), .ZN(new_n4223_));
  NOR2_X1    g03221(.A1(new_n4216_), .A2(new_n4223_), .ZN(new_n4224_));
  NAND2_X1   g03222(.A1(new_n4211_), .A2(\A[403] ), .ZN(new_n4225_));
  NAND2_X1   g03223(.A1(new_n4214_), .A2(\A[404] ), .ZN(new_n4226_));
  AOI21_X1   g03224(.A1(new_n4225_), .A2(new_n4226_), .B(\A[405] ), .ZN(new_n4227_));
  NOR2_X1    g03225(.A1(new_n4215_), .A2(new_n4212_), .ZN(new_n4228_));
  NOR2_X1    g03226(.A1(new_n4227_), .A2(new_n4228_), .ZN(new_n4229_));
  NOR2_X1    g03227(.A1(new_n4221_), .A2(\A[406] ), .ZN(new_n4230_));
  NOR2_X1    g03228(.A1(new_n4218_), .A2(\A[407] ), .ZN(new_n4231_));
  NOR2_X1    g03229(.A1(new_n4231_), .A2(new_n4230_), .ZN(new_n4232_));
  OAI21_X1   g03230(.A1(new_n4218_), .A2(\A[407] ), .B(\A[408] ), .ZN(new_n4233_));
  OAI22_X1   g03231(.A1(new_n4232_), .A2(\A[408] ), .B1(new_n4230_), .B2(new_n4233_), .ZN(new_n4234_));
  NOR2_X1    g03232(.A1(new_n4234_), .A2(new_n4229_), .ZN(new_n4235_));
  NOR2_X1    g03233(.A1(new_n4235_), .A2(new_n4224_), .ZN(new_n4236_));
  NOR2_X1    g03234(.A1(new_n4218_), .A2(new_n4221_), .ZN(new_n4237_));
  AOI21_X1   g03235(.A1(new_n4220_), .A2(\A[408] ), .B(new_n4237_), .ZN(new_n4238_));
  NAND2_X1   g03236(.A1(new_n4225_), .A2(new_n4226_), .ZN(new_n4239_));
  NAND2_X1   g03237(.A1(\A[403] ), .A2(\A[404] ), .ZN(new_n4240_));
  INV_X1     g03238(.I(new_n4240_), .ZN(new_n4241_));
  AOI21_X1   g03239(.A1(new_n4239_), .A2(\A[405] ), .B(new_n4241_), .ZN(new_n4242_));
  NAND2_X1   g03240(.A1(new_n4221_), .A2(\A[406] ), .ZN(new_n4243_));
  AOI21_X1   g03241(.A1(new_n4243_), .A2(new_n4219_), .B(\A[408] ), .ZN(new_n4244_));
  NOR3_X1    g03242(.A1(new_n4231_), .A2(new_n4230_), .A3(new_n4217_), .ZN(new_n4245_));
  OAI22_X1   g03243(.A1(new_n4244_), .A2(new_n4245_), .B1(new_n4227_), .B2(new_n4228_), .ZN(new_n4246_));
  NOR3_X1    g03244(.A1(new_n4246_), .A2(new_n4238_), .A3(new_n4242_), .ZN(new_n4247_));
  NOR2_X1    g03245(.A1(new_n4236_), .A2(new_n4247_), .ZN(new_n4248_));
  NAND2_X1   g03246(.A1(new_n4248_), .A2(new_n4210_), .ZN(new_n4249_));
  INV_X1     g03247(.I(new_n4173_), .ZN(new_n4250_));
  XOR2_X1    g03248(.A1(\A[412] ), .A2(\A[413] ), .Z(new_n4251_));
  AOI21_X1   g03249(.A1(new_n4251_), .A2(\A[414] ), .B(new_n4250_), .ZN(new_n4252_));
  INV_X1     g03250(.I(new_n4177_), .ZN(new_n4253_));
  XOR2_X1    g03251(.A1(\A[409] ), .A2(\A[410] ), .Z(new_n4254_));
  AOI21_X1   g03252(.A1(new_n4254_), .A2(\A[411] ), .B(new_n4253_), .ZN(new_n4255_));
  OAI22_X1   g03253(.A1(new_n4198_), .A2(new_n4199_), .B1(new_n4204_), .B2(new_n4206_), .ZN(new_n4256_));
  NOR3_X1    g03254(.A1(new_n4256_), .A2(new_n4252_), .A3(new_n4255_), .ZN(new_n4257_));
  NOR2_X1    g03255(.A1(new_n4203_), .A2(new_n4207_), .ZN(new_n4258_));
  NOR2_X1    g03256(.A1(new_n4200_), .A2(new_n4201_), .ZN(new_n4259_));
  NOR2_X1    g03257(.A1(new_n4259_), .A2(new_n4258_), .ZN(new_n4260_));
  NOR2_X1    g03258(.A1(new_n4260_), .A2(new_n4257_), .ZN(new_n4261_));
  NAND2_X1   g03259(.A1(new_n4234_), .A2(new_n4229_), .ZN(new_n4262_));
  NAND2_X1   g03260(.A1(new_n4216_), .A2(new_n4223_), .ZN(new_n4263_));
  NAND2_X1   g03261(.A1(new_n4262_), .A2(new_n4263_), .ZN(new_n4264_));
  INV_X1     g03262(.I(new_n4237_), .ZN(new_n4265_));
  OAI21_X1   g03263(.A1(new_n4232_), .A2(new_n4217_), .B(new_n4265_), .ZN(new_n4266_));
  INV_X1     g03264(.I(\A[405] ), .ZN(new_n4267_));
  OAI21_X1   g03265(.A1(new_n4213_), .A2(new_n4267_), .B(new_n4240_), .ZN(new_n4268_));
  NAND4_X1   g03266(.A1(new_n4234_), .A2(new_n4266_), .A3(new_n4216_), .A4(new_n4268_), .ZN(new_n4269_));
  NAND2_X1   g03267(.A1(new_n4264_), .A2(new_n4269_), .ZN(new_n4270_));
  NAND2_X1   g03268(.A1(new_n4261_), .A2(new_n4270_), .ZN(new_n4271_));
  NAND2_X1   g03269(.A1(new_n4249_), .A2(new_n4271_), .ZN(new_n4272_));
  INV_X1     g03270(.I(\A[402] ), .ZN(new_n4273_));
  INV_X1     g03271(.I(\A[400] ), .ZN(new_n4274_));
  INV_X1     g03272(.I(\A[401] ), .ZN(new_n4275_));
  NOR2_X1    g03273(.A1(new_n4274_), .A2(new_n4275_), .ZN(new_n4276_));
  INV_X1     g03274(.I(new_n4276_), .ZN(new_n4277_));
  NOR2_X1    g03275(.A1(new_n4274_), .A2(\A[401] ), .ZN(new_n4278_));
  NOR2_X1    g03276(.A1(new_n4275_), .A2(\A[400] ), .ZN(new_n4279_));
  NOR2_X1    g03277(.A1(new_n4278_), .A2(new_n4279_), .ZN(new_n4280_));
  OAI21_X1   g03278(.A1(new_n4280_), .A2(new_n4273_), .B(new_n4277_), .ZN(new_n4281_));
  INV_X1     g03279(.I(\A[399] ), .ZN(new_n4282_));
  INV_X1     g03280(.I(\A[397] ), .ZN(new_n4283_));
  INV_X1     g03281(.I(\A[398] ), .ZN(new_n4284_));
  NOR2_X1    g03282(.A1(new_n4283_), .A2(new_n4284_), .ZN(new_n4285_));
  INV_X1     g03283(.I(new_n4285_), .ZN(new_n4286_));
  NOR2_X1    g03284(.A1(new_n4283_), .A2(\A[398] ), .ZN(new_n4287_));
  NOR2_X1    g03285(.A1(new_n4284_), .A2(\A[397] ), .ZN(new_n4288_));
  NOR2_X1    g03286(.A1(new_n4287_), .A2(new_n4288_), .ZN(new_n4289_));
  OAI21_X1   g03287(.A1(new_n4289_), .A2(new_n4282_), .B(new_n4286_), .ZN(new_n4290_));
  XOR2_X1    g03288(.A1(\A[397] ), .A2(\A[398] ), .Z(new_n4291_));
  NAND2_X1   g03289(.A1(new_n4291_), .A2(new_n4282_), .ZN(new_n4292_));
  NAND2_X1   g03290(.A1(new_n4284_), .A2(\A[397] ), .ZN(new_n4293_));
  NAND2_X1   g03291(.A1(new_n4283_), .A2(\A[398] ), .ZN(new_n4294_));
  NAND3_X1   g03292(.A1(new_n4293_), .A2(new_n4294_), .A3(\A[399] ), .ZN(new_n4295_));
  OAI21_X1   g03293(.A1(new_n4278_), .A2(new_n4279_), .B(new_n4273_), .ZN(new_n4296_));
  NAND2_X1   g03294(.A1(new_n4274_), .A2(\A[401] ), .ZN(new_n4297_));
  AOI21_X1   g03295(.A1(\A[400] ), .A2(new_n4275_), .B(new_n4273_), .ZN(new_n4298_));
  NAND2_X1   g03296(.A1(new_n4298_), .A2(new_n4297_), .ZN(new_n4299_));
  AOI22_X1   g03297(.A1(new_n4292_), .A2(new_n4295_), .B1(new_n4296_), .B2(new_n4299_), .ZN(new_n4300_));
  NAND3_X1   g03298(.A1(new_n4300_), .A2(new_n4281_), .A3(new_n4290_), .ZN(new_n4301_));
  AOI21_X1   g03299(.A1(new_n4293_), .A2(new_n4294_), .B(\A[399] ), .ZN(new_n4302_));
  OAI21_X1   g03300(.A1(new_n4283_), .A2(\A[398] ), .B(\A[399] ), .ZN(new_n4303_));
  NOR2_X1    g03301(.A1(new_n4303_), .A2(new_n4288_), .ZN(new_n4304_));
  NOR2_X1    g03302(.A1(new_n4302_), .A2(new_n4304_), .ZN(new_n4305_));
  NAND2_X1   g03303(.A1(new_n4299_), .A2(new_n4296_), .ZN(new_n4306_));
  NAND2_X1   g03304(.A1(new_n4306_), .A2(new_n4305_), .ZN(new_n4307_));
  OAI21_X1   g03305(.A1(\A[399] ), .A2(new_n4289_), .B(new_n4295_), .ZN(new_n4308_));
  NAND2_X1   g03306(.A1(new_n4275_), .A2(\A[400] ), .ZN(new_n4309_));
  AOI21_X1   g03307(.A1(new_n4309_), .A2(new_n4297_), .B(\A[402] ), .ZN(new_n4310_));
  NOR3_X1    g03308(.A1(new_n4278_), .A2(new_n4279_), .A3(new_n4273_), .ZN(new_n4311_));
  NOR2_X1    g03309(.A1(new_n4310_), .A2(new_n4311_), .ZN(new_n4312_));
  NAND2_X1   g03310(.A1(new_n4308_), .A2(new_n4312_), .ZN(new_n4313_));
  NAND2_X1   g03311(.A1(new_n4313_), .A2(new_n4307_), .ZN(new_n4314_));
  NAND2_X1   g03312(.A1(new_n4314_), .A2(new_n4301_), .ZN(new_n4315_));
  INV_X1     g03313(.I(\A[393] ), .ZN(new_n4316_));
  XOR2_X1    g03314(.A1(\A[391] ), .A2(\A[392] ), .Z(new_n4317_));
  NAND2_X1   g03315(.A1(new_n4317_), .A2(new_n4316_), .ZN(new_n4318_));
  INV_X1     g03316(.I(\A[391] ), .ZN(new_n4319_));
  NAND2_X1   g03317(.A1(new_n4319_), .A2(\A[392] ), .ZN(new_n4320_));
  INV_X1     g03318(.I(\A[392] ), .ZN(new_n4321_));
  AOI21_X1   g03319(.A1(\A[391] ), .A2(new_n4321_), .B(new_n4316_), .ZN(new_n4322_));
  NAND2_X1   g03320(.A1(new_n4322_), .A2(new_n4320_), .ZN(new_n4323_));
  NAND2_X1   g03321(.A1(new_n4318_), .A2(new_n4323_), .ZN(new_n4324_));
  INV_X1     g03322(.I(\A[395] ), .ZN(new_n4325_));
  NAND2_X1   g03323(.A1(new_n4325_), .A2(\A[394] ), .ZN(new_n4326_));
  INV_X1     g03324(.I(\A[394] ), .ZN(new_n4327_));
  NAND2_X1   g03325(.A1(new_n4327_), .A2(\A[395] ), .ZN(new_n4328_));
  AOI21_X1   g03326(.A1(new_n4326_), .A2(new_n4328_), .B(\A[396] ), .ZN(new_n4329_));
  INV_X1     g03327(.I(\A[396] ), .ZN(new_n4330_));
  NOR2_X1    g03328(.A1(new_n4327_), .A2(\A[395] ), .ZN(new_n4331_));
  NOR2_X1    g03329(.A1(new_n4325_), .A2(\A[394] ), .ZN(new_n4332_));
  NOR3_X1    g03330(.A1(new_n4331_), .A2(new_n4332_), .A3(new_n4330_), .ZN(new_n4333_));
  NOR2_X1    g03331(.A1(new_n4329_), .A2(new_n4333_), .ZN(new_n4334_));
  NOR2_X1    g03332(.A1(new_n4324_), .A2(new_n4334_), .ZN(new_n4335_));
  AOI22_X1   g03333(.A1(new_n4317_), .A2(new_n4316_), .B1(new_n4320_), .B2(new_n4322_), .ZN(new_n4336_));
  OAI21_X1   g03334(.A1(new_n4331_), .A2(new_n4332_), .B(new_n4330_), .ZN(new_n4337_));
  NAND3_X1   g03335(.A1(new_n4326_), .A2(new_n4328_), .A3(\A[396] ), .ZN(new_n4338_));
  NAND2_X1   g03336(.A1(new_n4337_), .A2(new_n4338_), .ZN(new_n4339_));
  NOR2_X1    g03337(.A1(new_n4339_), .A2(new_n4336_), .ZN(new_n4340_));
  NOR2_X1    g03338(.A1(new_n4335_), .A2(new_n4340_), .ZN(new_n4341_));
  NAND2_X1   g03339(.A1(new_n4326_), .A2(new_n4328_), .ZN(new_n4342_));
  NOR2_X1    g03340(.A1(new_n4327_), .A2(new_n4325_), .ZN(new_n4343_));
  AOI21_X1   g03341(.A1(new_n4342_), .A2(\A[396] ), .B(new_n4343_), .ZN(new_n4344_));
  NOR2_X1    g03342(.A1(new_n4319_), .A2(new_n4321_), .ZN(new_n4345_));
  AOI21_X1   g03343(.A1(new_n4317_), .A2(\A[393] ), .B(new_n4345_), .ZN(new_n4346_));
  NOR2_X1    g03344(.A1(new_n4319_), .A2(\A[392] ), .ZN(new_n4347_));
  INV_X1     g03345(.I(new_n4347_), .ZN(new_n4348_));
  AOI21_X1   g03346(.A1(new_n4348_), .A2(new_n4320_), .B(\A[393] ), .ZN(new_n4349_));
  NOR2_X1    g03347(.A1(new_n4321_), .A2(\A[391] ), .ZN(new_n4350_));
  NOR3_X1    g03348(.A1(new_n4347_), .A2(new_n4350_), .A3(new_n4316_), .ZN(new_n4351_));
  OAI22_X1   g03349(.A1(new_n4349_), .A2(new_n4351_), .B1(new_n4329_), .B2(new_n4333_), .ZN(new_n4352_));
  NOR3_X1    g03350(.A1(new_n4352_), .A2(new_n4344_), .A3(new_n4346_), .ZN(new_n4353_));
  NOR2_X1    g03351(.A1(new_n4341_), .A2(new_n4353_), .ZN(new_n4354_));
  NOR2_X1    g03352(.A1(new_n4354_), .A2(new_n4315_), .ZN(new_n4355_));
  INV_X1     g03353(.I(new_n4355_), .ZN(new_n4356_));
  NAND2_X1   g03354(.A1(new_n4354_), .A2(new_n4315_), .ZN(new_n4357_));
  NAND3_X1   g03355(.A1(new_n4272_), .A2(new_n4356_), .A3(new_n4357_), .ZN(new_n4358_));
  NOR2_X1    g03356(.A1(new_n4261_), .A2(new_n4270_), .ZN(new_n4359_));
  NOR2_X1    g03357(.A1(new_n4248_), .A2(new_n4210_), .ZN(new_n4360_));
  NOR2_X1    g03358(.A1(new_n4360_), .A2(new_n4359_), .ZN(new_n4361_));
  XOR2_X1    g03359(.A1(\A[400] ), .A2(\A[401] ), .Z(new_n4362_));
  AOI21_X1   g03360(.A1(new_n4362_), .A2(\A[402] ), .B(new_n4276_), .ZN(new_n4363_));
  AOI21_X1   g03361(.A1(new_n4291_), .A2(\A[399] ), .B(new_n4285_), .ZN(new_n4364_));
  OAI22_X1   g03362(.A1(new_n4310_), .A2(new_n4311_), .B1(new_n4302_), .B2(new_n4304_), .ZN(new_n4365_));
  NOR3_X1    g03363(.A1(new_n4365_), .A2(new_n4363_), .A3(new_n4364_), .ZN(new_n4366_));
  NOR2_X1    g03364(.A1(new_n4308_), .A2(new_n4312_), .ZN(new_n4367_));
  NOR2_X1    g03365(.A1(new_n4306_), .A2(new_n4305_), .ZN(new_n4368_));
  NOR2_X1    g03366(.A1(new_n4367_), .A2(new_n4368_), .ZN(new_n4369_));
  NOR2_X1    g03367(.A1(new_n4369_), .A2(new_n4366_), .ZN(new_n4370_));
  NOR3_X1    g03368(.A1(new_n4370_), .A2(new_n4341_), .A3(new_n4353_), .ZN(new_n4371_));
  OAI21_X1   g03369(.A1(new_n4355_), .A2(new_n4371_), .B(new_n4361_), .ZN(new_n4372_));
  NAND2_X1   g03370(.A1(new_n4372_), .A2(new_n4358_), .ZN(new_n4373_));
  INV_X1     g03371(.I(\A[385] ), .ZN(new_n4374_));
  NAND2_X1   g03372(.A1(new_n4374_), .A2(\A[386] ), .ZN(new_n4375_));
  INV_X1     g03373(.I(\A[386] ), .ZN(new_n4376_));
  INV_X1     g03374(.I(\A[387] ), .ZN(new_n4377_));
  AOI21_X1   g03375(.A1(\A[385] ), .A2(new_n4376_), .B(new_n4377_), .ZN(new_n4378_));
  NAND2_X1   g03376(.A1(new_n4378_), .A2(new_n4375_), .ZN(new_n4379_));
  NOR2_X1    g03377(.A1(new_n4376_), .A2(\A[385] ), .ZN(new_n4380_));
  NOR2_X1    g03378(.A1(new_n4374_), .A2(\A[386] ), .ZN(new_n4381_));
  OAI21_X1   g03379(.A1(new_n4380_), .A2(new_n4381_), .B(new_n4377_), .ZN(new_n4382_));
  NAND2_X1   g03380(.A1(new_n4379_), .A2(new_n4382_), .ZN(new_n4383_));
  INV_X1     g03381(.I(\A[390] ), .ZN(new_n4384_));
  INV_X1     g03382(.I(\A[388] ), .ZN(new_n4385_));
  NAND2_X1   g03383(.A1(new_n4385_), .A2(\A[389] ), .ZN(new_n4386_));
  INV_X1     g03384(.I(\A[389] ), .ZN(new_n4387_));
  AOI21_X1   g03385(.A1(\A[388] ), .A2(new_n4387_), .B(new_n4384_), .ZN(new_n4388_));
  XOR2_X1    g03386(.A1(\A[388] ), .A2(\A[389] ), .Z(new_n4389_));
  AOI22_X1   g03387(.A1(new_n4389_), .A2(new_n4384_), .B1(new_n4386_), .B2(new_n4388_), .ZN(new_n4390_));
  XOR2_X1    g03388(.A1(new_n4383_), .A2(new_n4390_), .Z(new_n4391_));
  NAND2_X1   g03389(.A1(\A[388] ), .A2(\A[389] ), .ZN(new_n4392_));
  INV_X1     g03390(.I(new_n4392_), .ZN(new_n4393_));
  AOI21_X1   g03391(.A1(new_n4389_), .A2(\A[390] ), .B(new_n4393_), .ZN(new_n4394_));
  XOR2_X1    g03392(.A1(\A[385] ), .A2(\A[386] ), .Z(new_n4395_));
  NAND2_X1   g03393(.A1(\A[385] ), .A2(\A[386] ), .ZN(new_n4396_));
  INV_X1     g03394(.I(new_n4396_), .ZN(new_n4397_));
  AOI21_X1   g03395(.A1(new_n4395_), .A2(\A[387] ), .B(new_n4397_), .ZN(new_n4398_));
  NOR3_X1    g03396(.A1(new_n4380_), .A2(new_n4381_), .A3(new_n4377_), .ZN(new_n4399_));
  NAND2_X1   g03397(.A1(new_n4376_), .A2(\A[385] ), .ZN(new_n4400_));
  AOI21_X1   g03398(.A1(new_n4375_), .A2(new_n4400_), .B(\A[387] ), .ZN(new_n4401_));
  NOR2_X1    g03399(.A1(new_n4387_), .A2(\A[388] ), .ZN(new_n4402_));
  NOR2_X1    g03400(.A1(new_n4385_), .A2(\A[389] ), .ZN(new_n4403_));
  NOR3_X1    g03401(.A1(new_n4402_), .A2(new_n4403_), .A3(new_n4384_), .ZN(new_n4404_));
  NAND2_X1   g03402(.A1(new_n4387_), .A2(\A[388] ), .ZN(new_n4405_));
  AOI21_X1   g03403(.A1(new_n4386_), .A2(new_n4405_), .B(\A[390] ), .ZN(new_n4406_));
  OAI22_X1   g03404(.A1(new_n4399_), .A2(new_n4401_), .B1(new_n4406_), .B2(new_n4404_), .ZN(new_n4407_));
  NOR3_X1    g03405(.A1(new_n4407_), .A2(new_n4394_), .A3(new_n4398_), .ZN(new_n4408_));
  NOR2_X1    g03406(.A1(new_n4391_), .A2(new_n4408_), .ZN(new_n4409_));
  INV_X1     g03407(.I(\A[381] ), .ZN(new_n4410_));
  INV_X1     g03408(.I(\A[379] ), .ZN(new_n4411_));
  NAND2_X1   g03409(.A1(new_n4411_), .A2(\A[380] ), .ZN(new_n4412_));
  INV_X1     g03410(.I(\A[380] ), .ZN(new_n4413_));
  AOI21_X1   g03411(.A1(\A[379] ), .A2(new_n4413_), .B(new_n4410_), .ZN(new_n4414_));
  XOR2_X1    g03412(.A1(\A[379] ), .A2(\A[380] ), .Z(new_n4415_));
  AOI22_X1   g03413(.A1(new_n4415_), .A2(new_n4410_), .B1(new_n4412_), .B2(new_n4414_), .ZN(new_n4416_));
  INV_X1     g03414(.I(\A[382] ), .ZN(new_n4417_));
  NAND2_X1   g03415(.A1(new_n4417_), .A2(\A[383] ), .ZN(new_n4418_));
  INV_X1     g03416(.I(\A[383] ), .ZN(new_n4419_));
  INV_X1     g03417(.I(\A[384] ), .ZN(new_n4420_));
  AOI21_X1   g03418(.A1(\A[382] ), .A2(new_n4419_), .B(new_n4420_), .ZN(new_n4421_));
  NAND2_X1   g03419(.A1(new_n4421_), .A2(new_n4418_), .ZN(new_n4422_));
  NOR2_X1    g03420(.A1(new_n4419_), .A2(\A[382] ), .ZN(new_n4423_));
  NOR2_X1    g03421(.A1(new_n4417_), .A2(\A[383] ), .ZN(new_n4424_));
  OAI21_X1   g03422(.A1(new_n4423_), .A2(new_n4424_), .B(new_n4420_), .ZN(new_n4425_));
  NAND2_X1   g03423(.A1(new_n4422_), .A2(new_n4425_), .ZN(new_n4426_));
  NAND2_X1   g03424(.A1(new_n4426_), .A2(new_n4416_), .ZN(new_n4427_));
  NAND2_X1   g03425(.A1(new_n4414_), .A2(new_n4412_), .ZN(new_n4428_));
  NOR2_X1    g03426(.A1(new_n4413_), .A2(\A[379] ), .ZN(new_n4429_));
  NOR2_X1    g03427(.A1(new_n4411_), .A2(\A[380] ), .ZN(new_n4430_));
  OAI21_X1   g03428(.A1(new_n4429_), .A2(new_n4430_), .B(new_n4410_), .ZN(new_n4431_));
  NAND2_X1   g03429(.A1(new_n4428_), .A2(new_n4431_), .ZN(new_n4432_));
  XOR2_X1    g03430(.A1(\A[382] ), .A2(\A[383] ), .Z(new_n4433_));
  AOI22_X1   g03431(.A1(new_n4433_), .A2(new_n4420_), .B1(new_n4418_), .B2(new_n4421_), .ZN(new_n4434_));
  NAND2_X1   g03432(.A1(new_n4432_), .A2(new_n4434_), .ZN(new_n4435_));
  NAND2_X1   g03433(.A1(new_n4427_), .A2(new_n4435_), .ZN(new_n4436_));
  NOR2_X1    g03434(.A1(new_n4417_), .A2(new_n4419_), .ZN(new_n4437_));
  AOI21_X1   g03435(.A1(new_n4433_), .A2(\A[384] ), .B(new_n4437_), .ZN(new_n4438_));
  NOR2_X1    g03436(.A1(new_n4411_), .A2(new_n4413_), .ZN(new_n4439_));
  AOI21_X1   g03437(.A1(new_n4415_), .A2(\A[381] ), .B(new_n4439_), .ZN(new_n4440_));
  NOR4_X1    g03438(.A1(new_n4416_), .A2(new_n4434_), .A3(new_n4438_), .A4(new_n4440_), .ZN(new_n4441_));
  INV_X1     g03439(.I(new_n4441_), .ZN(new_n4442_));
  NAND2_X1   g03440(.A1(new_n4436_), .A2(new_n4442_), .ZN(new_n4443_));
  NOR2_X1    g03441(.A1(new_n4409_), .A2(new_n4443_), .ZN(new_n4444_));
  NOR2_X1    g03442(.A1(new_n4401_), .A2(new_n4399_), .ZN(new_n4445_));
  NAND2_X1   g03443(.A1(new_n4388_), .A2(new_n4386_), .ZN(new_n4446_));
  OAI21_X1   g03444(.A1(new_n4402_), .A2(new_n4403_), .B(new_n4384_), .ZN(new_n4447_));
  NAND2_X1   g03445(.A1(new_n4446_), .A2(new_n4447_), .ZN(new_n4448_));
  NAND2_X1   g03446(.A1(new_n4445_), .A2(new_n4448_), .ZN(new_n4449_));
  NAND2_X1   g03447(.A1(new_n4383_), .A2(new_n4390_), .ZN(new_n4450_));
  NAND2_X1   g03448(.A1(new_n4449_), .A2(new_n4450_), .ZN(new_n4451_));
  NOR2_X1    g03449(.A1(new_n4402_), .A2(new_n4403_), .ZN(new_n4452_));
  OAI21_X1   g03450(.A1(new_n4452_), .A2(new_n4384_), .B(new_n4392_), .ZN(new_n4453_));
  NOR2_X1    g03451(.A1(new_n4380_), .A2(new_n4381_), .ZN(new_n4454_));
  OAI21_X1   g03452(.A1(new_n4454_), .A2(new_n4377_), .B(new_n4396_), .ZN(new_n4455_));
  AOI22_X1   g03453(.A1(new_n4379_), .A2(new_n4382_), .B1(new_n4446_), .B2(new_n4447_), .ZN(new_n4456_));
  NAND3_X1   g03454(.A1(new_n4456_), .A2(new_n4453_), .A3(new_n4455_), .ZN(new_n4457_));
  NAND2_X1   g03455(.A1(new_n4451_), .A2(new_n4457_), .ZN(new_n4458_));
  NOR2_X1    g03456(.A1(new_n4432_), .A2(new_n4434_), .ZN(new_n4459_));
  NOR2_X1    g03457(.A1(new_n4426_), .A2(new_n4416_), .ZN(new_n4460_));
  NOR2_X1    g03458(.A1(new_n4459_), .A2(new_n4460_), .ZN(new_n4461_));
  NOR2_X1    g03459(.A1(new_n4461_), .A2(new_n4441_), .ZN(new_n4462_));
  NOR2_X1    g03460(.A1(new_n4462_), .A2(new_n4458_), .ZN(new_n4463_));
  NOR2_X1    g03461(.A1(new_n4444_), .A2(new_n4463_), .ZN(new_n4464_));
  INV_X1     g03462(.I(\A[373] ), .ZN(new_n4465_));
  NAND2_X1   g03463(.A1(new_n4465_), .A2(\A[374] ), .ZN(new_n4466_));
  INV_X1     g03464(.I(\A[374] ), .ZN(new_n4467_));
  INV_X1     g03465(.I(\A[375] ), .ZN(new_n4468_));
  AOI21_X1   g03466(.A1(\A[373] ), .A2(new_n4467_), .B(new_n4468_), .ZN(new_n4469_));
  NAND2_X1   g03467(.A1(new_n4469_), .A2(new_n4466_), .ZN(new_n4470_));
  NOR2_X1    g03468(.A1(new_n4467_), .A2(\A[373] ), .ZN(new_n4471_));
  NOR2_X1    g03469(.A1(new_n4465_), .A2(\A[374] ), .ZN(new_n4472_));
  OAI21_X1   g03470(.A1(new_n4471_), .A2(new_n4472_), .B(new_n4468_), .ZN(new_n4473_));
  NAND2_X1   g03471(.A1(new_n4470_), .A2(new_n4473_), .ZN(new_n4474_));
  INV_X1     g03472(.I(\A[378] ), .ZN(new_n4475_));
  INV_X1     g03473(.I(\A[377] ), .ZN(new_n4476_));
  NOR2_X1    g03474(.A1(new_n4476_), .A2(\A[376] ), .ZN(new_n4477_));
  INV_X1     g03475(.I(\A[376] ), .ZN(new_n4478_));
  NOR2_X1    g03476(.A1(new_n4478_), .A2(\A[377] ), .ZN(new_n4479_));
  NOR3_X1    g03477(.A1(new_n4477_), .A2(new_n4479_), .A3(new_n4475_), .ZN(new_n4480_));
  NAND2_X1   g03478(.A1(new_n4478_), .A2(\A[377] ), .ZN(new_n4481_));
  NAND2_X1   g03479(.A1(new_n4476_), .A2(\A[376] ), .ZN(new_n4482_));
  AOI21_X1   g03480(.A1(new_n4481_), .A2(new_n4482_), .B(\A[378] ), .ZN(new_n4483_));
  NOR2_X1    g03481(.A1(new_n4483_), .A2(new_n4480_), .ZN(new_n4484_));
  NOR2_X1    g03482(.A1(new_n4484_), .A2(new_n4474_), .ZN(new_n4485_));
  NOR3_X1    g03483(.A1(new_n4471_), .A2(new_n4472_), .A3(new_n4468_), .ZN(new_n4486_));
  NAND2_X1   g03484(.A1(new_n4467_), .A2(\A[373] ), .ZN(new_n4487_));
  AOI21_X1   g03485(.A1(new_n4466_), .A2(new_n4487_), .B(\A[375] ), .ZN(new_n4488_));
  NOR2_X1    g03486(.A1(new_n4488_), .A2(new_n4486_), .ZN(new_n4489_));
  NAND3_X1   g03487(.A1(new_n4481_), .A2(new_n4482_), .A3(\A[378] ), .ZN(new_n4490_));
  OAI21_X1   g03488(.A1(new_n4477_), .A2(new_n4479_), .B(new_n4475_), .ZN(new_n4491_));
  NAND2_X1   g03489(.A1(new_n4491_), .A2(new_n4490_), .ZN(new_n4492_));
  NOR2_X1    g03490(.A1(new_n4489_), .A2(new_n4492_), .ZN(new_n4493_));
  NOR2_X1    g03491(.A1(new_n4485_), .A2(new_n4493_), .ZN(new_n4494_));
  NAND2_X1   g03492(.A1(new_n4481_), .A2(new_n4482_), .ZN(new_n4495_));
  NOR2_X1    g03493(.A1(new_n4478_), .A2(new_n4476_), .ZN(new_n4496_));
  AOI21_X1   g03494(.A1(new_n4495_), .A2(\A[378] ), .B(new_n4496_), .ZN(new_n4497_));
  NAND2_X1   g03495(.A1(new_n4466_), .A2(new_n4487_), .ZN(new_n4498_));
  NOR2_X1    g03496(.A1(new_n4465_), .A2(new_n4467_), .ZN(new_n4499_));
  AOI21_X1   g03497(.A1(new_n4498_), .A2(\A[375] ), .B(new_n4499_), .ZN(new_n4500_));
  OAI22_X1   g03498(.A1(new_n4486_), .A2(new_n4488_), .B1(new_n4483_), .B2(new_n4480_), .ZN(new_n4501_));
  NOR3_X1    g03499(.A1(new_n4501_), .A2(new_n4497_), .A3(new_n4500_), .ZN(new_n4502_));
  NOR2_X1    g03500(.A1(new_n4494_), .A2(new_n4502_), .ZN(new_n4503_));
  INV_X1     g03501(.I(\A[369] ), .ZN(new_n4504_));
  INV_X1     g03502(.I(\A[368] ), .ZN(new_n4505_));
  NOR2_X1    g03503(.A1(new_n4505_), .A2(\A[367] ), .ZN(new_n4506_));
  INV_X1     g03504(.I(\A[367] ), .ZN(new_n4507_));
  NOR2_X1    g03505(.A1(new_n4507_), .A2(\A[368] ), .ZN(new_n4508_));
  NOR3_X1    g03506(.A1(new_n4506_), .A2(new_n4508_), .A3(new_n4504_), .ZN(new_n4509_));
  NAND2_X1   g03507(.A1(new_n4507_), .A2(\A[368] ), .ZN(new_n4510_));
  NAND2_X1   g03508(.A1(new_n4505_), .A2(\A[367] ), .ZN(new_n4511_));
  AOI21_X1   g03509(.A1(new_n4510_), .A2(new_n4511_), .B(\A[369] ), .ZN(new_n4512_));
  NOR2_X1    g03510(.A1(new_n4512_), .A2(new_n4509_), .ZN(new_n4513_));
  INV_X1     g03511(.I(\A[370] ), .ZN(new_n4514_));
  NAND2_X1   g03512(.A1(new_n4514_), .A2(\A[371] ), .ZN(new_n4515_));
  INV_X1     g03513(.I(\A[371] ), .ZN(new_n4516_));
  INV_X1     g03514(.I(\A[372] ), .ZN(new_n4517_));
  AOI21_X1   g03515(.A1(\A[370] ), .A2(new_n4516_), .B(new_n4517_), .ZN(new_n4518_));
  NAND2_X1   g03516(.A1(new_n4518_), .A2(new_n4515_), .ZN(new_n4519_));
  NOR2_X1    g03517(.A1(new_n4516_), .A2(\A[370] ), .ZN(new_n4520_));
  NOR2_X1    g03518(.A1(new_n4514_), .A2(\A[371] ), .ZN(new_n4521_));
  OAI21_X1   g03519(.A1(new_n4520_), .A2(new_n4521_), .B(new_n4517_), .ZN(new_n4522_));
  NAND2_X1   g03520(.A1(new_n4519_), .A2(new_n4522_), .ZN(new_n4523_));
  NAND2_X1   g03521(.A1(new_n4513_), .A2(new_n4523_), .ZN(new_n4524_));
  AOI21_X1   g03522(.A1(\A[367] ), .A2(new_n4505_), .B(new_n4504_), .ZN(new_n4525_));
  NAND2_X1   g03523(.A1(new_n4525_), .A2(new_n4510_), .ZN(new_n4526_));
  OAI21_X1   g03524(.A1(new_n4506_), .A2(new_n4508_), .B(new_n4504_), .ZN(new_n4527_));
  NAND2_X1   g03525(.A1(new_n4526_), .A2(new_n4527_), .ZN(new_n4528_));
  XOR2_X1    g03526(.A1(\A[370] ), .A2(\A[371] ), .Z(new_n4529_));
  AOI22_X1   g03527(.A1(new_n4529_), .A2(new_n4517_), .B1(new_n4515_), .B2(new_n4518_), .ZN(new_n4530_));
  NAND2_X1   g03528(.A1(new_n4528_), .A2(new_n4530_), .ZN(new_n4531_));
  NAND2_X1   g03529(.A1(new_n4524_), .A2(new_n4531_), .ZN(new_n4532_));
  NOR2_X1    g03530(.A1(new_n4520_), .A2(new_n4521_), .ZN(new_n4533_));
  NOR2_X1    g03531(.A1(new_n4514_), .A2(new_n4516_), .ZN(new_n4534_));
  INV_X1     g03532(.I(new_n4534_), .ZN(new_n4535_));
  OAI21_X1   g03533(.A1(new_n4533_), .A2(new_n4517_), .B(new_n4535_), .ZN(new_n4536_));
  NOR2_X1    g03534(.A1(new_n4506_), .A2(new_n4508_), .ZN(new_n4537_));
  NOR2_X1    g03535(.A1(new_n4507_), .A2(new_n4505_), .ZN(new_n4538_));
  INV_X1     g03536(.I(new_n4538_), .ZN(new_n4539_));
  OAI21_X1   g03537(.A1(new_n4537_), .A2(new_n4504_), .B(new_n4539_), .ZN(new_n4540_));
  AOI22_X1   g03538(.A1(new_n4526_), .A2(new_n4527_), .B1(new_n4519_), .B2(new_n4522_), .ZN(new_n4541_));
  NAND3_X1   g03539(.A1(new_n4541_), .A2(new_n4536_), .A3(new_n4540_), .ZN(new_n4542_));
  NAND2_X1   g03540(.A1(new_n4532_), .A2(new_n4542_), .ZN(new_n4543_));
  NOR2_X1    g03541(.A1(new_n4503_), .A2(new_n4543_), .ZN(new_n4544_));
  NOR2_X1    g03542(.A1(new_n4528_), .A2(new_n4530_), .ZN(new_n4545_));
  NOR2_X1    g03543(.A1(new_n4513_), .A2(new_n4523_), .ZN(new_n4546_));
  NOR2_X1    g03544(.A1(new_n4546_), .A2(new_n4545_), .ZN(new_n4547_));
  AOI21_X1   g03545(.A1(new_n4529_), .A2(\A[372] ), .B(new_n4534_), .ZN(new_n4548_));
  NAND2_X1   g03546(.A1(new_n4510_), .A2(new_n4511_), .ZN(new_n4549_));
  AOI21_X1   g03547(.A1(new_n4549_), .A2(\A[369] ), .B(new_n4538_), .ZN(new_n4550_));
  NOR3_X1    g03548(.A1(new_n4520_), .A2(new_n4521_), .A3(new_n4517_), .ZN(new_n4551_));
  NAND2_X1   g03549(.A1(new_n4516_), .A2(\A[370] ), .ZN(new_n4552_));
  AOI21_X1   g03550(.A1(new_n4515_), .A2(new_n4552_), .B(\A[372] ), .ZN(new_n4553_));
  OAI22_X1   g03551(.A1(new_n4509_), .A2(new_n4512_), .B1(new_n4553_), .B2(new_n4551_), .ZN(new_n4554_));
  NOR3_X1    g03552(.A1(new_n4554_), .A2(new_n4548_), .A3(new_n4550_), .ZN(new_n4555_));
  NOR2_X1    g03553(.A1(new_n4547_), .A2(new_n4555_), .ZN(new_n4556_));
  NOR3_X1    g03554(.A1(new_n4556_), .A2(new_n4494_), .A3(new_n4502_), .ZN(new_n4557_));
  OAI21_X1   g03555(.A1(new_n4544_), .A2(new_n4557_), .B(new_n4464_), .ZN(new_n4558_));
  NOR2_X1    g03556(.A1(new_n4557_), .A2(new_n4544_), .ZN(new_n4559_));
  OAI21_X1   g03557(.A1(new_n4444_), .A2(new_n4463_), .B(new_n4559_), .ZN(new_n4560_));
  NAND2_X1   g03558(.A1(new_n4558_), .A2(new_n4560_), .ZN(new_n4561_));
  XOR2_X1    g03559(.A1(new_n4561_), .A2(new_n4373_), .Z(new_n4562_));
  INV_X1     g03560(.I(\A[462] ), .ZN(new_n4563_));
  NAND2_X1   g03561(.A1(\A[460] ), .A2(\A[461] ), .ZN(new_n4564_));
  INV_X1     g03562(.I(\A[460] ), .ZN(new_n4565_));
  NOR2_X1    g03563(.A1(new_n4565_), .A2(\A[461] ), .ZN(new_n4566_));
  INV_X1     g03564(.I(\A[461] ), .ZN(new_n4567_));
  NOR2_X1    g03565(.A1(new_n4567_), .A2(\A[460] ), .ZN(new_n4568_));
  NOR2_X1    g03566(.A1(new_n4566_), .A2(new_n4568_), .ZN(new_n4569_));
  OAI21_X1   g03567(.A1(new_n4569_), .A2(new_n4563_), .B(new_n4564_), .ZN(new_n4570_));
  INV_X1     g03568(.I(\A[459] ), .ZN(new_n4571_));
  NAND2_X1   g03569(.A1(\A[457] ), .A2(\A[458] ), .ZN(new_n4572_));
  XNOR2_X1   g03570(.A1(\A[457] ), .A2(\A[458] ), .ZN(new_n4573_));
  OAI21_X1   g03571(.A1(new_n4573_), .A2(new_n4571_), .B(new_n4572_), .ZN(new_n4574_));
  INV_X1     g03572(.I(\A[457] ), .ZN(new_n4575_));
  NOR2_X1    g03573(.A1(new_n4575_), .A2(\A[458] ), .ZN(new_n4576_));
  INV_X1     g03574(.I(\A[458] ), .ZN(new_n4577_));
  NOR2_X1    g03575(.A1(new_n4577_), .A2(\A[457] ), .ZN(new_n4578_));
  OAI21_X1   g03576(.A1(new_n4576_), .A2(new_n4578_), .B(new_n4571_), .ZN(new_n4579_));
  NAND2_X1   g03577(.A1(new_n4575_), .A2(\A[458] ), .ZN(new_n4580_));
  AOI21_X1   g03578(.A1(\A[457] ), .A2(new_n4577_), .B(new_n4571_), .ZN(new_n4581_));
  NAND2_X1   g03579(.A1(new_n4581_), .A2(new_n4580_), .ZN(new_n4582_));
  OAI21_X1   g03580(.A1(new_n4566_), .A2(new_n4568_), .B(new_n4563_), .ZN(new_n4583_));
  NAND2_X1   g03581(.A1(new_n4567_), .A2(\A[460] ), .ZN(new_n4584_));
  NAND2_X1   g03582(.A1(new_n4565_), .A2(\A[461] ), .ZN(new_n4585_));
  NAND3_X1   g03583(.A1(new_n4584_), .A2(new_n4585_), .A3(\A[462] ), .ZN(new_n4586_));
  AOI22_X1   g03584(.A1(new_n4579_), .A2(new_n4582_), .B1(new_n4583_), .B2(new_n4586_), .ZN(new_n4587_));
  NAND3_X1   g03585(.A1(new_n4587_), .A2(new_n4570_), .A3(new_n4574_), .ZN(new_n4588_));
  NAND2_X1   g03586(.A1(new_n4582_), .A2(new_n4579_), .ZN(new_n4589_));
  AOI21_X1   g03587(.A1(new_n4584_), .A2(new_n4585_), .B(\A[462] ), .ZN(new_n4590_));
  NOR3_X1    g03588(.A1(new_n4566_), .A2(new_n4568_), .A3(new_n4563_), .ZN(new_n4591_));
  NOR2_X1    g03589(.A1(new_n4590_), .A2(new_n4591_), .ZN(new_n4592_));
  NAND2_X1   g03590(.A1(new_n4592_), .A2(new_n4589_), .ZN(new_n4593_));
  XOR2_X1    g03591(.A1(\A[457] ), .A2(\A[458] ), .Z(new_n4594_));
  AOI22_X1   g03592(.A1(new_n4594_), .A2(new_n4571_), .B1(new_n4580_), .B2(new_n4581_), .ZN(new_n4595_));
  NAND2_X1   g03593(.A1(new_n4583_), .A2(new_n4586_), .ZN(new_n4596_));
  NAND2_X1   g03594(.A1(new_n4596_), .A2(new_n4595_), .ZN(new_n4597_));
  NAND2_X1   g03595(.A1(new_n4593_), .A2(new_n4597_), .ZN(new_n4598_));
  NAND2_X1   g03596(.A1(new_n4598_), .A2(new_n4588_), .ZN(new_n4599_));
  NAND2_X1   g03597(.A1(\A[454] ), .A2(\A[455] ), .ZN(new_n4600_));
  INV_X1     g03598(.I(new_n4600_), .ZN(new_n4601_));
  XOR2_X1    g03599(.A1(\A[454] ), .A2(\A[455] ), .Z(new_n4602_));
  AOI21_X1   g03600(.A1(new_n4602_), .A2(\A[456] ), .B(new_n4601_), .ZN(new_n4603_));
  NAND2_X1   g03601(.A1(\A[451] ), .A2(\A[452] ), .ZN(new_n4604_));
  INV_X1     g03602(.I(new_n4604_), .ZN(new_n4605_));
  XOR2_X1    g03603(.A1(\A[451] ), .A2(\A[452] ), .Z(new_n4606_));
  AOI21_X1   g03604(.A1(new_n4606_), .A2(\A[453] ), .B(new_n4605_), .ZN(new_n4607_));
  INV_X1     g03605(.I(\A[452] ), .ZN(new_n4608_));
  NAND2_X1   g03606(.A1(new_n4608_), .A2(\A[451] ), .ZN(new_n4609_));
  INV_X1     g03607(.I(\A[451] ), .ZN(new_n4610_));
  NAND2_X1   g03608(.A1(new_n4610_), .A2(\A[452] ), .ZN(new_n4611_));
  AOI21_X1   g03609(.A1(new_n4609_), .A2(new_n4611_), .B(\A[453] ), .ZN(new_n4612_));
  INV_X1     g03610(.I(\A[453] ), .ZN(new_n4613_));
  NOR2_X1    g03611(.A1(new_n4610_), .A2(\A[452] ), .ZN(new_n4614_));
  NOR2_X1    g03612(.A1(new_n4608_), .A2(\A[451] ), .ZN(new_n4615_));
  NOR3_X1    g03613(.A1(new_n4614_), .A2(new_n4615_), .A3(new_n4613_), .ZN(new_n4616_));
  INV_X1     g03614(.I(\A[455] ), .ZN(new_n4617_));
  NAND2_X1   g03615(.A1(new_n4617_), .A2(\A[454] ), .ZN(new_n4618_));
  INV_X1     g03616(.I(\A[454] ), .ZN(new_n4619_));
  NAND2_X1   g03617(.A1(new_n4619_), .A2(\A[455] ), .ZN(new_n4620_));
  AOI21_X1   g03618(.A1(new_n4618_), .A2(new_n4620_), .B(\A[456] ), .ZN(new_n4621_));
  NOR2_X1    g03619(.A1(new_n4617_), .A2(\A[454] ), .ZN(new_n4622_));
  OAI21_X1   g03620(.A1(new_n4619_), .A2(\A[455] ), .B(\A[456] ), .ZN(new_n4623_));
  NOR2_X1    g03621(.A1(new_n4623_), .A2(new_n4622_), .ZN(new_n4624_));
  OAI22_X1   g03622(.A1(new_n4612_), .A2(new_n4616_), .B1(new_n4621_), .B2(new_n4624_), .ZN(new_n4625_));
  NOR3_X1    g03623(.A1(new_n4625_), .A2(new_n4603_), .A3(new_n4607_), .ZN(new_n4626_));
  OAI21_X1   g03624(.A1(new_n4614_), .A2(new_n4615_), .B(new_n4613_), .ZN(new_n4627_));
  AOI21_X1   g03625(.A1(\A[451] ), .A2(new_n4608_), .B(new_n4613_), .ZN(new_n4628_));
  NAND2_X1   g03626(.A1(new_n4628_), .A2(new_n4611_), .ZN(new_n4629_));
  NAND2_X1   g03627(.A1(new_n4629_), .A2(new_n4627_), .ZN(new_n4630_));
  NOR2_X1    g03628(.A1(new_n4621_), .A2(new_n4624_), .ZN(new_n4631_));
  NOR2_X1    g03629(.A1(new_n4630_), .A2(new_n4631_), .ZN(new_n4632_));
  AOI22_X1   g03630(.A1(new_n4606_), .A2(new_n4613_), .B1(new_n4611_), .B2(new_n4628_), .ZN(new_n4633_));
  INV_X1     g03631(.I(\A[456] ), .ZN(new_n4634_));
  NOR2_X1    g03632(.A1(new_n4619_), .A2(\A[455] ), .ZN(new_n4635_));
  OAI21_X1   g03633(.A1(new_n4635_), .A2(new_n4622_), .B(new_n4634_), .ZN(new_n4636_));
  NAND3_X1   g03634(.A1(new_n4618_), .A2(new_n4620_), .A3(\A[456] ), .ZN(new_n4637_));
  NAND2_X1   g03635(.A1(new_n4636_), .A2(new_n4637_), .ZN(new_n4638_));
  NOR2_X1    g03636(.A1(new_n4638_), .A2(new_n4633_), .ZN(new_n4639_));
  NOR2_X1    g03637(.A1(new_n4632_), .A2(new_n4639_), .ZN(new_n4640_));
  NOR2_X1    g03638(.A1(new_n4640_), .A2(new_n4626_), .ZN(new_n4641_));
  NOR2_X1    g03639(.A1(new_n4641_), .A2(new_n4599_), .ZN(new_n4642_));
  INV_X1     g03640(.I(new_n4564_), .ZN(new_n4643_));
  XOR2_X1    g03641(.A1(\A[460] ), .A2(\A[461] ), .Z(new_n4644_));
  AOI21_X1   g03642(.A1(new_n4644_), .A2(\A[462] ), .B(new_n4643_), .ZN(new_n4645_));
  INV_X1     g03643(.I(new_n4572_), .ZN(new_n4646_));
  AOI21_X1   g03644(.A1(new_n4594_), .A2(\A[459] ), .B(new_n4646_), .ZN(new_n4647_));
  NAND2_X1   g03645(.A1(new_n4577_), .A2(\A[457] ), .ZN(new_n4648_));
  AOI21_X1   g03646(.A1(new_n4648_), .A2(new_n4580_), .B(\A[459] ), .ZN(new_n4649_));
  NOR3_X1    g03647(.A1(new_n4576_), .A2(new_n4578_), .A3(new_n4571_), .ZN(new_n4650_));
  OAI22_X1   g03648(.A1(new_n4649_), .A2(new_n4650_), .B1(new_n4590_), .B2(new_n4591_), .ZN(new_n4651_));
  NOR3_X1    g03649(.A1(new_n4651_), .A2(new_n4645_), .A3(new_n4647_), .ZN(new_n4652_));
  NOR2_X1    g03650(.A1(new_n4596_), .A2(new_n4595_), .ZN(new_n4653_));
  NOR2_X1    g03651(.A1(new_n4592_), .A2(new_n4589_), .ZN(new_n4654_));
  NOR2_X1    g03652(.A1(new_n4654_), .A2(new_n4653_), .ZN(new_n4655_));
  NOR2_X1    g03653(.A1(new_n4655_), .A2(new_n4652_), .ZN(new_n4656_));
  XNOR2_X1   g03654(.A1(\A[454] ), .A2(\A[455] ), .ZN(new_n4657_));
  OAI21_X1   g03655(.A1(new_n4657_), .A2(new_n4634_), .B(new_n4600_), .ZN(new_n4658_));
  XNOR2_X1   g03656(.A1(\A[451] ), .A2(\A[452] ), .ZN(new_n4659_));
  OAI21_X1   g03657(.A1(new_n4659_), .A2(new_n4613_), .B(new_n4604_), .ZN(new_n4660_));
  AOI22_X1   g03658(.A1(new_n4627_), .A2(new_n4629_), .B1(new_n4636_), .B2(new_n4637_), .ZN(new_n4661_));
  NAND3_X1   g03659(.A1(new_n4661_), .A2(new_n4658_), .A3(new_n4660_), .ZN(new_n4662_));
  NAND2_X1   g03660(.A1(new_n4638_), .A2(new_n4633_), .ZN(new_n4663_));
  NAND2_X1   g03661(.A1(new_n4630_), .A2(new_n4631_), .ZN(new_n4664_));
  NAND2_X1   g03662(.A1(new_n4664_), .A2(new_n4663_), .ZN(new_n4665_));
  NAND2_X1   g03663(.A1(new_n4665_), .A2(new_n4662_), .ZN(new_n4666_));
  NOR2_X1    g03664(.A1(new_n4656_), .A2(new_n4666_), .ZN(new_n4667_));
  NOR2_X1    g03665(.A1(new_n4642_), .A2(new_n4667_), .ZN(new_n4668_));
  INV_X1     g03666(.I(\A[448] ), .ZN(new_n4669_));
  INV_X1     g03667(.I(\A[449] ), .ZN(new_n4670_));
  NOR2_X1    g03668(.A1(new_n4669_), .A2(new_n4670_), .ZN(new_n4671_));
  XOR2_X1    g03669(.A1(\A[448] ), .A2(\A[449] ), .Z(new_n4672_));
  AOI21_X1   g03670(.A1(new_n4672_), .A2(\A[450] ), .B(new_n4671_), .ZN(new_n4673_));
  INV_X1     g03671(.I(\A[445] ), .ZN(new_n4674_));
  INV_X1     g03672(.I(\A[446] ), .ZN(new_n4675_));
  NOR2_X1    g03673(.A1(new_n4674_), .A2(new_n4675_), .ZN(new_n4676_));
  XOR2_X1    g03674(.A1(\A[445] ), .A2(\A[446] ), .Z(new_n4677_));
  AOI21_X1   g03675(.A1(new_n4677_), .A2(\A[447] ), .B(new_n4676_), .ZN(new_n4678_));
  NAND2_X1   g03676(.A1(new_n4675_), .A2(\A[445] ), .ZN(new_n4679_));
  NAND2_X1   g03677(.A1(new_n4674_), .A2(\A[446] ), .ZN(new_n4680_));
  AOI21_X1   g03678(.A1(new_n4679_), .A2(new_n4680_), .B(\A[447] ), .ZN(new_n4681_));
  NOR2_X1    g03679(.A1(new_n4675_), .A2(\A[445] ), .ZN(new_n4682_));
  OAI21_X1   g03680(.A1(new_n4674_), .A2(\A[446] ), .B(\A[447] ), .ZN(new_n4683_));
  NOR2_X1    g03681(.A1(new_n4683_), .A2(new_n4682_), .ZN(new_n4684_));
  NAND2_X1   g03682(.A1(new_n4670_), .A2(\A[448] ), .ZN(new_n4685_));
  NAND2_X1   g03683(.A1(new_n4669_), .A2(\A[449] ), .ZN(new_n4686_));
  AOI21_X1   g03684(.A1(new_n4685_), .A2(new_n4686_), .B(\A[450] ), .ZN(new_n4687_));
  INV_X1     g03685(.I(\A[450] ), .ZN(new_n4688_));
  NOR2_X1    g03686(.A1(new_n4669_), .A2(\A[449] ), .ZN(new_n4689_));
  NOR2_X1    g03687(.A1(new_n4670_), .A2(\A[448] ), .ZN(new_n4690_));
  NOR3_X1    g03688(.A1(new_n4689_), .A2(new_n4690_), .A3(new_n4688_), .ZN(new_n4691_));
  OAI22_X1   g03689(.A1(new_n4687_), .A2(new_n4691_), .B1(new_n4681_), .B2(new_n4684_), .ZN(new_n4692_));
  NOR3_X1    g03690(.A1(new_n4692_), .A2(new_n4673_), .A3(new_n4678_), .ZN(new_n4693_));
  NOR2_X1    g03691(.A1(new_n4681_), .A2(new_n4684_), .ZN(new_n4694_));
  OAI21_X1   g03692(.A1(new_n4689_), .A2(new_n4690_), .B(new_n4688_), .ZN(new_n4695_));
  NAND3_X1   g03693(.A1(new_n4685_), .A2(new_n4686_), .A3(\A[450] ), .ZN(new_n4696_));
  NAND2_X1   g03694(.A1(new_n4695_), .A2(new_n4696_), .ZN(new_n4697_));
  NOR2_X1    g03695(.A1(new_n4697_), .A2(new_n4694_), .ZN(new_n4698_));
  NOR2_X1    g03696(.A1(new_n4674_), .A2(\A[446] ), .ZN(new_n4699_));
  NOR2_X1    g03697(.A1(new_n4699_), .A2(new_n4682_), .ZN(new_n4700_));
  NAND3_X1   g03698(.A1(new_n4679_), .A2(new_n4680_), .A3(\A[447] ), .ZN(new_n4701_));
  OAI21_X1   g03699(.A1(\A[447] ), .A2(new_n4700_), .B(new_n4701_), .ZN(new_n4702_));
  NOR2_X1    g03700(.A1(new_n4687_), .A2(new_n4691_), .ZN(new_n4703_));
  NOR2_X1    g03701(.A1(new_n4702_), .A2(new_n4703_), .ZN(new_n4704_));
  NOR2_X1    g03702(.A1(new_n4704_), .A2(new_n4698_), .ZN(new_n4705_));
  NOR2_X1    g03703(.A1(new_n4705_), .A2(new_n4693_), .ZN(new_n4706_));
  INV_X1     g03704(.I(\A[444] ), .ZN(new_n4707_));
  INV_X1     g03705(.I(\A[442] ), .ZN(new_n4708_));
  INV_X1     g03706(.I(\A[443] ), .ZN(new_n4709_));
  NOR2_X1    g03707(.A1(new_n4708_), .A2(new_n4709_), .ZN(new_n4710_));
  INV_X1     g03708(.I(new_n4710_), .ZN(new_n4711_));
  NOR2_X1    g03709(.A1(new_n4708_), .A2(\A[443] ), .ZN(new_n4712_));
  NOR2_X1    g03710(.A1(new_n4709_), .A2(\A[442] ), .ZN(new_n4713_));
  NOR2_X1    g03711(.A1(new_n4712_), .A2(new_n4713_), .ZN(new_n4714_));
  OAI21_X1   g03712(.A1(new_n4714_), .A2(new_n4707_), .B(new_n4711_), .ZN(new_n4715_));
  INV_X1     g03713(.I(\A[441] ), .ZN(new_n4716_));
  INV_X1     g03714(.I(\A[439] ), .ZN(new_n4717_));
  INV_X1     g03715(.I(\A[440] ), .ZN(new_n4718_));
  NOR2_X1    g03716(.A1(new_n4717_), .A2(new_n4718_), .ZN(new_n4719_));
  INV_X1     g03717(.I(new_n4719_), .ZN(new_n4720_));
  NOR2_X1    g03718(.A1(new_n4717_), .A2(\A[440] ), .ZN(new_n4721_));
  NOR2_X1    g03719(.A1(new_n4718_), .A2(\A[439] ), .ZN(new_n4722_));
  NOR2_X1    g03720(.A1(new_n4721_), .A2(new_n4722_), .ZN(new_n4723_));
  OAI21_X1   g03721(.A1(new_n4723_), .A2(new_n4716_), .B(new_n4720_), .ZN(new_n4724_));
  XOR2_X1    g03722(.A1(\A[439] ), .A2(\A[440] ), .Z(new_n4725_));
  NAND2_X1   g03723(.A1(new_n4725_), .A2(new_n4716_), .ZN(new_n4726_));
  NAND2_X1   g03724(.A1(new_n4718_), .A2(\A[439] ), .ZN(new_n4727_));
  NAND2_X1   g03725(.A1(new_n4717_), .A2(\A[440] ), .ZN(new_n4728_));
  NAND3_X1   g03726(.A1(new_n4727_), .A2(new_n4728_), .A3(\A[441] ), .ZN(new_n4729_));
  OAI21_X1   g03727(.A1(new_n4712_), .A2(new_n4713_), .B(new_n4707_), .ZN(new_n4730_));
  NAND2_X1   g03728(.A1(new_n4709_), .A2(\A[442] ), .ZN(new_n4731_));
  NAND2_X1   g03729(.A1(new_n4708_), .A2(\A[443] ), .ZN(new_n4732_));
  NAND3_X1   g03730(.A1(new_n4731_), .A2(new_n4732_), .A3(\A[444] ), .ZN(new_n4733_));
  AOI22_X1   g03731(.A1(new_n4726_), .A2(new_n4729_), .B1(new_n4730_), .B2(new_n4733_), .ZN(new_n4734_));
  NAND3_X1   g03732(.A1(new_n4734_), .A2(new_n4715_), .A3(new_n4724_), .ZN(new_n4735_));
  NOR3_X1    g03733(.A1(new_n4721_), .A2(new_n4722_), .A3(new_n4716_), .ZN(new_n4736_));
  AOI21_X1   g03734(.A1(new_n4716_), .A2(new_n4725_), .B(new_n4736_), .ZN(new_n4737_));
  NAND2_X1   g03735(.A1(new_n4730_), .A2(new_n4733_), .ZN(new_n4738_));
  NAND2_X1   g03736(.A1(new_n4737_), .A2(new_n4738_), .ZN(new_n4739_));
  NAND2_X1   g03737(.A1(new_n4726_), .A2(new_n4729_), .ZN(new_n4740_));
  XOR2_X1    g03738(.A1(\A[442] ), .A2(\A[443] ), .Z(new_n4741_));
  NOR3_X1    g03739(.A1(new_n4712_), .A2(new_n4713_), .A3(new_n4707_), .ZN(new_n4742_));
  AOI21_X1   g03740(.A1(new_n4707_), .A2(new_n4741_), .B(new_n4742_), .ZN(new_n4743_));
  NAND2_X1   g03741(.A1(new_n4740_), .A2(new_n4743_), .ZN(new_n4744_));
  NAND2_X1   g03742(.A1(new_n4744_), .A2(new_n4739_), .ZN(new_n4745_));
  NAND2_X1   g03743(.A1(new_n4745_), .A2(new_n4735_), .ZN(new_n4746_));
  NOR2_X1    g03744(.A1(new_n4746_), .A2(new_n4706_), .ZN(new_n4747_));
  INV_X1     g03745(.I(new_n4671_), .ZN(new_n4748_));
  NOR2_X1    g03746(.A1(new_n4689_), .A2(new_n4690_), .ZN(new_n4749_));
  OAI21_X1   g03747(.A1(new_n4749_), .A2(new_n4688_), .B(new_n4748_), .ZN(new_n4750_));
  INV_X1     g03748(.I(\A[447] ), .ZN(new_n4751_));
  INV_X1     g03749(.I(new_n4676_), .ZN(new_n4752_));
  OAI21_X1   g03750(.A1(new_n4700_), .A2(new_n4751_), .B(new_n4752_), .ZN(new_n4753_));
  NAND2_X1   g03751(.A1(new_n4677_), .A2(new_n4751_), .ZN(new_n4754_));
  AOI22_X1   g03752(.A1(new_n4754_), .A2(new_n4701_), .B1(new_n4695_), .B2(new_n4696_), .ZN(new_n4755_));
  NAND3_X1   g03753(.A1(new_n4755_), .A2(new_n4750_), .A3(new_n4753_), .ZN(new_n4756_));
  NAND2_X1   g03754(.A1(new_n4702_), .A2(new_n4703_), .ZN(new_n4757_));
  NAND2_X1   g03755(.A1(new_n4697_), .A2(new_n4694_), .ZN(new_n4758_));
  NAND2_X1   g03756(.A1(new_n4757_), .A2(new_n4758_), .ZN(new_n4759_));
  NAND2_X1   g03757(.A1(new_n4759_), .A2(new_n4756_), .ZN(new_n4760_));
  AOI21_X1   g03758(.A1(new_n4741_), .A2(\A[444] ), .B(new_n4710_), .ZN(new_n4761_));
  AOI21_X1   g03759(.A1(new_n4725_), .A2(\A[441] ), .B(new_n4719_), .ZN(new_n4762_));
  NOR4_X1    g03760(.A1(new_n4737_), .A2(new_n4743_), .A3(new_n4761_), .A4(new_n4762_), .ZN(new_n4763_));
  NOR2_X1    g03761(.A1(new_n4740_), .A2(new_n4743_), .ZN(new_n4764_));
  NOR2_X1    g03762(.A1(new_n4737_), .A2(new_n4738_), .ZN(new_n4765_));
  NOR2_X1    g03763(.A1(new_n4764_), .A2(new_n4765_), .ZN(new_n4766_));
  NOR2_X1    g03764(.A1(new_n4766_), .A2(new_n4763_), .ZN(new_n4767_));
  NOR2_X1    g03765(.A1(new_n4767_), .A2(new_n4760_), .ZN(new_n4768_));
  NOR3_X1    g03766(.A1(new_n4668_), .A2(new_n4747_), .A3(new_n4768_), .ZN(new_n4769_));
  NOR2_X1    g03767(.A1(new_n4768_), .A2(new_n4747_), .ZN(new_n4770_));
  NOR3_X1    g03768(.A1(new_n4770_), .A2(new_n4642_), .A3(new_n4667_), .ZN(new_n4771_));
  NOR2_X1    g03769(.A1(new_n4771_), .A2(new_n4769_), .ZN(new_n4772_));
  INV_X1     g03770(.I(\A[435] ), .ZN(new_n4773_));
  INV_X1     g03771(.I(\A[433] ), .ZN(new_n4774_));
  NOR2_X1    g03772(.A1(new_n4774_), .A2(\A[434] ), .ZN(new_n4775_));
  INV_X1     g03773(.I(\A[434] ), .ZN(new_n4776_));
  NOR2_X1    g03774(.A1(new_n4776_), .A2(\A[433] ), .ZN(new_n4777_));
  OAI21_X1   g03775(.A1(new_n4775_), .A2(new_n4777_), .B(new_n4773_), .ZN(new_n4778_));
  NAND2_X1   g03776(.A1(new_n4776_), .A2(\A[433] ), .ZN(new_n4779_));
  NAND2_X1   g03777(.A1(new_n4774_), .A2(\A[434] ), .ZN(new_n4780_));
  NAND3_X1   g03778(.A1(new_n4779_), .A2(new_n4780_), .A3(\A[435] ), .ZN(new_n4781_));
  NAND2_X1   g03779(.A1(new_n4778_), .A2(new_n4781_), .ZN(new_n4782_));
  INV_X1     g03780(.I(\A[438] ), .ZN(new_n4783_));
  INV_X1     g03781(.I(\A[436] ), .ZN(new_n4784_));
  NAND2_X1   g03782(.A1(new_n4784_), .A2(\A[437] ), .ZN(new_n4785_));
  XOR2_X1    g03783(.A1(\A[436] ), .A2(\A[437] ), .Z(new_n4786_));
  INV_X1     g03784(.I(\A[437] ), .ZN(new_n4787_));
  AOI21_X1   g03785(.A1(\A[436] ), .A2(new_n4787_), .B(new_n4783_), .ZN(new_n4788_));
  AOI22_X1   g03786(.A1(new_n4786_), .A2(new_n4783_), .B1(new_n4785_), .B2(new_n4788_), .ZN(new_n4789_));
  NOR2_X1    g03787(.A1(new_n4782_), .A2(new_n4789_), .ZN(new_n4790_));
  AOI21_X1   g03788(.A1(new_n4779_), .A2(new_n4780_), .B(\A[435] ), .ZN(new_n4791_));
  NOR3_X1    g03789(.A1(new_n4775_), .A2(new_n4777_), .A3(new_n4773_), .ZN(new_n4792_));
  NOR2_X1    g03790(.A1(new_n4791_), .A2(new_n4792_), .ZN(new_n4793_));
  NOR2_X1    g03791(.A1(new_n4784_), .A2(\A[437] ), .ZN(new_n4794_));
  NOR2_X1    g03792(.A1(new_n4787_), .A2(\A[436] ), .ZN(new_n4795_));
  OAI21_X1   g03793(.A1(new_n4794_), .A2(new_n4795_), .B(new_n4783_), .ZN(new_n4796_));
  NAND2_X1   g03794(.A1(new_n4788_), .A2(new_n4785_), .ZN(new_n4797_));
  NAND2_X1   g03795(.A1(new_n4797_), .A2(new_n4796_), .ZN(new_n4798_));
  NOR2_X1    g03796(.A1(new_n4793_), .A2(new_n4798_), .ZN(new_n4799_));
  NOR2_X1    g03797(.A1(new_n4799_), .A2(new_n4790_), .ZN(new_n4800_));
  NOR2_X1    g03798(.A1(new_n4784_), .A2(new_n4787_), .ZN(new_n4801_));
  AOI21_X1   g03799(.A1(new_n4786_), .A2(\A[438] ), .B(new_n4801_), .ZN(new_n4802_));
  XOR2_X1    g03800(.A1(\A[433] ), .A2(\A[434] ), .Z(new_n4803_));
  NAND2_X1   g03801(.A1(\A[433] ), .A2(\A[434] ), .ZN(new_n4804_));
  INV_X1     g03802(.I(new_n4804_), .ZN(new_n4805_));
  AOI21_X1   g03803(.A1(new_n4803_), .A2(\A[435] ), .B(new_n4805_), .ZN(new_n4806_));
  NAND2_X1   g03804(.A1(new_n4787_), .A2(\A[436] ), .ZN(new_n4807_));
  AOI21_X1   g03805(.A1(new_n4807_), .A2(new_n4785_), .B(\A[438] ), .ZN(new_n4808_));
  NOR3_X1    g03806(.A1(new_n4794_), .A2(new_n4795_), .A3(new_n4783_), .ZN(new_n4809_));
  OAI22_X1   g03807(.A1(new_n4808_), .A2(new_n4809_), .B1(new_n4791_), .B2(new_n4792_), .ZN(new_n4810_));
  NOR3_X1    g03808(.A1(new_n4810_), .A2(new_n4802_), .A3(new_n4806_), .ZN(new_n4811_));
  NOR2_X1    g03809(.A1(new_n4800_), .A2(new_n4811_), .ZN(new_n4812_));
  INV_X1     g03810(.I(\A[429] ), .ZN(new_n4813_));
  XOR2_X1    g03811(.A1(\A[427] ), .A2(\A[428] ), .Z(new_n4814_));
  INV_X1     g03812(.I(\A[428] ), .ZN(new_n4815_));
  NOR2_X1    g03813(.A1(new_n4815_), .A2(\A[427] ), .ZN(new_n4816_));
  INV_X1     g03814(.I(\A[427] ), .ZN(new_n4817_));
  OAI21_X1   g03815(.A1(new_n4817_), .A2(\A[428] ), .B(\A[429] ), .ZN(new_n4818_));
  NOR2_X1    g03816(.A1(new_n4818_), .A2(new_n4816_), .ZN(new_n4819_));
  AOI21_X1   g03817(.A1(new_n4813_), .A2(new_n4814_), .B(new_n4819_), .ZN(new_n4820_));
  INV_X1     g03818(.I(\A[432] ), .ZN(new_n4821_));
  INV_X1     g03819(.I(\A[430] ), .ZN(new_n4822_));
  NOR2_X1    g03820(.A1(new_n4822_), .A2(\A[431] ), .ZN(new_n4823_));
  INV_X1     g03821(.I(\A[431] ), .ZN(new_n4824_));
  NOR2_X1    g03822(.A1(new_n4824_), .A2(\A[430] ), .ZN(new_n4825_));
  OAI21_X1   g03823(.A1(new_n4823_), .A2(new_n4825_), .B(new_n4821_), .ZN(new_n4826_));
  NAND2_X1   g03824(.A1(new_n4822_), .A2(\A[431] ), .ZN(new_n4827_));
  AOI21_X1   g03825(.A1(\A[430] ), .A2(new_n4824_), .B(new_n4821_), .ZN(new_n4828_));
  NAND2_X1   g03826(.A1(new_n4828_), .A2(new_n4827_), .ZN(new_n4829_));
  NAND2_X1   g03827(.A1(new_n4829_), .A2(new_n4826_), .ZN(new_n4830_));
  NAND2_X1   g03828(.A1(new_n4820_), .A2(new_n4830_), .ZN(new_n4831_));
  NOR2_X1    g03829(.A1(new_n4817_), .A2(\A[428] ), .ZN(new_n4832_));
  NOR2_X1    g03830(.A1(new_n4832_), .A2(new_n4816_), .ZN(new_n4833_));
  OAI22_X1   g03831(.A1(new_n4833_), .A2(\A[429] ), .B1(new_n4816_), .B2(new_n4818_), .ZN(new_n4834_));
  XOR2_X1    g03832(.A1(\A[430] ), .A2(\A[431] ), .Z(new_n4835_));
  AOI22_X1   g03833(.A1(new_n4835_), .A2(new_n4821_), .B1(new_n4827_), .B2(new_n4828_), .ZN(new_n4836_));
  NAND2_X1   g03834(.A1(new_n4834_), .A2(new_n4836_), .ZN(new_n4837_));
  NAND2_X1   g03835(.A1(new_n4831_), .A2(new_n4837_), .ZN(new_n4838_));
  NOR2_X1    g03836(.A1(new_n4822_), .A2(new_n4824_), .ZN(new_n4839_));
  AOI21_X1   g03837(.A1(new_n4835_), .A2(\A[432] ), .B(new_n4839_), .ZN(new_n4840_));
  NOR2_X1    g03838(.A1(new_n4817_), .A2(new_n4815_), .ZN(new_n4841_));
  AOI21_X1   g03839(.A1(new_n4814_), .A2(\A[429] ), .B(new_n4841_), .ZN(new_n4842_));
  NOR4_X1    g03840(.A1(new_n4820_), .A2(new_n4836_), .A3(new_n4840_), .A4(new_n4842_), .ZN(new_n4843_));
  INV_X1     g03841(.I(new_n4843_), .ZN(new_n4844_));
  NAND2_X1   g03842(.A1(new_n4844_), .A2(new_n4838_), .ZN(new_n4845_));
  NAND2_X1   g03843(.A1(new_n4845_), .A2(new_n4812_), .ZN(new_n4846_));
  NAND2_X1   g03844(.A1(new_n4793_), .A2(new_n4798_), .ZN(new_n4847_));
  NAND2_X1   g03845(.A1(new_n4782_), .A2(new_n4789_), .ZN(new_n4848_));
  NAND2_X1   g03846(.A1(new_n4847_), .A2(new_n4848_), .ZN(new_n4849_));
  NOR2_X1    g03847(.A1(new_n4794_), .A2(new_n4795_), .ZN(new_n4850_));
  INV_X1     g03848(.I(new_n4801_), .ZN(new_n4851_));
  OAI21_X1   g03849(.A1(new_n4850_), .A2(new_n4783_), .B(new_n4851_), .ZN(new_n4852_));
  XNOR2_X1   g03850(.A1(\A[433] ), .A2(\A[434] ), .ZN(new_n4853_));
  OAI21_X1   g03851(.A1(new_n4853_), .A2(new_n4773_), .B(new_n4804_), .ZN(new_n4854_));
  AOI22_X1   g03852(.A1(new_n4796_), .A2(new_n4797_), .B1(new_n4778_), .B2(new_n4781_), .ZN(new_n4855_));
  NAND3_X1   g03853(.A1(new_n4855_), .A2(new_n4852_), .A3(new_n4854_), .ZN(new_n4856_));
  NAND2_X1   g03854(.A1(new_n4849_), .A2(new_n4856_), .ZN(new_n4857_));
  NOR2_X1    g03855(.A1(new_n4834_), .A2(new_n4836_), .ZN(new_n4858_));
  NOR2_X1    g03856(.A1(new_n4820_), .A2(new_n4830_), .ZN(new_n4859_));
  NOR2_X1    g03857(.A1(new_n4859_), .A2(new_n4858_), .ZN(new_n4860_));
  NOR2_X1    g03858(.A1(new_n4860_), .A2(new_n4843_), .ZN(new_n4861_));
  NAND2_X1   g03859(.A1(new_n4861_), .A2(new_n4857_), .ZN(new_n4862_));
  NAND2_X1   g03860(.A1(new_n4846_), .A2(new_n4862_), .ZN(new_n4863_));
  INV_X1     g03861(.I(\A[421] ), .ZN(new_n4864_));
  NAND2_X1   g03862(.A1(new_n4864_), .A2(\A[422] ), .ZN(new_n4865_));
  INV_X1     g03863(.I(\A[423] ), .ZN(new_n4866_));
  NOR2_X1    g03864(.A1(new_n4864_), .A2(\A[422] ), .ZN(new_n4867_));
  NOR2_X1    g03865(.A1(new_n4867_), .A2(new_n4866_), .ZN(new_n4868_));
  NAND2_X1   g03866(.A1(new_n4868_), .A2(new_n4865_), .ZN(new_n4869_));
  INV_X1     g03867(.I(\A[422] ), .ZN(new_n4870_));
  NOR2_X1    g03868(.A1(new_n4870_), .A2(\A[421] ), .ZN(new_n4871_));
  OAI21_X1   g03869(.A1(new_n4871_), .A2(new_n4867_), .B(new_n4866_), .ZN(new_n4872_));
  NAND2_X1   g03870(.A1(new_n4869_), .A2(new_n4872_), .ZN(new_n4873_));
  INV_X1     g03871(.I(\A[426] ), .ZN(new_n4874_));
  INV_X1     g03872(.I(\A[425] ), .ZN(new_n4875_));
  NOR2_X1    g03873(.A1(new_n4875_), .A2(\A[424] ), .ZN(new_n4876_));
  INV_X1     g03874(.I(\A[424] ), .ZN(new_n4877_));
  NOR2_X1    g03875(.A1(new_n4877_), .A2(\A[425] ), .ZN(new_n4878_));
  NOR3_X1    g03876(.A1(new_n4876_), .A2(new_n4878_), .A3(new_n4874_), .ZN(new_n4879_));
  NAND2_X1   g03877(.A1(new_n4877_), .A2(\A[425] ), .ZN(new_n4880_));
  NAND2_X1   g03878(.A1(new_n4875_), .A2(\A[424] ), .ZN(new_n4881_));
  AOI21_X1   g03879(.A1(new_n4880_), .A2(new_n4881_), .B(\A[426] ), .ZN(new_n4882_));
  NOR2_X1    g03880(.A1(new_n4882_), .A2(new_n4879_), .ZN(new_n4883_));
  NOR2_X1    g03881(.A1(new_n4873_), .A2(new_n4883_), .ZN(new_n4884_));
  NOR3_X1    g03882(.A1(new_n4871_), .A2(new_n4867_), .A3(new_n4866_), .ZN(new_n4885_));
  NAND2_X1   g03883(.A1(new_n4870_), .A2(\A[421] ), .ZN(new_n4886_));
  AOI21_X1   g03884(.A1(new_n4865_), .A2(new_n4886_), .B(\A[423] ), .ZN(new_n4887_));
  NOR2_X1    g03885(.A1(new_n4887_), .A2(new_n4885_), .ZN(new_n4888_));
  NAND3_X1   g03886(.A1(new_n4880_), .A2(new_n4881_), .A3(\A[426] ), .ZN(new_n4889_));
  OAI21_X1   g03887(.A1(new_n4876_), .A2(new_n4878_), .B(new_n4874_), .ZN(new_n4890_));
  NAND2_X1   g03888(.A1(new_n4890_), .A2(new_n4889_), .ZN(new_n4891_));
  NOR2_X1    g03889(.A1(new_n4888_), .A2(new_n4891_), .ZN(new_n4892_));
  NOR2_X1    g03890(.A1(new_n4884_), .A2(new_n4892_), .ZN(new_n4893_));
  NAND2_X1   g03891(.A1(new_n4880_), .A2(new_n4881_), .ZN(new_n4894_));
  NOR2_X1    g03892(.A1(new_n4877_), .A2(new_n4875_), .ZN(new_n4895_));
  AOI21_X1   g03893(.A1(new_n4894_), .A2(\A[426] ), .B(new_n4895_), .ZN(new_n4896_));
  XOR2_X1    g03894(.A1(\A[421] ), .A2(\A[422] ), .Z(new_n4897_));
  NOR2_X1    g03895(.A1(new_n4864_), .A2(new_n4870_), .ZN(new_n4898_));
  AOI21_X1   g03896(.A1(new_n4897_), .A2(\A[423] ), .B(new_n4898_), .ZN(new_n4899_));
  OAI22_X1   g03897(.A1(new_n4885_), .A2(new_n4887_), .B1(new_n4882_), .B2(new_n4879_), .ZN(new_n4900_));
  NOR3_X1    g03898(.A1(new_n4900_), .A2(new_n4896_), .A3(new_n4899_), .ZN(new_n4901_));
  NOR2_X1    g03899(.A1(new_n4893_), .A2(new_n4901_), .ZN(new_n4902_));
  INV_X1     g03900(.I(\A[417] ), .ZN(new_n4903_));
  INV_X1     g03901(.I(\A[415] ), .ZN(new_n4904_));
  NAND2_X1   g03902(.A1(new_n4904_), .A2(\A[416] ), .ZN(new_n4905_));
  NOR2_X1    g03903(.A1(new_n4904_), .A2(\A[416] ), .ZN(new_n4906_));
  NOR2_X1    g03904(.A1(new_n4906_), .A2(new_n4903_), .ZN(new_n4907_));
  INV_X1     g03905(.I(\A[416] ), .ZN(new_n4908_));
  NAND2_X1   g03906(.A1(new_n4908_), .A2(\A[415] ), .ZN(new_n4909_));
  NAND2_X1   g03907(.A1(new_n4905_), .A2(new_n4909_), .ZN(new_n4910_));
  AOI22_X1   g03908(.A1(new_n4910_), .A2(new_n4903_), .B1(new_n4907_), .B2(new_n4905_), .ZN(new_n4911_));
  INV_X1     g03909(.I(\A[418] ), .ZN(new_n4912_));
  NAND2_X1   g03910(.A1(new_n4912_), .A2(\A[419] ), .ZN(new_n4913_));
  INV_X1     g03911(.I(\A[419] ), .ZN(new_n4914_));
  INV_X1     g03912(.I(\A[420] ), .ZN(new_n4915_));
  AOI21_X1   g03913(.A1(\A[418] ), .A2(new_n4914_), .B(new_n4915_), .ZN(new_n4916_));
  NAND2_X1   g03914(.A1(new_n4916_), .A2(new_n4913_), .ZN(new_n4917_));
  NOR2_X1    g03915(.A1(new_n4914_), .A2(\A[418] ), .ZN(new_n4918_));
  NOR2_X1    g03916(.A1(new_n4912_), .A2(\A[419] ), .ZN(new_n4919_));
  OAI21_X1   g03917(.A1(new_n4918_), .A2(new_n4919_), .B(new_n4915_), .ZN(new_n4920_));
  NAND2_X1   g03918(.A1(new_n4917_), .A2(new_n4920_), .ZN(new_n4921_));
  NAND2_X1   g03919(.A1(new_n4911_), .A2(new_n4921_), .ZN(new_n4922_));
  NAND2_X1   g03920(.A1(new_n4907_), .A2(new_n4905_), .ZN(new_n4923_));
  NOR2_X1    g03921(.A1(new_n4908_), .A2(\A[415] ), .ZN(new_n4924_));
  OAI21_X1   g03922(.A1(new_n4924_), .A2(new_n4906_), .B(new_n4903_), .ZN(new_n4925_));
  NAND2_X1   g03923(.A1(new_n4923_), .A2(new_n4925_), .ZN(new_n4926_));
  NAND2_X1   g03924(.A1(new_n4914_), .A2(\A[418] ), .ZN(new_n4927_));
  NAND2_X1   g03925(.A1(new_n4913_), .A2(new_n4927_), .ZN(new_n4928_));
  AOI22_X1   g03926(.A1(new_n4928_), .A2(new_n4915_), .B1(new_n4913_), .B2(new_n4916_), .ZN(new_n4929_));
  NAND2_X1   g03927(.A1(new_n4926_), .A2(new_n4929_), .ZN(new_n4930_));
  NAND2_X1   g03928(.A1(new_n4930_), .A2(new_n4922_), .ZN(new_n4931_));
  NOR2_X1    g03929(.A1(new_n4918_), .A2(new_n4919_), .ZN(new_n4932_));
  NOR2_X1    g03930(.A1(new_n4912_), .A2(new_n4914_), .ZN(new_n4933_));
  INV_X1     g03931(.I(new_n4933_), .ZN(new_n4934_));
  OAI21_X1   g03932(.A1(new_n4932_), .A2(new_n4915_), .B(new_n4934_), .ZN(new_n4935_));
  NOR2_X1    g03933(.A1(new_n4924_), .A2(new_n4906_), .ZN(new_n4936_));
  NOR2_X1    g03934(.A1(new_n4904_), .A2(new_n4908_), .ZN(new_n4937_));
  INV_X1     g03935(.I(new_n4937_), .ZN(new_n4938_));
  OAI21_X1   g03936(.A1(new_n4936_), .A2(new_n4903_), .B(new_n4938_), .ZN(new_n4939_));
  AOI22_X1   g03937(.A1(new_n4923_), .A2(new_n4925_), .B1(new_n4920_), .B2(new_n4917_), .ZN(new_n4940_));
  NAND3_X1   g03938(.A1(new_n4940_), .A2(new_n4935_), .A3(new_n4939_), .ZN(new_n4941_));
  NAND2_X1   g03939(.A1(new_n4931_), .A2(new_n4941_), .ZN(new_n4942_));
  NOR2_X1    g03940(.A1(new_n4902_), .A2(new_n4942_), .ZN(new_n4943_));
  NAND2_X1   g03941(.A1(new_n4888_), .A2(new_n4891_), .ZN(new_n4944_));
  NAND2_X1   g03942(.A1(new_n4873_), .A2(new_n4883_), .ZN(new_n4945_));
  NAND2_X1   g03943(.A1(new_n4945_), .A2(new_n4944_), .ZN(new_n4946_));
  NOR2_X1    g03944(.A1(new_n4876_), .A2(new_n4878_), .ZN(new_n4947_));
  INV_X1     g03945(.I(new_n4895_), .ZN(new_n4948_));
  OAI21_X1   g03946(.A1(new_n4947_), .A2(new_n4874_), .B(new_n4948_), .ZN(new_n4949_));
  NOR2_X1    g03947(.A1(new_n4871_), .A2(new_n4867_), .ZN(new_n4950_));
  INV_X1     g03948(.I(new_n4898_), .ZN(new_n4951_));
  OAI21_X1   g03949(.A1(new_n4950_), .A2(new_n4866_), .B(new_n4951_), .ZN(new_n4952_));
  AOI22_X1   g03950(.A1(new_n4869_), .A2(new_n4872_), .B1(new_n4890_), .B2(new_n4889_), .ZN(new_n4953_));
  NAND3_X1   g03951(.A1(new_n4953_), .A2(new_n4949_), .A3(new_n4952_), .ZN(new_n4954_));
  NAND2_X1   g03952(.A1(new_n4946_), .A2(new_n4954_), .ZN(new_n4955_));
  XOR2_X1    g03953(.A1(new_n4911_), .A2(new_n4921_), .Z(new_n4956_));
  AOI21_X1   g03954(.A1(new_n4928_), .A2(\A[420] ), .B(new_n4933_), .ZN(new_n4957_));
  AOI21_X1   g03955(.A1(new_n4910_), .A2(\A[417] ), .B(new_n4937_), .ZN(new_n4958_));
  NOR4_X1    g03956(.A1(new_n4911_), .A2(new_n4929_), .A3(new_n4957_), .A4(new_n4958_), .ZN(new_n4959_));
  NOR2_X1    g03957(.A1(new_n4956_), .A2(new_n4959_), .ZN(new_n4960_));
  NOR2_X1    g03958(.A1(new_n4960_), .A2(new_n4955_), .ZN(new_n4961_));
  NOR2_X1    g03959(.A1(new_n4961_), .A2(new_n4943_), .ZN(new_n4962_));
  NAND2_X1   g03960(.A1(new_n4962_), .A2(new_n4863_), .ZN(new_n4963_));
  NOR2_X1    g03961(.A1(new_n4861_), .A2(new_n4857_), .ZN(new_n4964_));
  NOR2_X1    g03962(.A1(new_n4845_), .A2(new_n4812_), .ZN(new_n4965_));
  NOR2_X1    g03963(.A1(new_n4965_), .A2(new_n4964_), .ZN(new_n4966_));
  NAND2_X1   g03964(.A1(new_n4960_), .A2(new_n4955_), .ZN(new_n4967_));
  NAND2_X1   g03965(.A1(new_n4902_), .A2(new_n4942_), .ZN(new_n4968_));
  NAND2_X1   g03966(.A1(new_n4967_), .A2(new_n4968_), .ZN(new_n4969_));
  NAND2_X1   g03967(.A1(new_n4969_), .A2(new_n4966_), .ZN(new_n4970_));
  NAND2_X1   g03968(.A1(new_n4963_), .A2(new_n4970_), .ZN(new_n4971_));
  XNOR2_X1   g03969(.A1(new_n4772_), .A2(new_n4971_), .ZN(new_n4972_));
  XNOR2_X1   g03970(.A1(new_n4562_), .A2(new_n4972_), .ZN(new_n4973_));
  INV_X1     g03971(.I(\A[366] ), .ZN(new_n4974_));
  NAND2_X1   g03972(.A1(\A[364] ), .A2(\A[365] ), .ZN(new_n4975_));
  XNOR2_X1   g03973(.A1(\A[364] ), .A2(\A[365] ), .ZN(new_n4976_));
  OAI21_X1   g03974(.A1(new_n4976_), .A2(new_n4974_), .B(new_n4975_), .ZN(new_n4977_));
  INV_X1     g03975(.I(\A[363] ), .ZN(new_n4978_));
  NAND2_X1   g03976(.A1(\A[361] ), .A2(\A[362] ), .ZN(new_n4979_));
  XNOR2_X1   g03977(.A1(\A[361] ), .A2(\A[362] ), .ZN(new_n4980_));
  OAI21_X1   g03978(.A1(new_n4980_), .A2(new_n4978_), .B(new_n4979_), .ZN(new_n4981_));
  INV_X1     g03979(.I(\A[361] ), .ZN(new_n4982_));
  NOR2_X1    g03980(.A1(new_n4982_), .A2(\A[362] ), .ZN(new_n4983_));
  INV_X1     g03981(.I(\A[362] ), .ZN(new_n4984_));
  NOR2_X1    g03982(.A1(new_n4984_), .A2(\A[361] ), .ZN(new_n4985_));
  OAI21_X1   g03983(.A1(new_n4983_), .A2(new_n4985_), .B(new_n4978_), .ZN(new_n4986_));
  NAND2_X1   g03984(.A1(new_n4984_), .A2(\A[361] ), .ZN(new_n4987_));
  NAND2_X1   g03985(.A1(new_n4982_), .A2(\A[362] ), .ZN(new_n4988_));
  NAND3_X1   g03986(.A1(new_n4987_), .A2(new_n4988_), .A3(\A[363] ), .ZN(new_n4989_));
  INV_X1     g03987(.I(\A[364] ), .ZN(new_n4990_));
  NOR2_X1    g03988(.A1(new_n4990_), .A2(\A[365] ), .ZN(new_n4991_));
  INV_X1     g03989(.I(\A[365] ), .ZN(new_n4992_));
  NOR2_X1    g03990(.A1(new_n4992_), .A2(\A[364] ), .ZN(new_n4993_));
  OAI21_X1   g03991(.A1(new_n4991_), .A2(new_n4993_), .B(new_n4974_), .ZN(new_n4994_));
  NAND2_X1   g03992(.A1(new_n4992_), .A2(\A[364] ), .ZN(new_n4995_));
  NAND2_X1   g03993(.A1(new_n4990_), .A2(\A[365] ), .ZN(new_n4996_));
  NAND3_X1   g03994(.A1(new_n4995_), .A2(new_n4996_), .A3(\A[366] ), .ZN(new_n4997_));
  AOI22_X1   g03995(.A1(new_n4986_), .A2(new_n4989_), .B1(new_n4994_), .B2(new_n4997_), .ZN(new_n4998_));
  NAND3_X1   g03996(.A1(new_n4998_), .A2(new_n4977_), .A3(new_n4981_), .ZN(new_n4999_));
  NAND2_X1   g03997(.A1(new_n4986_), .A2(new_n4989_), .ZN(new_n5000_));
  XOR2_X1    g03998(.A1(\A[364] ), .A2(\A[365] ), .Z(new_n5001_));
  AOI21_X1   g03999(.A1(\A[364] ), .A2(new_n4992_), .B(new_n4974_), .ZN(new_n5002_));
  AOI22_X1   g04000(.A1(new_n5001_), .A2(new_n4974_), .B1(new_n4996_), .B2(new_n5002_), .ZN(new_n5003_));
  NAND2_X1   g04001(.A1(new_n5000_), .A2(new_n5003_), .ZN(new_n5004_));
  AOI21_X1   g04002(.A1(new_n4987_), .A2(new_n4988_), .B(\A[363] ), .ZN(new_n5005_));
  NOR3_X1    g04003(.A1(new_n4983_), .A2(new_n4985_), .A3(new_n4978_), .ZN(new_n5006_));
  NOR2_X1    g04004(.A1(new_n5005_), .A2(new_n5006_), .ZN(new_n5007_));
  NAND2_X1   g04005(.A1(new_n4994_), .A2(new_n4997_), .ZN(new_n5008_));
  NAND2_X1   g04006(.A1(new_n5007_), .A2(new_n5008_), .ZN(new_n5009_));
  NAND2_X1   g04007(.A1(new_n5009_), .A2(new_n5004_), .ZN(new_n5010_));
  NAND2_X1   g04008(.A1(new_n5010_), .A2(new_n4999_), .ZN(new_n5011_));
  NAND2_X1   g04009(.A1(\A[358] ), .A2(\A[359] ), .ZN(new_n5012_));
  INV_X1     g04010(.I(new_n5012_), .ZN(new_n5013_));
  XOR2_X1    g04011(.A1(\A[358] ), .A2(\A[359] ), .Z(new_n5014_));
  AOI21_X1   g04012(.A1(new_n5014_), .A2(\A[360] ), .B(new_n5013_), .ZN(new_n5015_));
  NAND2_X1   g04013(.A1(\A[355] ), .A2(\A[356] ), .ZN(new_n5016_));
  INV_X1     g04014(.I(new_n5016_), .ZN(new_n5017_));
  XOR2_X1    g04015(.A1(\A[355] ), .A2(\A[356] ), .Z(new_n5018_));
  AOI21_X1   g04016(.A1(new_n5018_), .A2(\A[357] ), .B(new_n5017_), .ZN(new_n5019_));
  INV_X1     g04017(.I(\A[356] ), .ZN(new_n5020_));
  NAND2_X1   g04018(.A1(new_n5020_), .A2(\A[355] ), .ZN(new_n5021_));
  INV_X1     g04019(.I(\A[355] ), .ZN(new_n5022_));
  NAND2_X1   g04020(.A1(new_n5022_), .A2(\A[356] ), .ZN(new_n5023_));
  AOI21_X1   g04021(.A1(new_n5021_), .A2(new_n5023_), .B(\A[357] ), .ZN(new_n5024_));
  INV_X1     g04022(.I(\A[357] ), .ZN(new_n5025_));
  NOR2_X1    g04023(.A1(new_n5022_), .A2(\A[356] ), .ZN(new_n5026_));
  NOR2_X1    g04024(.A1(new_n5020_), .A2(\A[355] ), .ZN(new_n5027_));
  NOR3_X1    g04025(.A1(new_n5026_), .A2(new_n5027_), .A3(new_n5025_), .ZN(new_n5028_));
  INV_X1     g04026(.I(\A[359] ), .ZN(new_n5029_));
  NAND2_X1   g04027(.A1(new_n5029_), .A2(\A[358] ), .ZN(new_n5030_));
  INV_X1     g04028(.I(\A[358] ), .ZN(new_n5031_));
  NAND2_X1   g04029(.A1(new_n5031_), .A2(\A[359] ), .ZN(new_n5032_));
  AOI21_X1   g04030(.A1(new_n5030_), .A2(new_n5032_), .B(\A[360] ), .ZN(new_n5033_));
  INV_X1     g04031(.I(\A[360] ), .ZN(new_n5034_));
  NOR2_X1    g04032(.A1(new_n5031_), .A2(\A[359] ), .ZN(new_n5035_));
  NOR2_X1    g04033(.A1(new_n5029_), .A2(\A[358] ), .ZN(new_n5036_));
  NOR3_X1    g04034(.A1(new_n5035_), .A2(new_n5036_), .A3(new_n5034_), .ZN(new_n5037_));
  OAI22_X1   g04035(.A1(new_n5024_), .A2(new_n5028_), .B1(new_n5033_), .B2(new_n5037_), .ZN(new_n5038_));
  NOR3_X1    g04036(.A1(new_n5038_), .A2(new_n5015_), .A3(new_n5019_), .ZN(new_n5039_));
  XNOR2_X1   g04037(.A1(\A[355] ), .A2(\A[356] ), .ZN(new_n5040_));
  NAND2_X1   g04038(.A1(new_n5021_), .A2(\A[357] ), .ZN(new_n5041_));
  OAI22_X1   g04039(.A1(\A[357] ), .A2(new_n5040_), .B1(new_n5041_), .B2(new_n5027_), .ZN(new_n5042_));
  NOR2_X1    g04040(.A1(new_n5033_), .A2(new_n5037_), .ZN(new_n5043_));
  NOR2_X1    g04041(.A1(new_n5042_), .A2(new_n5043_), .ZN(new_n5044_));
  AOI21_X1   g04042(.A1(\A[355] ), .A2(new_n5020_), .B(new_n5025_), .ZN(new_n5045_));
  AOI22_X1   g04043(.A1(new_n5018_), .A2(new_n5025_), .B1(new_n5023_), .B2(new_n5045_), .ZN(new_n5046_));
  NOR2_X1    g04044(.A1(new_n5035_), .A2(new_n5036_), .ZN(new_n5047_));
  OAI21_X1   g04045(.A1(new_n5031_), .A2(\A[359] ), .B(\A[360] ), .ZN(new_n5048_));
  OAI22_X1   g04046(.A1(new_n5047_), .A2(\A[360] ), .B1(new_n5036_), .B2(new_n5048_), .ZN(new_n5049_));
  NOR2_X1    g04047(.A1(new_n5049_), .A2(new_n5046_), .ZN(new_n5050_));
  NOR2_X1    g04048(.A1(new_n5044_), .A2(new_n5050_), .ZN(new_n5051_));
  NOR2_X1    g04049(.A1(new_n5051_), .A2(new_n5039_), .ZN(new_n5052_));
  NOR2_X1    g04050(.A1(new_n5052_), .A2(new_n5011_), .ZN(new_n5053_));
  INV_X1     g04051(.I(new_n4975_), .ZN(new_n5054_));
  AOI21_X1   g04052(.A1(new_n5001_), .A2(\A[366] ), .B(new_n5054_), .ZN(new_n5055_));
  INV_X1     g04053(.I(new_n4979_), .ZN(new_n5056_));
  XOR2_X1    g04054(.A1(\A[361] ), .A2(\A[362] ), .Z(new_n5057_));
  AOI21_X1   g04055(.A1(new_n5057_), .A2(\A[363] ), .B(new_n5056_), .ZN(new_n5058_));
  AOI21_X1   g04056(.A1(new_n4995_), .A2(new_n4996_), .B(\A[366] ), .ZN(new_n5059_));
  NOR3_X1    g04057(.A1(new_n4991_), .A2(new_n4993_), .A3(new_n4974_), .ZN(new_n5060_));
  OAI22_X1   g04058(.A1(new_n5005_), .A2(new_n5006_), .B1(new_n5059_), .B2(new_n5060_), .ZN(new_n5061_));
  NOR3_X1    g04059(.A1(new_n5061_), .A2(new_n5055_), .A3(new_n5058_), .ZN(new_n5062_));
  NOR2_X1    g04060(.A1(new_n5007_), .A2(new_n5008_), .ZN(new_n5063_));
  NOR2_X1    g04061(.A1(new_n5000_), .A2(new_n5003_), .ZN(new_n5064_));
  NOR2_X1    g04062(.A1(new_n5063_), .A2(new_n5064_), .ZN(new_n5065_));
  NOR2_X1    g04063(.A1(new_n5065_), .A2(new_n5062_), .ZN(new_n5066_));
  OAI21_X1   g04064(.A1(new_n5047_), .A2(new_n5034_), .B(new_n5012_), .ZN(new_n5067_));
  OAI21_X1   g04065(.A1(new_n5040_), .A2(new_n5025_), .B(new_n5016_), .ZN(new_n5068_));
  NAND4_X1   g04066(.A1(new_n5042_), .A2(new_n5049_), .A3(new_n5067_), .A4(new_n5068_), .ZN(new_n5069_));
  NAND2_X1   g04067(.A1(new_n5049_), .A2(new_n5046_), .ZN(new_n5070_));
  NAND2_X1   g04068(.A1(new_n5042_), .A2(new_n5043_), .ZN(new_n5071_));
  NAND2_X1   g04069(.A1(new_n5071_), .A2(new_n5070_), .ZN(new_n5072_));
  NAND2_X1   g04070(.A1(new_n5072_), .A2(new_n5069_), .ZN(new_n5073_));
  NOR2_X1    g04071(.A1(new_n5073_), .A2(new_n5066_), .ZN(new_n5074_));
  NOR2_X1    g04072(.A1(new_n5074_), .A2(new_n5053_), .ZN(new_n5075_));
  INV_X1     g04073(.I(\A[354] ), .ZN(new_n5076_));
  INV_X1     g04074(.I(\A[352] ), .ZN(new_n5077_));
  INV_X1     g04075(.I(\A[353] ), .ZN(new_n5078_));
  NOR2_X1    g04076(.A1(new_n5077_), .A2(new_n5078_), .ZN(new_n5079_));
  INV_X1     g04077(.I(new_n5079_), .ZN(new_n5080_));
  NOR2_X1    g04078(.A1(new_n5077_), .A2(\A[353] ), .ZN(new_n5081_));
  NOR2_X1    g04079(.A1(new_n5078_), .A2(\A[352] ), .ZN(new_n5082_));
  NOR2_X1    g04080(.A1(new_n5081_), .A2(new_n5082_), .ZN(new_n5083_));
  OAI21_X1   g04081(.A1(new_n5083_), .A2(new_n5076_), .B(new_n5080_), .ZN(new_n5084_));
  INV_X1     g04082(.I(\A[351] ), .ZN(new_n5085_));
  INV_X1     g04083(.I(\A[349] ), .ZN(new_n5086_));
  INV_X1     g04084(.I(\A[350] ), .ZN(new_n5087_));
  NOR2_X1    g04085(.A1(new_n5086_), .A2(new_n5087_), .ZN(new_n5088_));
  INV_X1     g04086(.I(new_n5088_), .ZN(new_n5089_));
  NOR2_X1    g04087(.A1(new_n5086_), .A2(\A[350] ), .ZN(new_n5090_));
  NOR2_X1    g04088(.A1(new_n5087_), .A2(\A[349] ), .ZN(new_n5091_));
  NOR2_X1    g04089(.A1(new_n5090_), .A2(new_n5091_), .ZN(new_n5092_));
  OAI21_X1   g04090(.A1(new_n5092_), .A2(new_n5085_), .B(new_n5089_), .ZN(new_n5093_));
  XOR2_X1    g04091(.A1(\A[349] ), .A2(\A[350] ), .Z(new_n5094_));
  NAND2_X1   g04092(.A1(new_n5094_), .A2(new_n5085_), .ZN(new_n5095_));
  NAND2_X1   g04093(.A1(new_n5087_), .A2(\A[349] ), .ZN(new_n5096_));
  NAND2_X1   g04094(.A1(new_n5086_), .A2(\A[350] ), .ZN(new_n5097_));
  NAND3_X1   g04095(.A1(new_n5096_), .A2(new_n5097_), .A3(\A[351] ), .ZN(new_n5098_));
  OAI21_X1   g04096(.A1(new_n5081_), .A2(new_n5082_), .B(new_n5076_), .ZN(new_n5099_));
  NAND2_X1   g04097(.A1(new_n5077_), .A2(\A[353] ), .ZN(new_n5100_));
  AOI21_X1   g04098(.A1(\A[352] ), .A2(new_n5078_), .B(new_n5076_), .ZN(new_n5101_));
  NAND2_X1   g04099(.A1(new_n5101_), .A2(new_n5100_), .ZN(new_n5102_));
  AOI22_X1   g04100(.A1(new_n5095_), .A2(new_n5098_), .B1(new_n5099_), .B2(new_n5102_), .ZN(new_n5103_));
  NAND3_X1   g04101(.A1(new_n5103_), .A2(new_n5084_), .A3(new_n5093_), .ZN(new_n5104_));
  OAI21_X1   g04102(.A1(new_n5086_), .A2(\A[350] ), .B(\A[351] ), .ZN(new_n5105_));
  OAI22_X1   g04103(.A1(new_n5092_), .A2(\A[351] ), .B1(new_n5091_), .B2(new_n5105_), .ZN(new_n5106_));
  XOR2_X1    g04104(.A1(\A[352] ), .A2(\A[353] ), .Z(new_n5107_));
  AOI22_X1   g04105(.A1(new_n5107_), .A2(new_n5076_), .B1(new_n5100_), .B2(new_n5101_), .ZN(new_n5108_));
  NAND2_X1   g04106(.A1(new_n5106_), .A2(new_n5108_), .ZN(new_n5109_));
  AOI21_X1   g04107(.A1(new_n5096_), .A2(new_n5097_), .B(\A[351] ), .ZN(new_n5110_));
  NOR2_X1    g04108(.A1(new_n5105_), .A2(new_n5091_), .ZN(new_n5111_));
  NOR2_X1    g04109(.A1(new_n5110_), .A2(new_n5111_), .ZN(new_n5112_));
  NAND2_X1   g04110(.A1(new_n5102_), .A2(new_n5099_), .ZN(new_n5113_));
  NAND2_X1   g04111(.A1(new_n5113_), .A2(new_n5112_), .ZN(new_n5114_));
  NAND2_X1   g04112(.A1(new_n5109_), .A2(new_n5114_), .ZN(new_n5115_));
  NAND2_X1   g04113(.A1(new_n5115_), .A2(new_n5104_), .ZN(new_n5116_));
  INV_X1     g04114(.I(\A[348] ), .ZN(new_n5117_));
  INV_X1     g04115(.I(\A[346] ), .ZN(new_n5118_));
  INV_X1     g04116(.I(\A[347] ), .ZN(new_n5119_));
  NOR2_X1    g04117(.A1(new_n5118_), .A2(new_n5119_), .ZN(new_n5120_));
  INV_X1     g04118(.I(new_n5120_), .ZN(new_n5121_));
  NOR2_X1    g04119(.A1(new_n5118_), .A2(\A[347] ), .ZN(new_n5122_));
  NOR2_X1    g04120(.A1(new_n5119_), .A2(\A[346] ), .ZN(new_n5123_));
  NOR2_X1    g04121(.A1(new_n5122_), .A2(new_n5123_), .ZN(new_n5124_));
  OAI21_X1   g04122(.A1(new_n5124_), .A2(new_n5117_), .B(new_n5121_), .ZN(new_n5125_));
  INV_X1     g04123(.I(\A[345] ), .ZN(new_n5126_));
  NAND2_X1   g04124(.A1(\A[343] ), .A2(\A[344] ), .ZN(new_n5127_));
  XNOR2_X1   g04125(.A1(\A[343] ), .A2(\A[344] ), .ZN(new_n5128_));
  OAI21_X1   g04126(.A1(new_n5128_), .A2(new_n5126_), .B(new_n5127_), .ZN(new_n5129_));
  INV_X1     g04127(.I(\A[344] ), .ZN(new_n5130_));
  NOR2_X1    g04128(.A1(new_n5130_), .A2(\A[343] ), .ZN(new_n5131_));
  INV_X1     g04129(.I(\A[343] ), .ZN(new_n5132_));
  OAI21_X1   g04130(.A1(new_n5132_), .A2(\A[344] ), .B(\A[345] ), .ZN(new_n5133_));
  OAI22_X1   g04131(.A1(new_n5128_), .A2(\A[345] ), .B1(new_n5131_), .B2(new_n5133_), .ZN(new_n5134_));
  OAI21_X1   g04132(.A1(new_n5118_), .A2(\A[347] ), .B(\A[348] ), .ZN(new_n5135_));
  OAI22_X1   g04133(.A1(new_n5124_), .A2(\A[348] ), .B1(new_n5123_), .B2(new_n5135_), .ZN(new_n5136_));
  NAND4_X1   g04134(.A1(new_n5136_), .A2(new_n5125_), .A3(new_n5134_), .A4(new_n5129_), .ZN(new_n5137_));
  INV_X1     g04135(.I(new_n5137_), .ZN(new_n5138_));
  NAND2_X1   g04136(.A1(new_n5119_), .A2(\A[346] ), .ZN(new_n5139_));
  NAND2_X1   g04137(.A1(new_n5118_), .A2(\A[347] ), .ZN(new_n5140_));
  AOI21_X1   g04138(.A1(new_n5139_), .A2(new_n5140_), .B(\A[348] ), .ZN(new_n5141_));
  NOR3_X1    g04139(.A1(new_n5122_), .A2(new_n5123_), .A3(new_n5117_), .ZN(new_n5142_));
  NOR2_X1    g04140(.A1(new_n5141_), .A2(new_n5142_), .ZN(new_n5143_));
  NOR2_X1    g04141(.A1(new_n5143_), .A2(new_n5134_), .ZN(new_n5144_));
  XOR2_X1    g04142(.A1(\A[343] ), .A2(\A[344] ), .Z(new_n5145_));
  NOR2_X1    g04143(.A1(new_n5133_), .A2(new_n5131_), .ZN(new_n5146_));
  AOI21_X1   g04144(.A1(new_n5126_), .A2(new_n5145_), .B(new_n5146_), .ZN(new_n5147_));
  NOR2_X1    g04145(.A1(new_n5147_), .A2(new_n5136_), .ZN(new_n5148_));
  NOR2_X1    g04146(.A1(new_n5148_), .A2(new_n5144_), .ZN(new_n5149_));
  NOR2_X1    g04147(.A1(new_n5149_), .A2(new_n5138_), .ZN(new_n5150_));
  NAND2_X1   g04148(.A1(new_n5150_), .A2(new_n5116_), .ZN(new_n5151_));
  AOI21_X1   g04149(.A1(new_n5107_), .A2(\A[354] ), .B(new_n5079_), .ZN(new_n5152_));
  AOI21_X1   g04150(.A1(new_n5094_), .A2(\A[351] ), .B(new_n5088_), .ZN(new_n5153_));
  NAND2_X1   g04151(.A1(new_n5078_), .A2(\A[352] ), .ZN(new_n5154_));
  AOI21_X1   g04152(.A1(new_n5154_), .A2(new_n5100_), .B(\A[354] ), .ZN(new_n5155_));
  NOR3_X1    g04153(.A1(new_n5081_), .A2(new_n5082_), .A3(new_n5076_), .ZN(new_n5156_));
  OAI22_X1   g04154(.A1(new_n5155_), .A2(new_n5156_), .B1(new_n5110_), .B2(new_n5111_), .ZN(new_n5157_));
  NOR3_X1    g04155(.A1(new_n5157_), .A2(new_n5152_), .A3(new_n5153_), .ZN(new_n5158_));
  NOR2_X1    g04156(.A1(new_n5113_), .A2(new_n5112_), .ZN(new_n5159_));
  NOR2_X1    g04157(.A1(new_n5106_), .A2(new_n5108_), .ZN(new_n5160_));
  NOR2_X1    g04158(.A1(new_n5160_), .A2(new_n5159_), .ZN(new_n5161_));
  NOR2_X1    g04159(.A1(new_n5161_), .A2(new_n5158_), .ZN(new_n5162_));
  NAND2_X1   g04160(.A1(new_n5147_), .A2(new_n5136_), .ZN(new_n5163_));
  NAND2_X1   g04161(.A1(new_n5143_), .A2(new_n5134_), .ZN(new_n5164_));
  NAND2_X1   g04162(.A1(new_n5163_), .A2(new_n5164_), .ZN(new_n5165_));
  NAND2_X1   g04163(.A1(new_n5165_), .A2(new_n5137_), .ZN(new_n5166_));
  NAND2_X1   g04164(.A1(new_n5162_), .A2(new_n5166_), .ZN(new_n5167_));
  NAND2_X1   g04165(.A1(new_n5151_), .A2(new_n5167_), .ZN(new_n5168_));
  NOR2_X1    g04166(.A1(new_n5168_), .A2(new_n5075_), .ZN(new_n5169_));
  NAND2_X1   g04167(.A1(new_n5073_), .A2(new_n5066_), .ZN(new_n5170_));
  NAND2_X1   g04168(.A1(new_n5052_), .A2(new_n5011_), .ZN(new_n5171_));
  NAND2_X1   g04169(.A1(new_n5170_), .A2(new_n5171_), .ZN(new_n5172_));
  NOR2_X1    g04170(.A1(new_n5162_), .A2(new_n5166_), .ZN(new_n5173_));
  NOR2_X1    g04171(.A1(new_n5150_), .A2(new_n5116_), .ZN(new_n5174_));
  NOR2_X1    g04172(.A1(new_n5174_), .A2(new_n5173_), .ZN(new_n5175_));
  NOR2_X1    g04173(.A1(new_n5175_), .A2(new_n5172_), .ZN(new_n5176_));
  NOR2_X1    g04174(.A1(new_n5169_), .A2(new_n5176_), .ZN(new_n5177_));
  INV_X1     g04175(.I(\A[337] ), .ZN(new_n5178_));
  NOR2_X1    g04176(.A1(new_n5178_), .A2(\A[338] ), .ZN(new_n5179_));
  INV_X1     g04177(.I(\A[338] ), .ZN(new_n5180_));
  NOR2_X1    g04178(.A1(new_n5180_), .A2(\A[337] ), .ZN(new_n5181_));
  NOR2_X1    g04179(.A1(new_n5179_), .A2(new_n5181_), .ZN(new_n5182_));
  NAND2_X1   g04180(.A1(new_n5180_), .A2(\A[337] ), .ZN(new_n5183_));
  NAND2_X1   g04181(.A1(new_n5178_), .A2(\A[338] ), .ZN(new_n5184_));
  NAND3_X1   g04182(.A1(new_n5183_), .A2(new_n5184_), .A3(\A[339] ), .ZN(new_n5185_));
  OAI21_X1   g04183(.A1(\A[339] ), .A2(new_n5182_), .B(new_n5185_), .ZN(new_n5186_));
  INV_X1     g04184(.I(\A[341] ), .ZN(new_n5187_));
  NAND2_X1   g04185(.A1(new_n5187_), .A2(\A[340] ), .ZN(new_n5188_));
  INV_X1     g04186(.I(\A[340] ), .ZN(new_n5189_));
  NAND2_X1   g04187(.A1(new_n5189_), .A2(\A[341] ), .ZN(new_n5190_));
  AOI21_X1   g04188(.A1(new_n5188_), .A2(new_n5190_), .B(\A[342] ), .ZN(new_n5191_));
  INV_X1     g04189(.I(\A[342] ), .ZN(new_n5192_));
  NOR2_X1    g04190(.A1(new_n5189_), .A2(\A[341] ), .ZN(new_n5193_));
  NOR2_X1    g04191(.A1(new_n5187_), .A2(\A[340] ), .ZN(new_n5194_));
  NOR3_X1    g04192(.A1(new_n5193_), .A2(new_n5194_), .A3(new_n5192_), .ZN(new_n5195_));
  NOR2_X1    g04193(.A1(new_n5191_), .A2(new_n5195_), .ZN(new_n5196_));
  NOR2_X1    g04194(.A1(new_n5186_), .A2(new_n5196_), .ZN(new_n5197_));
  AOI21_X1   g04195(.A1(new_n5183_), .A2(new_n5184_), .B(\A[339] ), .ZN(new_n5198_));
  OAI21_X1   g04196(.A1(new_n5178_), .A2(\A[338] ), .B(\A[339] ), .ZN(new_n5199_));
  NOR2_X1    g04197(.A1(new_n5199_), .A2(new_n5181_), .ZN(new_n5200_));
  NOR2_X1    g04198(.A1(new_n5198_), .A2(new_n5200_), .ZN(new_n5201_));
  OAI21_X1   g04199(.A1(new_n5193_), .A2(new_n5194_), .B(new_n5192_), .ZN(new_n5202_));
  NAND3_X1   g04200(.A1(new_n5188_), .A2(new_n5190_), .A3(\A[342] ), .ZN(new_n5203_));
  NAND2_X1   g04201(.A1(new_n5202_), .A2(new_n5203_), .ZN(new_n5204_));
  NOR2_X1    g04202(.A1(new_n5204_), .A2(new_n5201_), .ZN(new_n5205_));
  NOR2_X1    g04203(.A1(new_n5197_), .A2(new_n5205_), .ZN(new_n5206_));
  XOR2_X1    g04204(.A1(\A[340] ), .A2(\A[341] ), .Z(new_n5207_));
  NOR2_X1    g04205(.A1(new_n5189_), .A2(new_n5187_), .ZN(new_n5208_));
  AOI21_X1   g04206(.A1(new_n5207_), .A2(\A[342] ), .B(new_n5208_), .ZN(new_n5209_));
  XOR2_X1    g04207(.A1(\A[337] ), .A2(\A[338] ), .Z(new_n5210_));
  NAND2_X1   g04208(.A1(\A[337] ), .A2(\A[338] ), .ZN(new_n5211_));
  INV_X1     g04209(.I(new_n5211_), .ZN(new_n5212_));
  AOI21_X1   g04210(.A1(new_n5210_), .A2(\A[339] ), .B(new_n5212_), .ZN(new_n5213_));
  OAI22_X1   g04211(.A1(new_n5191_), .A2(new_n5195_), .B1(new_n5198_), .B2(new_n5200_), .ZN(new_n5214_));
  NOR3_X1    g04212(.A1(new_n5214_), .A2(new_n5209_), .A3(new_n5213_), .ZN(new_n5215_));
  NOR2_X1    g04213(.A1(new_n5206_), .A2(new_n5215_), .ZN(new_n5216_));
  INV_X1     g04214(.I(\A[332] ), .ZN(new_n5217_));
  NAND2_X1   g04215(.A1(new_n5217_), .A2(\A[331] ), .ZN(new_n5218_));
  INV_X1     g04216(.I(\A[331] ), .ZN(new_n5219_));
  NAND2_X1   g04217(.A1(new_n5219_), .A2(\A[332] ), .ZN(new_n5220_));
  AOI21_X1   g04218(.A1(new_n5218_), .A2(new_n5220_), .B(\A[333] ), .ZN(new_n5221_));
  INV_X1     g04219(.I(\A[333] ), .ZN(new_n5222_));
  NOR2_X1    g04220(.A1(new_n5219_), .A2(\A[332] ), .ZN(new_n5223_));
  NOR2_X1    g04221(.A1(new_n5217_), .A2(\A[331] ), .ZN(new_n5224_));
  NOR3_X1    g04222(.A1(new_n5223_), .A2(new_n5224_), .A3(new_n5222_), .ZN(new_n5225_));
  NOR2_X1    g04223(.A1(new_n5221_), .A2(new_n5225_), .ZN(new_n5226_));
  INV_X1     g04224(.I(\A[336] ), .ZN(new_n5227_));
  INV_X1     g04225(.I(\A[334] ), .ZN(new_n5228_));
  NOR2_X1    g04226(.A1(new_n5228_), .A2(\A[335] ), .ZN(new_n5229_));
  INV_X1     g04227(.I(\A[335] ), .ZN(new_n5230_));
  NOR2_X1    g04228(.A1(new_n5230_), .A2(\A[334] ), .ZN(new_n5231_));
  OAI21_X1   g04229(.A1(new_n5229_), .A2(new_n5231_), .B(new_n5227_), .ZN(new_n5232_));
  NAND2_X1   g04230(.A1(new_n5228_), .A2(\A[335] ), .ZN(new_n5233_));
  AOI21_X1   g04231(.A1(\A[334] ), .A2(new_n5230_), .B(new_n5227_), .ZN(new_n5234_));
  NAND2_X1   g04232(.A1(new_n5234_), .A2(new_n5233_), .ZN(new_n5235_));
  NAND2_X1   g04233(.A1(new_n5235_), .A2(new_n5232_), .ZN(new_n5236_));
  NAND2_X1   g04234(.A1(new_n5226_), .A2(new_n5236_), .ZN(new_n5237_));
  XOR2_X1    g04235(.A1(\A[331] ), .A2(\A[332] ), .Z(new_n5238_));
  NAND2_X1   g04236(.A1(new_n5238_), .A2(new_n5222_), .ZN(new_n5239_));
  NAND3_X1   g04237(.A1(new_n5218_), .A2(new_n5220_), .A3(\A[333] ), .ZN(new_n5240_));
  NAND2_X1   g04238(.A1(new_n5239_), .A2(new_n5240_), .ZN(new_n5241_));
  NAND2_X1   g04239(.A1(new_n5230_), .A2(\A[334] ), .ZN(new_n5242_));
  AOI21_X1   g04240(.A1(new_n5242_), .A2(new_n5233_), .B(\A[336] ), .ZN(new_n5243_));
  NOR3_X1    g04241(.A1(new_n5229_), .A2(new_n5231_), .A3(new_n5227_), .ZN(new_n5244_));
  NOR2_X1    g04242(.A1(new_n5243_), .A2(new_n5244_), .ZN(new_n5245_));
  NAND2_X1   g04243(.A1(new_n5241_), .A2(new_n5245_), .ZN(new_n5246_));
  NAND2_X1   g04244(.A1(new_n5246_), .A2(new_n5237_), .ZN(new_n5247_));
  XOR2_X1    g04245(.A1(\A[334] ), .A2(\A[335] ), .Z(new_n5248_));
  NAND2_X1   g04246(.A1(\A[334] ), .A2(\A[335] ), .ZN(new_n5249_));
  INV_X1     g04247(.I(new_n5249_), .ZN(new_n5250_));
  AOI21_X1   g04248(.A1(new_n5248_), .A2(\A[336] ), .B(new_n5250_), .ZN(new_n5251_));
  NOR2_X1    g04249(.A1(new_n5219_), .A2(new_n5217_), .ZN(new_n5252_));
  AOI21_X1   g04250(.A1(new_n5238_), .A2(\A[333] ), .B(new_n5252_), .ZN(new_n5253_));
  OAI22_X1   g04251(.A1(new_n5221_), .A2(new_n5225_), .B1(new_n5243_), .B2(new_n5244_), .ZN(new_n5254_));
  NOR3_X1    g04252(.A1(new_n5254_), .A2(new_n5251_), .A3(new_n5253_), .ZN(new_n5255_));
  INV_X1     g04253(.I(new_n5255_), .ZN(new_n5256_));
  NAND2_X1   g04254(.A1(new_n5256_), .A2(new_n5247_), .ZN(new_n5257_));
  NAND2_X1   g04255(.A1(new_n5257_), .A2(new_n5216_), .ZN(new_n5258_));
  NAND2_X1   g04256(.A1(new_n5204_), .A2(new_n5201_), .ZN(new_n5259_));
  NAND2_X1   g04257(.A1(new_n5186_), .A2(new_n5196_), .ZN(new_n5260_));
  NAND2_X1   g04258(.A1(new_n5260_), .A2(new_n5259_), .ZN(new_n5261_));
  NOR2_X1    g04259(.A1(new_n5193_), .A2(new_n5194_), .ZN(new_n5262_));
  INV_X1     g04260(.I(new_n5208_), .ZN(new_n5263_));
  OAI21_X1   g04261(.A1(new_n5262_), .A2(new_n5192_), .B(new_n5263_), .ZN(new_n5264_));
  INV_X1     g04262(.I(\A[339] ), .ZN(new_n5265_));
  OAI21_X1   g04263(.A1(new_n5182_), .A2(new_n5265_), .B(new_n5211_), .ZN(new_n5266_));
  NAND2_X1   g04264(.A1(new_n5210_), .A2(new_n5265_), .ZN(new_n5267_));
  AOI22_X1   g04265(.A1(new_n5267_), .A2(new_n5185_), .B1(new_n5202_), .B2(new_n5203_), .ZN(new_n5268_));
  NAND3_X1   g04266(.A1(new_n5268_), .A2(new_n5264_), .A3(new_n5266_), .ZN(new_n5269_));
  NAND2_X1   g04267(.A1(new_n5261_), .A2(new_n5269_), .ZN(new_n5270_));
  NOR2_X1    g04268(.A1(new_n5241_), .A2(new_n5245_), .ZN(new_n5271_));
  NOR2_X1    g04269(.A1(new_n5226_), .A2(new_n5236_), .ZN(new_n5272_));
  NOR2_X1    g04270(.A1(new_n5271_), .A2(new_n5272_), .ZN(new_n5273_));
  NOR2_X1    g04271(.A1(new_n5273_), .A2(new_n5255_), .ZN(new_n5274_));
  NAND2_X1   g04272(.A1(new_n5274_), .A2(new_n5270_), .ZN(new_n5275_));
  NAND2_X1   g04273(.A1(new_n5258_), .A2(new_n5275_), .ZN(new_n5276_));
  INV_X1     g04274(.I(\A[327] ), .ZN(new_n5277_));
  INV_X1     g04275(.I(\A[326] ), .ZN(new_n5278_));
  NOR2_X1    g04276(.A1(new_n5278_), .A2(\A[325] ), .ZN(new_n5279_));
  INV_X1     g04277(.I(\A[325] ), .ZN(new_n5280_));
  NOR2_X1    g04278(.A1(new_n5280_), .A2(\A[326] ), .ZN(new_n5281_));
  NOR3_X1    g04279(.A1(new_n5279_), .A2(new_n5281_), .A3(new_n5277_), .ZN(new_n5282_));
  NAND2_X1   g04280(.A1(new_n5280_), .A2(\A[326] ), .ZN(new_n5283_));
  NAND2_X1   g04281(.A1(new_n5278_), .A2(\A[325] ), .ZN(new_n5284_));
  AOI21_X1   g04282(.A1(new_n5283_), .A2(new_n5284_), .B(\A[327] ), .ZN(new_n5285_));
  NOR2_X1    g04283(.A1(new_n5285_), .A2(new_n5282_), .ZN(new_n5286_));
  INV_X1     g04284(.I(\A[328] ), .ZN(new_n5287_));
  NAND2_X1   g04285(.A1(new_n5287_), .A2(\A[329] ), .ZN(new_n5288_));
  INV_X1     g04286(.I(\A[329] ), .ZN(new_n5289_));
  NAND2_X1   g04287(.A1(new_n5289_), .A2(\A[328] ), .ZN(new_n5290_));
  NAND3_X1   g04288(.A1(new_n5288_), .A2(new_n5290_), .A3(\A[330] ), .ZN(new_n5291_));
  INV_X1     g04289(.I(\A[330] ), .ZN(new_n5292_));
  NOR2_X1    g04290(.A1(new_n5289_), .A2(\A[328] ), .ZN(new_n5293_));
  NOR2_X1    g04291(.A1(new_n5287_), .A2(\A[329] ), .ZN(new_n5294_));
  OAI21_X1   g04292(.A1(new_n5293_), .A2(new_n5294_), .B(new_n5292_), .ZN(new_n5295_));
  NAND2_X1   g04293(.A1(new_n5295_), .A2(new_n5291_), .ZN(new_n5296_));
  NAND2_X1   g04294(.A1(new_n5286_), .A2(new_n5296_), .ZN(new_n5297_));
  INV_X1     g04295(.I(new_n5282_), .ZN(new_n5298_));
  OAI21_X1   g04296(.A1(new_n5279_), .A2(new_n5281_), .B(new_n5277_), .ZN(new_n5299_));
  NAND2_X1   g04297(.A1(new_n5298_), .A2(new_n5299_), .ZN(new_n5300_));
  NOR3_X1    g04298(.A1(new_n5293_), .A2(new_n5294_), .A3(new_n5292_), .ZN(new_n5301_));
  AOI21_X1   g04299(.A1(new_n5288_), .A2(new_n5290_), .B(\A[330] ), .ZN(new_n5302_));
  NOR2_X1    g04300(.A1(new_n5302_), .A2(new_n5301_), .ZN(new_n5303_));
  NAND2_X1   g04301(.A1(new_n5300_), .A2(new_n5303_), .ZN(new_n5304_));
  NAND2_X1   g04302(.A1(new_n5304_), .A2(new_n5297_), .ZN(new_n5305_));
  NAND2_X1   g04303(.A1(new_n5288_), .A2(new_n5290_), .ZN(new_n5306_));
  NOR2_X1    g04304(.A1(new_n5287_), .A2(new_n5289_), .ZN(new_n5307_));
  AOI21_X1   g04305(.A1(new_n5306_), .A2(\A[330] ), .B(new_n5307_), .ZN(new_n5308_));
  NAND2_X1   g04306(.A1(new_n5283_), .A2(new_n5284_), .ZN(new_n5309_));
  NOR2_X1    g04307(.A1(new_n5280_), .A2(new_n5278_), .ZN(new_n5310_));
  AOI21_X1   g04308(.A1(new_n5309_), .A2(\A[327] ), .B(new_n5310_), .ZN(new_n5311_));
  OAI22_X1   g04309(.A1(new_n5282_), .A2(new_n5285_), .B1(new_n5302_), .B2(new_n5301_), .ZN(new_n5312_));
  NOR3_X1    g04310(.A1(new_n5312_), .A2(new_n5308_), .A3(new_n5311_), .ZN(new_n5313_));
  INV_X1     g04311(.I(new_n5313_), .ZN(new_n5314_));
  NAND2_X1   g04312(.A1(new_n5314_), .A2(new_n5305_), .ZN(new_n5315_));
  INV_X1     g04313(.I(\A[321] ), .ZN(new_n5316_));
  INV_X1     g04314(.I(\A[320] ), .ZN(new_n5317_));
  NOR2_X1    g04315(.A1(new_n5317_), .A2(\A[319] ), .ZN(new_n5318_));
  INV_X1     g04316(.I(\A[319] ), .ZN(new_n5319_));
  NOR2_X1    g04317(.A1(new_n5319_), .A2(\A[320] ), .ZN(new_n5320_));
  NOR3_X1    g04318(.A1(new_n5318_), .A2(new_n5320_), .A3(new_n5316_), .ZN(new_n5321_));
  NAND2_X1   g04319(.A1(new_n5319_), .A2(\A[320] ), .ZN(new_n5322_));
  NAND2_X1   g04320(.A1(new_n5317_), .A2(\A[319] ), .ZN(new_n5323_));
  AOI21_X1   g04321(.A1(new_n5322_), .A2(new_n5323_), .B(\A[321] ), .ZN(new_n5324_));
  NOR2_X1    g04322(.A1(new_n5324_), .A2(new_n5321_), .ZN(new_n5325_));
  INV_X1     g04323(.I(\A[323] ), .ZN(new_n5326_));
  NOR2_X1    g04324(.A1(new_n5326_), .A2(\A[322] ), .ZN(new_n5327_));
  NAND2_X1   g04325(.A1(new_n5326_), .A2(\A[322] ), .ZN(new_n5328_));
  NAND2_X1   g04326(.A1(new_n5328_), .A2(\A[324] ), .ZN(new_n5329_));
  INV_X1     g04327(.I(\A[322] ), .ZN(new_n5330_));
  NOR2_X1    g04328(.A1(new_n5330_), .A2(\A[323] ), .ZN(new_n5331_));
  NOR2_X1    g04329(.A1(new_n5327_), .A2(new_n5331_), .ZN(new_n5332_));
  OAI22_X1   g04330(.A1(new_n5332_), .A2(\A[324] ), .B1(new_n5329_), .B2(new_n5327_), .ZN(new_n5333_));
  XOR2_X1    g04331(.A1(new_n5333_), .A2(new_n5325_), .Z(new_n5334_));
  XOR2_X1    g04332(.A1(\A[322] ), .A2(\A[323] ), .Z(new_n5335_));
  NOR2_X1    g04333(.A1(new_n5330_), .A2(new_n5326_), .ZN(new_n5336_));
  AOI21_X1   g04334(.A1(new_n5335_), .A2(\A[324] ), .B(new_n5336_), .ZN(new_n5337_));
  NAND2_X1   g04335(.A1(new_n5322_), .A2(new_n5323_), .ZN(new_n5338_));
  NOR2_X1    g04336(.A1(new_n5319_), .A2(new_n5317_), .ZN(new_n5339_));
  AOI21_X1   g04337(.A1(new_n5338_), .A2(\A[321] ), .B(new_n5339_), .ZN(new_n5340_));
  INV_X1     g04338(.I(\A[324] ), .ZN(new_n5341_));
  NOR3_X1    g04339(.A1(new_n5327_), .A2(new_n5331_), .A3(new_n5341_), .ZN(new_n5342_));
  NAND2_X1   g04340(.A1(new_n5330_), .A2(\A[323] ), .ZN(new_n5343_));
  AOI21_X1   g04341(.A1(new_n5343_), .A2(new_n5328_), .B(\A[324] ), .ZN(new_n5344_));
  OAI22_X1   g04342(.A1(new_n5321_), .A2(new_n5324_), .B1(new_n5344_), .B2(new_n5342_), .ZN(new_n5345_));
  NOR3_X1    g04343(.A1(new_n5345_), .A2(new_n5337_), .A3(new_n5340_), .ZN(new_n5346_));
  NOR2_X1    g04344(.A1(new_n5334_), .A2(new_n5346_), .ZN(new_n5347_));
  NAND2_X1   g04345(.A1(new_n5315_), .A2(new_n5347_), .ZN(new_n5348_));
  NOR2_X1    g04346(.A1(new_n5300_), .A2(new_n5303_), .ZN(new_n5349_));
  NOR2_X1    g04347(.A1(new_n5286_), .A2(new_n5296_), .ZN(new_n5350_));
  NOR2_X1    g04348(.A1(new_n5349_), .A2(new_n5350_), .ZN(new_n5351_));
  NOR2_X1    g04349(.A1(new_n5351_), .A2(new_n5313_), .ZN(new_n5352_));
  NAND2_X1   g04350(.A1(new_n5333_), .A2(new_n5325_), .ZN(new_n5353_));
  OR2_X2     g04351(.A1(new_n5324_), .A2(new_n5321_), .Z(new_n5354_));
  NOR2_X1    g04352(.A1(new_n5344_), .A2(new_n5342_), .ZN(new_n5355_));
  NAND2_X1   g04353(.A1(new_n5354_), .A2(new_n5355_), .ZN(new_n5356_));
  NAND2_X1   g04354(.A1(new_n5356_), .A2(new_n5353_), .ZN(new_n5357_));
  INV_X1     g04355(.I(new_n5336_), .ZN(new_n5358_));
  OAI21_X1   g04356(.A1(new_n5332_), .A2(new_n5341_), .B(new_n5358_), .ZN(new_n5359_));
  NOR2_X1    g04357(.A1(new_n5318_), .A2(new_n5320_), .ZN(new_n5360_));
  INV_X1     g04358(.I(new_n5339_), .ZN(new_n5361_));
  OAI21_X1   g04359(.A1(new_n5360_), .A2(new_n5316_), .B(new_n5361_), .ZN(new_n5362_));
  NAND4_X1   g04360(.A1(new_n5354_), .A2(new_n5333_), .A3(new_n5359_), .A4(new_n5362_), .ZN(new_n5363_));
  NAND2_X1   g04361(.A1(new_n5357_), .A2(new_n5363_), .ZN(new_n5364_));
  NAND2_X1   g04362(.A1(new_n5352_), .A2(new_n5364_), .ZN(new_n5365_));
  NAND3_X1   g04363(.A1(new_n5276_), .A2(new_n5348_), .A3(new_n5365_), .ZN(new_n5366_));
  NAND2_X1   g04364(.A1(new_n5348_), .A2(new_n5365_), .ZN(new_n5367_));
  NAND3_X1   g04365(.A1(new_n5367_), .A2(new_n5258_), .A3(new_n5275_), .ZN(new_n5368_));
  NAND2_X1   g04366(.A1(new_n5368_), .A2(new_n5366_), .ZN(new_n5369_));
  XOR2_X1    g04367(.A1(new_n5369_), .A2(new_n5177_), .Z(new_n5370_));
  INV_X1     g04368(.I(\A[315] ), .ZN(new_n5371_));
  INV_X1     g04369(.I(\A[314] ), .ZN(new_n5372_));
  NOR2_X1    g04370(.A1(new_n5372_), .A2(\A[313] ), .ZN(new_n5373_));
  INV_X1     g04371(.I(\A[313] ), .ZN(new_n5374_));
  NOR2_X1    g04372(.A1(new_n5374_), .A2(\A[314] ), .ZN(new_n5375_));
  NOR3_X1    g04373(.A1(new_n5373_), .A2(new_n5375_), .A3(new_n5371_), .ZN(new_n5376_));
  NAND2_X1   g04374(.A1(new_n5374_), .A2(\A[314] ), .ZN(new_n5377_));
  NAND2_X1   g04375(.A1(new_n5372_), .A2(\A[313] ), .ZN(new_n5378_));
  AOI21_X1   g04376(.A1(new_n5377_), .A2(new_n5378_), .B(\A[315] ), .ZN(new_n5379_));
  NOR2_X1    g04377(.A1(new_n5379_), .A2(new_n5376_), .ZN(new_n5380_));
  INV_X1     g04378(.I(\A[316] ), .ZN(new_n5381_));
  NAND2_X1   g04379(.A1(new_n5381_), .A2(\A[317] ), .ZN(new_n5382_));
  INV_X1     g04380(.I(\A[317] ), .ZN(new_n5383_));
  NAND2_X1   g04381(.A1(new_n5383_), .A2(\A[316] ), .ZN(new_n5384_));
  NAND3_X1   g04382(.A1(new_n5382_), .A2(new_n5384_), .A3(\A[318] ), .ZN(new_n5385_));
  INV_X1     g04383(.I(\A[318] ), .ZN(new_n5386_));
  NOR2_X1    g04384(.A1(new_n5383_), .A2(\A[316] ), .ZN(new_n5387_));
  NOR2_X1    g04385(.A1(new_n5381_), .A2(\A[317] ), .ZN(new_n5388_));
  OAI21_X1   g04386(.A1(new_n5387_), .A2(new_n5388_), .B(new_n5386_), .ZN(new_n5389_));
  NAND2_X1   g04387(.A1(new_n5389_), .A2(new_n5385_), .ZN(new_n5390_));
  NAND2_X1   g04388(.A1(new_n5380_), .A2(new_n5390_), .ZN(new_n5391_));
  AOI21_X1   g04389(.A1(\A[313] ), .A2(new_n5372_), .B(new_n5371_), .ZN(new_n5392_));
  NAND2_X1   g04390(.A1(new_n5392_), .A2(new_n5377_), .ZN(new_n5393_));
  OAI21_X1   g04391(.A1(new_n5373_), .A2(new_n5375_), .B(new_n5371_), .ZN(new_n5394_));
  NAND2_X1   g04392(.A1(new_n5393_), .A2(new_n5394_), .ZN(new_n5395_));
  NOR3_X1    g04393(.A1(new_n5387_), .A2(new_n5388_), .A3(new_n5386_), .ZN(new_n5396_));
  AOI21_X1   g04394(.A1(new_n5382_), .A2(new_n5384_), .B(\A[318] ), .ZN(new_n5397_));
  NOR2_X1    g04395(.A1(new_n5397_), .A2(new_n5396_), .ZN(new_n5398_));
  NAND2_X1   g04396(.A1(new_n5398_), .A2(new_n5395_), .ZN(new_n5399_));
  NAND2_X1   g04397(.A1(new_n5399_), .A2(new_n5391_), .ZN(new_n5400_));
  NOR2_X1    g04398(.A1(new_n5387_), .A2(new_n5388_), .ZN(new_n5401_));
  NOR2_X1    g04399(.A1(new_n5381_), .A2(new_n5383_), .ZN(new_n5402_));
  INV_X1     g04400(.I(new_n5402_), .ZN(new_n5403_));
  OAI21_X1   g04401(.A1(new_n5401_), .A2(new_n5386_), .B(new_n5403_), .ZN(new_n5404_));
  NOR2_X1    g04402(.A1(new_n5373_), .A2(new_n5375_), .ZN(new_n5405_));
  NOR2_X1    g04403(.A1(new_n5374_), .A2(new_n5372_), .ZN(new_n5406_));
  INV_X1     g04404(.I(new_n5406_), .ZN(new_n5407_));
  OAI21_X1   g04405(.A1(new_n5405_), .A2(new_n5371_), .B(new_n5407_), .ZN(new_n5408_));
  AOI22_X1   g04406(.A1(new_n5393_), .A2(new_n5394_), .B1(new_n5389_), .B2(new_n5385_), .ZN(new_n5409_));
  NAND3_X1   g04407(.A1(new_n5409_), .A2(new_n5404_), .A3(new_n5408_), .ZN(new_n5410_));
  NAND2_X1   g04408(.A1(new_n5400_), .A2(new_n5410_), .ZN(new_n5411_));
  INV_X1     g04409(.I(\A[307] ), .ZN(new_n5412_));
  NAND2_X1   g04410(.A1(new_n5412_), .A2(\A[308] ), .ZN(new_n5413_));
  INV_X1     g04411(.I(\A[308] ), .ZN(new_n5414_));
  INV_X1     g04412(.I(\A[309] ), .ZN(new_n5415_));
  AOI21_X1   g04413(.A1(\A[307] ), .A2(new_n5414_), .B(new_n5415_), .ZN(new_n5416_));
  NAND2_X1   g04414(.A1(new_n5416_), .A2(new_n5413_), .ZN(new_n5417_));
  NOR2_X1    g04415(.A1(new_n5414_), .A2(\A[307] ), .ZN(new_n5418_));
  NOR2_X1    g04416(.A1(new_n5412_), .A2(\A[308] ), .ZN(new_n5419_));
  OAI21_X1   g04417(.A1(new_n5418_), .A2(new_n5419_), .B(new_n5415_), .ZN(new_n5420_));
  NAND2_X1   g04418(.A1(new_n5417_), .A2(new_n5420_), .ZN(new_n5421_));
  INV_X1     g04419(.I(\A[312] ), .ZN(new_n5422_));
  INV_X1     g04420(.I(\A[310] ), .ZN(new_n5423_));
  NAND2_X1   g04421(.A1(new_n5423_), .A2(\A[311] ), .ZN(new_n5424_));
  INV_X1     g04422(.I(\A[311] ), .ZN(new_n5425_));
  AOI21_X1   g04423(.A1(\A[310] ), .A2(new_n5425_), .B(new_n5422_), .ZN(new_n5426_));
  XOR2_X1    g04424(.A1(\A[310] ), .A2(\A[311] ), .Z(new_n5427_));
  AOI22_X1   g04425(.A1(new_n5427_), .A2(new_n5422_), .B1(new_n5424_), .B2(new_n5426_), .ZN(new_n5428_));
  XOR2_X1    g04426(.A1(new_n5421_), .A2(new_n5428_), .Z(new_n5429_));
  NAND2_X1   g04427(.A1(new_n5414_), .A2(\A[307] ), .ZN(new_n5430_));
  NAND2_X1   g04428(.A1(new_n5413_), .A2(new_n5430_), .ZN(new_n5431_));
  AOI22_X1   g04429(.A1(new_n5431_), .A2(new_n5415_), .B1(new_n5413_), .B2(new_n5416_), .ZN(new_n5432_));
  NOR2_X1    g04430(.A1(new_n5423_), .A2(new_n5425_), .ZN(new_n5433_));
  AOI21_X1   g04431(.A1(new_n5427_), .A2(\A[312] ), .B(new_n5433_), .ZN(new_n5434_));
  NOR2_X1    g04432(.A1(new_n5412_), .A2(new_n5414_), .ZN(new_n5435_));
  AOI21_X1   g04433(.A1(new_n5431_), .A2(\A[309] ), .B(new_n5435_), .ZN(new_n5436_));
  NOR4_X1    g04434(.A1(new_n5432_), .A2(new_n5436_), .A3(new_n5428_), .A4(new_n5434_), .ZN(new_n5437_));
  NOR2_X1    g04435(.A1(new_n5429_), .A2(new_n5437_), .ZN(new_n5438_));
  NAND2_X1   g04436(.A1(new_n5438_), .A2(new_n5411_), .ZN(new_n5439_));
  NOR2_X1    g04437(.A1(new_n5398_), .A2(new_n5395_), .ZN(new_n5440_));
  NOR2_X1    g04438(.A1(new_n5380_), .A2(new_n5390_), .ZN(new_n5441_));
  NOR2_X1    g04439(.A1(new_n5440_), .A2(new_n5441_), .ZN(new_n5442_));
  NAND2_X1   g04440(.A1(new_n5382_), .A2(new_n5384_), .ZN(new_n5443_));
  AOI21_X1   g04441(.A1(new_n5443_), .A2(\A[318] ), .B(new_n5402_), .ZN(new_n5444_));
  XOR2_X1    g04442(.A1(\A[313] ), .A2(\A[314] ), .Z(new_n5445_));
  AOI21_X1   g04443(.A1(new_n5445_), .A2(\A[315] ), .B(new_n5406_), .ZN(new_n5446_));
  OAI22_X1   g04444(.A1(new_n5376_), .A2(new_n5379_), .B1(new_n5397_), .B2(new_n5396_), .ZN(new_n5447_));
  NOR3_X1    g04445(.A1(new_n5447_), .A2(new_n5444_), .A3(new_n5446_), .ZN(new_n5448_));
  NOR2_X1    g04446(.A1(new_n5442_), .A2(new_n5448_), .ZN(new_n5449_));
  NAND2_X1   g04447(.A1(new_n5426_), .A2(new_n5424_), .ZN(new_n5450_));
  NOR2_X1    g04448(.A1(new_n5425_), .A2(\A[310] ), .ZN(new_n5451_));
  NOR2_X1    g04449(.A1(new_n5423_), .A2(\A[311] ), .ZN(new_n5452_));
  OAI21_X1   g04450(.A1(new_n5451_), .A2(new_n5452_), .B(new_n5422_), .ZN(new_n5453_));
  NAND2_X1   g04451(.A1(new_n5450_), .A2(new_n5453_), .ZN(new_n5454_));
  NAND2_X1   g04452(.A1(new_n5432_), .A2(new_n5454_), .ZN(new_n5455_));
  NAND2_X1   g04453(.A1(new_n5421_), .A2(new_n5428_), .ZN(new_n5456_));
  NAND2_X1   g04454(.A1(new_n5455_), .A2(new_n5456_), .ZN(new_n5457_));
  NOR2_X1    g04455(.A1(new_n5451_), .A2(new_n5452_), .ZN(new_n5458_));
  INV_X1     g04456(.I(new_n5433_), .ZN(new_n5459_));
  OAI21_X1   g04457(.A1(new_n5458_), .A2(new_n5422_), .B(new_n5459_), .ZN(new_n5460_));
  NOR2_X1    g04458(.A1(new_n5418_), .A2(new_n5419_), .ZN(new_n5461_));
  INV_X1     g04459(.I(new_n5435_), .ZN(new_n5462_));
  OAI21_X1   g04460(.A1(new_n5461_), .A2(new_n5415_), .B(new_n5462_), .ZN(new_n5463_));
  AOI22_X1   g04461(.A1(new_n5417_), .A2(new_n5420_), .B1(new_n5450_), .B2(new_n5453_), .ZN(new_n5464_));
  NAND3_X1   g04462(.A1(new_n5464_), .A2(new_n5460_), .A3(new_n5463_), .ZN(new_n5465_));
  NAND2_X1   g04463(.A1(new_n5457_), .A2(new_n5465_), .ZN(new_n5466_));
  NAND2_X1   g04464(.A1(new_n5449_), .A2(new_n5466_), .ZN(new_n5467_));
  INV_X1     g04465(.I(\A[303] ), .ZN(new_n5468_));
  INV_X1     g04466(.I(\A[302] ), .ZN(new_n5469_));
  NOR2_X1    g04467(.A1(new_n5469_), .A2(\A[301] ), .ZN(new_n5470_));
  INV_X1     g04468(.I(\A[301] ), .ZN(new_n5471_));
  NOR2_X1    g04469(.A1(new_n5471_), .A2(\A[302] ), .ZN(new_n5472_));
  NOR3_X1    g04470(.A1(new_n5470_), .A2(new_n5472_), .A3(new_n5468_), .ZN(new_n5473_));
  NAND2_X1   g04471(.A1(new_n5471_), .A2(\A[302] ), .ZN(new_n5474_));
  NAND2_X1   g04472(.A1(new_n5469_), .A2(\A[301] ), .ZN(new_n5475_));
  AOI21_X1   g04473(.A1(new_n5474_), .A2(new_n5475_), .B(\A[303] ), .ZN(new_n5476_));
  NOR2_X1    g04474(.A1(new_n5476_), .A2(new_n5473_), .ZN(new_n5477_));
  INV_X1     g04475(.I(\A[304] ), .ZN(new_n5478_));
  NAND2_X1   g04476(.A1(new_n5478_), .A2(\A[305] ), .ZN(new_n5479_));
  INV_X1     g04477(.I(\A[305] ), .ZN(new_n5480_));
  NAND2_X1   g04478(.A1(new_n5480_), .A2(\A[304] ), .ZN(new_n5481_));
  NAND3_X1   g04479(.A1(new_n5479_), .A2(new_n5481_), .A3(\A[306] ), .ZN(new_n5482_));
  INV_X1     g04480(.I(\A[306] ), .ZN(new_n5483_));
  NOR2_X1    g04481(.A1(new_n5480_), .A2(\A[304] ), .ZN(new_n5484_));
  NOR2_X1    g04482(.A1(new_n5478_), .A2(\A[305] ), .ZN(new_n5485_));
  OAI21_X1   g04483(.A1(new_n5484_), .A2(new_n5485_), .B(new_n5483_), .ZN(new_n5486_));
  NAND2_X1   g04484(.A1(new_n5486_), .A2(new_n5482_), .ZN(new_n5487_));
  NAND2_X1   g04485(.A1(new_n5477_), .A2(new_n5487_), .ZN(new_n5488_));
  AOI21_X1   g04486(.A1(\A[301] ), .A2(new_n5469_), .B(new_n5468_), .ZN(new_n5489_));
  NAND2_X1   g04487(.A1(new_n5489_), .A2(new_n5474_), .ZN(new_n5490_));
  OAI21_X1   g04488(.A1(new_n5470_), .A2(new_n5472_), .B(new_n5468_), .ZN(new_n5491_));
  NAND2_X1   g04489(.A1(new_n5490_), .A2(new_n5491_), .ZN(new_n5492_));
  NOR3_X1    g04490(.A1(new_n5484_), .A2(new_n5485_), .A3(new_n5483_), .ZN(new_n5493_));
  AOI21_X1   g04491(.A1(new_n5479_), .A2(new_n5481_), .B(\A[306] ), .ZN(new_n5494_));
  NOR2_X1    g04492(.A1(new_n5494_), .A2(new_n5493_), .ZN(new_n5495_));
  NAND2_X1   g04493(.A1(new_n5495_), .A2(new_n5492_), .ZN(new_n5496_));
  NAND2_X1   g04494(.A1(new_n5496_), .A2(new_n5488_), .ZN(new_n5497_));
  NOR2_X1    g04495(.A1(new_n5484_), .A2(new_n5485_), .ZN(new_n5498_));
  NOR2_X1    g04496(.A1(new_n5478_), .A2(new_n5480_), .ZN(new_n5499_));
  INV_X1     g04497(.I(new_n5499_), .ZN(new_n5500_));
  OAI21_X1   g04498(.A1(new_n5498_), .A2(new_n5483_), .B(new_n5500_), .ZN(new_n5501_));
  NOR2_X1    g04499(.A1(new_n5470_), .A2(new_n5472_), .ZN(new_n5502_));
  NOR2_X1    g04500(.A1(new_n5471_), .A2(new_n5469_), .ZN(new_n5503_));
  INV_X1     g04501(.I(new_n5503_), .ZN(new_n5504_));
  OAI21_X1   g04502(.A1(new_n5502_), .A2(new_n5468_), .B(new_n5504_), .ZN(new_n5505_));
  AOI22_X1   g04503(.A1(new_n5490_), .A2(new_n5491_), .B1(new_n5486_), .B2(new_n5482_), .ZN(new_n5506_));
  NAND3_X1   g04504(.A1(new_n5506_), .A2(new_n5501_), .A3(new_n5505_), .ZN(new_n5507_));
  NAND2_X1   g04505(.A1(new_n5497_), .A2(new_n5507_), .ZN(new_n5508_));
  INV_X1     g04506(.I(\A[295] ), .ZN(new_n5509_));
  NAND2_X1   g04507(.A1(new_n5509_), .A2(\A[296] ), .ZN(new_n5510_));
  INV_X1     g04508(.I(\A[296] ), .ZN(new_n5511_));
  INV_X1     g04509(.I(\A[297] ), .ZN(new_n5512_));
  AOI21_X1   g04510(.A1(\A[295] ), .A2(new_n5511_), .B(new_n5512_), .ZN(new_n5513_));
  NAND2_X1   g04511(.A1(new_n5513_), .A2(new_n5510_), .ZN(new_n5514_));
  NOR2_X1    g04512(.A1(new_n5511_), .A2(\A[295] ), .ZN(new_n5515_));
  NOR2_X1    g04513(.A1(new_n5509_), .A2(\A[296] ), .ZN(new_n5516_));
  OAI21_X1   g04514(.A1(new_n5515_), .A2(new_n5516_), .B(new_n5512_), .ZN(new_n5517_));
  NAND2_X1   g04515(.A1(new_n5514_), .A2(new_n5517_), .ZN(new_n5518_));
  INV_X1     g04516(.I(\A[300] ), .ZN(new_n5519_));
  INV_X1     g04517(.I(\A[299] ), .ZN(new_n5520_));
  NOR2_X1    g04518(.A1(new_n5520_), .A2(\A[298] ), .ZN(new_n5521_));
  INV_X1     g04519(.I(\A[298] ), .ZN(new_n5522_));
  NOR2_X1    g04520(.A1(new_n5522_), .A2(\A[299] ), .ZN(new_n5523_));
  NOR3_X1    g04521(.A1(new_n5521_), .A2(new_n5523_), .A3(new_n5519_), .ZN(new_n5524_));
  NAND2_X1   g04522(.A1(new_n5522_), .A2(\A[299] ), .ZN(new_n5525_));
  NAND2_X1   g04523(.A1(new_n5520_), .A2(\A[298] ), .ZN(new_n5526_));
  AOI21_X1   g04524(.A1(new_n5525_), .A2(new_n5526_), .B(\A[300] ), .ZN(new_n5527_));
  NOR2_X1    g04525(.A1(new_n5527_), .A2(new_n5524_), .ZN(new_n5528_));
  NOR2_X1    g04526(.A1(new_n5528_), .A2(new_n5518_), .ZN(new_n5529_));
  NOR3_X1    g04527(.A1(new_n5515_), .A2(new_n5516_), .A3(new_n5512_), .ZN(new_n5530_));
  NAND2_X1   g04528(.A1(new_n5511_), .A2(\A[295] ), .ZN(new_n5531_));
  AOI21_X1   g04529(.A1(new_n5510_), .A2(new_n5531_), .B(\A[297] ), .ZN(new_n5532_));
  NOR2_X1    g04530(.A1(new_n5532_), .A2(new_n5530_), .ZN(new_n5533_));
  NAND3_X1   g04531(.A1(new_n5525_), .A2(new_n5526_), .A3(\A[300] ), .ZN(new_n5534_));
  OAI21_X1   g04532(.A1(new_n5521_), .A2(new_n5523_), .B(new_n5519_), .ZN(new_n5535_));
  NAND2_X1   g04533(.A1(new_n5535_), .A2(new_n5534_), .ZN(new_n5536_));
  NOR2_X1    g04534(.A1(new_n5533_), .A2(new_n5536_), .ZN(new_n5537_));
  NOR2_X1    g04535(.A1(new_n5529_), .A2(new_n5537_), .ZN(new_n5538_));
  NAND2_X1   g04536(.A1(new_n5525_), .A2(new_n5526_), .ZN(new_n5539_));
  NOR2_X1    g04537(.A1(new_n5522_), .A2(new_n5520_), .ZN(new_n5540_));
  AOI21_X1   g04538(.A1(new_n5539_), .A2(\A[300] ), .B(new_n5540_), .ZN(new_n5541_));
  NAND2_X1   g04539(.A1(new_n5510_), .A2(new_n5531_), .ZN(new_n5542_));
  NOR2_X1    g04540(.A1(new_n5509_), .A2(new_n5511_), .ZN(new_n5543_));
  AOI21_X1   g04541(.A1(new_n5542_), .A2(\A[297] ), .B(new_n5543_), .ZN(new_n5544_));
  OAI22_X1   g04542(.A1(new_n5530_), .A2(new_n5532_), .B1(new_n5527_), .B2(new_n5524_), .ZN(new_n5545_));
  NOR3_X1    g04543(.A1(new_n5545_), .A2(new_n5541_), .A3(new_n5544_), .ZN(new_n5546_));
  NOR2_X1    g04544(.A1(new_n5538_), .A2(new_n5546_), .ZN(new_n5547_));
  NAND2_X1   g04545(.A1(new_n5547_), .A2(new_n5508_), .ZN(new_n5548_));
  NOR2_X1    g04546(.A1(new_n5495_), .A2(new_n5492_), .ZN(new_n5549_));
  NOR2_X1    g04547(.A1(new_n5477_), .A2(new_n5487_), .ZN(new_n5550_));
  NOR2_X1    g04548(.A1(new_n5549_), .A2(new_n5550_), .ZN(new_n5551_));
  NAND2_X1   g04549(.A1(new_n5479_), .A2(new_n5481_), .ZN(new_n5552_));
  AOI21_X1   g04550(.A1(new_n5552_), .A2(\A[306] ), .B(new_n5499_), .ZN(new_n5553_));
  NAND2_X1   g04551(.A1(new_n5474_), .A2(new_n5475_), .ZN(new_n5554_));
  AOI21_X1   g04552(.A1(new_n5554_), .A2(\A[303] ), .B(new_n5503_), .ZN(new_n5555_));
  OAI22_X1   g04553(.A1(new_n5473_), .A2(new_n5476_), .B1(new_n5494_), .B2(new_n5493_), .ZN(new_n5556_));
  NOR3_X1    g04554(.A1(new_n5556_), .A2(new_n5553_), .A3(new_n5555_), .ZN(new_n5557_));
  NOR2_X1    g04555(.A1(new_n5551_), .A2(new_n5557_), .ZN(new_n5558_));
  XOR2_X1    g04556(.A1(new_n5518_), .A2(new_n5536_), .Z(new_n5559_));
  INV_X1     g04557(.I(new_n5546_), .ZN(new_n5560_));
  NAND2_X1   g04558(.A1(new_n5560_), .A2(new_n5559_), .ZN(new_n5561_));
  NAND2_X1   g04559(.A1(new_n5561_), .A2(new_n5558_), .ZN(new_n5562_));
  NAND2_X1   g04560(.A1(new_n5562_), .A2(new_n5548_), .ZN(new_n5563_));
  NAND3_X1   g04561(.A1(new_n5563_), .A2(new_n5439_), .A3(new_n5467_), .ZN(new_n5564_));
  NAND2_X1   g04562(.A1(new_n5439_), .A2(new_n5467_), .ZN(new_n5565_));
  NAND3_X1   g04563(.A1(new_n5565_), .A2(new_n5548_), .A3(new_n5562_), .ZN(new_n5566_));
  NAND2_X1   g04564(.A1(new_n5564_), .A2(new_n5566_), .ZN(new_n5567_));
  INV_X1     g04565(.I(\A[290] ), .ZN(new_n5568_));
  NOR2_X1    g04566(.A1(new_n5568_), .A2(\A[289] ), .ZN(new_n5569_));
  INV_X1     g04567(.I(\A[289] ), .ZN(new_n5570_));
  OAI21_X1   g04568(.A1(new_n5570_), .A2(\A[290] ), .B(\A[291] ), .ZN(new_n5571_));
  NOR2_X1    g04569(.A1(new_n5571_), .A2(new_n5569_), .ZN(new_n5572_));
  NAND2_X1   g04570(.A1(new_n5570_), .A2(\A[290] ), .ZN(new_n5573_));
  NAND2_X1   g04571(.A1(new_n5568_), .A2(\A[289] ), .ZN(new_n5574_));
  AOI21_X1   g04572(.A1(new_n5573_), .A2(new_n5574_), .B(\A[291] ), .ZN(new_n5575_));
  NOR2_X1    g04573(.A1(new_n5575_), .A2(new_n5572_), .ZN(new_n5576_));
  INV_X1     g04574(.I(\A[292] ), .ZN(new_n5577_));
  NAND2_X1   g04575(.A1(new_n5577_), .A2(\A[293] ), .ZN(new_n5578_));
  INV_X1     g04576(.I(\A[293] ), .ZN(new_n5579_));
  INV_X1     g04577(.I(\A[294] ), .ZN(new_n5580_));
  AOI21_X1   g04578(.A1(\A[292] ), .A2(new_n5579_), .B(new_n5580_), .ZN(new_n5581_));
  NAND2_X1   g04579(.A1(new_n5581_), .A2(new_n5578_), .ZN(new_n5582_));
  NOR2_X1    g04580(.A1(new_n5579_), .A2(\A[292] ), .ZN(new_n5583_));
  NOR2_X1    g04581(.A1(new_n5577_), .A2(\A[293] ), .ZN(new_n5584_));
  OAI21_X1   g04582(.A1(new_n5583_), .A2(new_n5584_), .B(new_n5580_), .ZN(new_n5585_));
  NAND2_X1   g04583(.A1(new_n5582_), .A2(new_n5585_), .ZN(new_n5586_));
  NAND2_X1   g04584(.A1(new_n5586_), .A2(new_n5576_), .ZN(new_n5587_));
  NAND3_X1   g04585(.A1(new_n5573_), .A2(new_n5574_), .A3(\A[291] ), .ZN(new_n5588_));
  INV_X1     g04586(.I(\A[291] ), .ZN(new_n5589_));
  NOR2_X1    g04587(.A1(new_n5570_), .A2(\A[290] ), .ZN(new_n5590_));
  OAI21_X1   g04588(.A1(new_n5569_), .A2(new_n5590_), .B(new_n5589_), .ZN(new_n5591_));
  NAND2_X1   g04589(.A1(new_n5591_), .A2(new_n5588_), .ZN(new_n5592_));
  XOR2_X1    g04590(.A1(\A[292] ), .A2(\A[293] ), .Z(new_n5593_));
  AOI22_X1   g04591(.A1(new_n5593_), .A2(new_n5580_), .B1(new_n5578_), .B2(new_n5581_), .ZN(new_n5594_));
  NAND2_X1   g04592(.A1(new_n5592_), .A2(new_n5594_), .ZN(new_n5595_));
  NAND2_X1   g04593(.A1(new_n5587_), .A2(new_n5595_), .ZN(new_n5596_));
  NOR2_X1    g04594(.A1(new_n5583_), .A2(new_n5584_), .ZN(new_n5597_));
  NOR2_X1    g04595(.A1(new_n5577_), .A2(new_n5579_), .ZN(new_n5598_));
  INV_X1     g04596(.I(new_n5598_), .ZN(new_n5599_));
  OAI21_X1   g04597(.A1(new_n5597_), .A2(new_n5580_), .B(new_n5599_), .ZN(new_n5600_));
  XNOR2_X1   g04598(.A1(\A[289] ), .A2(\A[290] ), .ZN(new_n5601_));
  NAND2_X1   g04599(.A1(\A[289] ), .A2(\A[290] ), .ZN(new_n5602_));
  OAI21_X1   g04600(.A1(new_n5601_), .A2(new_n5589_), .B(new_n5602_), .ZN(new_n5603_));
  AOI22_X1   g04601(.A1(new_n5582_), .A2(new_n5585_), .B1(new_n5591_), .B2(new_n5588_), .ZN(new_n5604_));
  NAND3_X1   g04602(.A1(new_n5604_), .A2(new_n5600_), .A3(new_n5603_), .ZN(new_n5605_));
  NAND2_X1   g04603(.A1(new_n5596_), .A2(new_n5605_), .ZN(new_n5606_));
  INV_X1     g04604(.I(\A[283] ), .ZN(new_n5607_));
  NAND2_X1   g04605(.A1(new_n5607_), .A2(\A[284] ), .ZN(new_n5608_));
  INV_X1     g04606(.I(\A[284] ), .ZN(new_n5609_));
  INV_X1     g04607(.I(\A[285] ), .ZN(new_n5610_));
  AOI21_X1   g04608(.A1(\A[283] ), .A2(new_n5609_), .B(new_n5610_), .ZN(new_n5611_));
  NAND2_X1   g04609(.A1(new_n5611_), .A2(new_n5608_), .ZN(new_n5612_));
  NOR2_X1    g04610(.A1(new_n5609_), .A2(\A[283] ), .ZN(new_n5613_));
  NOR2_X1    g04611(.A1(new_n5607_), .A2(\A[284] ), .ZN(new_n5614_));
  OAI21_X1   g04612(.A1(new_n5613_), .A2(new_n5614_), .B(new_n5610_), .ZN(new_n5615_));
  NAND2_X1   g04613(.A1(new_n5612_), .A2(new_n5615_), .ZN(new_n5616_));
  INV_X1     g04614(.I(\A[288] ), .ZN(new_n5617_));
  INV_X1     g04615(.I(\A[287] ), .ZN(new_n5618_));
  NOR2_X1    g04616(.A1(new_n5618_), .A2(\A[286] ), .ZN(new_n5619_));
  INV_X1     g04617(.I(\A[286] ), .ZN(new_n5620_));
  NOR2_X1    g04618(.A1(new_n5620_), .A2(\A[287] ), .ZN(new_n5621_));
  NOR3_X1    g04619(.A1(new_n5619_), .A2(new_n5621_), .A3(new_n5617_), .ZN(new_n5622_));
  NAND2_X1   g04620(.A1(new_n5620_), .A2(\A[287] ), .ZN(new_n5623_));
  NAND2_X1   g04621(.A1(new_n5618_), .A2(\A[286] ), .ZN(new_n5624_));
  AOI21_X1   g04622(.A1(new_n5623_), .A2(new_n5624_), .B(\A[288] ), .ZN(new_n5625_));
  NOR2_X1    g04623(.A1(new_n5625_), .A2(new_n5622_), .ZN(new_n5626_));
  NOR2_X1    g04624(.A1(new_n5626_), .A2(new_n5616_), .ZN(new_n5627_));
  NOR3_X1    g04625(.A1(new_n5613_), .A2(new_n5614_), .A3(new_n5610_), .ZN(new_n5628_));
  NAND2_X1   g04626(.A1(new_n5609_), .A2(\A[283] ), .ZN(new_n5629_));
  AOI21_X1   g04627(.A1(new_n5608_), .A2(new_n5629_), .B(\A[285] ), .ZN(new_n5630_));
  NOR2_X1    g04628(.A1(new_n5630_), .A2(new_n5628_), .ZN(new_n5631_));
  NAND3_X1   g04629(.A1(new_n5623_), .A2(new_n5624_), .A3(\A[288] ), .ZN(new_n5632_));
  OAI21_X1   g04630(.A1(new_n5619_), .A2(new_n5621_), .B(new_n5617_), .ZN(new_n5633_));
  NAND2_X1   g04631(.A1(new_n5633_), .A2(new_n5632_), .ZN(new_n5634_));
  NOR2_X1    g04632(.A1(new_n5631_), .A2(new_n5634_), .ZN(new_n5635_));
  NOR2_X1    g04633(.A1(new_n5627_), .A2(new_n5635_), .ZN(new_n5636_));
  XOR2_X1    g04634(.A1(\A[286] ), .A2(\A[287] ), .Z(new_n5637_));
  NOR2_X1    g04635(.A1(new_n5620_), .A2(new_n5618_), .ZN(new_n5638_));
  AOI21_X1   g04636(.A1(new_n5637_), .A2(\A[288] ), .B(new_n5638_), .ZN(new_n5639_));
  XOR2_X1    g04637(.A1(\A[283] ), .A2(\A[284] ), .Z(new_n5640_));
  NAND2_X1   g04638(.A1(\A[283] ), .A2(\A[284] ), .ZN(new_n5641_));
  INV_X1     g04639(.I(new_n5641_), .ZN(new_n5642_));
  AOI21_X1   g04640(.A1(new_n5640_), .A2(\A[285] ), .B(new_n5642_), .ZN(new_n5643_));
  OAI22_X1   g04641(.A1(new_n5628_), .A2(new_n5630_), .B1(new_n5625_), .B2(new_n5622_), .ZN(new_n5644_));
  NOR3_X1    g04642(.A1(new_n5644_), .A2(new_n5639_), .A3(new_n5643_), .ZN(new_n5645_));
  NOR2_X1    g04643(.A1(new_n5636_), .A2(new_n5645_), .ZN(new_n5646_));
  NAND2_X1   g04644(.A1(new_n5646_), .A2(new_n5606_), .ZN(new_n5647_));
  NAND2_X1   g04645(.A1(new_n5631_), .A2(new_n5634_), .ZN(new_n5648_));
  NAND2_X1   g04646(.A1(new_n5626_), .A2(new_n5616_), .ZN(new_n5649_));
  NAND2_X1   g04647(.A1(new_n5649_), .A2(new_n5648_), .ZN(new_n5650_));
  NOR2_X1    g04648(.A1(new_n5619_), .A2(new_n5621_), .ZN(new_n5651_));
  INV_X1     g04649(.I(new_n5638_), .ZN(new_n5652_));
  OAI21_X1   g04650(.A1(new_n5651_), .A2(new_n5617_), .B(new_n5652_), .ZN(new_n5653_));
  NOR2_X1    g04651(.A1(new_n5613_), .A2(new_n5614_), .ZN(new_n5654_));
  OAI21_X1   g04652(.A1(new_n5654_), .A2(new_n5610_), .B(new_n5641_), .ZN(new_n5655_));
  AOI22_X1   g04653(.A1(new_n5612_), .A2(new_n5615_), .B1(new_n5633_), .B2(new_n5632_), .ZN(new_n5656_));
  NAND3_X1   g04654(.A1(new_n5656_), .A2(new_n5653_), .A3(new_n5655_), .ZN(new_n5657_));
  NAND2_X1   g04655(.A1(new_n5650_), .A2(new_n5657_), .ZN(new_n5658_));
  NAND3_X1   g04656(.A1(new_n5658_), .A2(new_n5596_), .A3(new_n5605_), .ZN(new_n5659_));
  INV_X1     g04657(.I(\A[278] ), .ZN(new_n5660_));
  NOR2_X1    g04658(.A1(new_n5660_), .A2(\A[277] ), .ZN(new_n5661_));
  NAND2_X1   g04659(.A1(new_n5660_), .A2(\A[277] ), .ZN(new_n5662_));
  NAND2_X1   g04660(.A1(new_n5662_), .A2(\A[279] ), .ZN(new_n5663_));
  NOR2_X1    g04661(.A1(new_n5663_), .A2(new_n5661_), .ZN(new_n5664_));
  INV_X1     g04662(.I(\A[277] ), .ZN(new_n5665_));
  NAND2_X1   g04663(.A1(new_n5665_), .A2(\A[278] ), .ZN(new_n5666_));
  AOI21_X1   g04664(.A1(new_n5666_), .A2(new_n5662_), .B(\A[279] ), .ZN(new_n5667_));
  NOR2_X1    g04665(.A1(new_n5664_), .A2(new_n5667_), .ZN(new_n5668_));
  INV_X1     g04666(.I(\A[280] ), .ZN(new_n5669_));
  NAND2_X1   g04667(.A1(new_n5669_), .A2(\A[281] ), .ZN(new_n5670_));
  INV_X1     g04668(.I(\A[281] ), .ZN(new_n5671_));
  NAND2_X1   g04669(.A1(new_n5671_), .A2(\A[280] ), .ZN(new_n5672_));
  NAND3_X1   g04670(.A1(new_n5670_), .A2(new_n5672_), .A3(\A[282] ), .ZN(new_n5673_));
  INV_X1     g04671(.I(\A[282] ), .ZN(new_n5674_));
  NOR2_X1    g04672(.A1(new_n5671_), .A2(\A[280] ), .ZN(new_n5675_));
  NOR2_X1    g04673(.A1(new_n5669_), .A2(\A[281] ), .ZN(new_n5676_));
  OAI21_X1   g04674(.A1(new_n5675_), .A2(new_n5676_), .B(new_n5674_), .ZN(new_n5677_));
  NAND2_X1   g04675(.A1(new_n5677_), .A2(new_n5673_), .ZN(new_n5678_));
  NAND2_X1   g04676(.A1(new_n5668_), .A2(new_n5678_), .ZN(new_n5679_));
  NAND3_X1   g04677(.A1(new_n5666_), .A2(new_n5662_), .A3(\A[279] ), .ZN(new_n5680_));
  INV_X1     g04678(.I(\A[279] ), .ZN(new_n5681_));
  NOR2_X1    g04679(.A1(new_n5665_), .A2(\A[278] ), .ZN(new_n5682_));
  OAI21_X1   g04680(.A1(new_n5661_), .A2(new_n5682_), .B(new_n5681_), .ZN(new_n5683_));
  NAND2_X1   g04681(.A1(new_n5683_), .A2(new_n5680_), .ZN(new_n5684_));
  NOR3_X1    g04682(.A1(new_n5675_), .A2(new_n5676_), .A3(new_n5674_), .ZN(new_n5685_));
  AOI21_X1   g04683(.A1(new_n5670_), .A2(new_n5672_), .B(\A[282] ), .ZN(new_n5686_));
  NOR2_X1    g04684(.A1(new_n5686_), .A2(new_n5685_), .ZN(new_n5687_));
  NAND2_X1   g04685(.A1(new_n5687_), .A2(new_n5684_), .ZN(new_n5688_));
  NAND2_X1   g04686(.A1(new_n5679_), .A2(new_n5688_), .ZN(new_n5689_));
  NOR2_X1    g04687(.A1(new_n5675_), .A2(new_n5676_), .ZN(new_n5690_));
  NOR2_X1    g04688(.A1(new_n5669_), .A2(new_n5671_), .ZN(new_n5691_));
  INV_X1     g04689(.I(new_n5691_), .ZN(new_n5692_));
  OAI21_X1   g04690(.A1(new_n5690_), .A2(new_n5674_), .B(new_n5692_), .ZN(new_n5693_));
  NOR2_X1    g04691(.A1(new_n5661_), .A2(new_n5682_), .ZN(new_n5694_));
  NOR2_X1    g04692(.A1(new_n5665_), .A2(new_n5660_), .ZN(new_n5695_));
  INV_X1     g04693(.I(new_n5695_), .ZN(new_n5696_));
  OAI21_X1   g04694(.A1(new_n5694_), .A2(new_n5681_), .B(new_n5696_), .ZN(new_n5697_));
  AOI22_X1   g04695(.A1(new_n5680_), .A2(new_n5683_), .B1(new_n5677_), .B2(new_n5673_), .ZN(new_n5698_));
  NAND3_X1   g04696(.A1(new_n5698_), .A2(new_n5693_), .A3(new_n5697_), .ZN(new_n5699_));
  NAND2_X1   g04697(.A1(new_n5689_), .A2(new_n5699_), .ZN(new_n5700_));
  INV_X1     g04698(.I(\A[272] ), .ZN(new_n5701_));
  NOR2_X1    g04699(.A1(new_n5701_), .A2(\A[271] ), .ZN(new_n5702_));
  NAND2_X1   g04700(.A1(new_n5701_), .A2(\A[271] ), .ZN(new_n5703_));
  NAND2_X1   g04701(.A1(new_n5703_), .A2(\A[273] ), .ZN(new_n5704_));
  INV_X1     g04702(.I(\A[271] ), .ZN(new_n5705_));
  NOR2_X1    g04703(.A1(new_n5705_), .A2(\A[272] ), .ZN(new_n5706_));
  NOR2_X1    g04704(.A1(new_n5702_), .A2(new_n5706_), .ZN(new_n5707_));
  OAI22_X1   g04705(.A1(new_n5707_), .A2(\A[273] ), .B1(new_n5704_), .B2(new_n5702_), .ZN(new_n5708_));
  INV_X1     g04706(.I(\A[276] ), .ZN(new_n5709_));
  INV_X1     g04707(.I(\A[275] ), .ZN(new_n5710_));
  NOR2_X1    g04708(.A1(new_n5710_), .A2(\A[274] ), .ZN(new_n5711_));
  INV_X1     g04709(.I(\A[274] ), .ZN(new_n5712_));
  NOR2_X1    g04710(.A1(new_n5712_), .A2(\A[275] ), .ZN(new_n5713_));
  NOR3_X1    g04711(.A1(new_n5711_), .A2(new_n5713_), .A3(new_n5709_), .ZN(new_n5714_));
  NAND2_X1   g04712(.A1(new_n5712_), .A2(\A[275] ), .ZN(new_n5715_));
  NAND2_X1   g04713(.A1(new_n5710_), .A2(\A[274] ), .ZN(new_n5716_));
  AOI21_X1   g04714(.A1(new_n5715_), .A2(new_n5716_), .B(\A[276] ), .ZN(new_n5717_));
  NOR2_X1    g04715(.A1(new_n5717_), .A2(new_n5714_), .ZN(new_n5718_));
  NOR2_X1    g04716(.A1(new_n5708_), .A2(new_n5718_), .ZN(new_n5719_));
  NOR2_X1    g04717(.A1(new_n5704_), .A2(new_n5702_), .ZN(new_n5720_));
  NAND2_X1   g04718(.A1(new_n5705_), .A2(\A[272] ), .ZN(new_n5721_));
  AOI21_X1   g04719(.A1(new_n5721_), .A2(new_n5703_), .B(\A[273] ), .ZN(new_n5722_));
  NOR2_X1    g04720(.A1(new_n5720_), .A2(new_n5722_), .ZN(new_n5723_));
  NAND2_X1   g04721(.A1(new_n5716_), .A2(\A[276] ), .ZN(new_n5724_));
  NOR2_X1    g04722(.A1(new_n5711_), .A2(new_n5713_), .ZN(new_n5725_));
  OAI22_X1   g04723(.A1(new_n5725_), .A2(\A[276] ), .B1(new_n5724_), .B2(new_n5711_), .ZN(new_n5726_));
  NOR2_X1    g04724(.A1(new_n5723_), .A2(new_n5726_), .ZN(new_n5727_));
  NOR2_X1    g04725(.A1(new_n5727_), .A2(new_n5719_), .ZN(new_n5728_));
  NOR2_X1    g04726(.A1(new_n5712_), .A2(new_n5710_), .ZN(new_n5729_));
  INV_X1     g04727(.I(new_n5729_), .ZN(new_n5730_));
  OAI21_X1   g04728(.A1(new_n5725_), .A2(new_n5709_), .B(new_n5730_), .ZN(new_n5731_));
  INV_X1     g04729(.I(\A[273] ), .ZN(new_n5732_));
  NOR2_X1    g04730(.A1(new_n5705_), .A2(new_n5701_), .ZN(new_n5733_));
  INV_X1     g04731(.I(new_n5733_), .ZN(new_n5734_));
  OAI21_X1   g04732(.A1(new_n5707_), .A2(new_n5732_), .B(new_n5734_), .ZN(new_n5735_));
  NAND4_X1   g04733(.A1(new_n5708_), .A2(new_n5726_), .A3(new_n5731_), .A4(new_n5735_), .ZN(new_n5736_));
  INV_X1     g04734(.I(new_n5736_), .ZN(new_n5737_));
  NOR2_X1    g04735(.A1(new_n5737_), .A2(new_n5728_), .ZN(new_n5738_));
  NAND2_X1   g04736(.A1(new_n5738_), .A2(new_n5700_), .ZN(new_n5739_));
  NAND2_X1   g04737(.A1(new_n5723_), .A2(new_n5726_), .ZN(new_n5740_));
  NAND2_X1   g04738(.A1(new_n5708_), .A2(new_n5718_), .ZN(new_n5741_));
  NAND2_X1   g04739(.A1(new_n5740_), .A2(new_n5741_), .ZN(new_n5742_));
  NAND2_X1   g04740(.A1(new_n5742_), .A2(new_n5736_), .ZN(new_n5743_));
  NAND3_X1   g04741(.A1(new_n5743_), .A2(new_n5689_), .A3(new_n5699_), .ZN(new_n5744_));
  NAND2_X1   g04742(.A1(new_n5739_), .A2(new_n5744_), .ZN(new_n5745_));
  NAND3_X1   g04743(.A1(new_n5745_), .A2(new_n5647_), .A3(new_n5659_), .ZN(new_n5746_));
  NAND2_X1   g04744(.A1(new_n5659_), .A2(new_n5647_), .ZN(new_n5747_));
  NAND3_X1   g04745(.A1(new_n5747_), .A2(new_n5739_), .A3(new_n5744_), .ZN(new_n5748_));
  NAND2_X1   g04746(.A1(new_n5746_), .A2(new_n5748_), .ZN(new_n5749_));
  XOR2_X1    g04747(.A1(new_n5567_), .A2(new_n5749_), .Z(new_n5750_));
  XOR2_X1    g04748(.A1(new_n5370_), .A2(new_n5750_), .Z(new_n5751_));
  XNOR2_X1   g04749(.A1(new_n4973_), .A2(new_n5751_), .ZN(new_n5752_));
  INV_X1     g04750(.I(\A[222] ), .ZN(new_n5753_));
  NAND2_X1   g04751(.A1(\A[220] ), .A2(\A[221] ), .ZN(new_n5754_));
  XNOR2_X1   g04752(.A1(\A[220] ), .A2(\A[221] ), .ZN(new_n5755_));
  OAI21_X1   g04753(.A1(new_n5755_), .A2(new_n5753_), .B(new_n5754_), .ZN(new_n5756_));
  INV_X1     g04754(.I(\A[219] ), .ZN(new_n5757_));
  NAND2_X1   g04755(.A1(\A[217] ), .A2(\A[218] ), .ZN(new_n5758_));
  XNOR2_X1   g04756(.A1(\A[217] ), .A2(\A[218] ), .ZN(new_n5759_));
  OAI21_X1   g04757(.A1(new_n5759_), .A2(new_n5757_), .B(new_n5758_), .ZN(new_n5760_));
  INV_X1     g04758(.I(\A[217] ), .ZN(new_n5761_));
  NOR2_X1    g04759(.A1(new_n5761_), .A2(\A[218] ), .ZN(new_n5762_));
  INV_X1     g04760(.I(\A[218] ), .ZN(new_n5763_));
  NOR2_X1    g04761(.A1(new_n5763_), .A2(\A[217] ), .ZN(new_n5764_));
  OAI21_X1   g04762(.A1(new_n5762_), .A2(new_n5764_), .B(new_n5757_), .ZN(new_n5765_));
  NAND2_X1   g04763(.A1(new_n5763_), .A2(\A[217] ), .ZN(new_n5766_));
  NAND2_X1   g04764(.A1(new_n5761_), .A2(\A[218] ), .ZN(new_n5767_));
  NAND3_X1   g04765(.A1(new_n5766_), .A2(new_n5767_), .A3(\A[219] ), .ZN(new_n5768_));
  INV_X1     g04766(.I(\A[220] ), .ZN(new_n5769_));
  NOR2_X1    g04767(.A1(new_n5769_), .A2(\A[221] ), .ZN(new_n5770_));
  INV_X1     g04768(.I(\A[221] ), .ZN(new_n5771_));
  NOR2_X1    g04769(.A1(new_n5771_), .A2(\A[220] ), .ZN(new_n5772_));
  OAI21_X1   g04770(.A1(new_n5770_), .A2(new_n5772_), .B(new_n5753_), .ZN(new_n5773_));
  NAND2_X1   g04771(.A1(new_n5771_), .A2(\A[220] ), .ZN(new_n5774_));
  NAND2_X1   g04772(.A1(new_n5769_), .A2(\A[221] ), .ZN(new_n5775_));
  NAND3_X1   g04773(.A1(new_n5774_), .A2(new_n5775_), .A3(\A[222] ), .ZN(new_n5776_));
  AOI22_X1   g04774(.A1(new_n5765_), .A2(new_n5768_), .B1(new_n5773_), .B2(new_n5776_), .ZN(new_n5777_));
  NAND3_X1   g04775(.A1(new_n5777_), .A2(new_n5756_), .A3(new_n5760_), .ZN(new_n5778_));
  AOI21_X1   g04776(.A1(new_n5766_), .A2(new_n5767_), .B(\A[219] ), .ZN(new_n5779_));
  OAI21_X1   g04777(.A1(new_n5761_), .A2(\A[218] ), .B(\A[219] ), .ZN(new_n5780_));
  NOR2_X1    g04778(.A1(new_n5780_), .A2(new_n5764_), .ZN(new_n5781_));
  NOR2_X1    g04779(.A1(new_n5779_), .A2(new_n5781_), .ZN(new_n5782_));
  NAND2_X1   g04780(.A1(new_n5773_), .A2(new_n5776_), .ZN(new_n5783_));
  NAND2_X1   g04781(.A1(new_n5783_), .A2(new_n5782_), .ZN(new_n5784_));
  NAND2_X1   g04782(.A1(new_n5765_), .A2(new_n5768_), .ZN(new_n5785_));
  AOI21_X1   g04783(.A1(new_n5774_), .A2(new_n5775_), .B(\A[222] ), .ZN(new_n5786_));
  OAI21_X1   g04784(.A1(new_n5769_), .A2(\A[221] ), .B(\A[222] ), .ZN(new_n5787_));
  NOR2_X1    g04785(.A1(new_n5787_), .A2(new_n5772_), .ZN(new_n5788_));
  NOR2_X1    g04786(.A1(new_n5786_), .A2(new_n5788_), .ZN(new_n5789_));
  NAND2_X1   g04787(.A1(new_n5785_), .A2(new_n5789_), .ZN(new_n5790_));
  NAND2_X1   g04788(.A1(new_n5784_), .A2(new_n5790_), .ZN(new_n5791_));
  NAND2_X1   g04789(.A1(new_n5791_), .A2(new_n5778_), .ZN(new_n5792_));
  INV_X1     g04790(.I(\A[213] ), .ZN(new_n5793_));
  INV_X1     g04791(.I(\A[211] ), .ZN(new_n5794_));
  NOR2_X1    g04792(.A1(new_n5794_), .A2(\A[212] ), .ZN(new_n5795_));
  INV_X1     g04793(.I(\A[212] ), .ZN(new_n5796_));
  NOR2_X1    g04794(.A1(new_n5796_), .A2(\A[211] ), .ZN(new_n5797_));
  OAI21_X1   g04795(.A1(new_n5795_), .A2(new_n5797_), .B(new_n5793_), .ZN(new_n5798_));
  NAND2_X1   g04796(.A1(new_n5796_), .A2(\A[211] ), .ZN(new_n5799_));
  NAND2_X1   g04797(.A1(new_n5794_), .A2(\A[212] ), .ZN(new_n5800_));
  NAND3_X1   g04798(.A1(new_n5799_), .A2(new_n5800_), .A3(\A[213] ), .ZN(new_n5801_));
  NAND2_X1   g04799(.A1(new_n5798_), .A2(new_n5801_), .ZN(new_n5802_));
  INV_X1     g04800(.I(\A[215] ), .ZN(new_n5803_));
  NAND2_X1   g04801(.A1(new_n5803_), .A2(\A[214] ), .ZN(new_n5804_));
  INV_X1     g04802(.I(\A[214] ), .ZN(new_n5805_));
  NAND2_X1   g04803(.A1(new_n5805_), .A2(\A[215] ), .ZN(new_n5806_));
  AOI21_X1   g04804(.A1(new_n5804_), .A2(new_n5806_), .B(\A[216] ), .ZN(new_n5807_));
  NOR2_X1    g04805(.A1(new_n5803_), .A2(\A[214] ), .ZN(new_n5808_));
  OAI21_X1   g04806(.A1(new_n5805_), .A2(\A[215] ), .B(\A[216] ), .ZN(new_n5809_));
  NOR2_X1    g04807(.A1(new_n5809_), .A2(new_n5808_), .ZN(new_n5810_));
  NOR2_X1    g04808(.A1(new_n5807_), .A2(new_n5810_), .ZN(new_n5811_));
  NOR2_X1    g04809(.A1(new_n5802_), .A2(new_n5811_), .ZN(new_n5812_));
  AOI21_X1   g04810(.A1(new_n5799_), .A2(new_n5800_), .B(\A[213] ), .ZN(new_n5813_));
  OAI21_X1   g04811(.A1(new_n5794_), .A2(\A[212] ), .B(\A[213] ), .ZN(new_n5814_));
  NOR2_X1    g04812(.A1(new_n5814_), .A2(new_n5797_), .ZN(new_n5815_));
  NOR2_X1    g04813(.A1(new_n5813_), .A2(new_n5815_), .ZN(new_n5816_));
  INV_X1     g04814(.I(\A[216] ), .ZN(new_n5817_));
  NOR2_X1    g04815(.A1(new_n5805_), .A2(\A[215] ), .ZN(new_n5818_));
  OAI21_X1   g04816(.A1(new_n5818_), .A2(new_n5808_), .B(new_n5817_), .ZN(new_n5819_));
  NAND3_X1   g04817(.A1(new_n5804_), .A2(new_n5806_), .A3(\A[216] ), .ZN(new_n5820_));
  NAND2_X1   g04818(.A1(new_n5819_), .A2(new_n5820_), .ZN(new_n5821_));
  NOR2_X1    g04819(.A1(new_n5821_), .A2(new_n5816_), .ZN(new_n5822_));
  NOR2_X1    g04820(.A1(new_n5812_), .A2(new_n5822_), .ZN(new_n5823_));
  XOR2_X1    g04821(.A1(\A[214] ), .A2(\A[215] ), .Z(new_n5824_));
  NAND2_X1   g04822(.A1(\A[214] ), .A2(\A[215] ), .ZN(new_n5825_));
  INV_X1     g04823(.I(new_n5825_), .ZN(new_n5826_));
  AOI21_X1   g04824(.A1(new_n5824_), .A2(\A[216] ), .B(new_n5826_), .ZN(new_n5827_));
  XOR2_X1    g04825(.A1(\A[211] ), .A2(\A[212] ), .Z(new_n5828_));
  NOR2_X1    g04826(.A1(new_n5794_), .A2(new_n5796_), .ZN(new_n5829_));
  AOI21_X1   g04827(.A1(new_n5828_), .A2(\A[213] ), .B(new_n5829_), .ZN(new_n5830_));
  OAI22_X1   g04828(.A1(new_n5813_), .A2(new_n5815_), .B1(new_n5807_), .B2(new_n5810_), .ZN(new_n5831_));
  NOR3_X1    g04829(.A1(new_n5831_), .A2(new_n5827_), .A3(new_n5830_), .ZN(new_n5832_));
  NOR2_X1    g04830(.A1(new_n5823_), .A2(new_n5832_), .ZN(new_n5833_));
  NAND2_X1   g04831(.A1(new_n5833_), .A2(new_n5792_), .ZN(new_n5834_));
  INV_X1     g04832(.I(new_n5754_), .ZN(new_n5835_));
  XOR2_X1    g04833(.A1(\A[220] ), .A2(\A[221] ), .Z(new_n5836_));
  AOI21_X1   g04834(.A1(new_n5836_), .A2(\A[222] ), .B(new_n5835_), .ZN(new_n5837_));
  INV_X1     g04835(.I(new_n5758_), .ZN(new_n5838_));
  XOR2_X1    g04836(.A1(\A[217] ), .A2(\A[218] ), .Z(new_n5839_));
  AOI21_X1   g04837(.A1(new_n5839_), .A2(\A[219] ), .B(new_n5838_), .ZN(new_n5840_));
  OAI22_X1   g04838(.A1(new_n5779_), .A2(new_n5781_), .B1(new_n5786_), .B2(new_n5788_), .ZN(new_n5841_));
  NOR3_X1    g04839(.A1(new_n5841_), .A2(new_n5837_), .A3(new_n5840_), .ZN(new_n5842_));
  NOR2_X1    g04840(.A1(new_n5785_), .A2(new_n5789_), .ZN(new_n5843_));
  NOR2_X1    g04841(.A1(new_n5783_), .A2(new_n5782_), .ZN(new_n5844_));
  NOR2_X1    g04842(.A1(new_n5843_), .A2(new_n5844_), .ZN(new_n5845_));
  NOR2_X1    g04843(.A1(new_n5845_), .A2(new_n5842_), .ZN(new_n5846_));
  NAND2_X1   g04844(.A1(new_n5821_), .A2(new_n5816_), .ZN(new_n5847_));
  NAND2_X1   g04845(.A1(new_n5802_), .A2(new_n5811_), .ZN(new_n5848_));
  NAND2_X1   g04846(.A1(new_n5847_), .A2(new_n5848_), .ZN(new_n5849_));
  XNOR2_X1   g04847(.A1(\A[214] ), .A2(\A[215] ), .ZN(new_n5850_));
  OAI21_X1   g04848(.A1(new_n5850_), .A2(new_n5817_), .B(new_n5825_), .ZN(new_n5851_));
  NOR2_X1    g04849(.A1(new_n5795_), .A2(new_n5797_), .ZN(new_n5852_));
  INV_X1     g04850(.I(new_n5829_), .ZN(new_n5853_));
  OAI21_X1   g04851(.A1(new_n5852_), .A2(new_n5793_), .B(new_n5853_), .ZN(new_n5854_));
  AOI22_X1   g04852(.A1(new_n5798_), .A2(new_n5801_), .B1(new_n5819_), .B2(new_n5820_), .ZN(new_n5855_));
  NAND3_X1   g04853(.A1(new_n5855_), .A2(new_n5851_), .A3(new_n5854_), .ZN(new_n5856_));
  NAND2_X1   g04854(.A1(new_n5849_), .A2(new_n5856_), .ZN(new_n5857_));
  NAND2_X1   g04855(.A1(new_n5846_), .A2(new_n5857_), .ZN(new_n5858_));
  NAND2_X1   g04856(.A1(new_n5834_), .A2(new_n5858_), .ZN(new_n5859_));
  INV_X1     g04857(.I(\A[208] ), .ZN(new_n5860_));
  INV_X1     g04858(.I(\A[209] ), .ZN(new_n5861_));
  NOR2_X1    g04859(.A1(new_n5860_), .A2(new_n5861_), .ZN(new_n5862_));
  XOR2_X1    g04860(.A1(\A[208] ), .A2(\A[209] ), .Z(new_n5863_));
  AOI21_X1   g04861(.A1(new_n5863_), .A2(\A[210] ), .B(new_n5862_), .ZN(new_n5864_));
  INV_X1     g04862(.I(\A[205] ), .ZN(new_n5865_));
  INV_X1     g04863(.I(\A[206] ), .ZN(new_n5866_));
  NOR2_X1    g04864(.A1(new_n5865_), .A2(new_n5866_), .ZN(new_n5867_));
  XOR2_X1    g04865(.A1(\A[205] ), .A2(\A[206] ), .Z(new_n5868_));
  AOI21_X1   g04866(.A1(new_n5868_), .A2(\A[207] ), .B(new_n5867_), .ZN(new_n5869_));
  NAND2_X1   g04867(.A1(new_n5866_), .A2(\A[205] ), .ZN(new_n5870_));
  NAND2_X1   g04868(.A1(new_n5865_), .A2(\A[206] ), .ZN(new_n5871_));
  AOI21_X1   g04869(.A1(new_n5870_), .A2(new_n5871_), .B(\A[207] ), .ZN(new_n5872_));
  NOR2_X1    g04870(.A1(new_n5866_), .A2(\A[205] ), .ZN(new_n5873_));
  OAI21_X1   g04871(.A1(new_n5865_), .A2(\A[206] ), .B(\A[207] ), .ZN(new_n5874_));
  NOR2_X1    g04872(.A1(new_n5874_), .A2(new_n5873_), .ZN(new_n5875_));
  NAND2_X1   g04873(.A1(new_n5861_), .A2(\A[208] ), .ZN(new_n5876_));
  NAND2_X1   g04874(.A1(new_n5860_), .A2(\A[209] ), .ZN(new_n5877_));
  AOI21_X1   g04875(.A1(new_n5876_), .A2(new_n5877_), .B(\A[210] ), .ZN(new_n5878_));
  INV_X1     g04876(.I(\A[210] ), .ZN(new_n5879_));
  NOR2_X1    g04877(.A1(new_n5860_), .A2(\A[209] ), .ZN(new_n5880_));
  NOR2_X1    g04878(.A1(new_n5861_), .A2(\A[208] ), .ZN(new_n5881_));
  NOR3_X1    g04879(.A1(new_n5880_), .A2(new_n5881_), .A3(new_n5879_), .ZN(new_n5882_));
  OAI22_X1   g04880(.A1(new_n5878_), .A2(new_n5882_), .B1(new_n5872_), .B2(new_n5875_), .ZN(new_n5883_));
  NOR3_X1    g04881(.A1(new_n5883_), .A2(new_n5864_), .A3(new_n5869_), .ZN(new_n5884_));
  NOR2_X1    g04882(.A1(new_n5865_), .A2(\A[206] ), .ZN(new_n5885_));
  NOR2_X1    g04883(.A1(new_n5885_), .A2(new_n5873_), .ZN(new_n5886_));
  OAI22_X1   g04884(.A1(new_n5886_), .A2(\A[207] ), .B1(new_n5873_), .B2(new_n5874_), .ZN(new_n5887_));
  AOI21_X1   g04885(.A1(\A[208] ), .A2(new_n5861_), .B(new_n5879_), .ZN(new_n5888_));
  AOI22_X1   g04886(.A1(new_n5863_), .A2(new_n5879_), .B1(new_n5877_), .B2(new_n5888_), .ZN(new_n5889_));
  NOR2_X1    g04887(.A1(new_n5887_), .A2(new_n5889_), .ZN(new_n5890_));
  NOR2_X1    g04888(.A1(new_n5872_), .A2(new_n5875_), .ZN(new_n5891_));
  OAI21_X1   g04889(.A1(new_n5880_), .A2(new_n5881_), .B(new_n5879_), .ZN(new_n5892_));
  NAND2_X1   g04890(.A1(new_n5888_), .A2(new_n5877_), .ZN(new_n5893_));
  NAND2_X1   g04891(.A1(new_n5893_), .A2(new_n5892_), .ZN(new_n5894_));
  NOR2_X1    g04892(.A1(new_n5894_), .A2(new_n5891_), .ZN(new_n5895_));
  NOR2_X1    g04893(.A1(new_n5890_), .A2(new_n5895_), .ZN(new_n5896_));
  NOR2_X1    g04894(.A1(new_n5896_), .A2(new_n5884_), .ZN(new_n5897_));
  INV_X1     g04895(.I(\A[200] ), .ZN(new_n5898_));
  NAND2_X1   g04896(.A1(new_n5898_), .A2(\A[199] ), .ZN(new_n5899_));
  INV_X1     g04897(.I(\A[199] ), .ZN(new_n5900_));
  NAND2_X1   g04898(.A1(new_n5900_), .A2(\A[200] ), .ZN(new_n5901_));
  AOI21_X1   g04899(.A1(new_n5899_), .A2(new_n5901_), .B(\A[201] ), .ZN(new_n5902_));
  INV_X1     g04900(.I(\A[201] ), .ZN(new_n5903_));
  NOR2_X1    g04901(.A1(new_n5900_), .A2(\A[200] ), .ZN(new_n5904_));
  NOR2_X1    g04902(.A1(new_n5898_), .A2(\A[199] ), .ZN(new_n5905_));
  NOR3_X1    g04903(.A1(new_n5904_), .A2(new_n5905_), .A3(new_n5903_), .ZN(new_n5906_));
  NOR2_X1    g04904(.A1(new_n5902_), .A2(new_n5906_), .ZN(new_n5907_));
  INV_X1     g04905(.I(\A[204] ), .ZN(new_n5908_));
  INV_X1     g04906(.I(\A[202] ), .ZN(new_n5909_));
  NOR2_X1    g04907(.A1(new_n5909_), .A2(\A[203] ), .ZN(new_n5910_));
  INV_X1     g04908(.I(\A[203] ), .ZN(new_n5911_));
  NOR2_X1    g04909(.A1(new_n5911_), .A2(\A[202] ), .ZN(new_n5912_));
  OAI21_X1   g04910(.A1(new_n5910_), .A2(new_n5912_), .B(new_n5908_), .ZN(new_n5913_));
  NAND2_X1   g04911(.A1(new_n5911_), .A2(\A[202] ), .ZN(new_n5914_));
  NAND2_X1   g04912(.A1(new_n5909_), .A2(\A[203] ), .ZN(new_n5915_));
  NAND3_X1   g04913(.A1(new_n5914_), .A2(new_n5915_), .A3(\A[204] ), .ZN(new_n5916_));
  NAND2_X1   g04914(.A1(new_n5913_), .A2(new_n5916_), .ZN(new_n5917_));
  NAND2_X1   g04915(.A1(new_n5907_), .A2(new_n5917_), .ZN(new_n5918_));
  XOR2_X1    g04916(.A1(\A[199] ), .A2(\A[200] ), .Z(new_n5919_));
  NAND2_X1   g04917(.A1(new_n5919_), .A2(new_n5903_), .ZN(new_n5920_));
  AOI21_X1   g04918(.A1(\A[199] ), .A2(new_n5898_), .B(new_n5903_), .ZN(new_n5921_));
  NAND2_X1   g04919(.A1(new_n5921_), .A2(new_n5901_), .ZN(new_n5922_));
  NAND2_X1   g04920(.A1(new_n5920_), .A2(new_n5922_), .ZN(new_n5923_));
  AOI21_X1   g04921(.A1(new_n5914_), .A2(new_n5915_), .B(\A[204] ), .ZN(new_n5924_));
  NOR3_X1    g04922(.A1(new_n5910_), .A2(new_n5912_), .A3(new_n5908_), .ZN(new_n5925_));
  NOR2_X1    g04923(.A1(new_n5924_), .A2(new_n5925_), .ZN(new_n5926_));
  NAND2_X1   g04924(.A1(new_n5923_), .A2(new_n5926_), .ZN(new_n5927_));
  NAND2_X1   g04925(.A1(new_n5927_), .A2(new_n5918_), .ZN(new_n5928_));
  NOR2_X1    g04926(.A1(new_n5910_), .A2(new_n5912_), .ZN(new_n5929_));
  NOR2_X1    g04927(.A1(new_n5909_), .A2(new_n5911_), .ZN(new_n5930_));
  INV_X1     g04928(.I(new_n5930_), .ZN(new_n5931_));
  OAI21_X1   g04929(.A1(new_n5929_), .A2(new_n5908_), .B(new_n5931_), .ZN(new_n5932_));
  NOR2_X1    g04930(.A1(new_n5904_), .A2(new_n5905_), .ZN(new_n5933_));
  NOR2_X1    g04931(.A1(new_n5900_), .A2(new_n5898_), .ZN(new_n5934_));
  INV_X1     g04932(.I(new_n5934_), .ZN(new_n5935_));
  OAI21_X1   g04933(.A1(new_n5933_), .A2(new_n5903_), .B(new_n5935_), .ZN(new_n5936_));
  AOI22_X1   g04934(.A1(new_n5920_), .A2(new_n5922_), .B1(new_n5913_), .B2(new_n5916_), .ZN(new_n5937_));
  NAND3_X1   g04935(.A1(new_n5937_), .A2(new_n5932_), .A3(new_n5936_), .ZN(new_n5938_));
  NAND2_X1   g04936(.A1(new_n5928_), .A2(new_n5938_), .ZN(new_n5939_));
  NAND2_X1   g04937(.A1(new_n5939_), .A2(new_n5897_), .ZN(new_n5940_));
  INV_X1     g04938(.I(new_n5862_), .ZN(new_n5941_));
  NOR2_X1    g04939(.A1(new_n5880_), .A2(new_n5881_), .ZN(new_n5942_));
  OAI21_X1   g04940(.A1(new_n5942_), .A2(new_n5879_), .B(new_n5941_), .ZN(new_n5943_));
  INV_X1     g04941(.I(\A[207] ), .ZN(new_n5944_));
  INV_X1     g04942(.I(new_n5867_), .ZN(new_n5945_));
  OAI21_X1   g04943(.A1(new_n5886_), .A2(new_n5944_), .B(new_n5945_), .ZN(new_n5946_));
  NAND2_X1   g04944(.A1(new_n5868_), .A2(new_n5944_), .ZN(new_n5947_));
  NAND3_X1   g04945(.A1(new_n5870_), .A2(new_n5871_), .A3(\A[207] ), .ZN(new_n5948_));
  AOI22_X1   g04946(.A1(new_n5947_), .A2(new_n5948_), .B1(new_n5892_), .B2(new_n5893_), .ZN(new_n5949_));
  NAND3_X1   g04947(.A1(new_n5949_), .A2(new_n5943_), .A3(new_n5946_), .ZN(new_n5950_));
  NAND2_X1   g04948(.A1(new_n5894_), .A2(new_n5891_), .ZN(new_n5951_));
  NAND2_X1   g04949(.A1(new_n5887_), .A2(new_n5889_), .ZN(new_n5952_));
  NAND2_X1   g04950(.A1(new_n5952_), .A2(new_n5951_), .ZN(new_n5953_));
  NAND2_X1   g04951(.A1(new_n5953_), .A2(new_n5950_), .ZN(new_n5954_));
  XOR2_X1    g04952(.A1(new_n5907_), .A2(new_n5917_), .Z(new_n5955_));
  XOR2_X1    g04953(.A1(\A[202] ), .A2(\A[203] ), .Z(new_n5956_));
  AOI21_X1   g04954(.A1(new_n5956_), .A2(\A[204] ), .B(new_n5930_), .ZN(new_n5957_));
  AOI21_X1   g04955(.A1(new_n5919_), .A2(\A[201] ), .B(new_n5934_), .ZN(new_n5958_));
  OAI22_X1   g04956(.A1(new_n5902_), .A2(new_n5906_), .B1(new_n5924_), .B2(new_n5925_), .ZN(new_n5959_));
  NOR3_X1    g04957(.A1(new_n5959_), .A2(new_n5957_), .A3(new_n5958_), .ZN(new_n5960_));
  NOR2_X1    g04958(.A1(new_n5955_), .A2(new_n5960_), .ZN(new_n5961_));
  NAND2_X1   g04959(.A1(new_n5961_), .A2(new_n5954_), .ZN(new_n5962_));
  NAND3_X1   g04960(.A1(new_n5859_), .A2(new_n5940_), .A3(new_n5962_), .ZN(new_n5963_));
  NAND2_X1   g04961(.A1(new_n5962_), .A2(new_n5940_), .ZN(new_n5964_));
  NAND3_X1   g04962(.A1(new_n5964_), .A2(new_n5834_), .A3(new_n5858_), .ZN(new_n5965_));
  NAND2_X1   g04963(.A1(new_n5965_), .A2(new_n5963_), .ZN(new_n5966_));
  INV_X1     g04964(.I(\A[195] ), .ZN(new_n5967_));
  INV_X1     g04965(.I(\A[193] ), .ZN(new_n5968_));
  NAND2_X1   g04966(.A1(new_n5968_), .A2(\A[194] ), .ZN(new_n5969_));
  INV_X1     g04967(.I(\A[194] ), .ZN(new_n5970_));
  AOI21_X1   g04968(.A1(\A[193] ), .A2(new_n5970_), .B(new_n5967_), .ZN(new_n5971_));
  XOR2_X1    g04969(.A1(\A[193] ), .A2(\A[194] ), .Z(new_n5972_));
  AOI22_X1   g04970(.A1(new_n5972_), .A2(new_n5967_), .B1(new_n5969_), .B2(new_n5971_), .ZN(new_n5973_));
  INV_X1     g04971(.I(\A[196] ), .ZN(new_n5974_));
  NAND2_X1   g04972(.A1(new_n5974_), .A2(\A[197] ), .ZN(new_n5975_));
  INV_X1     g04973(.I(\A[197] ), .ZN(new_n5976_));
  INV_X1     g04974(.I(\A[198] ), .ZN(new_n5977_));
  AOI21_X1   g04975(.A1(\A[196] ), .A2(new_n5976_), .B(new_n5977_), .ZN(new_n5978_));
  NAND2_X1   g04976(.A1(new_n5978_), .A2(new_n5975_), .ZN(new_n5979_));
  NOR2_X1    g04977(.A1(new_n5976_), .A2(\A[196] ), .ZN(new_n5980_));
  NOR2_X1    g04978(.A1(new_n5974_), .A2(\A[197] ), .ZN(new_n5981_));
  OAI21_X1   g04979(.A1(new_n5980_), .A2(new_n5981_), .B(new_n5977_), .ZN(new_n5982_));
  NAND2_X1   g04980(.A1(new_n5979_), .A2(new_n5982_), .ZN(new_n5983_));
  NAND2_X1   g04981(.A1(new_n5983_), .A2(new_n5973_), .ZN(new_n5984_));
  NAND2_X1   g04982(.A1(new_n5971_), .A2(new_n5969_), .ZN(new_n5985_));
  NOR2_X1    g04983(.A1(new_n5970_), .A2(\A[193] ), .ZN(new_n5986_));
  NOR2_X1    g04984(.A1(new_n5968_), .A2(\A[194] ), .ZN(new_n5987_));
  OAI21_X1   g04985(.A1(new_n5986_), .A2(new_n5987_), .B(new_n5967_), .ZN(new_n5988_));
  NAND2_X1   g04986(.A1(new_n5985_), .A2(new_n5988_), .ZN(new_n5989_));
  XOR2_X1    g04987(.A1(\A[196] ), .A2(\A[197] ), .Z(new_n5990_));
  AOI22_X1   g04988(.A1(new_n5990_), .A2(new_n5977_), .B1(new_n5975_), .B2(new_n5978_), .ZN(new_n5991_));
  NAND2_X1   g04989(.A1(new_n5989_), .A2(new_n5991_), .ZN(new_n5992_));
  NAND2_X1   g04990(.A1(new_n5984_), .A2(new_n5992_), .ZN(new_n5993_));
  NOR2_X1    g04991(.A1(new_n5980_), .A2(new_n5981_), .ZN(new_n5994_));
  NOR2_X1    g04992(.A1(new_n5974_), .A2(new_n5976_), .ZN(new_n5995_));
  INV_X1     g04993(.I(new_n5995_), .ZN(new_n5996_));
  OAI21_X1   g04994(.A1(new_n5994_), .A2(new_n5977_), .B(new_n5996_), .ZN(new_n5997_));
  NOR2_X1    g04995(.A1(new_n5986_), .A2(new_n5987_), .ZN(new_n5998_));
  NAND2_X1   g04996(.A1(\A[193] ), .A2(\A[194] ), .ZN(new_n5999_));
  OAI21_X1   g04997(.A1(new_n5998_), .A2(new_n5967_), .B(new_n5999_), .ZN(new_n6000_));
  AOI22_X1   g04998(.A1(new_n5985_), .A2(new_n5988_), .B1(new_n5979_), .B2(new_n5982_), .ZN(new_n6001_));
  NAND3_X1   g04999(.A1(new_n6001_), .A2(new_n5997_), .A3(new_n6000_), .ZN(new_n6002_));
  NAND2_X1   g05000(.A1(new_n5993_), .A2(new_n6002_), .ZN(new_n6003_));
  INV_X1     g05001(.I(\A[187] ), .ZN(new_n6004_));
  NAND2_X1   g05002(.A1(new_n6004_), .A2(\A[188] ), .ZN(new_n6005_));
  INV_X1     g05003(.I(\A[188] ), .ZN(new_n6006_));
  INV_X1     g05004(.I(\A[189] ), .ZN(new_n6007_));
  AOI21_X1   g05005(.A1(\A[187] ), .A2(new_n6006_), .B(new_n6007_), .ZN(new_n6008_));
  NAND2_X1   g05006(.A1(new_n6008_), .A2(new_n6005_), .ZN(new_n6009_));
  NOR2_X1    g05007(.A1(new_n6006_), .A2(\A[187] ), .ZN(new_n6010_));
  NOR2_X1    g05008(.A1(new_n6004_), .A2(\A[188] ), .ZN(new_n6011_));
  OAI21_X1   g05009(.A1(new_n6010_), .A2(new_n6011_), .B(new_n6007_), .ZN(new_n6012_));
  NAND2_X1   g05010(.A1(new_n6009_), .A2(new_n6012_), .ZN(new_n6013_));
  INV_X1     g05011(.I(\A[192] ), .ZN(new_n6014_));
  INV_X1     g05012(.I(\A[191] ), .ZN(new_n6015_));
  NOR2_X1    g05013(.A1(new_n6015_), .A2(\A[190] ), .ZN(new_n6016_));
  INV_X1     g05014(.I(\A[190] ), .ZN(new_n6017_));
  NOR2_X1    g05015(.A1(new_n6017_), .A2(\A[191] ), .ZN(new_n6018_));
  NOR3_X1    g05016(.A1(new_n6016_), .A2(new_n6018_), .A3(new_n6014_), .ZN(new_n6019_));
  NAND2_X1   g05017(.A1(new_n6017_), .A2(\A[191] ), .ZN(new_n6020_));
  NAND2_X1   g05018(.A1(new_n6015_), .A2(\A[190] ), .ZN(new_n6021_));
  AOI21_X1   g05019(.A1(new_n6020_), .A2(new_n6021_), .B(\A[192] ), .ZN(new_n6022_));
  NOR2_X1    g05020(.A1(new_n6022_), .A2(new_n6019_), .ZN(new_n6023_));
  NOR2_X1    g05021(.A1(new_n6023_), .A2(new_n6013_), .ZN(new_n6024_));
  NOR3_X1    g05022(.A1(new_n6010_), .A2(new_n6011_), .A3(new_n6007_), .ZN(new_n6025_));
  NAND2_X1   g05023(.A1(new_n6006_), .A2(\A[187] ), .ZN(new_n6026_));
  AOI21_X1   g05024(.A1(new_n6005_), .A2(new_n6026_), .B(\A[189] ), .ZN(new_n6027_));
  NOR2_X1    g05025(.A1(new_n6027_), .A2(new_n6025_), .ZN(new_n6028_));
  NAND3_X1   g05026(.A1(new_n6020_), .A2(new_n6021_), .A3(\A[192] ), .ZN(new_n6029_));
  OAI21_X1   g05027(.A1(new_n6016_), .A2(new_n6018_), .B(new_n6014_), .ZN(new_n6030_));
  NAND2_X1   g05028(.A1(new_n6030_), .A2(new_n6029_), .ZN(new_n6031_));
  NOR2_X1    g05029(.A1(new_n6028_), .A2(new_n6031_), .ZN(new_n6032_));
  NOR2_X1    g05030(.A1(new_n6024_), .A2(new_n6032_), .ZN(new_n6033_));
  NAND2_X1   g05031(.A1(new_n6020_), .A2(new_n6021_), .ZN(new_n6034_));
  NOR2_X1    g05032(.A1(new_n6017_), .A2(new_n6015_), .ZN(new_n6035_));
  AOI21_X1   g05033(.A1(new_n6034_), .A2(\A[192] ), .B(new_n6035_), .ZN(new_n6036_));
  NAND2_X1   g05034(.A1(new_n6005_), .A2(new_n6026_), .ZN(new_n6037_));
  NOR2_X1    g05035(.A1(new_n6004_), .A2(new_n6006_), .ZN(new_n6038_));
  AOI21_X1   g05036(.A1(new_n6037_), .A2(\A[189] ), .B(new_n6038_), .ZN(new_n6039_));
  OAI22_X1   g05037(.A1(new_n6025_), .A2(new_n6027_), .B1(new_n6022_), .B2(new_n6019_), .ZN(new_n6040_));
  NOR3_X1    g05038(.A1(new_n6040_), .A2(new_n6036_), .A3(new_n6039_), .ZN(new_n6041_));
  NOR2_X1    g05039(.A1(new_n6033_), .A2(new_n6041_), .ZN(new_n6042_));
  NAND2_X1   g05040(.A1(new_n6042_), .A2(new_n6003_), .ZN(new_n6043_));
  NOR2_X1    g05041(.A1(new_n5989_), .A2(new_n5991_), .ZN(new_n6044_));
  NOR2_X1    g05042(.A1(new_n5983_), .A2(new_n5973_), .ZN(new_n6045_));
  NOR2_X1    g05043(.A1(new_n6044_), .A2(new_n6045_), .ZN(new_n6046_));
  AOI21_X1   g05044(.A1(new_n5990_), .A2(\A[198] ), .B(new_n5995_), .ZN(new_n6047_));
  INV_X1     g05045(.I(new_n5999_), .ZN(new_n6048_));
  AOI21_X1   g05046(.A1(new_n5972_), .A2(\A[195] ), .B(new_n6048_), .ZN(new_n6049_));
  NOR3_X1    g05047(.A1(new_n5986_), .A2(new_n5987_), .A3(new_n5967_), .ZN(new_n6050_));
  NAND2_X1   g05048(.A1(new_n5970_), .A2(\A[193] ), .ZN(new_n6051_));
  AOI21_X1   g05049(.A1(new_n5969_), .A2(new_n6051_), .B(\A[195] ), .ZN(new_n6052_));
  NOR3_X1    g05050(.A1(new_n5980_), .A2(new_n5981_), .A3(new_n5977_), .ZN(new_n6053_));
  NAND2_X1   g05051(.A1(new_n5976_), .A2(\A[196] ), .ZN(new_n6054_));
  AOI21_X1   g05052(.A1(new_n5975_), .A2(new_n6054_), .B(\A[198] ), .ZN(new_n6055_));
  OAI22_X1   g05053(.A1(new_n6050_), .A2(new_n6052_), .B1(new_n6055_), .B2(new_n6053_), .ZN(new_n6056_));
  NOR3_X1    g05054(.A1(new_n6056_), .A2(new_n6047_), .A3(new_n6049_), .ZN(new_n6057_));
  NOR2_X1    g05055(.A1(new_n6046_), .A2(new_n6057_), .ZN(new_n6058_));
  NAND2_X1   g05056(.A1(new_n6028_), .A2(new_n6031_), .ZN(new_n6059_));
  NAND2_X1   g05057(.A1(new_n6023_), .A2(new_n6013_), .ZN(new_n6060_));
  NAND2_X1   g05058(.A1(new_n6060_), .A2(new_n6059_), .ZN(new_n6061_));
  NOR2_X1    g05059(.A1(new_n6016_), .A2(new_n6018_), .ZN(new_n6062_));
  INV_X1     g05060(.I(new_n6035_), .ZN(new_n6063_));
  OAI21_X1   g05061(.A1(new_n6062_), .A2(new_n6014_), .B(new_n6063_), .ZN(new_n6064_));
  NOR2_X1    g05062(.A1(new_n6010_), .A2(new_n6011_), .ZN(new_n6065_));
  INV_X1     g05063(.I(new_n6038_), .ZN(new_n6066_));
  OAI21_X1   g05064(.A1(new_n6065_), .A2(new_n6007_), .B(new_n6066_), .ZN(new_n6067_));
  AOI22_X1   g05065(.A1(new_n6009_), .A2(new_n6012_), .B1(new_n6030_), .B2(new_n6029_), .ZN(new_n6068_));
  NAND3_X1   g05066(.A1(new_n6068_), .A2(new_n6064_), .A3(new_n6067_), .ZN(new_n6069_));
  NAND2_X1   g05067(.A1(new_n6061_), .A2(new_n6069_), .ZN(new_n6070_));
  NAND2_X1   g05068(.A1(new_n6070_), .A2(new_n6058_), .ZN(new_n6071_));
  INV_X1     g05069(.I(\A[183] ), .ZN(new_n6072_));
  INV_X1     g05070(.I(\A[182] ), .ZN(new_n6073_));
  NOR2_X1    g05071(.A1(new_n6073_), .A2(\A[181] ), .ZN(new_n6074_));
  INV_X1     g05072(.I(\A[181] ), .ZN(new_n6075_));
  NOR2_X1    g05073(.A1(new_n6075_), .A2(\A[182] ), .ZN(new_n6076_));
  NOR3_X1    g05074(.A1(new_n6074_), .A2(new_n6076_), .A3(new_n6072_), .ZN(new_n6077_));
  NAND2_X1   g05075(.A1(new_n6075_), .A2(\A[182] ), .ZN(new_n6078_));
  NAND2_X1   g05076(.A1(new_n6073_), .A2(\A[181] ), .ZN(new_n6079_));
  AOI21_X1   g05077(.A1(new_n6078_), .A2(new_n6079_), .B(\A[183] ), .ZN(new_n6080_));
  NOR2_X1    g05078(.A1(new_n6080_), .A2(new_n6077_), .ZN(new_n6081_));
  INV_X1     g05079(.I(\A[184] ), .ZN(new_n6082_));
  NAND2_X1   g05080(.A1(new_n6082_), .A2(\A[185] ), .ZN(new_n6083_));
  INV_X1     g05081(.I(\A[185] ), .ZN(new_n6084_));
  NAND2_X1   g05082(.A1(new_n6084_), .A2(\A[184] ), .ZN(new_n6085_));
  NAND3_X1   g05083(.A1(new_n6083_), .A2(new_n6085_), .A3(\A[186] ), .ZN(new_n6086_));
  INV_X1     g05084(.I(\A[186] ), .ZN(new_n6087_));
  NOR2_X1    g05085(.A1(new_n6084_), .A2(\A[184] ), .ZN(new_n6088_));
  NOR2_X1    g05086(.A1(new_n6082_), .A2(\A[185] ), .ZN(new_n6089_));
  OAI21_X1   g05087(.A1(new_n6088_), .A2(new_n6089_), .B(new_n6087_), .ZN(new_n6090_));
  NAND2_X1   g05088(.A1(new_n6090_), .A2(new_n6086_), .ZN(new_n6091_));
  NAND2_X1   g05089(.A1(new_n6081_), .A2(new_n6091_), .ZN(new_n6092_));
  AOI21_X1   g05090(.A1(\A[181] ), .A2(new_n6073_), .B(new_n6072_), .ZN(new_n6093_));
  NAND2_X1   g05091(.A1(new_n6093_), .A2(new_n6078_), .ZN(new_n6094_));
  OAI21_X1   g05092(.A1(new_n6074_), .A2(new_n6076_), .B(new_n6072_), .ZN(new_n6095_));
  NAND2_X1   g05093(.A1(new_n6094_), .A2(new_n6095_), .ZN(new_n6096_));
  NOR3_X1    g05094(.A1(new_n6088_), .A2(new_n6089_), .A3(new_n6087_), .ZN(new_n6097_));
  AOI21_X1   g05095(.A1(new_n6083_), .A2(new_n6085_), .B(\A[186] ), .ZN(new_n6098_));
  NOR2_X1    g05096(.A1(new_n6098_), .A2(new_n6097_), .ZN(new_n6099_));
  NAND2_X1   g05097(.A1(new_n6099_), .A2(new_n6096_), .ZN(new_n6100_));
  NAND2_X1   g05098(.A1(new_n6100_), .A2(new_n6092_), .ZN(new_n6101_));
  NOR2_X1    g05099(.A1(new_n6088_), .A2(new_n6089_), .ZN(new_n6102_));
  NOR2_X1    g05100(.A1(new_n6082_), .A2(new_n6084_), .ZN(new_n6103_));
  INV_X1     g05101(.I(new_n6103_), .ZN(new_n6104_));
  OAI21_X1   g05102(.A1(new_n6102_), .A2(new_n6087_), .B(new_n6104_), .ZN(new_n6105_));
  NOR2_X1    g05103(.A1(new_n6074_), .A2(new_n6076_), .ZN(new_n6106_));
  NOR2_X1    g05104(.A1(new_n6075_), .A2(new_n6073_), .ZN(new_n6107_));
  INV_X1     g05105(.I(new_n6107_), .ZN(new_n6108_));
  OAI21_X1   g05106(.A1(new_n6106_), .A2(new_n6072_), .B(new_n6108_), .ZN(new_n6109_));
  AOI22_X1   g05107(.A1(new_n6094_), .A2(new_n6095_), .B1(new_n6090_), .B2(new_n6086_), .ZN(new_n6110_));
  NAND3_X1   g05108(.A1(new_n6110_), .A2(new_n6105_), .A3(new_n6109_), .ZN(new_n6111_));
  NAND2_X1   g05109(.A1(new_n6101_), .A2(new_n6111_), .ZN(new_n6112_));
  INV_X1     g05110(.I(\A[175] ), .ZN(new_n6113_));
  NAND2_X1   g05111(.A1(new_n6113_), .A2(\A[176] ), .ZN(new_n6114_));
  INV_X1     g05112(.I(\A[176] ), .ZN(new_n6115_));
  INV_X1     g05113(.I(\A[177] ), .ZN(new_n6116_));
  AOI21_X1   g05114(.A1(\A[175] ), .A2(new_n6115_), .B(new_n6116_), .ZN(new_n6117_));
  NAND2_X1   g05115(.A1(new_n6117_), .A2(new_n6114_), .ZN(new_n6118_));
  NOR2_X1    g05116(.A1(new_n6115_), .A2(\A[175] ), .ZN(new_n6119_));
  NOR2_X1    g05117(.A1(new_n6113_), .A2(\A[176] ), .ZN(new_n6120_));
  OAI21_X1   g05118(.A1(new_n6119_), .A2(new_n6120_), .B(new_n6116_), .ZN(new_n6121_));
  NAND2_X1   g05119(.A1(new_n6118_), .A2(new_n6121_), .ZN(new_n6122_));
  INV_X1     g05120(.I(\A[180] ), .ZN(new_n6123_));
  INV_X1     g05121(.I(\A[179] ), .ZN(new_n6124_));
  NOR2_X1    g05122(.A1(new_n6124_), .A2(\A[178] ), .ZN(new_n6125_));
  INV_X1     g05123(.I(\A[178] ), .ZN(new_n6126_));
  NOR2_X1    g05124(.A1(new_n6126_), .A2(\A[179] ), .ZN(new_n6127_));
  NOR3_X1    g05125(.A1(new_n6125_), .A2(new_n6127_), .A3(new_n6123_), .ZN(new_n6128_));
  NAND2_X1   g05126(.A1(new_n6126_), .A2(\A[179] ), .ZN(new_n6129_));
  NAND2_X1   g05127(.A1(new_n6124_), .A2(\A[178] ), .ZN(new_n6130_));
  AOI21_X1   g05128(.A1(new_n6129_), .A2(new_n6130_), .B(\A[180] ), .ZN(new_n6131_));
  NOR2_X1    g05129(.A1(new_n6131_), .A2(new_n6128_), .ZN(new_n6132_));
  NOR2_X1    g05130(.A1(new_n6132_), .A2(new_n6122_), .ZN(new_n6133_));
  NOR3_X1    g05131(.A1(new_n6119_), .A2(new_n6120_), .A3(new_n6116_), .ZN(new_n6134_));
  NAND2_X1   g05132(.A1(new_n6115_), .A2(\A[175] ), .ZN(new_n6135_));
  AOI21_X1   g05133(.A1(new_n6114_), .A2(new_n6135_), .B(\A[177] ), .ZN(new_n6136_));
  NOR2_X1    g05134(.A1(new_n6136_), .A2(new_n6134_), .ZN(new_n6137_));
  NAND3_X1   g05135(.A1(new_n6129_), .A2(new_n6130_), .A3(\A[180] ), .ZN(new_n6138_));
  OAI21_X1   g05136(.A1(new_n6125_), .A2(new_n6127_), .B(new_n6123_), .ZN(new_n6139_));
  NAND2_X1   g05137(.A1(new_n6139_), .A2(new_n6138_), .ZN(new_n6140_));
  NOR2_X1    g05138(.A1(new_n6137_), .A2(new_n6140_), .ZN(new_n6141_));
  NOR2_X1    g05139(.A1(new_n6133_), .A2(new_n6141_), .ZN(new_n6142_));
  NAND2_X1   g05140(.A1(new_n6129_), .A2(new_n6130_), .ZN(new_n6143_));
  NOR2_X1    g05141(.A1(new_n6126_), .A2(new_n6124_), .ZN(new_n6144_));
  AOI21_X1   g05142(.A1(new_n6143_), .A2(\A[180] ), .B(new_n6144_), .ZN(new_n6145_));
  NAND2_X1   g05143(.A1(new_n6114_), .A2(new_n6135_), .ZN(new_n6146_));
  NOR2_X1    g05144(.A1(new_n6113_), .A2(new_n6115_), .ZN(new_n6147_));
  AOI21_X1   g05145(.A1(new_n6146_), .A2(\A[177] ), .B(new_n6147_), .ZN(new_n6148_));
  OAI22_X1   g05146(.A1(new_n6134_), .A2(new_n6136_), .B1(new_n6131_), .B2(new_n6128_), .ZN(new_n6149_));
  NOR3_X1    g05147(.A1(new_n6149_), .A2(new_n6145_), .A3(new_n6148_), .ZN(new_n6150_));
  NOR2_X1    g05148(.A1(new_n6142_), .A2(new_n6150_), .ZN(new_n6151_));
  NAND2_X1   g05149(.A1(new_n6151_), .A2(new_n6112_), .ZN(new_n6152_));
  NOR2_X1    g05150(.A1(new_n6099_), .A2(new_n6096_), .ZN(new_n6153_));
  NOR2_X1    g05151(.A1(new_n6081_), .A2(new_n6091_), .ZN(new_n6154_));
  NOR2_X1    g05152(.A1(new_n6153_), .A2(new_n6154_), .ZN(new_n6155_));
  NAND2_X1   g05153(.A1(new_n6083_), .A2(new_n6085_), .ZN(new_n6156_));
  AOI21_X1   g05154(.A1(new_n6156_), .A2(\A[186] ), .B(new_n6103_), .ZN(new_n6157_));
  NAND2_X1   g05155(.A1(new_n6078_), .A2(new_n6079_), .ZN(new_n6158_));
  AOI21_X1   g05156(.A1(new_n6158_), .A2(\A[183] ), .B(new_n6107_), .ZN(new_n6159_));
  OAI22_X1   g05157(.A1(new_n6077_), .A2(new_n6080_), .B1(new_n6098_), .B2(new_n6097_), .ZN(new_n6160_));
  NOR3_X1    g05158(.A1(new_n6160_), .A2(new_n6157_), .A3(new_n6159_), .ZN(new_n6161_));
  NOR2_X1    g05159(.A1(new_n6155_), .A2(new_n6161_), .ZN(new_n6162_));
  INV_X1     g05160(.I(new_n6151_), .ZN(new_n6163_));
  NAND2_X1   g05161(.A1(new_n6163_), .A2(new_n6162_), .ZN(new_n6164_));
  NAND2_X1   g05162(.A1(new_n6164_), .A2(new_n6152_), .ZN(new_n6165_));
  NAND3_X1   g05163(.A1(new_n6165_), .A2(new_n6043_), .A3(new_n6071_), .ZN(new_n6166_));
  NAND2_X1   g05164(.A1(new_n6071_), .A2(new_n6043_), .ZN(new_n6167_));
  NAND3_X1   g05165(.A1(new_n6167_), .A2(new_n6152_), .A3(new_n6164_), .ZN(new_n6168_));
  NAND2_X1   g05166(.A1(new_n6166_), .A2(new_n6168_), .ZN(new_n6169_));
  XOR2_X1    g05167(.A1(new_n6169_), .A2(new_n5966_), .Z(new_n6170_));
  INV_X1     g05168(.I(\A[270] ), .ZN(new_n6171_));
  INV_X1     g05169(.I(\A[268] ), .ZN(new_n6172_));
  INV_X1     g05170(.I(\A[269] ), .ZN(new_n6173_));
  NOR2_X1    g05171(.A1(new_n6172_), .A2(new_n6173_), .ZN(new_n6174_));
  INV_X1     g05172(.I(new_n6174_), .ZN(new_n6175_));
  NOR2_X1    g05173(.A1(new_n6172_), .A2(\A[269] ), .ZN(new_n6176_));
  NOR2_X1    g05174(.A1(new_n6173_), .A2(\A[268] ), .ZN(new_n6177_));
  NOR2_X1    g05175(.A1(new_n6176_), .A2(new_n6177_), .ZN(new_n6178_));
  OAI21_X1   g05176(.A1(new_n6178_), .A2(new_n6171_), .B(new_n6175_), .ZN(new_n6179_));
  INV_X1     g05177(.I(\A[267] ), .ZN(new_n6180_));
  NAND2_X1   g05178(.A1(\A[265] ), .A2(\A[266] ), .ZN(new_n6181_));
  XNOR2_X1   g05179(.A1(\A[265] ), .A2(\A[266] ), .ZN(new_n6182_));
  OAI21_X1   g05180(.A1(new_n6182_), .A2(new_n6180_), .B(new_n6181_), .ZN(new_n6183_));
  INV_X1     g05181(.I(\A[265] ), .ZN(new_n6184_));
  NOR2_X1    g05182(.A1(new_n6184_), .A2(\A[266] ), .ZN(new_n6185_));
  INV_X1     g05183(.I(\A[266] ), .ZN(new_n6186_));
  NOR2_X1    g05184(.A1(new_n6186_), .A2(\A[265] ), .ZN(new_n6187_));
  OAI21_X1   g05185(.A1(new_n6185_), .A2(new_n6187_), .B(new_n6180_), .ZN(new_n6188_));
  NAND2_X1   g05186(.A1(new_n6186_), .A2(\A[265] ), .ZN(new_n6189_));
  NAND2_X1   g05187(.A1(new_n6184_), .A2(\A[266] ), .ZN(new_n6190_));
  NAND3_X1   g05188(.A1(new_n6189_), .A2(new_n6190_), .A3(\A[267] ), .ZN(new_n6191_));
  OAI21_X1   g05189(.A1(new_n6176_), .A2(new_n6177_), .B(new_n6171_), .ZN(new_n6192_));
  NAND2_X1   g05190(.A1(new_n6173_), .A2(\A[268] ), .ZN(new_n6193_));
  NAND2_X1   g05191(.A1(new_n6172_), .A2(\A[269] ), .ZN(new_n6194_));
  NAND3_X1   g05192(.A1(new_n6193_), .A2(new_n6194_), .A3(\A[270] ), .ZN(new_n6195_));
  AOI22_X1   g05193(.A1(new_n6188_), .A2(new_n6191_), .B1(new_n6192_), .B2(new_n6195_), .ZN(new_n6196_));
  NAND3_X1   g05194(.A1(new_n6196_), .A2(new_n6179_), .A3(new_n6183_), .ZN(new_n6197_));
  NAND2_X1   g05195(.A1(new_n6188_), .A2(new_n6191_), .ZN(new_n6198_));
  AOI21_X1   g05196(.A1(new_n6193_), .A2(new_n6194_), .B(\A[270] ), .ZN(new_n6199_));
  OAI21_X1   g05197(.A1(new_n6172_), .A2(\A[269] ), .B(\A[270] ), .ZN(new_n6200_));
  NOR2_X1    g05198(.A1(new_n6200_), .A2(new_n6177_), .ZN(new_n6201_));
  NOR2_X1    g05199(.A1(new_n6199_), .A2(new_n6201_), .ZN(new_n6202_));
  NAND2_X1   g05200(.A1(new_n6198_), .A2(new_n6202_), .ZN(new_n6203_));
  AOI21_X1   g05201(.A1(new_n6189_), .A2(new_n6190_), .B(\A[267] ), .ZN(new_n6204_));
  NOR3_X1    g05202(.A1(new_n6185_), .A2(new_n6187_), .A3(new_n6180_), .ZN(new_n6205_));
  NOR2_X1    g05203(.A1(new_n6204_), .A2(new_n6205_), .ZN(new_n6206_));
  NAND2_X1   g05204(.A1(new_n6192_), .A2(new_n6195_), .ZN(new_n6207_));
  NAND2_X1   g05205(.A1(new_n6206_), .A2(new_n6207_), .ZN(new_n6208_));
  NAND2_X1   g05206(.A1(new_n6208_), .A2(new_n6203_), .ZN(new_n6209_));
  NAND2_X1   g05207(.A1(new_n6209_), .A2(new_n6197_), .ZN(new_n6210_));
  INV_X1     g05208(.I(\A[264] ), .ZN(new_n6211_));
  NAND2_X1   g05209(.A1(\A[262] ), .A2(\A[263] ), .ZN(new_n6212_));
  XNOR2_X1   g05210(.A1(\A[262] ), .A2(\A[263] ), .ZN(new_n6213_));
  OAI21_X1   g05211(.A1(new_n6213_), .A2(new_n6211_), .B(new_n6212_), .ZN(new_n6214_));
  INV_X1     g05212(.I(\A[261] ), .ZN(new_n6215_));
  NAND2_X1   g05213(.A1(\A[259] ), .A2(\A[260] ), .ZN(new_n6216_));
  XNOR2_X1   g05214(.A1(\A[259] ), .A2(\A[260] ), .ZN(new_n6217_));
  OAI21_X1   g05215(.A1(new_n6217_), .A2(new_n6215_), .B(new_n6216_), .ZN(new_n6218_));
  INV_X1     g05216(.I(\A[260] ), .ZN(new_n6219_));
  NOR2_X1    g05217(.A1(new_n6219_), .A2(\A[259] ), .ZN(new_n6220_));
  INV_X1     g05218(.I(\A[259] ), .ZN(new_n6221_));
  OAI21_X1   g05219(.A1(new_n6221_), .A2(\A[260] ), .B(\A[261] ), .ZN(new_n6222_));
  OAI22_X1   g05220(.A1(new_n6217_), .A2(\A[261] ), .B1(new_n6220_), .B2(new_n6222_), .ZN(new_n6223_));
  INV_X1     g05221(.I(\A[263] ), .ZN(new_n6224_));
  NOR2_X1    g05222(.A1(new_n6224_), .A2(\A[262] ), .ZN(new_n6225_));
  INV_X1     g05223(.I(\A[262] ), .ZN(new_n6226_));
  OAI21_X1   g05224(.A1(new_n6226_), .A2(\A[263] ), .B(\A[264] ), .ZN(new_n6227_));
  OAI22_X1   g05225(.A1(new_n6213_), .A2(\A[264] ), .B1(new_n6225_), .B2(new_n6227_), .ZN(new_n6228_));
  NAND4_X1   g05226(.A1(new_n6228_), .A2(new_n6223_), .A3(new_n6214_), .A4(new_n6218_), .ZN(new_n6229_));
  INV_X1     g05227(.I(new_n6229_), .ZN(new_n6230_));
  NAND2_X1   g05228(.A1(new_n6226_), .A2(\A[263] ), .ZN(new_n6231_));
  XOR2_X1    g05229(.A1(\A[262] ), .A2(\A[263] ), .Z(new_n6232_));
  AOI21_X1   g05230(.A1(\A[262] ), .A2(new_n6224_), .B(new_n6211_), .ZN(new_n6233_));
  AOI22_X1   g05231(.A1(new_n6232_), .A2(new_n6211_), .B1(new_n6231_), .B2(new_n6233_), .ZN(new_n6234_));
  XOR2_X1    g05232(.A1(new_n6223_), .A2(new_n6234_), .Z(new_n6235_));
  NOR2_X1    g05233(.A1(new_n6235_), .A2(new_n6230_), .ZN(new_n6236_));
  NOR2_X1    g05234(.A1(new_n6236_), .A2(new_n6210_), .ZN(new_n6237_));
  XOR2_X1    g05235(.A1(\A[268] ), .A2(\A[269] ), .Z(new_n6238_));
  AOI21_X1   g05236(.A1(new_n6238_), .A2(\A[270] ), .B(new_n6174_), .ZN(new_n6239_));
  INV_X1     g05237(.I(new_n6181_), .ZN(new_n6240_));
  XOR2_X1    g05238(.A1(\A[265] ), .A2(\A[266] ), .Z(new_n6241_));
  AOI21_X1   g05239(.A1(new_n6241_), .A2(\A[267] ), .B(new_n6240_), .ZN(new_n6242_));
  OAI22_X1   g05240(.A1(new_n6204_), .A2(new_n6205_), .B1(new_n6199_), .B2(new_n6201_), .ZN(new_n6243_));
  NOR3_X1    g05241(.A1(new_n6243_), .A2(new_n6239_), .A3(new_n6242_), .ZN(new_n6244_));
  NOR2_X1    g05242(.A1(new_n6206_), .A2(new_n6207_), .ZN(new_n6245_));
  NOR2_X1    g05243(.A1(new_n6198_), .A2(new_n6202_), .ZN(new_n6246_));
  NOR2_X1    g05244(.A1(new_n6245_), .A2(new_n6246_), .ZN(new_n6247_));
  NOR2_X1    g05245(.A1(new_n6247_), .A2(new_n6244_), .ZN(new_n6248_));
  NAND2_X1   g05246(.A1(new_n6219_), .A2(\A[259] ), .ZN(new_n6249_));
  NAND2_X1   g05247(.A1(new_n6221_), .A2(\A[260] ), .ZN(new_n6250_));
  AOI21_X1   g05248(.A1(new_n6249_), .A2(new_n6250_), .B(\A[261] ), .ZN(new_n6251_));
  NOR2_X1    g05249(.A1(new_n6222_), .A2(new_n6220_), .ZN(new_n6252_));
  NOR2_X1    g05250(.A1(new_n6251_), .A2(new_n6252_), .ZN(new_n6253_));
  NAND2_X1   g05251(.A1(new_n6228_), .A2(new_n6253_), .ZN(new_n6254_));
  NAND2_X1   g05252(.A1(new_n6223_), .A2(new_n6234_), .ZN(new_n6255_));
  NAND2_X1   g05253(.A1(new_n6254_), .A2(new_n6255_), .ZN(new_n6256_));
  NAND2_X1   g05254(.A1(new_n6256_), .A2(new_n6229_), .ZN(new_n6257_));
  NOR2_X1    g05255(.A1(new_n6248_), .A2(new_n6257_), .ZN(new_n6258_));
  NOR2_X1    g05256(.A1(new_n6237_), .A2(new_n6258_), .ZN(new_n6259_));
  INV_X1     g05257(.I(\A[258] ), .ZN(new_n6260_));
  INV_X1     g05258(.I(\A[256] ), .ZN(new_n6261_));
  INV_X1     g05259(.I(\A[257] ), .ZN(new_n6262_));
  NOR2_X1    g05260(.A1(new_n6261_), .A2(new_n6262_), .ZN(new_n6263_));
  INV_X1     g05261(.I(new_n6263_), .ZN(new_n6264_));
  NOR2_X1    g05262(.A1(new_n6261_), .A2(\A[257] ), .ZN(new_n6265_));
  NOR2_X1    g05263(.A1(new_n6262_), .A2(\A[256] ), .ZN(new_n6266_));
  NOR2_X1    g05264(.A1(new_n6265_), .A2(new_n6266_), .ZN(new_n6267_));
  OAI21_X1   g05265(.A1(new_n6267_), .A2(new_n6260_), .B(new_n6264_), .ZN(new_n6268_));
  INV_X1     g05266(.I(\A[255] ), .ZN(new_n6269_));
  INV_X1     g05267(.I(\A[253] ), .ZN(new_n6270_));
  INV_X1     g05268(.I(\A[254] ), .ZN(new_n6271_));
  NOR2_X1    g05269(.A1(new_n6270_), .A2(new_n6271_), .ZN(new_n6272_));
  INV_X1     g05270(.I(new_n6272_), .ZN(new_n6273_));
  NOR2_X1    g05271(.A1(new_n6270_), .A2(\A[254] ), .ZN(new_n6274_));
  NOR2_X1    g05272(.A1(new_n6271_), .A2(\A[253] ), .ZN(new_n6275_));
  NOR2_X1    g05273(.A1(new_n6274_), .A2(new_n6275_), .ZN(new_n6276_));
  OAI21_X1   g05274(.A1(new_n6276_), .A2(new_n6269_), .B(new_n6273_), .ZN(new_n6277_));
  OAI21_X1   g05275(.A1(new_n6274_), .A2(new_n6275_), .B(new_n6269_), .ZN(new_n6278_));
  NAND2_X1   g05276(.A1(new_n6271_), .A2(\A[253] ), .ZN(new_n6279_));
  NAND2_X1   g05277(.A1(new_n6270_), .A2(\A[254] ), .ZN(new_n6280_));
  NAND3_X1   g05278(.A1(new_n6279_), .A2(new_n6280_), .A3(\A[255] ), .ZN(new_n6281_));
  OAI21_X1   g05279(.A1(new_n6265_), .A2(new_n6266_), .B(new_n6260_), .ZN(new_n6282_));
  NAND2_X1   g05280(.A1(new_n6262_), .A2(\A[256] ), .ZN(new_n6283_));
  NAND2_X1   g05281(.A1(new_n6261_), .A2(\A[257] ), .ZN(new_n6284_));
  NAND3_X1   g05282(.A1(new_n6283_), .A2(new_n6284_), .A3(\A[258] ), .ZN(new_n6285_));
  AOI22_X1   g05283(.A1(new_n6278_), .A2(new_n6281_), .B1(new_n6282_), .B2(new_n6285_), .ZN(new_n6286_));
  NAND3_X1   g05284(.A1(new_n6286_), .A2(new_n6268_), .A3(new_n6277_), .ZN(new_n6287_));
  NAND2_X1   g05285(.A1(new_n6278_), .A2(new_n6281_), .ZN(new_n6288_));
  AOI21_X1   g05286(.A1(new_n6283_), .A2(new_n6284_), .B(\A[258] ), .ZN(new_n6289_));
  NOR3_X1    g05287(.A1(new_n6265_), .A2(new_n6266_), .A3(new_n6260_), .ZN(new_n6290_));
  NOR2_X1    g05288(.A1(new_n6289_), .A2(new_n6290_), .ZN(new_n6291_));
  NAND2_X1   g05289(.A1(new_n6291_), .A2(new_n6288_), .ZN(new_n6292_));
  AOI21_X1   g05290(.A1(new_n6279_), .A2(new_n6280_), .B(\A[255] ), .ZN(new_n6293_));
  NOR3_X1    g05291(.A1(new_n6274_), .A2(new_n6275_), .A3(new_n6269_), .ZN(new_n6294_));
  NOR2_X1    g05292(.A1(new_n6293_), .A2(new_n6294_), .ZN(new_n6295_));
  NAND2_X1   g05293(.A1(new_n6282_), .A2(new_n6285_), .ZN(new_n6296_));
  NAND2_X1   g05294(.A1(new_n6295_), .A2(new_n6296_), .ZN(new_n6297_));
  NAND2_X1   g05295(.A1(new_n6297_), .A2(new_n6292_), .ZN(new_n6298_));
  NAND2_X1   g05296(.A1(new_n6298_), .A2(new_n6287_), .ZN(new_n6299_));
  INV_X1     g05297(.I(\A[252] ), .ZN(new_n6300_));
  INV_X1     g05298(.I(\A[250] ), .ZN(new_n6301_));
  INV_X1     g05299(.I(\A[251] ), .ZN(new_n6302_));
  NOR2_X1    g05300(.A1(new_n6301_), .A2(new_n6302_), .ZN(new_n6303_));
  INV_X1     g05301(.I(new_n6303_), .ZN(new_n6304_));
  NOR2_X1    g05302(.A1(new_n6301_), .A2(\A[251] ), .ZN(new_n6305_));
  NOR2_X1    g05303(.A1(new_n6302_), .A2(\A[250] ), .ZN(new_n6306_));
  NOR2_X1    g05304(.A1(new_n6305_), .A2(new_n6306_), .ZN(new_n6307_));
  OAI21_X1   g05305(.A1(new_n6307_), .A2(new_n6300_), .B(new_n6304_), .ZN(new_n6308_));
  INV_X1     g05306(.I(\A[249] ), .ZN(new_n6309_));
  INV_X1     g05307(.I(\A[247] ), .ZN(new_n6310_));
  INV_X1     g05308(.I(\A[248] ), .ZN(new_n6311_));
  NOR2_X1    g05309(.A1(new_n6310_), .A2(new_n6311_), .ZN(new_n6312_));
  INV_X1     g05310(.I(new_n6312_), .ZN(new_n6313_));
  NOR2_X1    g05311(.A1(new_n6310_), .A2(\A[248] ), .ZN(new_n6314_));
  NOR2_X1    g05312(.A1(new_n6311_), .A2(\A[247] ), .ZN(new_n6315_));
  NOR2_X1    g05313(.A1(new_n6314_), .A2(new_n6315_), .ZN(new_n6316_));
  OAI21_X1   g05314(.A1(new_n6316_), .A2(new_n6309_), .B(new_n6313_), .ZN(new_n6317_));
  NAND2_X1   g05315(.A1(new_n6311_), .A2(\A[247] ), .ZN(new_n6318_));
  NAND2_X1   g05316(.A1(new_n6318_), .A2(\A[249] ), .ZN(new_n6319_));
  OAI22_X1   g05317(.A1(new_n6316_), .A2(\A[249] ), .B1(new_n6319_), .B2(new_n6315_), .ZN(new_n6320_));
  NAND2_X1   g05318(.A1(new_n6302_), .A2(\A[250] ), .ZN(new_n6321_));
  NAND2_X1   g05319(.A1(new_n6321_), .A2(\A[252] ), .ZN(new_n6322_));
  OAI22_X1   g05320(.A1(new_n6307_), .A2(\A[252] ), .B1(new_n6322_), .B2(new_n6306_), .ZN(new_n6323_));
  NAND4_X1   g05321(.A1(new_n6323_), .A2(new_n6320_), .A3(new_n6308_), .A4(new_n6317_), .ZN(new_n6324_));
  NAND2_X1   g05322(.A1(new_n6310_), .A2(\A[248] ), .ZN(new_n6325_));
  AOI21_X1   g05323(.A1(new_n6318_), .A2(new_n6325_), .B(\A[249] ), .ZN(new_n6326_));
  NOR3_X1    g05324(.A1(new_n6314_), .A2(new_n6315_), .A3(new_n6309_), .ZN(new_n6327_));
  NOR2_X1    g05325(.A1(new_n6326_), .A2(new_n6327_), .ZN(new_n6328_));
  NAND2_X1   g05326(.A1(new_n6323_), .A2(new_n6328_), .ZN(new_n6329_));
  NAND2_X1   g05327(.A1(new_n6301_), .A2(\A[251] ), .ZN(new_n6330_));
  AOI21_X1   g05328(.A1(new_n6321_), .A2(new_n6330_), .B(\A[252] ), .ZN(new_n6331_));
  NOR3_X1    g05329(.A1(new_n6305_), .A2(new_n6306_), .A3(new_n6300_), .ZN(new_n6332_));
  NOR2_X1    g05330(.A1(new_n6331_), .A2(new_n6332_), .ZN(new_n6333_));
  NAND2_X1   g05331(.A1(new_n6320_), .A2(new_n6333_), .ZN(new_n6334_));
  NAND2_X1   g05332(.A1(new_n6329_), .A2(new_n6334_), .ZN(new_n6335_));
  NAND3_X1   g05333(.A1(new_n6299_), .A2(new_n6324_), .A3(new_n6335_), .ZN(new_n6336_));
  XOR2_X1    g05334(.A1(\A[256] ), .A2(\A[257] ), .Z(new_n6337_));
  AOI21_X1   g05335(.A1(new_n6337_), .A2(\A[258] ), .B(new_n6263_), .ZN(new_n6338_));
  NAND2_X1   g05336(.A1(new_n6279_), .A2(new_n6280_), .ZN(new_n6339_));
  AOI21_X1   g05337(.A1(new_n6339_), .A2(\A[255] ), .B(new_n6272_), .ZN(new_n6340_));
  OAI22_X1   g05338(.A1(new_n6293_), .A2(new_n6294_), .B1(new_n6289_), .B2(new_n6290_), .ZN(new_n6341_));
  NOR3_X1    g05339(.A1(new_n6341_), .A2(new_n6338_), .A3(new_n6340_), .ZN(new_n6342_));
  NOR2_X1    g05340(.A1(new_n6295_), .A2(new_n6296_), .ZN(new_n6343_));
  NOR2_X1    g05341(.A1(new_n6291_), .A2(new_n6288_), .ZN(new_n6344_));
  NOR2_X1    g05342(.A1(new_n6343_), .A2(new_n6344_), .ZN(new_n6345_));
  NOR2_X1    g05343(.A1(new_n6345_), .A2(new_n6342_), .ZN(new_n6346_));
  NAND2_X1   g05344(.A1(new_n6335_), .A2(new_n6324_), .ZN(new_n6347_));
  NAND2_X1   g05345(.A1(new_n6347_), .A2(new_n6346_), .ZN(new_n6348_));
  NAND2_X1   g05346(.A1(new_n6348_), .A2(new_n6336_), .ZN(new_n6349_));
  NOR2_X1    g05347(.A1(new_n6349_), .A2(new_n6259_), .ZN(new_n6350_));
  NAND2_X1   g05348(.A1(new_n6248_), .A2(new_n6257_), .ZN(new_n6351_));
  NAND2_X1   g05349(.A1(new_n6236_), .A2(new_n6210_), .ZN(new_n6352_));
  NAND2_X1   g05350(.A1(new_n6352_), .A2(new_n6351_), .ZN(new_n6353_));
  NOR2_X1    g05351(.A1(new_n6347_), .A2(new_n6346_), .ZN(new_n6354_));
  AOI21_X1   g05352(.A1(new_n6324_), .A2(new_n6335_), .B(new_n6299_), .ZN(new_n6355_));
  NOR2_X1    g05353(.A1(new_n6355_), .A2(new_n6354_), .ZN(new_n6356_));
  NOR2_X1    g05354(.A1(new_n6356_), .A2(new_n6353_), .ZN(new_n6357_));
  NOR2_X1    g05355(.A1(new_n6357_), .A2(new_n6350_), .ZN(new_n6358_));
  INV_X1     g05356(.I(\A[243] ), .ZN(new_n6359_));
  XOR2_X1    g05357(.A1(\A[241] ), .A2(\A[242] ), .Z(new_n6360_));
  NAND2_X1   g05358(.A1(new_n6360_), .A2(new_n6359_), .ZN(new_n6361_));
  INV_X1     g05359(.I(\A[242] ), .ZN(new_n6362_));
  NAND2_X1   g05360(.A1(new_n6362_), .A2(\A[241] ), .ZN(new_n6363_));
  INV_X1     g05361(.I(\A[241] ), .ZN(new_n6364_));
  NAND2_X1   g05362(.A1(new_n6364_), .A2(\A[242] ), .ZN(new_n6365_));
  NAND3_X1   g05363(.A1(new_n6363_), .A2(new_n6365_), .A3(\A[243] ), .ZN(new_n6366_));
  NAND2_X1   g05364(.A1(new_n6361_), .A2(new_n6366_), .ZN(new_n6367_));
  INV_X1     g05365(.I(\A[245] ), .ZN(new_n6368_));
  NAND2_X1   g05366(.A1(new_n6368_), .A2(\A[244] ), .ZN(new_n6369_));
  INV_X1     g05367(.I(\A[244] ), .ZN(new_n6370_));
  NAND2_X1   g05368(.A1(new_n6370_), .A2(\A[245] ), .ZN(new_n6371_));
  AOI21_X1   g05369(.A1(new_n6369_), .A2(new_n6371_), .B(\A[246] ), .ZN(new_n6372_));
  INV_X1     g05370(.I(\A[246] ), .ZN(new_n6373_));
  NOR2_X1    g05371(.A1(new_n6370_), .A2(\A[245] ), .ZN(new_n6374_));
  NOR2_X1    g05372(.A1(new_n6368_), .A2(\A[244] ), .ZN(new_n6375_));
  NOR3_X1    g05373(.A1(new_n6374_), .A2(new_n6375_), .A3(new_n6373_), .ZN(new_n6376_));
  NOR2_X1    g05374(.A1(new_n6372_), .A2(new_n6376_), .ZN(new_n6377_));
  NOR2_X1    g05375(.A1(new_n6367_), .A2(new_n6377_), .ZN(new_n6378_));
  AOI21_X1   g05376(.A1(new_n6363_), .A2(new_n6365_), .B(\A[243] ), .ZN(new_n6379_));
  NOR2_X1    g05377(.A1(new_n6362_), .A2(\A[241] ), .ZN(new_n6380_));
  OAI21_X1   g05378(.A1(new_n6364_), .A2(\A[242] ), .B(\A[243] ), .ZN(new_n6381_));
  NOR2_X1    g05379(.A1(new_n6381_), .A2(new_n6380_), .ZN(new_n6382_));
  NOR2_X1    g05380(.A1(new_n6379_), .A2(new_n6382_), .ZN(new_n6383_));
  OAI21_X1   g05381(.A1(new_n6374_), .A2(new_n6375_), .B(new_n6373_), .ZN(new_n6384_));
  NAND3_X1   g05382(.A1(new_n6369_), .A2(new_n6371_), .A3(\A[246] ), .ZN(new_n6385_));
  NAND2_X1   g05383(.A1(new_n6384_), .A2(new_n6385_), .ZN(new_n6386_));
  NOR2_X1    g05384(.A1(new_n6386_), .A2(new_n6383_), .ZN(new_n6387_));
  NOR2_X1    g05385(.A1(new_n6378_), .A2(new_n6387_), .ZN(new_n6388_));
  XOR2_X1    g05386(.A1(\A[244] ), .A2(\A[245] ), .Z(new_n6389_));
  NOR2_X1    g05387(.A1(new_n6370_), .A2(new_n6368_), .ZN(new_n6390_));
  AOI21_X1   g05388(.A1(new_n6389_), .A2(\A[246] ), .B(new_n6390_), .ZN(new_n6391_));
  NOR2_X1    g05389(.A1(new_n6364_), .A2(new_n6362_), .ZN(new_n6392_));
  AOI21_X1   g05390(.A1(new_n6360_), .A2(\A[243] ), .B(new_n6392_), .ZN(new_n6393_));
  OAI22_X1   g05391(.A1(new_n6372_), .A2(new_n6376_), .B1(new_n6379_), .B2(new_n6382_), .ZN(new_n6394_));
  NOR3_X1    g05392(.A1(new_n6394_), .A2(new_n6391_), .A3(new_n6393_), .ZN(new_n6395_));
  NOR2_X1    g05393(.A1(new_n6388_), .A2(new_n6395_), .ZN(new_n6396_));
  INV_X1     g05394(.I(\A[236] ), .ZN(new_n6397_));
  NAND2_X1   g05395(.A1(new_n6397_), .A2(\A[235] ), .ZN(new_n6398_));
  INV_X1     g05396(.I(\A[235] ), .ZN(new_n6399_));
  NAND2_X1   g05397(.A1(new_n6399_), .A2(\A[236] ), .ZN(new_n6400_));
  AOI21_X1   g05398(.A1(new_n6398_), .A2(new_n6400_), .B(\A[237] ), .ZN(new_n6401_));
  NOR2_X1    g05399(.A1(new_n6397_), .A2(\A[235] ), .ZN(new_n6402_));
  OAI21_X1   g05400(.A1(new_n6399_), .A2(\A[236] ), .B(\A[237] ), .ZN(new_n6403_));
  NOR2_X1    g05401(.A1(new_n6403_), .A2(new_n6402_), .ZN(new_n6404_));
  NOR2_X1    g05402(.A1(new_n6401_), .A2(new_n6404_), .ZN(new_n6405_));
  INV_X1     g05403(.I(\A[240] ), .ZN(new_n6406_));
  INV_X1     g05404(.I(\A[238] ), .ZN(new_n6407_));
  NAND2_X1   g05405(.A1(new_n6407_), .A2(\A[239] ), .ZN(new_n6408_));
  XOR2_X1    g05406(.A1(\A[238] ), .A2(\A[239] ), .Z(new_n6409_));
  INV_X1     g05407(.I(\A[239] ), .ZN(new_n6410_));
  AOI21_X1   g05408(.A1(\A[238] ), .A2(new_n6410_), .B(new_n6406_), .ZN(new_n6411_));
  AOI22_X1   g05409(.A1(new_n6409_), .A2(new_n6406_), .B1(new_n6408_), .B2(new_n6411_), .ZN(new_n6412_));
  XOR2_X1    g05410(.A1(new_n6405_), .A2(new_n6412_), .Z(new_n6413_));
  NOR2_X1    g05411(.A1(new_n6407_), .A2(\A[239] ), .ZN(new_n6414_));
  NOR2_X1    g05412(.A1(new_n6410_), .A2(\A[238] ), .ZN(new_n6415_));
  NOR2_X1    g05413(.A1(new_n6414_), .A2(new_n6415_), .ZN(new_n6416_));
  NOR2_X1    g05414(.A1(new_n6407_), .A2(new_n6410_), .ZN(new_n6417_));
  INV_X1     g05415(.I(new_n6417_), .ZN(new_n6418_));
  OAI21_X1   g05416(.A1(new_n6416_), .A2(new_n6406_), .B(new_n6418_), .ZN(new_n6419_));
  INV_X1     g05417(.I(\A[237] ), .ZN(new_n6420_));
  NOR2_X1    g05418(.A1(new_n6399_), .A2(\A[236] ), .ZN(new_n6421_));
  NOR2_X1    g05419(.A1(new_n6421_), .A2(new_n6402_), .ZN(new_n6422_));
  NOR2_X1    g05420(.A1(new_n6399_), .A2(new_n6397_), .ZN(new_n6423_));
  INV_X1     g05421(.I(new_n6423_), .ZN(new_n6424_));
  OAI21_X1   g05422(.A1(new_n6422_), .A2(new_n6420_), .B(new_n6424_), .ZN(new_n6425_));
  XOR2_X1    g05423(.A1(\A[235] ), .A2(\A[236] ), .Z(new_n6426_));
  NAND2_X1   g05424(.A1(new_n6426_), .A2(new_n6420_), .ZN(new_n6427_));
  NAND3_X1   g05425(.A1(new_n6398_), .A2(new_n6400_), .A3(\A[237] ), .ZN(new_n6428_));
  OAI21_X1   g05426(.A1(new_n6414_), .A2(new_n6415_), .B(new_n6406_), .ZN(new_n6429_));
  NAND2_X1   g05427(.A1(new_n6411_), .A2(new_n6408_), .ZN(new_n6430_));
  AOI22_X1   g05428(.A1(new_n6427_), .A2(new_n6428_), .B1(new_n6429_), .B2(new_n6430_), .ZN(new_n6431_));
  NAND3_X1   g05429(.A1(new_n6431_), .A2(new_n6419_), .A3(new_n6425_), .ZN(new_n6432_));
  NAND2_X1   g05430(.A1(new_n6413_), .A2(new_n6432_), .ZN(new_n6433_));
  NAND2_X1   g05431(.A1(new_n6433_), .A2(new_n6396_), .ZN(new_n6434_));
  NAND2_X1   g05432(.A1(new_n6386_), .A2(new_n6383_), .ZN(new_n6435_));
  NAND2_X1   g05433(.A1(new_n6367_), .A2(new_n6377_), .ZN(new_n6436_));
  NAND2_X1   g05434(.A1(new_n6436_), .A2(new_n6435_), .ZN(new_n6437_));
  NOR2_X1    g05435(.A1(new_n6374_), .A2(new_n6375_), .ZN(new_n6438_));
  INV_X1     g05436(.I(new_n6390_), .ZN(new_n6439_));
  OAI21_X1   g05437(.A1(new_n6438_), .A2(new_n6373_), .B(new_n6439_), .ZN(new_n6440_));
  NOR2_X1    g05438(.A1(new_n6364_), .A2(\A[242] ), .ZN(new_n6441_));
  NOR2_X1    g05439(.A1(new_n6441_), .A2(new_n6380_), .ZN(new_n6442_));
  INV_X1     g05440(.I(new_n6392_), .ZN(new_n6443_));
  OAI21_X1   g05441(.A1(new_n6442_), .A2(new_n6359_), .B(new_n6443_), .ZN(new_n6444_));
  AOI22_X1   g05442(.A1(new_n6361_), .A2(new_n6366_), .B1(new_n6384_), .B2(new_n6385_), .ZN(new_n6445_));
  NAND3_X1   g05443(.A1(new_n6445_), .A2(new_n6440_), .A3(new_n6444_), .ZN(new_n6446_));
  NAND2_X1   g05444(.A1(new_n6437_), .A2(new_n6446_), .ZN(new_n6447_));
  NAND2_X1   g05445(.A1(new_n6427_), .A2(new_n6428_), .ZN(new_n6448_));
  NOR2_X1    g05446(.A1(new_n6448_), .A2(new_n6412_), .ZN(new_n6449_));
  NAND2_X1   g05447(.A1(new_n6430_), .A2(new_n6429_), .ZN(new_n6450_));
  NOR2_X1    g05448(.A1(new_n6450_), .A2(new_n6405_), .ZN(new_n6451_));
  NOR2_X1    g05449(.A1(new_n6449_), .A2(new_n6451_), .ZN(new_n6452_));
  AOI21_X1   g05450(.A1(new_n6409_), .A2(\A[240] ), .B(new_n6417_), .ZN(new_n6453_));
  AOI21_X1   g05451(.A1(new_n6426_), .A2(\A[237] ), .B(new_n6423_), .ZN(new_n6454_));
  INV_X1     g05452(.I(new_n6414_), .ZN(new_n6455_));
  AOI21_X1   g05453(.A1(new_n6455_), .A2(new_n6408_), .B(\A[240] ), .ZN(new_n6456_));
  NOR3_X1    g05454(.A1(new_n6414_), .A2(new_n6415_), .A3(new_n6406_), .ZN(new_n6457_));
  OAI22_X1   g05455(.A1(new_n6456_), .A2(new_n6457_), .B1(new_n6401_), .B2(new_n6404_), .ZN(new_n6458_));
  NOR3_X1    g05456(.A1(new_n6458_), .A2(new_n6453_), .A3(new_n6454_), .ZN(new_n6459_));
  NOR2_X1    g05457(.A1(new_n6452_), .A2(new_n6459_), .ZN(new_n6460_));
  NAND2_X1   g05458(.A1(new_n6460_), .A2(new_n6447_), .ZN(new_n6461_));
  NAND2_X1   g05459(.A1(new_n6434_), .A2(new_n6461_), .ZN(new_n6462_));
  INV_X1     g05460(.I(\A[229] ), .ZN(new_n6463_));
  NAND2_X1   g05461(.A1(new_n6463_), .A2(\A[230] ), .ZN(new_n6464_));
  INV_X1     g05462(.I(\A[230] ), .ZN(new_n6465_));
  NAND2_X1   g05463(.A1(new_n6465_), .A2(\A[229] ), .ZN(new_n6466_));
  NAND3_X1   g05464(.A1(new_n6464_), .A2(new_n6466_), .A3(\A[231] ), .ZN(new_n6467_));
  INV_X1     g05465(.I(\A[231] ), .ZN(new_n6468_));
  NOR2_X1    g05466(.A1(new_n6465_), .A2(\A[229] ), .ZN(new_n6469_));
  NOR2_X1    g05467(.A1(new_n6463_), .A2(\A[230] ), .ZN(new_n6470_));
  OAI21_X1   g05468(.A1(new_n6469_), .A2(new_n6470_), .B(new_n6468_), .ZN(new_n6471_));
  NAND2_X1   g05469(.A1(new_n6471_), .A2(new_n6467_), .ZN(new_n6472_));
  INV_X1     g05470(.I(\A[234] ), .ZN(new_n6473_));
  INV_X1     g05471(.I(\A[233] ), .ZN(new_n6474_));
  NOR2_X1    g05472(.A1(new_n6474_), .A2(\A[232] ), .ZN(new_n6475_));
  INV_X1     g05473(.I(\A[232] ), .ZN(new_n6476_));
  NOR2_X1    g05474(.A1(new_n6476_), .A2(\A[233] ), .ZN(new_n6477_));
  NOR3_X1    g05475(.A1(new_n6475_), .A2(new_n6477_), .A3(new_n6473_), .ZN(new_n6478_));
  NAND2_X1   g05476(.A1(new_n6476_), .A2(\A[233] ), .ZN(new_n6479_));
  NAND2_X1   g05477(.A1(new_n6474_), .A2(\A[232] ), .ZN(new_n6480_));
  AOI21_X1   g05478(.A1(new_n6479_), .A2(new_n6480_), .B(\A[234] ), .ZN(new_n6481_));
  NOR2_X1    g05479(.A1(new_n6481_), .A2(new_n6478_), .ZN(new_n6482_));
  NOR2_X1    g05480(.A1(new_n6482_), .A2(new_n6472_), .ZN(new_n6483_));
  INV_X1     g05481(.I(new_n6467_), .ZN(new_n6484_));
  AOI21_X1   g05482(.A1(new_n6464_), .A2(new_n6466_), .B(\A[231] ), .ZN(new_n6485_));
  NOR2_X1    g05483(.A1(new_n6484_), .A2(new_n6485_), .ZN(new_n6486_));
  NAND3_X1   g05484(.A1(new_n6479_), .A2(new_n6480_), .A3(\A[234] ), .ZN(new_n6487_));
  OAI21_X1   g05485(.A1(new_n6475_), .A2(new_n6477_), .B(new_n6473_), .ZN(new_n6488_));
  NAND2_X1   g05486(.A1(new_n6488_), .A2(new_n6487_), .ZN(new_n6489_));
  NOR2_X1    g05487(.A1(new_n6486_), .A2(new_n6489_), .ZN(new_n6490_));
  NOR2_X1    g05488(.A1(new_n6490_), .A2(new_n6483_), .ZN(new_n6491_));
  NAND2_X1   g05489(.A1(new_n6479_), .A2(new_n6480_), .ZN(new_n6492_));
  NOR2_X1    g05490(.A1(new_n6476_), .A2(new_n6474_), .ZN(new_n6493_));
  AOI21_X1   g05491(.A1(new_n6492_), .A2(\A[234] ), .B(new_n6493_), .ZN(new_n6494_));
  NAND2_X1   g05492(.A1(new_n6464_), .A2(new_n6466_), .ZN(new_n6495_));
  NOR2_X1    g05493(.A1(new_n6463_), .A2(new_n6465_), .ZN(new_n6496_));
  AOI21_X1   g05494(.A1(new_n6495_), .A2(\A[231] ), .B(new_n6496_), .ZN(new_n6497_));
  NAND2_X1   g05495(.A1(new_n6472_), .A2(new_n6489_), .ZN(new_n6498_));
  NOR3_X1    g05496(.A1(new_n6498_), .A2(new_n6494_), .A3(new_n6497_), .ZN(new_n6499_));
  NOR2_X1    g05497(.A1(new_n6491_), .A2(new_n6499_), .ZN(new_n6500_));
  INV_X1     g05498(.I(\A[225] ), .ZN(new_n6501_));
  INV_X1     g05499(.I(\A[223] ), .ZN(new_n6502_));
  NAND2_X1   g05500(.A1(new_n6502_), .A2(\A[224] ), .ZN(new_n6503_));
  INV_X1     g05501(.I(\A[224] ), .ZN(new_n6504_));
  AOI21_X1   g05502(.A1(\A[223] ), .A2(new_n6504_), .B(new_n6501_), .ZN(new_n6505_));
  NAND2_X1   g05503(.A1(new_n6504_), .A2(\A[223] ), .ZN(new_n6506_));
  NAND2_X1   g05504(.A1(new_n6503_), .A2(new_n6506_), .ZN(new_n6507_));
  AOI22_X1   g05505(.A1(new_n6507_), .A2(new_n6501_), .B1(new_n6503_), .B2(new_n6505_), .ZN(new_n6508_));
  INV_X1     g05506(.I(\A[226] ), .ZN(new_n6509_));
  NAND2_X1   g05507(.A1(new_n6509_), .A2(\A[227] ), .ZN(new_n6510_));
  INV_X1     g05508(.I(\A[227] ), .ZN(new_n6511_));
  NAND2_X1   g05509(.A1(new_n6511_), .A2(\A[226] ), .ZN(new_n6512_));
  NAND3_X1   g05510(.A1(new_n6510_), .A2(new_n6512_), .A3(\A[228] ), .ZN(new_n6513_));
  INV_X1     g05511(.I(\A[228] ), .ZN(new_n6514_));
  NOR2_X1    g05512(.A1(new_n6511_), .A2(\A[226] ), .ZN(new_n6515_));
  NOR2_X1    g05513(.A1(new_n6509_), .A2(\A[227] ), .ZN(new_n6516_));
  OAI21_X1   g05514(.A1(new_n6515_), .A2(new_n6516_), .B(new_n6514_), .ZN(new_n6517_));
  NAND2_X1   g05515(.A1(new_n6517_), .A2(new_n6513_), .ZN(new_n6518_));
  NAND2_X1   g05516(.A1(new_n6508_), .A2(new_n6518_), .ZN(new_n6519_));
  NAND2_X1   g05517(.A1(new_n6505_), .A2(new_n6503_), .ZN(new_n6520_));
  NOR2_X1    g05518(.A1(new_n6504_), .A2(\A[223] ), .ZN(new_n6521_));
  NOR2_X1    g05519(.A1(new_n6502_), .A2(\A[224] ), .ZN(new_n6522_));
  OAI21_X1   g05520(.A1(new_n6521_), .A2(new_n6522_), .B(new_n6501_), .ZN(new_n6523_));
  NAND2_X1   g05521(.A1(new_n6520_), .A2(new_n6523_), .ZN(new_n6524_));
  NOR3_X1    g05522(.A1(new_n6515_), .A2(new_n6516_), .A3(new_n6514_), .ZN(new_n6525_));
  NAND2_X1   g05523(.A1(new_n6510_), .A2(new_n6512_), .ZN(new_n6526_));
  AOI21_X1   g05524(.A1(new_n6514_), .A2(new_n6526_), .B(new_n6525_), .ZN(new_n6527_));
  NAND2_X1   g05525(.A1(new_n6527_), .A2(new_n6524_), .ZN(new_n6528_));
  NAND2_X1   g05526(.A1(new_n6528_), .A2(new_n6519_), .ZN(new_n6529_));
  NOR2_X1    g05527(.A1(new_n6515_), .A2(new_n6516_), .ZN(new_n6530_));
  NOR2_X1    g05528(.A1(new_n6509_), .A2(new_n6511_), .ZN(new_n6531_));
  INV_X1     g05529(.I(new_n6531_), .ZN(new_n6532_));
  OAI21_X1   g05530(.A1(new_n6530_), .A2(new_n6514_), .B(new_n6532_), .ZN(new_n6533_));
  NOR2_X1    g05531(.A1(new_n6521_), .A2(new_n6522_), .ZN(new_n6534_));
  NOR2_X1    g05532(.A1(new_n6502_), .A2(new_n6504_), .ZN(new_n6535_));
  INV_X1     g05533(.I(new_n6535_), .ZN(new_n6536_));
  OAI21_X1   g05534(.A1(new_n6534_), .A2(new_n6501_), .B(new_n6536_), .ZN(new_n6537_));
  AOI22_X1   g05535(.A1(new_n6520_), .A2(new_n6523_), .B1(new_n6517_), .B2(new_n6513_), .ZN(new_n6538_));
  NAND3_X1   g05536(.A1(new_n6538_), .A2(new_n6533_), .A3(new_n6537_), .ZN(new_n6539_));
  NAND2_X1   g05537(.A1(new_n6529_), .A2(new_n6539_), .ZN(new_n6540_));
  NOR2_X1    g05538(.A1(new_n6500_), .A2(new_n6540_), .ZN(new_n6541_));
  XOR2_X1    g05539(.A1(new_n6472_), .A2(new_n6489_), .Z(new_n6542_));
  NOR2_X1    g05540(.A1(new_n6475_), .A2(new_n6477_), .ZN(new_n6543_));
  INV_X1     g05541(.I(new_n6493_), .ZN(new_n6544_));
  OAI21_X1   g05542(.A1(new_n6543_), .A2(new_n6473_), .B(new_n6544_), .ZN(new_n6545_));
  NOR2_X1    g05543(.A1(new_n6469_), .A2(new_n6470_), .ZN(new_n6546_));
  INV_X1     g05544(.I(new_n6496_), .ZN(new_n6547_));
  OAI21_X1   g05545(.A1(new_n6546_), .A2(new_n6468_), .B(new_n6547_), .ZN(new_n6548_));
  AOI22_X1   g05546(.A1(new_n6467_), .A2(new_n6471_), .B1(new_n6488_), .B2(new_n6487_), .ZN(new_n6549_));
  NAND3_X1   g05547(.A1(new_n6549_), .A2(new_n6545_), .A3(new_n6548_), .ZN(new_n6550_));
  NAND2_X1   g05548(.A1(new_n6542_), .A2(new_n6550_), .ZN(new_n6551_));
  NOR2_X1    g05549(.A1(new_n6527_), .A2(new_n6524_), .ZN(new_n6552_));
  NOR2_X1    g05550(.A1(new_n6508_), .A2(new_n6518_), .ZN(new_n6553_));
  NOR2_X1    g05551(.A1(new_n6552_), .A2(new_n6553_), .ZN(new_n6554_));
  AOI21_X1   g05552(.A1(new_n6526_), .A2(\A[228] ), .B(new_n6531_), .ZN(new_n6555_));
  AOI21_X1   g05553(.A1(new_n6507_), .A2(\A[225] ), .B(new_n6535_), .ZN(new_n6556_));
  NOR4_X1    g05554(.A1(new_n6527_), .A2(new_n6508_), .A3(new_n6555_), .A4(new_n6556_), .ZN(new_n6557_));
  NOR2_X1    g05555(.A1(new_n6554_), .A2(new_n6557_), .ZN(new_n6558_));
  NOR2_X1    g05556(.A1(new_n6551_), .A2(new_n6558_), .ZN(new_n6559_));
  NOR2_X1    g05557(.A1(new_n6559_), .A2(new_n6541_), .ZN(new_n6560_));
  NAND2_X1   g05558(.A1(new_n6560_), .A2(new_n6462_), .ZN(new_n6561_));
  NOR2_X1    g05559(.A1(new_n6460_), .A2(new_n6447_), .ZN(new_n6562_));
  NOR2_X1    g05560(.A1(new_n6433_), .A2(new_n6396_), .ZN(new_n6563_));
  NOR2_X1    g05561(.A1(new_n6563_), .A2(new_n6562_), .ZN(new_n6564_));
  NAND2_X1   g05562(.A1(new_n6551_), .A2(new_n6558_), .ZN(new_n6565_));
  NAND2_X1   g05563(.A1(new_n6500_), .A2(new_n6540_), .ZN(new_n6566_));
  NAND2_X1   g05564(.A1(new_n6565_), .A2(new_n6566_), .ZN(new_n6567_));
  NAND2_X1   g05565(.A1(new_n6567_), .A2(new_n6564_), .ZN(new_n6568_));
  NAND2_X1   g05566(.A1(new_n6568_), .A2(new_n6561_), .ZN(new_n6569_));
  XNOR2_X1   g05567(.A1(new_n6569_), .A2(new_n6358_), .ZN(new_n6570_));
  XNOR2_X1   g05568(.A1(new_n6170_), .A2(new_n6570_), .ZN(new_n6571_));
  INV_X1     g05569(.I(\A[171] ), .ZN(new_n6572_));
  INV_X1     g05570(.I(\A[170] ), .ZN(new_n6573_));
  NOR2_X1    g05571(.A1(new_n6573_), .A2(\A[169] ), .ZN(new_n6574_));
  INV_X1     g05572(.I(\A[169] ), .ZN(new_n6575_));
  NOR2_X1    g05573(.A1(new_n6575_), .A2(\A[170] ), .ZN(new_n6576_));
  NOR3_X1    g05574(.A1(new_n6574_), .A2(new_n6576_), .A3(new_n6572_), .ZN(new_n6577_));
  NAND2_X1   g05575(.A1(new_n6575_), .A2(\A[170] ), .ZN(new_n6578_));
  NAND2_X1   g05576(.A1(new_n6573_), .A2(\A[169] ), .ZN(new_n6579_));
  AOI21_X1   g05577(.A1(new_n6578_), .A2(new_n6579_), .B(\A[171] ), .ZN(new_n6580_));
  NOR2_X1    g05578(.A1(new_n6580_), .A2(new_n6577_), .ZN(new_n6581_));
  INV_X1     g05579(.I(\A[172] ), .ZN(new_n6582_));
  NAND2_X1   g05580(.A1(new_n6582_), .A2(\A[173] ), .ZN(new_n6583_));
  INV_X1     g05581(.I(\A[173] ), .ZN(new_n6584_));
  INV_X1     g05582(.I(\A[174] ), .ZN(new_n6585_));
  AOI21_X1   g05583(.A1(\A[172] ), .A2(new_n6584_), .B(new_n6585_), .ZN(new_n6586_));
  NAND2_X1   g05584(.A1(new_n6586_), .A2(new_n6583_), .ZN(new_n6587_));
  NOR2_X1    g05585(.A1(new_n6584_), .A2(\A[172] ), .ZN(new_n6588_));
  NOR2_X1    g05586(.A1(new_n6582_), .A2(\A[173] ), .ZN(new_n6589_));
  OAI21_X1   g05587(.A1(new_n6588_), .A2(new_n6589_), .B(new_n6585_), .ZN(new_n6590_));
  NAND2_X1   g05588(.A1(new_n6587_), .A2(new_n6590_), .ZN(new_n6591_));
  NAND2_X1   g05589(.A1(new_n6581_), .A2(new_n6591_), .ZN(new_n6592_));
  AOI21_X1   g05590(.A1(\A[169] ), .A2(new_n6573_), .B(new_n6572_), .ZN(new_n6593_));
  NAND2_X1   g05591(.A1(new_n6593_), .A2(new_n6578_), .ZN(new_n6594_));
  OAI21_X1   g05592(.A1(new_n6574_), .A2(new_n6576_), .B(new_n6572_), .ZN(new_n6595_));
  NAND2_X1   g05593(.A1(new_n6594_), .A2(new_n6595_), .ZN(new_n6596_));
  XOR2_X1    g05594(.A1(\A[172] ), .A2(\A[173] ), .Z(new_n6597_));
  AOI22_X1   g05595(.A1(new_n6597_), .A2(new_n6585_), .B1(new_n6583_), .B2(new_n6586_), .ZN(new_n6598_));
  NAND2_X1   g05596(.A1(new_n6596_), .A2(new_n6598_), .ZN(new_n6599_));
  NAND2_X1   g05597(.A1(new_n6592_), .A2(new_n6599_), .ZN(new_n6600_));
  NOR2_X1    g05598(.A1(new_n6588_), .A2(new_n6589_), .ZN(new_n6601_));
  NOR2_X1    g05599(.A1(new_n6582_), .A2(new_n6584_), .ZN(new_n6602_));
  INV_X1     g05600(.I(new_n6602_), .ZN(new_n6603_));
  OAI21_X1   g05601(.A1(new_n6601_), .A2(new_n6585_), .B(new_n6603_), .ZN(new_n6604_));
  NOR2_X1    g05602(.A1(new_n6574_), .A2(new_n6576_), .ZN(new_n6605_));
  NOR2_X1    g05603(.A1(new_n6575_), .A2(new_n6573_), .ZN(new_n6606_));
  INV_X1     g05604(.I(new_n6606_), .ZN(new_n6607_));
  OAI21_X1   g05605(.A1(new_n6605_), .A2(new_n6572_), .B(new_n6607_), .ZN(new_n6608_));
  AOI22_X1   g05606(.A1(new_n6594_), .A2(new_n6595_), .B1(new_n6587_), .B2(new_n6590_), .ZN(new_n6609_));
  NAND3_X1   g05607(.A1(new_n6609_), .A2(new_n6604_), .A3(new_n6608_), .ZN(new_n6610_));
  NAND2_X1   g05608(.A1(new_n6600_), .A2(new_n6610_), .ZN(new_n6611_));
  INV_X1     g05609(.I(\A[164] ), .ZN(new_n6612_));
  NOR2_X1    g05610(.A1(new_n6612_), .A2(\A[163] ), .ZN(new_n6613_));
  INV_X1     g05611(.I(new_n6613_), .ZN(new_n6614_));
  INV_X1     g05612(.I(\A[165] ), .ZN(new_n6615_));
  AOI21_X1   g05613(.A1(\A[163] ), .A2(new_n6612_), .B(new_n6615_), .ZN(new_n6616_));
  NAND2_X1   g05614(.A1(new_n6614_), .A2(new_n6616_), .ZN(new_n6617_));
  INV_X1     g05615(.I(\A[163] ), .ZN(new_n6618_));
  NOR2_X1    g05616(.A1(new_n6618_), .A2(\A[164] ), .ZN(new_n6619_));
  OAI21_X1   g05617(.A1(new_n6613_), .A2(new_n6619_), .B(new_n6615_), .ZN(new_n6620_));
  NAND2_X1   g05618(.A1(new_n6617_), .A2(new_n6620_), .ZN(new_n6621_));
  INV_X1     g05619(.I(\A[168] ), .ZN(new_n6622_));
  INV_X1     g05620(.I(\A[167] ), .ZN(new_n6623_));
  NOR2_X1    g05621(.A1(new_n6623_), .A2(\A[166] ), .ZN(new_n6624_));
  INV_X1     g05622(.I(\A[166] ), .ZN(new_n6625_));
  NOR2_X1    g05623(.A1(new_n6625_), .A2(\A[167] ), .ZN(new_n6626_));
  NOR3_X1    g05624(.A1(new_n6624_), .A2(new_n6626_), .A3(new_n6622_), .ZN(new_n6627_));
  NAND2_X1   g05625(.A1(new_n6625_), .A2(\A[167] ), .ZN(new_n6628_));
  NAND2_X1   g05626(.A1(new_n6623_), .A2(\A[166] ), .ZN(new_n6629_));
  AOI21_X1   g05627(.A1(new_n6628_), .A2(new_n6629_), .B(\A[168] ), .ZN(new_n6630_));
  NOR2_X1    g05628(.A1(new_n6630_), .A2(new_n6627_), .ZN(new_n6631_));
  NOR2_X1    g05629(.A1(new_n6621_), .A2(new_n6631_), .ZN(new_n6632_));
  XOR2_X1    g05630(.A1(\A[163] ), .A2(\A[164] ), .Z(new_n6633_));
  AOI22_X1   g05631(.A1(new_n6633_), .A2(new_n6615_), .B1(new_n6614_), .B2(new_n6616_), .ZN(new_n6634_));
  AOI21_X1   g05632(.A1(\A[166] ), .A2(new_n6623_), .B(new_n6622_), .ZN(new_n6635_));
  NAND2_X1   g05633(.A1(new_n6635_), .A2(new_n6628_), .ZN(new_n6636_));
  OAI21_X1   g05634(.A1(new_n6624_), .A2(new_n6626_), .B(new_n6622_), .ZN(new_n6637_));
  NAND2_X1   g05635(.A1(new_n6636_), .A2(new_n6637_), .ZN(new_n6638_));
  NOR2_X1    g05636(.A1(new_n6638_), .A2(new_n6634_), .ZN(new_n6639_));
  NOR2_X1    g05637(.A1(new_n6632_), .A2(new_n6639_), .ZN(new_n6640_));
  NAND2_X1   g05638(.A1(new_n6628_), .A2(new_n6629_), .ZN(new_n6641_));
  NOR2_X1    g05639(.A1(new_n6625_), .A2(new_n6623_), .ZN(new_n6642_));
  AOI21_X1   g05640(.A1(new_n6641_), .A2(\A[168] ), .B(new_n6642_), .ZN(new_n6643_));
  NOR2_X1    g05641(.A1(new_n6618_), .A2(new_n6612_), .ZN(new_n6644_));
  AOI21_X1   g05642(.A1(new_n6633_), .A2(\A[165] ), .B(new_n6644_), .ZN(new_n6645_));
  NOR3_X1    g05643(.A1(new_n6613_), .A2(new_n6619_), .A3(new_n6615_), .ZN(new_n6646_));
  NAND2_X1   g05644(.A1(new_n6612_), .A2(\A[163] ), .ZN(new_n6647_));
  AOI21_X1   g05645(.A1(new_n6614_), .A2(new_n6647_), .B(\A[165] ), .ZN(new_n6648_));
  OAI22_X1   g05646(.A1(new_n6648_), .A2(new_n6646_), .B1(new_n6627_), .B2(new_n6630_), .ZN(new_n6649_));
  NOR3_X1    g05647(.A1(new_n6649_), .A2(new_n6643_), .A3(new_n6645_), .ZN(new_n6650_));
  NOR2_X1    g05648(.A1(new_n6640_), .A2(new_n6650_), .ZN(new_n6651_));
  NAND2_X1   g05649(.A1(new_n6651_), .A2(new_n6611_), .ZN(new_n6652_));
  XOR2_X1    g05650(.A1(new_n6596_), .A2(new_n6598_), .Z(new_n6653_));
  AOI21_X1   g05651(.A1(new_n6597_), .A2(\A[174] ), .B(new_n6602_), .ZN(new_n6654_));
  XOR2_X1    g05652(.A1(\A[169] ), .A2(\A[170] ), .Z(new_n6655_));
  AOI21_X1   g05653(.A1(new_n6655_), .A2(\A[171] ), .B(new_n6606_), .ZN(new_n6656_));
  NOR3_X1    g05654(.A1(new_n6588_), .A2(new_n6589_), .A3(new_n6585_), .ZN(new_n6657_));
  NAND2_X1   g05655(.A1(new_n6584_), .A2(\A[172] ), .ZN(new_n6658_));
  AOI21_X1   g05656(.A1(new_n6583_), .A2(new_n6658_), .B(\A[174] ), .ZN(new_n6659_));
  OAI22_X1   g05657(.A1(new_n6577_), .A2(new_n6580_), .B1(new_n6659_), .B2(new_n6657_), .ZN(new_n6660_));
  NOR3_X1    g05658(.A1(new_n6660_), .A2(new_n6654_), .A3(new_n6656_), .ZN(new_n6661_));
  NOR2_X1    g05659(.A1(new_n6653_), .A2(new_n6661_), .ZN(new_n6662_));
  NAND2_X1   g05660(.A1(new_n6638_), .A2(new_n6634_), .ZN(new_n6663_));
  NAND2_X1   g05661(.A1(new_n6621_), .A2(new_n6631_), .ZN(new_n6664_));
  NAND2_X1   g05662(.A1(new_n6664_), .A2(new_n6663_), .ZN(new_n6665_));
  NOR2_X1    g05663(.A1(new_n6624_), .A2(new_n6626_), .ZN(new_n6666_));
  INV_X1     g05664(.I(new_n6642_), .ZN(new_n6667_));
  OAI21_X1   g05665(.A1(new_n6666_), .A2(new_n6622_), .B(new_n6667_), .ZN(new_n6668_));
  NOR2_X1    g05666(.A1(new_n6613_), .A2(new_n6619_), .ZN(new_n6669_));
  INV_X1     g05667(.I(new_n6644_), .ZN(new_n6670_));
  OAI21_X1   g05668(.A1(new_n6669_), .A2(new_n6615_), .B(new_n6670_), .ZN(new_n6671_));
  AOI22_X1   g05669(.A1(new_n6617_), .A2(new_n6620_), .B1(new_n6636_), .B2(new_n6637_), .ZN(new_n6672_));
  NAND3_X1   g05670(.A1(new_n6672_), .A2(new_n6668_), .A3(new_n6671_), .ZN(new_n6673_));
  NAND2_X1   g05671(.A1(new_n6665_), .A2(new_n6673_), .ZN(new_n6674_));
  NAND2_X1   g05672(.A1(new_n6662_), .A2(new_n6674_), .ZN(new_n6675_));
  INV_X1     g05673(.I(\A[159] ), .ZN(new_n6676_));
  INV_X1     g05674(.I(\A[158] ), .ZN(new_n6677_));
  NOR2_X1    g05675(.A1(new_n6677_), .A2(\A[157] ), .ZN(new_n6678_));
  INV_X1     g05676(.I(\A[157] ), .ZN(new_n6679_));
  NOR2_X1    g05677(.A1(new_n6679_), .A2(\A[158] ), .ZN(new_n6680_));
  NOR3_X1    g05678(.A1(new_n6678_), .A2(new_n6680_), .A3(new_n6676_), .ZN(new_n6681_));
  NAND2_X1   g05679(.A1(new_n6679_), .A2(\A[158] ), .ZN(new_n6682_));
  NAND2_X1   g05680(.A1(new_n6677_), .A2(\A[157] ), .ZN(new_n6683_));
  AOI21_X1   g05681(.A1(new_n6682_), .A2(new_n6683_), .B(\A[159] ), .ZN(new_n6684_));
  NOR2_X1    g05682(.A1(new_n6684_), .A2(new_n6681_), .ZN(new_n6685_));
  INV_X1     g05683(.I(\A[160] ), .ZN(new_n6686_));
  NAND2_X1   g05684(.A1(new_n6686_), .A2(\A[161] ), .ZN(new_n6687_));
  INV_X1     g05685(.I(\A[161] ), .ZN(new_n6688_));
  NAND2_X1   g05686(.A1(new_n6688_), .A2(\A[160] ), .ZN(new_n6689_));
  NAND3_X1   g05687(.A1(new_n6687_), .A2(new_n6689_), .A3(\A[162] ), .ZN(new_n6690_));
  INV_X1     g05688(.I(\A[162] ), .ZN(new_n6691_));
  NOR2_X1    g05689(.A1(new_n6688_), .A2(\A[160] ), .ZN(new_n6692_));
  NOR2_X1    g05690(.A1(new_n6686_), .A2(\A[161] ), .ZN(new_n6693_));
  OAI21_X1   g05691(.A1(new_n6692_), .A2(new_n6693_), .B(new_n6691_), .ZN(new_n6694_));
  NAND2_X1   g05692(.A1(new_n6694_), .A2(new_n6690_), .ZN(new_n6695_));
  NAND2_X1   g05693(.A1(new_n6685_), .A2(new_n6695_), .ZN(new_n6696_));
  AOI21_X1   g05694(.A1(\A[157] ), .A2(new_n6677_), .B(new_n6676_), .ZN(new_n6697_));
  NAND2_X1   g05695(.A1(new_n6697_), .A2(new_n6682_), .ZN(new_n6698_));
  XOR2_X1    g05696(.A1(\A[157] ), .A2(\A[158] ), .Z(new_n6699_));
  NAND2_X1   g05697(.A1(new_n6699_), .A2(new_n6676_), .ZN(new_n6700_));
  NAND2_X1   g05698(.A1(new_n6700_), .A2(new_n6698_), .ZN(new_n6701_));
  NOR3_X1    g05699(.A1(new_n6692_), .A2(new_n6693_), .A3(new_n6691_), .ZN(new_n6702_));
  AOI21_X1   g05700(.A1(new_n6687_), .A2(new_n6689_), .B(\A[162] ), .ZN(new_n6703_));
  NOR2_X1    g05701(.A1(new_n6703_), .A2(new_n6702_), .ZN(new_n6704_));
  NAND2_X1   g05702(.A1(new_n6701_), .A2(new_n6704_), .ZN(new_n6705_));
  NAND2_X1   g05703(.A1(new_n6705_), .A2(new_n6696_), .ZN(new_n6706_));
  NOR2_X1    g05704(.A1(new_n6692_), .A2(new_n6693_), .ZN(new_n6707_));
  NOR2_X1    g05705(.A1(new_n6686_), .A2(new_n6688_), .ZN(new_n6708_));
  INV_X1     g05706(.I(new_n6708_), .ZN(new_n6709_));
  OAI21_X1   g05707(.A1(new_n6707_), .A2(new_n6691_), .B(new_n6709_), .ZN(new_n6710_));
  NOR2_X1    g05708(.A1(new_n6678_), .A2(new_n6680_), .ZN(new_n6711_));
  NOR2_X1    g05709(.A1(new_n6679_), .A2(new_n6677_), .ZN(new_n6712_));
  INV_X1     g05710(.I(new_n6712_), .ZN(new_n6713_));
  OAI21_X1   g05711(.A1(new_n6711_), .A2(new_n6676_), .B(new_n6713_), .ZN(new_n6714_));
  AOI22_X1   g05712(.A1(new_n6700_), .A2(new_n6698_), .B1(new_n6690_), .B2(new_n6694_), .ZN(new_n6715_));
  NAND3_X1   g05713(.A1(new_n6715_), .A2(new_n6710_), .A3(new_n6714_), .ZN(new_n6716_));
  NAND2_X1   g05714(.A1(new_n6706_), .A2(new_n6716_), .ZN(new_n6717_));
  INV_X1     g05715(.I(\A[152] ), .ZN(new_n6718_));
  NOR2_X1    g05716(.A1(new_n6718_), .A2(\A[151] ), .ZN(new_n6719_));
  NAND2_X1   g05717(.A1(new_n6718_), .A2(\A[151] ), .ZN(new_n6720_));
  NAND2_X1   g05718(.A1(new_n6720_), .A2(\A[153] ), .ZN(new_n6721_));
  INV_X1     g05719(.I(\A[151] ), .ZN(new_n6722_));
  NOR2_X1    g05720(.A1(new_n6722_), .A2(\A[152] ), .ZN(new_n6723_));
  NOR2_X1    g05721(.A1(new_n6719_), .A2(new_n6723_), .ZN(new_n6724_));
  OAI22_X1   g05722(.A1(new_n6724_), .A2(\A[153] ), .B1(new_n6721_), .B2(new_n6719_), .ZN(new_n6725_));
  INV_X1     g05723(.I(\A[156] ), .ZN(new_n6726_));
  INV_X1     g05724(.I(\A[155] ), .ZN(new_n6727_));
  NOR2_X1    g05725(.A1(new_n6727_), .A2(\A[154] ), .ZN(new_n6728_));
  INV_X1     g05726(.I(\A[154] ), .ZN(new_n6729_));
  NOR2_X1    g05727(.A1(new_n6729_), .A2(\A[155] ), .ZN(new_n6730_));
  NOR3_X1    g05728(.A1(new_n6728_), .A2(new_n6730_), .A3(new_n6726_), .ZN(new_n6731_));
  NAND2_X1   g05729(.A1(new_n6729_), .A2(\A[155] ), .ZN(new_n6732_));
  NAND2_X1   g05730(.A1(new_n6727_), .A2(\A[154] ), .ZN(new_n6733_));
  AOI21_X1   g05731(.A1(new_n6732_), .A2(new_n6733_), .B(\A[156] ), .ZN(new_n6734_));
  NOR2_X1    g05732(.A1(new_n6734_), .A2(new_n6731_), .ZN(new_n6735_));
  NOR2_X1    g05733(.A1(new_n6725_), .A2(new_n6735_), .ZN(new_n6736_));
  INV_X1     g05734(.I(\A[153] ), .ZN(new_n6737_));
  NOR3_X1    g05735(.A1(new_n6719_), .A2(new_n6723_), .A3(new_n6737_), .ZN(new_n6738_));
  NAND2_X1   g05736(.A1(new_n6722_), .A2(\A[152] ), .ZN(new_n6739_));
  AOI21_X1   g05737(.A1(new_n6739_), .A2(new_n6720_), .B(\A[153] ), .ZN(new_n6740_));
  NOR2_X1    g05738(.A1(new_n6740_), .A2(new_n6738_), .ZN(new_n6741_));
  AOI21_X1   g05739(.A1(\A[154] ), .A2(new_n6727_), .B(new_n6726_), .ZN(new_n6742_));
  NAND2_X1   g05740(.A1(new_n6742_), .A2(new_n6732_), .ZN(new_n6743_));
  NOR2_X1    g05741(.A1(new_n6728_), .A2(new_n6730_), .ZN(new_n6744_));
  OAI21_X1   g05742(.A1(\A[156] ), .A2(new_n6744_), .B(new_n6743_), .ZN(new_n6745_));
  NOR2_X1    g05743(.A1(new_n6745_), .A2(new_n6741_), .ZN(new_n6746_));
  NOR2_X1    g05744(.A1(new_n6746_), .A2(new_n6736_), .ZN(new_n6747_));
  XOR2_X1    g05745(.A1(\A[154] ), .A2(\A[155] ), .Z(new_n6748_));
  NOR2_X1    g05746(.A1(new_n6729_), .A2(new_n6727_), .ZN(new_n6749_));
  AOI21_X1   g05747(.A1(new_n6748_), .A2(\A[156] ), .B(new_n6749_), .ZN(new_n6750_));
  NAND2_X1   g05748(.A1(new_n6739_), .A2(new_n6720_), .ZN(new_n6751_));
  NOR2_X1    g05749(.A1(new_n6722_), .A2(new_n6718_), .ZN(new_n6752_));
  AOI21_X1   g05750(.A1(new_n6751_), .A2(\A[153] ), .B(new_n6752_), .ZN(new_n6753_));
  OAI22_X1   g05751(.A1(new_n6738_), .A2(new_n6740_), .B1(new_n6734_), .B2(new_n6731_), .ZN(new_n6754_));
  NOR3_X1    g05752(.A1(new_n6754_), .A2(new_n6750_), .A3(new_n6753_), .ZN(new_n6755_));
  NOR2_X1    g05753(.A1(new_n6747_), .A2(new_n6755_), .ZN(new_n6756_));
  NAND2_X1   g05754(.A1(new_n6756_), .A2(new_n6717_), .ZN(new_n6757_));
  INV_X1     g05755(.I(new_n6717_), .ZN(new_n6758_));
  NAND2_X1   g05756(.A1(new_n6745_), .A2(new_n6741_), .ZN(new_n6759_));
  NAND2_X1   g05757(.A1(new_n6725_), .A2(new_n6735_), .ZN(new_n6760_));
  NAND2_X1   g05758(.A1(new_n6759_), .A2(new_n6760_), .ZN(new_n6761_));
  INV_X1     g05759(.I(new_n6749_), .ZN(new_n6762_));
  OAI21_X1   g05760(.A1(new_n6744_), .A2(new_n6726_), .B(new_n6762_), .ZN(new_n6763_));
  INV_X1     g05761(.I(new_n6752_), .ZN(new_n6764_));
  OAI21_X1   g05762(.A1(new_n6724_), .A2(new_n6737_), .B(new_n6764_), .ZN(new_n6765_));
  NAND4_X1   g05763(.A1(new_n6745_), .A2(new_n6725_), .A3(new_n6763_), .A4(new_n6765_), .ZN(new_n6766_));
  NAND2_X1   g05764(.A1(new_n6761_), .A2(new_n6766_), .ZN(new_n6767_));
  NAND2_X1   g05765(.A1(new_n6758_), .A2(new_n6767_), .ZN(new_n6768_));
  NAND2_X1   g05766(.A1(new_n6768_), .A2(new_n6757_), .ZN(new_n6769_));
  NAND3_X1   g05767(.A1(new_n6769_), .A2(new_n6652_), .A3(new_n6675_), .ZN(new_n6770_));
  NAND2_X1   g05768(.A1(new_n6675_), .A2(new_n6652_), .ZN(new_n6771_));
  NAND3_X1   g05769(.A1(new_n6771_), .A2(new_n6757_), .A3(new_n6768_), .ZN(new_n6772_));
  NAND2_X1   g05770(.A1(new_n6770_), .A2(new_n6772_), .ZN(new_n6773_));
  INV_X1     g05771(.I(\A[145] ), .ZN(new_n6774_));
  NAND2_X1   g05772(.A1(new_n6774_), .A2(\A[146] ), .ZN(new_n6775_));
  INV_X1     g05773(.I(\A[146] ), .ZN(new_n6776_));
  NAND2_X1   g05774(.A1(new_n6776_), .A2(\A[145] ), .ZN(new_n6777_));
  NAND3_X1   g05775(.A1(new_n6775_), .A2(new_n6777_), .A3(\A[147] ), .ZN(new_n6778_));
  INV_X1     g05776(.I(\A[147] ), .ZN(new_n6779_));
  NOR2_X1    g05777(.A1(new_n6776_), .A2(\A[145] ), .ZN(new_n6780_));
  NOR2_X1    g05778(.A1(new_n6774_), .A2(\A[146] ), .ZN(new_n6781_));
  OAI21_X1   g05779(.A1(new_n6780_), .A2(new_n6781_), .B(new_n6779_), .ZN(new_n6782_));
  NAND2_X1   g05780(.A1(new_n6782_), .A2(new_n6778_), .ZN(new_n6783_));
  INV_X1     g05781(.I(\A[150] ), .ZN(new_n6784_));
  INV_X1     g05782(.I(\A[148] ), .ZN(new_n6785_));
  NAND2_X1   g05783(.A1(new_n6785_), .A2(\A[149] ), .ZN(new_n6786_));
  INV_X1     g05784(.I(\A[149] ), .ZN(new_n6787_));
  AOI21_X1   g05785(.A1(\A[148] ), .A2(new_n6787_), .B(new_n6784_), .ZN(new_n6788_));
  XOR2_X1    g05786(.A1(\A[148] ), .A2(\A[149] ), .Z(new_n6789_));
  AOI22_X1   g05787(.A1(new_n6789_), .A2(new_n6784_), .B1(new_n6786_), .B2(new_n6788_), .ZN(new_n6790_));
  NOR2_X1    g05788(.A1(new_n6783_), .A2(new_n6790_), .ZN(new_n6791_));
  NOR3_X1    g05789(.A1(new_n6780_), .A2(new_n6781_), .A3(new_n6779_), .ZN(new_n6792_));
  AOI21_X1   g05790(.A1(new_n6775_), .A2(new_n6777_), .B(\A[147] ), .ZN(new_n6793_));
  NOR2_X1    g05791(.A1(new_n6793_), .A2(new_n6792_), .ZN(new_n6794_));
  NAND2_X1   g05792(.A1(new_n6788_), .A2(new_n6786_), .ZN(new_n6795_));
  NOR2_X1    g05793(.A1(new_n6787_), .A2(\A[148] ), .ZN(new_n6796_));
  NOR2_X1    g05794(.A1(new_n6785_), .A2(\A[149] ), .ZN(new_n6797_));
  OAI21_X1   g05795(.A1(new_n6796_), .A2(new_n6797_), .B(new_n6784_), .ZN(new_n6798_));
  NAND2_X1   g05796(.A1(new_n6795_), .A2(new_n6798_), .ZN(new_n6799_));
  NOR2_X1    g05797(.A1(new_n6794_), .A2(new_n6799_), .ZN(new_n6800_));
  NOR2_X1    g05798(.A1(new_n6800_), .A2(new_n6791_), .ZN(new_n6801_));
  NOR2_X1    g05799(.A1(new_n6785_), .A2(new_n6787_), .ZN(new_n6802_));
  AOI21_X1   g05800(.A1(new_n6789_), .A2(\A[150] ), .B(new_n6802_), .ZN(new_n6803_));
  NAND2_X1   g05801(.A1(new_n6775_), .A2(new_n6777_), .ZN(new_n6804_));
  NAND2_X1   g05802(.A1(\A[145] ), .A2(\A[146] ), .ZN(new_n6805_));
  INV_X1     g05803(.I(new_n6805_), .ZN(new_n6806_));
  AOI21_X1   g05804(.A1(new_n6804_), .A2(\A[147] ), .B(new_n6806_), .ZN(new_n6807_));
  NOR3_X1    g05805(.A1(new_n6796_), .A2(new_n6797_), .A3(new_n6784_), .ZN(new_n6808_));
  NAND2_X1   g05806(.A1(new_n6787_), .A2(\A[148] ), .ZN(new_n6809_));
  AOI21_X1   g05807(.A1(new_n6786_), .A2(new_n6809_), .B(\A[150] ), .ZN(new_n6810_));
  OAI22_X1   g05808(.A1(new_n6808_), .A2(new_n6810_), .B1(new_n6793_), .B2(new_n6792_), .ZN(new_n6811_));
  NOR3_X1    g05809(.A1(new_n6811_), .A2(new_n6803_), .A3(new_n6807_), .ZN(new_n6812_));
  NOR2_X1    g05810(.A1(new_n6801_), .A2(new_n6812_), .ZN(new_n6813_));
  INV_X1     g05811(.I(\A[141] ), .ZN(new_n6814_));
  INV_X1     g05812(.I(\A[139] ), .ZN(new_n6815_));
  NAND2_X1   g05813(.A1(new_n6815_), .A2(\A[140] ), .ZN(new_n6816_));
  INV_X1     g05814(.I(\A[140] ), .ZN(new_n6817_));
  AOI21_X1   g05815(.A1(\A[139] ), .A2(new_n6817_), .B(new_n6814_), .ZN(new_n6818_));
  XOR2_X1    g05816(.A1(\A[139] ), .A2(\A[140] ), .Z(new_n6819_));
  AOI22_X1   g05817(.A1(new_n6819_), .A2(new_n6814_), .B1(new_n6816_), .B2(new_n6818_), .ZN(new_n6820_));
  INV_X1     g05818(.I(\A[142] ), .ZN(new_n6821_));
  NAND2_X1   g05819(.A1(new_n6821_), .A2(\A[143] ), .ZN(new_n6822_));
  INV_X1     g05820(.I(\A[143] ), .ZN(new_n6823_));
  NAND2_X1   g05821(.A1(new_n6823_), .A2(\A[142] ), .ZN(new_n6824_));
  NAND3_X1   g05822(.A1(new_n6822_), .A2(new_n6824_), .A3(\A[144] ), .ZN(new_n6825_));
  INV_X1     g05823(.I(\A[144] ), .ZN(new_n6826_));
  NOR2_X1    g05824(.A1(new_n6823_), .A2(\A[142] ), .ZN(new_n6827_));
  NOR2_X1    g05825(.A1(new_n6821_), .A2(\A[143] ), .ZN(new_n6828_));
  OAI21_X1   g05826(.A1(new_n6827_), .A2(new_n6828_), .B(new_n6826_), .ZN(new_n6829_));
  NAND2_X1   g05827(.A1(new_n6829_), .A2(new_n6825_), .ZN(new_n6830_));
  NAND2_X1   g05828(.A1(new_n6830_), .A2(new_n6820_), .ZN(new_n6831_));
  NAND2_X1   g05829(.A1(new_n6818_), .A2(new_n6816_), .ZN(new_n6832_));
  NOR2_X1    g05830(.A1(new_n6817_), .A2(\A[139] ), .ZN(new_n6833_));
  NOR2_X1    g05831(.A1(new_n6815_), .A2(\A[140] ), .ZN(new_n6834_));
  OAI21_X1   g05832(.A1(new_n6833_), .A2(new_n6834_), .B(new_n6814_), .ZN(new_n6835_));
  NAND2_X1   g05833(.A1(new_n6832_), .A2(new_n6835_), .ZN(new_n6836_));
  NOR3_X1    g05834(.A1(new_n6827_), .A2(new_n6828_), .A3(new_n6826_), .ZN(new_n6837_));
  AOI21_X1   g05835(.A1(new_n6822_), .A2(new_n6824_), .B(\A[144] ), .ZN(new_n6838_));
  NOR2_X1    g05836(.A1(new_n6838_), .A2(new_n6837_), .ZN(new_n6839_));
  NAND2_X1   g05837(.A1(new_n6839_), .A2(new_n6836_), .ZN(new_n6840_));
  NAND2_X1   g05838(.A1(new_n6840_), .A2(new_n6831_), .ZN(new_n6841_));
  NOR2_X1    g05839(.A1(new_n6827_), .A2(new_n6828_), .ZN(new_n6842_));
  NAND2_X1   g05840(.A1(\A[142] ), .A2(\A[143] ), .ZN(new_n6843_));
  OAI21_X1   g05841(.A1(new_n6842_), .A2(new_n6826_), .B(new_n6843_), .ZN(new_n6844_));
  NOR2_X1    g05842(.A1(new_n6833_), .A2(new_n6834_), .ZN(new_n6845_));
  NOR2_X1    g05843(.A1(new_n6815_), .A2(new_n6817_), .ZN(new_n6846_));
  INV_X1     g05844(.I(new_n6846_), .ZN(new_n6847_));
  OAI21_X1   g05845(.A1(new_n6845_), .A2(new_n6814_), .B(new_n6847_), .ZN(new_n6848_));
  AOI22_X1   g05846(.A1(new_n6832_), .A2(new_n6835_), .B1(new_n6829_), .B2(new_n6825_), .ZN(new_n6849_));
  NAND3_X1   g05847(.A1(new_n6849_), .A2(new_n6844_), .A3(new_n6848_), .ZN(new_n6850_));
  NAND2_X1   g05848(.A1(new_n6841_), .A2(new_n6850_), .ZN(new_n6851_));
  NOR2_X1    g05849(.A1(new_n6813_), .A2(new_n6851_), .ZN(new_n6852_));
  NAND2_X1   g05850(.A1(new_n6794_), .A2(new_n6799_), .ZN(new_n6853_));
  NAND2_X1   g05851(.A1(new_n6783_), .A2(new_n6790_), .ZN(new_n6854_));
  NAND2_X1   g05852(.A1(new_n6853_), .A2(new_n6854_), .ZN(new_n6855_));
  NOR2_X1    g05853(.A1(new_n6796_), .A2(new_n6797_), .ZN(new_n6856_));
  INV_X1     g05854(.I(new_n6802_), .ZN(new_n6857_));
  OAI21_X1   g05855(.A1(new_n6856_), .A2(new_n6784_), .B(new_n6857_), .ZN(new_n6858_));
  XNOR2_X1   g05856(.A1(\A[145] ), .A2(\A[146] ), .ZN(new_n6859_));
  OAI21_X1   g05857(.A1(new_n6859_), .A2(new_n6779_), .B(new_n6805_), .ZN(new_n6860_));
  AOI22_X1   g05858(.A1(new_n6795_), .A2(new_n6798_), .B1(new_n6782_), .B2(new_n6778_), .ZN(new_n6861_));
  NAND3_X1   g05859(.A1(new_n6861_), .A2(new_n6858_), .A3(new_n6860_), .ZN(new_n6862_));
  NAND2_X1   g05860(.A1(new_n6855_), .A2(new_n6862_), .ZN(new_n6863_));
  NOR2_X1    g05861(.A1(new_n6839_), .A2(new_n6836_), .ZN(new_n6864_));
  NOR2_X1    g05862(.A1(new_n6830_), .A2(new_n6820_), .ZN(new_n6865_));
  NOR2_X1    g05863(.A1(new_n6864_), .A2(new_n6865_), .ZN(new_n6866_));
  XOR2_X1    g05864(.A1(\A[142] ), .A2(\A[143] ), .Z(new_n6867_));
  INV_X1     g05865(.I(new_n6843_), .ZN(new_n6868_));
  AOI21_X1   g05866(.A1(new_n6867_), .A2(\A[144] ), .B(new_n6868_), .ZN(new_n6869_));
  AOI21_X1   g05867(.A1(new_n6819_), .A2(\A[141] ), .B(new_n6846_), .ZN(new_n6870_));
  NOR3_X1    g05868(.A1(new_n6833_), .A2(new_n6834_), .A3(new_n6814_), .ZN(new_n6871_));
  NAND2_X1   g05869(.A1(new_n6817_), .A2(\A[139] ), .ZN(new_n6872_));
  AOI21_X1   g05870(.A1(new_n6816_), .A2(new_n6872_), .B(\A[141] ), .ZN(new_n6873_));
  OAI22_X1   g05871(.A1(new_n6871_), .A2(new_n6873_), .B1(new_n6838_), .B2(new_n6837_), .ZN(new_n6874_));
  NOR3_X1    g05872(.A1(new_n6874_), .A2(new_n6869_), .A3(new_n6870_), .ZN(new_n6875_));
  NOR2_X1    g05873(.A1(new_n6866_), .A2(new_n6875_), .ZN(new_n6876_));
  NOR2_X1    g05874(.A1(new_n6876_), .A2(new_n6863_), .ZN(new_n6877_));
  NOR2_X1    g05875(.A1(new_n6852_), .A2(new_n6877_), .ZN(new_n6878_));
  INV_X1     g05876(.I(\A[133] ), .ZN(new_n6879_));
  NAND2_X1   g05877(.A1(new_n6879_), .A2(\A[134] ), .ZN(new_n6880_));
  INV_X1     g05878(.I(\A[134] ), .ZN(new_n6881_));
  NAND2_X1   g05879(.A1(new_n6881_), .A2(\A[133] ), .ZN(new_n6882_));
  NAND3_X1   g05880(.A1(new_n6880_), .A2(new_n6882_), .A3(\A[135] ), .ZN(new_n6883_));
  INV_X1     g05881(.I(new_n6883_), .ZN(new_n6884_));
  AOI21_X1   g05882(.A1(new_n6880_), .A2(new_n6882_), .B(\A[135] ), .ZN(new_n6885_));
  NOR2_X1    g05883(.A1(new_n6884_), .A2(new_n6885_), .ZN(new_n6886_));
  INV_X1     g05884(.I(\A[136] ), .ZN(new_n6887_));
  NAND2_X1   g05885(.A1(new_n6887_), .A2(\A[137] ), .ZN(new_n6888_));
  INV_X1     g05886(.I(\A[137] ), .ZN(new_n6889_));
  NAND2_X1   g05887(.A1(new_n6889_), .A2(\A[136] ), .ZN(new_n6890_));
  NAND3_X1   g05888(.A1(new_n6888_), .A2(new_n6890_), .A3(\A[138] ), .ZN(new_n6891_));
  INV_X1     g05889(.I(\A[138] ), .ZN(new_n6892_));
  NOR2_X1    g05890(.A1(new_n6889_), .A2(\A[136] ), .ZN(new_n6893_));
  NOR2_X1    g05891(.A1(new_n6887_), .A2(\A[137] ), .ZN(new_n6894_));
  OAI21_X1   g05892(.A1(new_n6893_), .A2(new_n6894_), .B(new_n6892_), .ZN(new_n6895_));
  NAND2_X1   g05893(.A1(new_n6895_), .A2(new_n6891_), .ZN(new_n6896_));
  NAND2_X1   g05894(.A1(new_n6886_), .A2(new_n6896_), .ZN(new_n6897_));
  INV_X1     g05895(.I(\A[135] ), .ZN(new_n6898_));
  NOR2_X1    g05896(.A1(new_n6881_), .A2(\A[133] ), .ZN(new_n6899_));
  NOR2_X1    g05897(.A1(new_n6879_), .A2(\A[134] ), .ZN(new_n6900_));
  OAI21_X1   g05898(.A1(new_n6899_), .A2(new_n6900_), .B(new_n6898_), .ZN(new_n6901_));
  NAND2_X1   g05899(.A1(new_n6901_), .A2(new_n6883_), .ZN(new_n6902_));
  NOR3_X1    g05900(.A1(new_n6893_), .A2(new_n6894_), .A3(new_n6892_), .ZN(new_n6903_));
  AOI21_X1   g05901(.A1(new_n6888_), .A2(new_n6890_), .B(\A[138] ), .ZN(new_n6904_));
  NOR2_X1    g05902(.A1(new_n6904_), .A2(new_n6903_), .ZN(new_n6905_));
  NAND2_X1   g05903(.A1(new_n6905_), .A2(new_n6902_), .ZN(new_n6906_));
  NAND2_X1   g05904(.A1(new_n6897_), .A2(new_n6906_), .ZN(new_n6907_));
  NOR2_X1    g05905(.A1(new_n6893_), .A2(new_n6894_), .ZN(new_n6908_));
  NOR2_X1    g05906(.A1(new_n6887_), .A2(new_n6889_), .ZN(new_n6909_));
  INV_X1     g05907(.I(new_n6909_), .ZN(new_n6910_));
  OAI21_X1   g05908(.A1(new_n6908_), .A2(new_n6892_), .B(new_n6910_), .ZN(new_n6911_));
  NOR2_X1    g05909(.A1(new_n6899_), .A2(new_n6900_), .ZN(new_n6912_));
  NOR2_X1    g05910(.A1(new_n6879_), .A2(new_n6881_), .ZN(new_n6913_));
  INV_X1     g05911(.I(new_n6913_), .ZN(new_n6914_));
  OAI21_X1   g05912(.A1(new_n6912_), .A2(new_n6898_), .B(new_n6914_), .ZN(new_n6915_));
  AOI22_X1   g05913(.A1(new_n6883_), .A2(new_n6901_), .B1(new_n6895_), .B2(new_n6891_), .ZN(new_n6916_));
  NAND3_X1   g05914(.A1(new_n6916_), .A2(new_n6911_), .A3(new_n6915_), .ZN(new_n6917_));
  NAND2_X1   g05915(.A1(new_n6907_), .A2(new_n6917_), .ZN(new_n6918_));
  INV_X1     g05916(.I(\A[128] ), .ZN(new_n6919_));
  NOR2_X1    g05917(.A1(new_n6919_), .A2(\A[127] ), .ZN(new_n6920_));
  INV_X1     g05918(.I(\A[127] ), .ZN(new_n6921_));
  OAI21_X1   g05919(.A1(new_n6921_), .A2(\A[128] ), .B(\A[129] ), .ZN(new_n6922_));
  NOR2_X1    g05920(.A1(new_n6921_), .A2(\A[128] ), .ZN(new_n6923_));
  NOR2_X1    g05921(.A1(new_n6920_), .A2(new_n6923_), .ZN(new_n6924_));
  OAI22_X1   g05922(.A1(new_n6924_), .A2(\A[129] ), .B1(new_n6920_), .B2(new_n6922_), .ZN(new_n6925_));
  INV_X1     g05923(.I(\A[132] ), .ZN(new_n6926_));
  INV_X1     g05924(.I(\A[131] ), .ZN(new_n6927_));
  NOR2_X1    g05925(.A1(new_n6927_), .A2(\A[130] ), .ZN(new_n6928_));
  INV_X1     g05926(.I(\A[130] ), .ZN(new_n6929_));
  NOR2_X1    g05927(.A1(new_n6929_), .A2(\A[131] ), .ZN(new_n6930_));
  NOR3_X1    g05928(.A1(new_n6928_), .A2(new_n6930_), .A3(new_n6926_), .ZN(new_n6931_));
  NAND2_X1   g05929(.A1(new_n6929_), .A2(\A[131] ), .ZN(new_n6932_));
  NAND2_X1   g05930(.A1(new_n6927_), .A2(\A[130] ), .ZN(new_n6933_));
  AOI21_X1   g05931(.A1(new_n6932_), .A2(new_n6933_), .B(\A[132] ), .ZN(new_n6934_));
  NOR2_X1    g05932(.A1(new_n6934_), .A2(new_n6931_), .ZN(new_n6935_));
  NOR2_X1    g05933(.A1(new_n6925_), .A2(new_n6935_), .ZN(new_n6936_));
  NOR2_X1    g05934(.A1(new_n6922_), .A2(new_n6920_), .ZN(new_n6937_));
  NAND2_X1   g05935(.A1(new_n6921_), .A2(\A[128] ), .ZN(new_n6938_));
  NAND2_X1   g05936(.A1(new_n6919_), .A2(\A[127] ), .ZN(new_n6939_));
  AOI21_X1   g05937(.A1(new_n6938_), .A2(new_n6939_), .B(\A[129] ), .ZN(new_n6940_));
  NOR2_X1    g05938(.A1(new_n6940_), .A2(new_n6937_), .ZN(new_n6941_));
  NAND2_X1   g05939(.A1(new_n6933_), .A2(\A[132] ), .ZN(new_n6942_));
  NOR2_X1    g05940(.A1(new_n6928_), .A2(new_n6930_), .ZN(new_n6943_));
  OAI22_X1   g05941(.A1(new_n6943_), .A2(\A[132] ), .B1(new_n6942_), .B2(new_n6928_), .ZN(new_n6944_));
  NOR2_X1    g05942(.A1(new_n6944_), .A2(new_n6941_), .ZN(new_n6945_));
  NOR2_X1    g05943(.A1(new_n6936_), .A2(new_n6945_), .ZN(new_n6946_));
  XOR2_X1    g05944(.A1(\A[130] ), .A2(\A[131] ), .Z(new_n6947_));
  NOR2_X1    g05945(.A1(new_n6929_), .A2(new_n6927_), .ZN(new_n6948_));
  AOI21_X1   g05946(.A1(new_n6947_), .A2(\A[132] ), .B(new_n6948_), .ZN(new_n6949_));
  XOR2_X1    g05947(.A1(\A[127] ), .A2(\A[128] ), .Z(new_n6950_));
  NOR2_X1    g05948(.A1(new_n6921_), .A2(new_n6919_), .ZN(new_n6951_));
  AOI21_X1   g05949(.A1(new_n6950_), .A2(\A[129] ), .B(new_n6951_), .ZN(new_n6952_));
  OAI22_X1   g05950(.A1(new_n6931_), .A2(new_n6934_), .B1(new_n6940_), .B2(new_n6937_), .ZN(new_n6953_));
  NOR3_X1    g05951(.A1(new_n6953_), .A2(new_n6949_), .A3(new_n6952_), .ZN(new_n6954_));
  NOR2_X1    g05952(.A1(new_n6946_), .A2(new_n6954_), .ZN(new_n6955_));
  NAND2_X1   g05953(.A1(new_n6918_), .A2(new_n6955_), .ZN(new_n6956_));
  NOR2_X1    g05954(.A1(new_n6905_), .A2(new_n6902_), .ZN(new_n6957_));
  NOR2_X1    g05955(.A1(new_n6886_), .A2(new_n6896_), .ZN(new_n6958_));
  NOR2_X1    g05956(.A1(new_n6958_), .A2(new_n6957_), .ZN(new_n6959_));
  INV_X1     g05957(.I(new_n6917_), .ZN(new_n6960_));
  NOR2_X1    g05958(.A1(new_n6959_), .A2(new_n6960_), .ZN(new_n6961_));
  NAND2_X1   g05959(.A1(new_n6944_), .A2(new_n6941_), .ZN(new_n6962_));
  NAND2_X1   g05960(.A1(new_n6925_), .A2(new_n6935_), .ZN(new_n6963_));
  NAND2_X1   g05961(.A1(new_n6963_), .A2(new_n6962_), .ZN(new_n6964_));
  INV_X1     g05962(.I(new_n6948_), .ZN(new_n6965_));
  OAI21_X1   g05963(.A1(new_n6943_), .A2(new_n6926_), .B(new_n6965_), .ZN(new_n6966_));
  INV_X1     g05964(.I(\A[129] ), .ZN(new_n6967_));
  INV_X1     g05965(.I(new_n6951_), .ZN(new_n6968_));
  OAI21_X1   g05966(.A1(new_n6924_), .A2(new_n6967_), .B(new_n6968_), .ZN(new_n6969_));
  NAND4_X1   g05967(.A1(new_n6944_), .A2(new_n6925_), .A3(new_n6966_), .A4(new_n6969_), .ZN(new_n6970_));
  NAND2_X1   g05968(.A1(new_n6964_), .A2(new_n6970_), .ZN(new_n6971_));
  NAND2_X1   g05969(.A1(new_n6961_), .A2(new_n6971_), .ZN(new_n6972_));
  NAND2_X1   g05970(.A1(new_n6972_), .A2(new_n6956_), .ZN(new_n6973_));
  NAND2_X1   g05971(.A1(new_n6973_), .A2(new_n6878_), .ZN(new_n6974_));
  NAND2_X1   g05972(.A1(new_n6876_), .A2(new_n6863_), .ZN(new_n6975_));
  NAND2_X1   g05973(.A1(new_n6813_), .A2(new_n6851_), .ZN(new_n6976_));
  NAND2_X1   g05974(.A1(new_n6976_), .A2(new_n6975_), .ZN(new_n6977_));
  NOR2_X1    g05975(.A1(new_n6961_), .A2(new_n6971_), .ZN(new_n6978_));
  NOR2_X1    g05976(.A1(new_n6918_), .A2(new_n6955_), .ZN(new_n6979_));
  NOR2_X1    g05977(.A1(new_n6978_), .A2(new_n6979_), .ZN(new_n6980_));
  NAND2_X1   g05978(.A1(new_n6980_), .A2(new_n6977_), .ZN(new_n6981_));
  NAND2_X1   g05979(.A1(new_n6974_), .A2(new_n6981_), .ZN(new_n6982_));
  XOR2_X1    g05980(.A1(new_n6773_), .A2(new_n6982_), .Z(new_n6983_));
  INV_X1     g05981(.I(\A[123] ), .ZN(new_n6984_));
  INV_X1     g05982(.I(\A[121] ), .ZN(new_n6985_));
  NAND2_X1   g05983(.A1(new_n6985_), .A2(\A[122] ), .ZN(new_n6986_));
  INV_X1     g05984(.I(\A[122] ), .ZN(new_n6987_));
  AOI21_X1   g05985(.A1(\A[121] ), .A2(new_n6987_), .B(new_n6984_), .ZN(new_n6988_));
  XOR2_X1    g05986(.A1(\A[121] ), .A2(\A[122] ), .Z(new_n6989_));
  AOI22_X1   g05987(.A1(new_n6989_), .A2(new_n6984_), .B1(new_n6986_), .B2(new_n6988_), .ZN(new_n6990_));
  INV_X1     g05988(.I(\A[124] ), .ZN(new_n6991_));
  NAND2_X1   g05989(.A1(new_n6991_), .A2(\A[125] ), .ZN(new_n6992_));
  INV_X1     g05990(.I(\A[125] ), .ZN(new_n6993_));
  INV_X1     g05991(.I(\A[126] ), .ZN(new_n6994_));
  AOI21_X1   g05992(.A1(\A[124] ), .A2(new_n6993_), .B(new_n6994_), .ZN(new_n6995_));
  NAND2_X1   g05993(.A1(new_n6995_), .A2(new_n6992_), .ZN(new_n6996_));
  NOR2_X1    g05994(.A1(new_n6993_), .A2(\A[124] ), .ZN(new_n6997_));
  NOR2_X1    g05995(.A1(new_n6991_), .A2(\A[125] ), .ZN(new_n6998_));
  OAI21_X1   g05996(.A1(new_n6997_), .A2(new_n6998_), .B(new_n6994_), .ZN(new_n6999_));
  NAND2_X1   g05997(.A1(new_n6996_), .A2(new_n6999_), .ZN(new_n7000_));
  NAND2_X1   g05998(.A1(new_n7000_), .A2(new_n6990_), .ZN(new_n7001_));
  NAND2_X1   g05999(.A1(new_n6988_), .A2(new_n6986_), .ZN(new_n7002_));
  NOR2_X1    g06000(.A1(new_n6987_), .A2(\A[121] ), .ZN(new_n7003_));
  NOR2_X1    g06001(.A1(new_n6985_), .A2(\A[122] ), .ZN(new_n7004_));
  OAI21_X1   g06002(.A1(new_n7003_), .A2(new_n7004_), .B(new_n6984_), .ZN(new_n7005_));
  NAND2_X1   g06003(.A1(new_n7002_), .A2(new_n7005_), .ZN(new_n7006_));
  XOR2_X1    g06004(.A1(\A[124] ), .A2(\A[125] ), .Z(new_n7007_));
  AOI22_X1   g06005(.A1(new_n7007_), .A2(new_n6994_), .B1(new_n6992_), .B2(new_n6995_), .ZN(new_n7008_));
  NAND2_X1   g06006(.A1(new_n7006_), .A2(new_n7008_), .ZN(new_n7009_));
  NAND2_X1   g06007(.A1(new_n7001_), .A2(new_n7009_), .ZN(new_n7010_));
  NOR2_X1    g06008(.A1(new_n6997_), .A2(new_n6998_), .ZN(new_n7011_));
  NAND2_X1   g06009(.A1(\A[124] ), .A2(\A[125] ), .ZN(new_n7012_));
  OAI21_X1   g06010(.A1(new_n7011_), .A2(new_n6994_), .B(new_n7012_), .ZN(new_n7013_));
  NOR2_X1    g06011(.A1(new_n7003_), .A2(new_n7004_), .ZN(new_n7014_));
  NAND2_X1   g06012(.A1(\A[121] ), .A2(\A[122] ), .ZN(new_n7015_));
  OAI21_X1   g06013(.A1(new_n7014_), .A2(new_n6984_), .B(new_n7015_), .ZN(new_n7016_));
  AOI22_X1   g06014(.A1(new_n7002_), .A2(new_n7005_), .B1(new_n6996_), .B2(new_n6999_), .ZN(new_n7017_));
  NAND3_X1   g06015(.A1(new_n7017_), .A2(new_n7013_), .A3(new_n7016_), .ZN(new_n7018_));
  NAND2_X1   g06016(.A1(new_n7010_), .A2(new_n7018_), .ZN(new_n7019_));
  INV_X1     g06017(.I(\A[115] ), .ZN(new_n7020_));
  NAND2_X1   g06018(.A1(new_n7020_), .A2(\A[116] ), .ZN(new_n7021_));
  INV_X1     g06019(.I(\A[116] ), .ZN(new_n7022_));
  INV_X1     g06020(.I(\A[117] ), .ZN(new_n7023_));
  AOI21_X1   g06021(.A1(\A[115] ), .A2(new_n7022_), .B(new_n7023_), .ZN(new_n7024_));
  NAND2_X1   g06022(.A1(new_n7024_), .A2(new_n7021_), .ZN(new_n7025_));
  NOR2_X1    g06023(.A1(new_n7022_), .A2(\A[115] ), .ZN(new_n7026_));
  NOR2_X1    g06024(.A1(new_n7020_), .A2(\A[116] ), .ZN(new_n7027_));
  OAI21_X1   g06025(.A1(new_n7026_), .A2(new_n7027_), .B(new_n7023_), .ZN(new_n7028_));
  NAND2_X1   g06026(.A1(new_n7025_), .A2(new_n7028_), .ZN(new_n7029_));
  INV_X1     g06027(.I(\A[119] ), .ZN(new_n7030_));
  NOR2_X1    g06028(.A1(new_n7030_), .A2(\A[118] ), .ZN(new_n7031_));
  INV_X1     g06029(.I(\A[118] ), .ZN(new_n7032_));
  OAI21_X1   g06030(.A1(new_n7032_), .A2(\A[119] ), .B(\A[120] ), .ZN(new_n7033_));
  NOR2_X1    g06031(.A1(new_n7033_), .A2(new_n7031_), .ZN(new_n7034_));
  NAND2_X1   g06032(.A1(new_n7032_), .A2(\A[119] ), .ZN(new_n7035_));
  NAND2_X1   g06033(.A1(new_n7030_), .A2(\A[118] ), .ZN(new_n7036_));
  AOI21_X1   g06034(.A1(new_n7035_), .A2(new_n7036_), .B(\A[120] ), .ZN(new_n7037_));
  NOR2_X1    g06035(.A1(new_n7037_), .A2(new_n7034_), .ZN(new_n7038_));
  NOR2_X1    g06036(.A1(new_n7029_), .A2(new_n7038_), .ZN(new_n7039_));
  XOR2_X1    g06037(.A1(\A[115] ), .A2(\A[116] ), .Z(new_n7040_));
  AOI22_X1   g06038(.A1(new_n7040_), .A2(new_n7023_), .B1(new_n7021_), .B2(new_n7024_), .ZN(new_n7041_));
  NAND3_X1   g06039(.A1(new_n7035_), .A2(new_n7036_), .A3(\A[120] ), .ZN(new_n7042_));
  INV_X1     g06040(.I(\A[120] ), .ZN(new_n7043_));
  NOR2_X1    g06041(.A1(new_n7032_), .A2(\A[119] ), .ZN(new_n7044_));
  OAI21_X1   g06042(.A1(new_n7031_), .A2(new_n7044_), .B(new_n7043_), .ZN(new_n7045_));
  NAND2_X1   g06043(.A1(new_n7045_), .A2(new_n7042_), .ZN(new_n7046_));
  NOR2_X1    g06044(.A1(new_n7046_), .A2(new_n7041_), .ZN(new_n7047_));
  NOR2_X1    g06045(.A1(new_n7039_), .A2(new_n7047_), .ZN(new_n7048_));
  NAND2_X1   g06046(.A1(new_n7035_), .A2(new_n7036_), .ZN(new_n7049_));
  NOR2_X1    g06047(.A1(new_n7032_), .A2(new_n7030_), .ZN(new_n7050_));
  AOI21_X1   g06048(.A1(new_n7049_), .A2(\A[120] ), .B(new_n7050_), .ZN(new_n7051_));
  NOR2_X1    g06049(.A1(new_n7020_), .A2(new_n7022_), .ZN(new_n7052_));
  AOI21_X1   g06050(.A1(new_n7040_), .A2(\A[117] ), .B(new_n7052_), .ZN(new_n7053_));
  NOR3_X1    g06051(.A1(new_n7026_), .A2(new_n7027_), .A3(new_n7023_), .ZN(new_n7054_));
  NAND2_X1   g06052(.A1(new_n7022_), .A2(\A[115] ), .ZN(new_n7055_));
  AOI21_X1   g06053(.A1(new_n7021_), .A2(new_n7055_), .B(\A[117] ), .ZN(new_n7056_));
  OAI22_X1   g06054(.A1(new_n7054_), .A2(new_n7056_), .B1(new_n7037_), .B2(new_n7034_), .ZN(new_n7057_));
  NOR3_X1    g06055(.A1(new_n7057_), .A2(new_n7051_), .A3(new_n7053_), .ZN(new_n7058_));
  NOR2_X1    g06056(.A1(new_n7048_), .A2(new_n7058_), .ZN(new_n7059_));
  NAND2_X1   g06057(.A1(new_n7059_), .A2(new_n7019_), .ZN(new_n7060_));
  NAND2_X1   g06058(.A1(new_n7046_), .A2(new_n7041_), .ZN(new_n7061_));
  NAND2_X1   g06059(.A1(new_n7029_), .A2(new_n7038_), .ZN(new_n7062_));
  NAND2_X1   g06060(.A1(new_n7062_), .A2(new_n7061_), .ZN(new_n7063_));
  NOR2_X1    g06061(.A1(new_n7031_), .A2(new_n7044_), .ZN(new_n7064_));
  INV_X1     g06062(.I(new_n7050_), .ZN(new_n7065_));
  OAI21_X1   g06063(.A1(new_n7064_), .A2(new_n7043_), .B(new_n7065_), .ZN(new_n7066_));
  NOR2_X1    g06064(.A1(new_n7026_), .A2(new_n7027_), .ZN(new_n7067_));
  INV_X1     g06065(.I(new_n7052_), .ZN(new_n7068_));
  OAI21_X1   g06066(.A1(new_n7067_), .A2(new_n7023_), .B(new_n7068_), .ZN(new_n7069_));
  AOI22_X1   g06067(.A1(new_n7025_), .A2(new_n7028_), .B1(new_n7045_), .B2(new_n7042_), .ZN(new_n7070_));
  NAND3_X1   g06068(.A1(new_n7070_), .A2(new_n7066_), .A3(new_n7069_), .ZN(new_n7071_));
  NAND2_X1   g06069(.A1(new_n7063_), .A2(new_n7071_), .ZN(new_n7072_));
  NAND3_X1   g06070(.A1(new_n7072_), .A2(new_n7010_), .A3(new_n7018_), .ZN(new_n7073_));
  INV_X1     g06071(.I(\A[111] ), .ZN(new_n7074_));
  INV_X1     g06072(.I(\A[109] ), .ZN(new_n7075_));
  NAND2_X1   g06073(.A1(new_n7075_), .A2(\A[110] ), .ZN(new_n7076_));
  INV_X1     g06074(.I(\A[110] ), .ZN(new_n7077_));
  AOI21_X1   g06075(.A1(\A[109] ), .A2(new_n7077_), .B(new_n7074_), .ZN(new_n7078_));
  XOR2_X1    g06076(.A1(\A[109] ), .A2(\A[110] ), .Z(new_n7079_));
  AOI22_X1   g06077(.A1(new_n7079_), .A2(new_n7074_), .B1(new_n7076_), .B2(new_n7078_), .ZN(new_n7080_));
  INV_X1     g06078(.I(\A[112] ), .ZN(new_n7081_));
  NAND2_X1   g06079(.A1(new_n7081_), .A2(\A[113] ), .ZN(new_n7082_));
  INV_X1     g06080(.I(\A[113] ), .ZN(new_n7083_));
  NAND2_X1   g06081(.A1(new_n7083_), .A2(\A[112] ), .ZN(new_n7084_));
  NAND3_X1   g06082(.A1(new_n7082_), .A2(new_n7084_), .A3(\A[114] ), .ZN(new_n7085_));
  INV_X1     g06083(.I(\A[114] ), .ZN(new_n7086_));
  NOR2_X1    g06084(.A1(new_n7083_), .A2(\A[112] ), .ZN(new_n7087_));
  NOR2_X1    g06085(.A1(new_n7081_), .A2(\A[113] ), .ZN(new_n7088_));
  OAI21_X1   g06086(.A1(new_n7087_), .A2(new_n7088_), .B(new_n7086_), .ZN(new_n7089_));
  NAND2_X1   g06087(.A1(new_n7089_), .A2(new_n7085_), .ZN(new_n7090_));
  NAND2_X1   g06088(.A1(new_n7090_), .A2(new_n7080_), .ZN(new_n7091_));
  NAND2_X1   g06089(.A1(new_n7078_), .A2(new_n7076_), .ZN(new_n7092_));
  NOR2_X1    g06090(.A1(new_n7077_), .A2(\A[109] ), .ZN(new_n7093_));
  NOR2_X1    g06091(.A1(new_n7075_), .A2(\A[110] ), .ZN(new_n7094_));
  OAI21_X1   g06092(.A1(new_n7093_), .A2(new_n7094_), .B(new_n7074_), .ZN(new_n7095_));
  NAND2_X1   g06093(.A1(new_n7092_), .A2(new_n7095_), .ZN(new_n7096_));
  OAI21_X1   g06094(.A1(new_n7081_), .A2(\A[113] ), .B(\A[114] ), .ZN(new_n7097_));
  NOR2_X1    g06095(.A1(new_n7097_), .A2(new_n7087_), .ZN(new_n7098_));
  AOI21_X1   g06096(.A1(new_n7082_), .A2(new_n7084_), .B(\A[114] ), .ZN(new_n7099_));
  NOR2_X1    g06097(.A1(new_n7099_), .A2(new_n7098_), .ZN(new_n7100_));
  NAND2_X1   g06098(.A1(new_n7096_), .A2(new_n7100_), .ZN(new_n7101_));
  NAND2_X1   g06099(.A1(new_n7101_), .A2(new_n7091_), .ZN(new_n7102_));
  NOR2_X1    g06100(.A1(new_n7087_), .A2(new_n7088_), .ZN(new_n7103_));
  NOR2_X1    g06101(.A1(new_n7081_), .A2(new_n7083_), .ZN(new_n7104_));
  INV_X1     g06102(.I(new_n7104_), .ZN(new_n7105_));
  OAI21_X1   g06103(.A1(new_n7103_), .A2(new_n7086_), .B(new_n7105_), .ZN(new_n7106_));
  NOR2_X1    g06104(.A1(new_n7093_), .A2(new_n7094_), .ZN(new_n7107_));
  NOR2_X1    g06105(.A1(new_n7075_), .A2(new_n7077_), .ZN(new_n7108_));
  INV_X1     g06106(.I(new_n7108_), .ZN(new_n7109_));
  OAI21_X1   g06107(.A1(new_n7107_), .A2(new_n7074_), .B(new_n7109_), .ZN(new_n7110_));
  AOI22_X1   g06108(.A1(new_n7092_), .A2(new_n7095_), .B1(new_n7089_), .B2(new_n7085_), .ZN(new_n7111_));
  NAND3_X1   g06109(.A1(new_n7111_), .A2(new_n7106_), .A3(new_n7110_), .ZN(new_n7112_));
  NAND2_X1   g06110(.A1(new_n7102_), .A2(new_n7112_), .ZN(new_n7113_));
  INV_X1     g06111(.I(\A[103] ), .ZN(new_n7114_));
  NAND2_X1   g06112(.A1(new_n7114_), .A2(\A[104] ), .ZN(new_n7115_));
  INV_X1     g06113(.I(\A[104] ), .ZN(new_n7116_));
  INV_X1     g06114(.I(\A[105] ), .ZN(new_n7117_));
  AOI21_X1   g06115(.A1(\A[103] ), .A2(new_n7116_), .B(new_n7117_), .ZN(new_n7118_));
  NAND2_X1   g06116(.A1(new_n7118_), .A2(new_n7115_), .ZN(new_n7119_));
  NOR2_X1    g06117(.A1(new_n7116_), .A2(\A[103] ), .ZN(new_n7120_));
  NOR2_X1    g06118(.A1(new_n7114_), .A2(\A[104] ), .ZN(new_n7121_));
  OAI21_X1   g06119(.A1(new_n7120_), .A2(new_n7121_), .B(new_n7117_), .ZN(new_n7122_));
  NAND2_X1   g06120(.A1(new_n7119_), .A2(new_n7122_), .ZN(new_n7123_));
  INV_X1     g06121(.I(\A[108] ), .ZN(new_n7124_));
  INV_X1     g06122(.I(\A[107] ), .ZN(new_n7125_));
  NOR2_X1    g06123(.A1(new_n7125_), .A2(\A[106] ), .ZN(new_n7126_));
  INV_X1     g06124(.I(\A[106] ), .ZN(new_n7127_));
  NOR2_X1    g06125(.A1(new_n7127_), .A2(\A[107] ), .ZN(new_n7128_));
  NOR3_X1    g06126(.A1(new_n7126_), .A2(new_n7128_), .A3(new_n7124_), .ZN(new_n7129_));
  NAND2_X1   g06127(.A1(new_n7127_), .A2(\A[107] ), .ZN(new_n7130_));
  NAND2_X1   g06128(.A1(new_n7125_), .A2(\A[106] ), .ZN(new_n7131_));
  AOI21_X1   g06129(.A1(new_n7130_), .A2(new_n7131_), .B(\A[108] ), .ZN(new_n7132_));
  NOR2_X1    g06130(.A1(new_n7132_), .A2(new_n7129_), .ZN(new_n7133_));
  NOR2_X1    g06131(.A1(new_n7133_), .A2(new_n7123_), .ZN(new_n7134_));
  NOR3_X1    g06132(.A1(new_n7120_), .A2(new_n7121_), .A3(new_n7117_), .ZN(new_n7135_));
  NAND2_X1   g06133(.A1(new_n7116_), .A2(\A[103] ), .ZN(new_n7136_));
  AOI21_X1   g06134(.A1(new_n7115_), .A2(new_n7136_), .B(\A[105] ), .ZN(new_n7137_));
  NOR2_X1    g06135(.A1(new_n7137_), .A2(new_n7135_), .ZN(new_n7138_));
  AOI21_X1   g06136(.A1(\A[106] ), .A2(new_n7125_), .B(new_n7124_), .ZN(new_n7139_));
  NAND2_X1   g06137(.A1(new_n7139_), .A2(new_n7130_), .ZN(new_n7140_));
  XOR2_X1    g06138(.A1(\A[106] ), .A2(\A[107] ), .Z(new_n7141_));
  NAND2_X1   g06139(.A1(new_n7141_), .A2(new_n7124_), .ZN(new_n7142_));
  NAND2_X1   g06140(.A1(new_n7142_), .A2(new_n7140_), .ZN(new_n7143_));
  NOR2_X1    g06141(.A1(new_n7143_), .A2(new_n7138_), .ZN(new_n7144_));
  NOR2_X1    g06142(.A1(new_n7144_), .A2(new_n7134_), .ZN(new_n7145_));
  NOR2_X1    g06143(.A1(new_n7127_), .A2(new_n7125_), .ZN(new_n7146_));
  AOI21_X1   g06144(.A1(new_n7141_), .A2(\A[108] ), .B(new_n7146_), .ZN(new_n7147_));
  NAND2_X1   g06145(.A1(new_n7115_), .A2(new_n7136_), .ZN(new_n7148_));
  NAND2_X1   g06146(.A1(\A[103] ), .A2(\A[104] ), .ZN(new_n7149_));
  INV_X1     g06147(.I(new_n7149_), .ZN(new_n7150_));
  AOI21_X1   g06148(.A1(new_n7148_), .A2(\A[105] ), .B(new_n7150_), .ZN(new_n7151_));
  OAI22_X1   g06149(.A1(new_n7135_), .A2(new_n7137_), .B1(new_n7132_), .B2(new_n7129_), .ZN(new_n7152_));
  NOR3_X1    g06150(.A1(new_n7152_), .A2(new_n7147_), .A3(new_n7151_), .ZN(new_n7153_));
  NOR2_X1    g06151(.A1(new_n7145_), .A2(new_n7153_), .ZN(new_n7154_));
  NAND2_X1   g06152(.A1(new_n7154_), .A2(new_n7113_), .ZN(new_n7155_));
  NAND2_X1   g06153(.A1(new_n7143_), .A2(new_n7138_), .ZN(new_n7156_));
  NAND2_X1   g06154(.A1(new_n7133_), .A2(new_n7123_), .ZN(new_n7157_));
  NAND2_X1   g06155(.A1(new_n7156_), .A2(new_n7157_), .ZN(new_n7158_));
  NOR2_X1    g06156(.A1(new_n7126_), .A2(new_n7128_), .ZN(new_n7159_));
  INV_X1     g06157(.I(new_n7146_), .ZN(new_n7160_));
  OAI21_X1   g06158(.A1(new_n7159_), .A2(new_n7124_), .B(new_n7160_), .ZN(new_n7161_));
  NOR2_X1    g06159(.A1(new_n7120_), .A2(new_n7121_), .ZN(new_n7162_));
  OAI21_X1   g06160(.A1(new_n7162_), .A2(new_n7117_), .B(new_n7149_), .ZN(new_n7163_));
  AOI22_X1   g06161(.A1(new_n7142_), .A2(new_n7140_), .B1(new_n7119_), .B2(new_n7122_), .ZN(new_n7164_));
  NAND3_X1   g06162(.A1(new_n7164_), .A2(new_n7161_), .A3(new_n7163_), .ZN(new_n7165_));
  NAND2_X1   g06163(.A1(new_n7158_), .A2(new_n7165_), .ZN(new_n7166_));
  NAND3_X1   g06164(.A1(new_n7166_), .A2(new_n7102_), .A3(new_n7112_), .ZN(new_n7167_));
  NAND2_X1   g06165(.A1(new_n7167_), .A2(new_n7155_), .ZN(new_n7168_));
  NAND3_X1   g06166(.A1(new_n7168_), .A2(new_n7060_), .A3(new_n7073_), .ZN(new_n7169_));
  NAND2_X1   g06167(.A1(new_n7060_), .A2(new_n7073_), .ZN(new_n7170_));
  NAND3_X1   g06168(.A1(new_n7170_), .A2(new_n7155_), .A3(new_n7167_), .ZN(new_n7171_));
  NAND2_X1   g06169(.A1(new_n7169_), .A2(new_n7171_), .ZN(new_n7172_));
  INV_X1     g06170(.I(\A[99] ), .ZN(new_n7173_));
  INV_X1     g06171(.I(\A[98] ), .ZN(new_n7174_));
  NOR2_X1    g06172(.A1(new_n7174_), .A2(\A[97] ), .ZN(new_n7175_));
  INV_X1     g06173(.I(\A[97] ), .ZN(new_n7176_));
  NOR2_X1    g06174(.A1(new_n7176_), .A2(\A[98] ), .ZN(new_n7177_));
  NOR3_X1    g06175(.A1(new_n7175_), .A2(new_n7177_), .A3(new_n7173_), .ZN(new_n7178_));
  NAND2_X1   g06176(.A1(new_n7176_), .A2(\A[98] ), .ZN(new_n7179_));
  NAND2_X1   g06177(.A1(new_n7174_), .A2(\A[97] ), .ZN(new_n7180_));
  AOI21_X1   g06178(.A1(new_n7179_), .A2(new_n7180_), .B(\A[99] ), .ZN(new_n7181_));
  NOR2_X1    g06179(.A1(new_n7181_), .A2(new_n7178_), .ZN(new_n7182_));
  INV_X1     g06180(.I(\A[100] ), .ZN(new_n7183_));
  NAND2_X1   g06181(.A1(new_n7183_), .A2(\A[101] ), .ZN(new_n7184_));
  INV_X1     g06182(.I(\A[101] ), .ZN(new_n7185_));
  NAND2_X1   g06183(.A1(new_n7185_), .A2(\A[100] ), .ZN(new_n7186_));
  NAND3_X1   g06184(.A1(new_n7184_), .A2(new_n7186_), .A3(\A[102] ), .ZN(new_n7187_));
  INV_X1     g06185(.I(\A[102] ), .ZN(new_n7188_));
  NOR2_X1    g06186(.A1(new_n7185_), .A2(\A[100] ), .ZN(new_n7189_));
  NOR2_X1    g06187(.A1(new_n7183_), .A2(\A[101] ), .ZN(new_n7190_));
  OAI21_X1   g06188(.A1(new_n7189_), .A2(new_n7190_), .B(new_n7188_), .ZN(new_n7191_));
  NAND2_X1   g06189(.A1(new_n7191_), .A2(new_n7187_), .ZN(new_n7192_));
  NAND2_X1   g06190(.A1(new_n7182_), .A2(new_n7192_), .ZN(new_n7193_));
  NAND3_X1   g06191(.A1(new_n7179_), .A2(new_n7180_), .A3(\A[99] ), .ZN(new_n7194_));
  OAI21_X1   g06192(.A1(new_n7175_), .A2(new_n7177_), .B(new_n7173_), .ZN(new_n7195_));
  NAND2_X1   g06193(.A1(new_n7195_), .A2(new_n7194_), .ZN(new_n7196_));
  AOI21_X1   g06194(.A1(\A[100] ), .A2(new_n7185_), .B(new_n7188_), .ZN(new_n7197_));
  XOR2_X1    g06195(.A1(\A[100] ), .A2(\A[101] ), .Z(new_n7198_));
  AOI22_X1   g06196(.A1(new_n7198_), .A2(new_n7188_), .B1(new_n7184_), .B2(new_n7197_), .ZN(new_n7199_));
  NAND2_X1   g06197(.A1(new_n7196_), .A2(new_n7199_), .ZN(new_n7200_));
  NAND2_X1   g06198(.A1(new_n7193_), .A2(new_n7200_), .ZN(new_n7201_));
  NOR2_X1    g06199(.A1(new_n7189_), .A2(new_n7190_), .ZN(new_n7202_));
  NOR2_X1    g06200(.A1(new_n7183_), .A2(new_n7185_), .ZN(new_n7203_));
  INV_X1     g06201(.I(new_n7203_), .ZN(new_n7204_));
  OAI21_X1   g06202(.A1(new_n7202_), .A2(new_n7188_), .B(new_n7204_), .ZN(new_n7205_));
  XNOR2_X1   g06203(.A1(\A[97] ), .A2(\A[98] ), .ZN(new_n7206_));
  NAND2_X1   g06204(.A1(\A[97] ), .A2(\A[98] ), .ZN(new_n7207_));
  OAI21_X1   g06205(.A1(new_n7206_), .A2(new_n7173_), .B(new_n7207_), .ZN(new_n7208_));
  AOI22_X1   g06206(.A1(new_n7194_), .A2(new_n7195_), .B1(new_n7191_), .B2(new_n7187_), .ZN(new_n7209_));
  NAND3_X1   g06207(.A1(new_n7209_), .A2(new_n7205_), .A3(new_n7208_), .ZN(new_n7210_));
  NAND2_X1   g06208(.A1(new_n7201_), .A2(new_n7210_), .ZN(new_n7211_));
  INV_X1     g06209(.I(\A[91] ), .ZN(new_n7212_));
  NAND2_X1   g06210(.A1(new_n7212_), .A2(\A[92] ), .ZN(new_n7213_));
  INV_X1     g06211(.I(\A[92] ), .ZN(new_n7214_));
  INV_X1     g06212(.I(\A[93] ), .ZN(new_n7215_));
  AOI21_X1   g06213(.A1(\A[91] ), .A2(new_n7214_), .B(new_n7215_), .ZN(new_n7216_));
  NAND2_X1   g06214(.A1(new_n7216_), .A2(new_n7213_), .ZN(new_n7217_));
  NOR2_X1    g06215(.A1(new_n7214_), .A2(\A[91] ), .ZN(new_n7218_));
  NOR2_X1    g06216(.A1(new_n7212_), .A2(\A[92] ), .ZN(new_n7219_));
  OAI21_X1   g06217(.A1(new_n7218_), .A2(new_n7219_), .B(new_n7215_), .ZN(new_n7220_));
  NAND2_X1   g06218(.A1(new_n7217_), .A2(new_n7220_), .ZN(new_n7221_));
  INV_X1     g06219(.I(\A[96] ), .ZN(new_n7222_));
  INV_X1     g06220(.I(\A[94] ), .ZN(new_n7223_));
  NAND2_X1   g06221(.A1(new_n7223_), .A2(\A[95] ), .ZN(new_n7224_));
  INV_X1     g06222(.I(\A[95] ), .ZN(new_n7225_));
  AOI21_X1   g06223(.A1(\A[94] ), .A2(new_n7225_), .B(new_n7222_), .ZN(new_n7226_));
  XOR2_X1    g06224(.A1(\A[94] ), .A2(\A[95] ), .Z(new_n7227_));
  AOI22_X1   g06225(.A1(new_n7227_), .A2(new_n7222_), .B1(new_n7224_), .B2(new_n7226_), .ZN(new_n7228_));
  NOR2_X1    g06226(.A1(new_n7221_), .A2(new_n7228_), .ZN(new_n7229_));
  XOR2_X1    g06227(.A1(\A[91] ), .A2(\A[92] ), .Z(new_n7230_));
  AOI22_X1   g06228(.A1(new_n7230_), .A2(new_n7215_), .B1(new_n7213_), .B2(new_n7216_), .ZN(new_n7231_));
  NAND2_X1   g06229(.A1(new_n7225_), .A2(\A[94] ), .ZN(new_n7232_));
  NAND3_X1   g06230(.A1(new_n7224_), .A2(new_n7232_), .A3(\A[96] ), .ZN(new_n7233_));
  NOR2_X1    g06231(.A1(new_n7225_), .A2(\A[94] ), .ZN(new_n7234_));
  NOR2_X1    g06232(.A1(new_n7223_), .A2(\A[95] ), .ZN(new_n7235_));
  OAI21_X1   g06233(.A1(new_n7234_), .A2(new_n7235_), .B(new_n7222_), .ZN(new_n7236_));
  NAND2_X1   g06234(.A1(new_n7236_), .A2(new_n7233_), .ZN(new_n7237_));
  NOR2_X1    g06235(.A1(new_n7237_), .A2(new_n7231_), .ZN(new_n7238_));
  NOR2_X1    g06236(.A1(new_n7229_), .A2(new_n7238_), .ZN(new_n7239_));
  NAND2_X1   g06237(.A1(\A[94] ), .A2(\A[95] ), .ZN(new_n7240_));
  INV_X1     g06238(.I(new_n7240_), .ZN(new_n7241_));
  AOI21_X1   g06239(.A1(new_n7227_), .A2(\A[96] ), .B(new_n7241_), .ZN(new_n7242_));
  NAND2_X1   g06240(.A1(\A[91] ), .A2(\A[92] ), .ZN(new_n7243_));
  INV_X1     g06241(.I(new_n7243_), .ZN(new_n7244_));
  AOI21_X1   g06242(.A1(new_n7230_), .A2(\A[93] ), .B(new_n7244_), .ZN(new_n7245_));
  NOR3_X1    g06243(.A1(new_n7218_), .A2(new_n7219_), .A3(new_n7215_), .ZN(new_n7246_));
  NAND2_X1   g06244(.A1(new_n7214_), .A2(\A[91] ), .ZN(new_n7247_));
  AOI21_X1   g06245(.A1(new_n7213_), .A2(new_n7247_), .B(\A[93] ), .ZN(new_n7248_));
  NOR3_X1    g06246(.A1(new_n7234_), .A2(new_n7235_), .A3(new_n7222_), .ZN(new_n7249_));
  AOI21_X1   g06247(.A1(new_n7224_), .A2(new_n7232_), .B(\A[96] ), .ZN(new_n7250_));
  OAI22_X1   g06248(.A1(new_n7246_), .A2(new_n7248_), .B1(new_n7250_), .B2(new_n7249_), .ZN(new_n7251_));
  NOR3_X1    g06249(.A1(new_n7251_), .A2(new_n7242_), .A3(new_n7245_), .ZN(new_n7252_));
  NOR2_X1    g06250(.A1(new_n7239_), .A2(new_n7252_), .ZN(new_n7253_));
  NAND2_X1   g06251(.A1(new_n7253_), .A2(new_n7211_), .ZN(new_n7254_));
  NOR2_X1    g06252(.A1(new_n7196_), .A2(new_n7199_), .ZN(new_n7255_));
  NOR2_X1    g06253(.A1(new_n7182_), .A2(new_n7192_), .ZN(new_n7256_));
  NOR2_X1    g06254(.A1(new_n7256_), .A2(new_n7255_), .ZN(new_n7257_));
  AOI21_X1   g06255(.A1(new_n7198_), .A2(\A[102] ), .B(new_n7203_), .ZN(new_n7258_));
  XOR2_X1    g06256(.A1(\A[97] ), .A2(\A[98] ), .Z(new_n7259_));
  INV_X1     g06257(.I(new_n7207_), .ZN(new_n7260_));
  AOI21_X1   g06258(.A1(new_n7259_), .A2(\A[99] ), .B(new_n7260_), .ZN(new_n7261_));
  NOR3_X1    g06259(.A1(new_n7189_), .A2(new_n7190_), .A3(new_n7188_), .ZN(new_n7262_));
  AOI21_X1   g06260(.A1(new_n7184_), .A2(new_n7186_), .B(\A[102] ), .ZN(new_n7263_));
  OAI22_X1   g06261(.A1(new_n7262_), .A2(new_n7263_), .B1(new_n7181_), .B2(new_n7178_), .ZN(new_n7264_));
  NOR3_X1    g06262(.A1(new_n7264_), .A2(new_n7258_), .A3(new_n7261_), .ZN(new_n7265_));
  NOR2_X1    g06263(.A1(new_n7257_), .A2(new_n7265_), .ZN(new_n7266_));
  NAND2_X1   g06264(.A1(new_n7237_), .A2(new_n7231_), .ZN(new_n7267_));
  NAND2_X1   g06265(.A1(new_n7221_), .A2(new_n7228_), .ZN(new_n7268_));
  NAND2_X1   g06266(.A1(new_n7268_), .A2(new_n7267_), .ZN(new_n7269_));
  XNOR2_X1   g06267(.A1(\A[94] ), .A2(\A[95] ), .ZN(new_n7270_));
  OAI21_X1   g06268(.A1(new_n7270_), .A2(new_n7222_), .B(new_n7240_), .ZN(new_n7271_));
  XNOR2_X1   g06269(.A1(\A[91] ), .A2(\A[92] ), .ZN(new_n7272_));
  OAI21_X1   g06270(.A1(new_n7272_), .A2(new_n7215_), .B(new_n7243_), .ZN(new_n7273_));
  AOI22_X1   g06271(.A1(new_n7217_), .A2(new_n7220_), .B1(new_n7236_), .B2(new_n7233_), .ZN(new_n7274_));
  NAND3_X1   g06272(.A1(new_n7274_), .A2(new_n7271_), .A3(new_n7273_), .ZN(new_n7275_));
  NAND2_X1   g06273(.A1(new_n7269_), .A2(new_n7275_), .ZN(new_n7276_));
  NAND2_X1   g06274(.A1(new_n7266_), .A2(new_n7276_), .ZN(new_n7277_));
  INV_X1     g06275(.I(\A[87] ), .ZN(new_n7278_));
  INV_X1     g06276(.I(\A[86] ), .ZN(new_n7279_));
  NOR2_X1    g06277(.A1(new_n7279_), .A2(\A[85] ), .ZN(new_n7280_));
  INV_X1     g06278(.I(\A[85] ), .ZN(new_n7281_));
  NOR2_X1    g06279(.A1(new_n7281_), .A2(\A[86] ), .ZN(new_n7282_));
  NOR3_X1    g06280(.A1(new_n7280_), .A2(new_n7282_), .A3(new_n7278_), .ZN(new_n7283_));
  NAND2_X1   g06281(.A1(new_n7281_), .A2(\A[86] ), .ZN(new_n7284_));
  NAND2_X1   g06282(.A1(new_n7279_), .A2(\A[85] ), .ZN(new_n7285_));
  AOI21_X1   g06283(.A1(new_n7284_), .A2(new_n7285_), .B(\A[87] ), .ZN(new_n7286_));
  NOR2_X1    g06284(.A1(new_n7286_), .A2(new_n7283_), .ZN(new_n7287_));
  INV_X1     g06285(.I(\A[88] ), .ZN(new_n7288_));
  NAND2_X1   g06286(.A1(new_n7288_), .A2(\A[89] ), .ZN(new_n7289_));
  INV_X1     g06287(.I(\A[89] ), .ZN(new_n7290_));
  NAND2_X1   g06288(.A1(new_n7290_), .A2(\A[88] ), .ZN(new_n7291_));
  NAND3_X1   g06289(.A1(new_n7289_), .A2(new_n7291_), .A3(\A[90] ), .ZN(new_n7292_));
  INV_X1     g06290(.I(\A[90] ), .ZN(new_n7293_));
  NOR2_X1    g06291(.A1(new_n7290_), .A2(\A[88] ), .ZN(new_n7294_));
  NOR2_X1    g06292(.A1(new_n7288_), .A2(\A[89] ), .ZN(new_n7295_));
  OAI21_X1   g06293(.A1(new_n7294_), .A2(new_n7295_), .B(new_n7293_), .ZN(new_n7296_));
  NAND2_X1   g06294(.A1(new_n7296_), .A2(new_n7292_), .ZN(new_n7297_));
  NAND2_X1   g06295(.A1(new_n7287_), .A2(new_n7297_), .ZN(new_n7298_));
  NAND3_X1   g06296(.A1(new_n7284_), .A2(new_n7285_), .A3(\A[87] ), .ZN(new_n7299_));
  OAI21_X1   g06297(.A1(new_n7280_), .A2(new_n7282_), .B(new_n7278_), .ZN(new_n7300_));
  NAND2_X1   g06298(.A1(new_n7300_), .A2(new_n7299_), .ZN(new_n7301_));
  NOR3_X1    g06299(.A1(new_n7294_), .A2(new_n7295_), .A3(new_n7293_), .ZN(new_n7302_));
  AOI21_X1   g06300(.A1(new_n7289_), .A2(new_n7291_), .B(\A[90] ), .ZN(new_n7303_));
  NOR2_X1    g06301(.A1(new_n7303_), .A2(new_n7302_), .ZN(new_n7304_));
  NAND2_X1   g06302(.A1(new_n7304_), .A2(new_n7301_), .ZN(new_n7305_));
  NAND2_X1   g06303(.A1(new_n7298_), .A2(new_n7305_), .ZN(new_n7306_));
  NOR2_X1    g06304(.A1(new_n7294_), .A2(new_n7295_), .ZN(new_n7307_));
  NOR2_X1    g06305(.A1(new_n7288_), .A2(new_n7290_), .ZN(new_n7308_));
  INV_X1     g06306(.I(new_n7308_), .ZN(new_n7309_));
  OAI21_X1   g06307(.A1(new_n7307_), .A2(new_n7293_), .B(new_n7309_), .ZN(new_n7310_));
  NOR2_X1    g06308(.A1(new_n7280_), .A2(new_n7282_), .ZN(new_n7311_));
  NOR2_X1    g06309(.A1(new_n7281_), .A2(new_n7279_), .ZN(new_n7312_));
  INV_X1     g06310(.I(new_n7312_), .ZN(new_n7313_));
  OAI21_X1   g06311(.A1(new_n7311_), .A2(new_n7278_), .B(new_n7313_), .ZN(new_n7314_));
  AOI22_X1   g06312(.A1(new_n7292_), .A2(new_n7296_), .B1(new_n7300_), .B2(new_n7299_), .ZN(new_n7315_));
  NAND3_X1   g06313(.A1(new_n7315_), .A2(new_n7310_), .A3(new_n7314_), .ZN(new_n7316_));
  NAND2_X1   g06314(.A1(new_n7306_), .A2(new_n7316_), .ZN(new_n7317_));
  INV_X1     g06315(.I(\A[79] ), .ZN(new_n7318_));
  NAND2_X1   g06316(.A1(new_n7318_), .A2(\A[80] ), .ZN(new_n7319_));
  INV_X1     g06317(.I(\A[80] ), .ZN(new_n7320_));
  NAND2_X1   g06318(.A1(new_n7320_), .A2(\A[79] ), .ZN(new_n7321_));
  NAND3_X1   g06319(.A1(new_n7319_), .A2(new_n7321_), .A3(\A[81] ), .ZN(new_n7322_));
  INV_X1     g06320(.I(\A[81] ), .ZN(new_n7323_));
  NOR2_X1    g06321(.A1(new_n7320_), .A2(\A[79] ), .ZN(new_n7324_));
  NOR2_X1    g06322(.A1(new_n7318_), .A2(\A[80] ), .ZN(new_n7325_));
  OAI21_X1   g06323(.A1(new_n7324_), .A2(new_n7325_), .B(new_n7323_), .ZN(new_n7326_));
  NAND2_X1   g06324(.A1(new_n7326_), .A2(new_n7322_), .ZN(new_n7327_));
  INV_X1     g06325(.I(\A[84] ), .ZN(new_n7328_));
  INV_X1     g06326(.I(\A[83] ), .ZN(new_n7329_));
  NOR2_X1    g06327(.A1(new_n7329_), .A2(\A[82] ), .ZN(new_n7330_));
  INV_X1     g06328(.I(\A[82] ), .ZN(new_n7331_));
  NOR2_X1    g06329(.A1(new_n7331_), .A2(\A[83] ), .ZN(new_n7332_));
  NOR3_X1    g06330(.A1(new_n7330_), .A2(new_n7332_), .A3(new_n7328_), .ZN(new_n7333_));
  NAND2_X1   g06331(.A1(new_n7331_), .A2(\A[83] ), .ZN(new_n7334_));
  NAND2_X1   g06332(.A1(new_n7329_), .A2(\A[82] ), .ZN(new_n7335_));
  AOI21_X1   g06333(.A1(new_n7334_), .A2(new_n7335_), .B(\A[84] ), .ZN(new_n7336_));
  NOR2_X1    g06334(.A1(new_n7336_), .A2(new_n7333_), .ZN(new_n7337_));
  NOR2_X1    g06335(.A1(new_n7337_), .A2(new_n7327_), .ZN(new_n7338_));
  OAI21_X1   g06336(.A1(new_n7318_), .A2(\A[80] ), .B(\A[81] ), .ZN(new_n7339_));
  NOR2_X1    g06337(.A1(new_n7339_), .A2(new_n7324_), .ZN(new_n7340_));
  AOI21_X1   g06338(.A1(new_n7319_), .A2(new_n7321_), .B(\A[81] ), .ZN(new_n7341_));
  NOR2_X1    g06339(.A1(new_n7341_), .A2(new_n7340_), .ZN(new_n7342_));
  NAND3_X1   g06340(.A1(new_n7334_), .A2(new_n7335_), .A3(\A[84] ), .ZN(new_n7343_));
  OAI21_X1   g06341(.A1(new_n7330_), .A2(new_n7332_), .B(new_n7328_), .ZN(new_n7344_));
  NAND2_X1   g06342(.A1(new_n7344_), .A2(new_n7343_), .ZN(new_n7345_));
  NOR2_X1    g06343(.A1(new_n7345_), .A2(new_n7342_), .ZN(new_n7346_));
  NOR2_X1    g06344(.A1(new_n7338_), .A2(new_n7346_), .ZN(new_n7347_));
  XOR2_X1    g06345(.A1(\A[82] ), .A2(\A[83] ), .Z(new_n7348_));
  NOR2_X1    g06346(.A1(new_n7331_), .A2(new_n7329_), .ZN(new_n7349_));
  AOI21_X1   g06347(.A1(new_n7348_), .A2(\A[84] ), .B(new_n7349_), .ZN(new_n7350_));
  XOR2_X1    g06348(.A1(\A[79] ), .A2(\A[80] ), .Z(new_n7351_));
  NAND2_X1   g06349(.A1(\A[79] ), .A2(\A[80] ), .ZN(new_n7352_));
  INV_X1     g06350(.I(new_n7352_), .ZN(new_n7353_));
  AOI21_X1   g06351(.A1(new_n7351_), .A2(\A[81] ), .B(new_n7353_), .ZN(new_n7354_));
  OAI22_X1   g06352(.A1(new_n7333_), .A2(new_n7336_), .B1(new_n7341_), .B2(new_n7340_), .ZN(new_n7355_));
  NOR3_X1    g06353(.A1(new_n7355_), .A2(new_n7350_), .A3(new_n7354_), .ZN(new_n7356_));
  NOR2_X1    g06354(.A1(new_n7347_), .A2(new_n7356_), .ZN(new_n7357_));
  NAND2_X1   g06355(.A1(new_n7357_), .A2(new_n7317_), .ZN(new_n7358_));
  NOR2_X1    g06356(.A1(new_n7304_), .A2(new_n7301_), .ZN(new_n7359_));
  NOR2_X1    g06357(.A1(new_n7287_), .A2(new_n7297_), .ZN(new_n7360_));
  NOR2_X1    g06358(.A1(new_n7360_), .A2(new_n7359_), .ZN(new_n7361_));
  INV_X1     g06359(.I(new_n7316_), .ZN(new_n7362_));
  NOR2_X1    g06360(.A1(new_n7362_), .A2(new_n7361_), .ZN(new_n7363_));
  NAND2_X1   g06361(.A1(new_n7345_), .A2(new_n7342_), .ZN(new_n7364_));
  NAND2_X1   g06362(.A1(new_n7337_), .A2(new_n7327_), .ZN(new_n7365_));
  NAND2_X1   g06363(.A1(new_n7365_), .A2(new_n7364_), .ZN(new_n7366_));
  NOR2_X1    g06364(.A1(new_n7330_), .A2(new_n7332_), .ZN(new_n7367_));
  INV_X1     g06365(.I(new_n7349_), .ZN(new_n7368_));
  OAI21_X1   g06366(.A1(new_n7367_), .A2(new_n7328_), .B(new_n7368_), .ZN(new_n7369_));
  XNOR2_X1   g06367(.A1(\A[79] ), .A2(\A[80] ), .ZN(new_n7370_));
  OAI21_X1   g06368(.A1(new_n7370_), .A2(new_n7323_), .B(new_n7352_), .ZN(new_n7371_));
  AOI22_X1   g06369(.A1(new_n7343_), .A2(new_n7344_), .B1(new_n7326_), .B2(new_n7322_), .ZN(new_n7372_));
  NAND3_X1   g06370(.A1(new_n7372_), .A2(new_n7369_), .A3(new_n7371_), .ZN(new_n7373_));
  NAND2_X1   g06371(.A1(new_n7366_), .A2(new_n7373_), .ZN(new_n7374_));
  NAND2_X1   g06372(.A1(new_n7363_), .A2(new_n7374_), .ZN(new_n7375_));
  NAND2_X1   g06373(.A1(new_n7375_), .A2(new_n7358_), .ZN(new_n7376_));
  NAND3_X1   g06374(.A1(new_n7376_), .A2(new_n7254_), .A3(new_n7277_), .ZN(new_n7377_));
  NAND2_X1   g06375(.A1(new_n7254_), .A2(new_n7277_), .ZN(new_n7378_));
  NAND3_X1   g06376(.A1(new_n7378_), .A2(new_n7358_), .A3(new_n7375_), .ZN(new_n7379_));
  NAND2_X1   g06377(.A1(new_n7377_), .A2(new_n7379_), .ZN(new_n7380_));
  XOR2_X1    g06378(.A1(new_n7380_), .A2(new_n7172_), .Z(new_n7381_));
  XNOR2_X1   g06379(.A1(new_n6983_), .A2(new_n7381_), .ZN(new_n7382_));
  XNOR2_X1   g06380(.A1(new_n6571_), .A2(new_n7382_), .ZN(new_n7383_));
  NOR2_X1    g06381(.A1(new_n7383_), .A2(new_n5752_), .ZN(new_n7384_));
  XOR2_X1    g06382(.A1(\A[274] ), .A2(\A[275] ), .Z(new_n7385_));
  AOI21_X1   g06383(.A1(new_n7385_), .A2(\A[276] ), .B(new_n5729_), .ZN(new_n7386_));
  NOR2_X1    g06384(.A1(new_n5735_), .A2(new_n7386_), .ZN(new_n7387_));
  XOR2_X1    g06385(.A1(\A[271] ), .A2(\A[272] ), .Z(new_n7388_));
  AOI21_X1   g06386(.A1(new_n7388_), .A2(\A[273] ), .B(new_n5733_), .ZN(new_n7389_));
  NOR2_X1    g06387(.A1(new_n5731_), .A2(new_n7389_), .ZN(new_n7390_));
  NOR2_X1    g06388(.A1(new_n7387_), .A2(new_n7390_), .ZN(new_n7391_));
  OAI22_X1   g06389(.A1(new_n5720_), .A2(new_n5722_), .B1(new_n5717_), .B2(new_n5714_), .ZN(new_n7392_));
  NOR2_X1    g06390(.A1(new_n7386_), .A2(new_n7389_), .ZN(new_n7393_));
  INV_X1     g06391(.I(new_n7393_), .ZN(new_n7394_));
  OAI21_X1   g06392(.A1(new_n7391_), .A2(new_n7392_), .B(new_n7394_), .ZN(new_n7395_));
  NAND2_X1   g06393(.A1(new_n5731_), .A2(new_n7389_), .ZN(new_n7396_));
  NAND2_X1   g06394(.A1(new_n5735_), .A2(new_n7386_), .ZN(new_n7397_));
  NAND4_X1   g06395(.A1(new_n7396_), .A2(new_n7397_), .A3(new_n5708_), .A4(new_n5726_), .ZN(new_n7398_));
  OAI21_X1   g06396(.A1(new_n7387_), .A2(new_n7390_), .B(new_n7392_), .ZN(new_n7399_));
  AOI22_X1   g06397(.A1(new_n7395_), .A2(new_n5742_), .B1(new_n7398_), .B2(new_n7399_), .ZN(new_n7400_));
  NAND2_X1   g06398(.A1(new_n5666_), .A2(new_n5662_), .ZN(new_n7401_));
  AOI21_X1   g06399(.A1(new_n7401_), .A2(\A[279] ), .B(new_n5695_), .ZN(new_n7402_));
  NAND2_X1   g06400(.A1(new_n5693_), .A2(new_n7402_), .ZN(new_n7403_));
  XOR2_X1    g06401(.A1(\A[280] ), .A2(\A[281] ), .Z(new_n7404_));
  AOI21_X1   g06402(.A1(new_n7404_), .A2(\A[282] ), .B(new_n5691_), .ZN(new_n7405_));
  NAND2_X1   g06403(.A1(new_n5697_), .A2(new_n7405_), .ZN(new_n7406_));
  NAND3_X1   g06404(.A1(new_n7403_), .A2(new_n7406_), .A3(new_n5698_), .ZN(new_n7407_));
  NOR2_X1    g06405(.A1(new_n5697_), .A2(new_n7405_), .ZN(new_n7408_));
  NOR2_X1    g06406(.A1(new_n5693_), .A2(new_n7402_), .ZN(new_n7409_));
  OAI22_X1   g06407(.A1(new_n5664_), .A2(new_n5667_), .B1(new_n5686_), .B2(new_n5685_), .ZN(new_n7410_));
  OAI21_X1   g06408(.A1(new_n7409_), .A2(new_n7408_), .B(new_n7410_), .ZN(new_n7411_));
  NAND2_X1   g06409(.A1(new_n7411_), .A2(new_n7407_), .ZN(new_n7412_));
  AOI22_X1   g06410(.A1(new_n5679_), .A2(new_n5688_), .B1(new_n5740_), .B2(new_n5741_), .ZN(new_n7413_));
  NAND3_X1   g06411(.A1(new_n7412_), .A2(new_n7413_), .A3(new_n5699_), .ZN(new_n7414_));
  XOR2_X1    g06412(.A1(new_n5687_), .A2(new_n5684_), .Z(new_n7415_));
  NAND2_X1   g06413(.A1(new_n7403_), .A2(new_n7406_), .ZN(new_n7416_));
  NOR2_X1    g06414(.A1(new_n7402_), .A2(new_n7405_), .ZN(new_n7417_));
  AOI21_X1   g06415(.A1(new_n7416_), .A2(new_n5698_), .B(new_n7417_), .ZN(new_n7418_));
  OAI21_X1   g06416(.A1(new_n7418_), .A2(new_n7415_), .B(new_n5736_), .ZN(new_n7419_));
  NOR2_X1    g06417(.A1(new_n7414_), .A2(new_n7419_), .ZN(new_n7420_));
  INV_X1     g06418(.I(new_n5699_), .ZN(new_n7421_));
  NOR4_X1    g06419(.A1(new_n7415_), .A2(new_n7421_), .A3(new_n5737_), .A4(new_n5728_), .ZN(new_n7422_));
  OAI21_X1   g06420(.A1(new_n7409_), .A2(new_n7408_), .B(new_n5698_), .ZN(new_n7423_));
  INV_X1     g06421(.I(new_n7417_), .ZN(new_n7424_));
  NAND2_X1   g06422(.A1(new_n7423_), .A2(new_n7424_), .ZN(new_n7425_));
  AOI22_X1   g06423(.A1(new_n7425_), .A2(new_n5689_), .B1(new_n7407_), .B2(new_n7411_), .ZN(new_n7426_));
  NOR2_X1    g06424(.A1(new_n7426_), .A2(new_n7422_), .ZN(new_n7427_));
  OAI21_X1   g06425(.A1(new_n7427_), .A2(new_n7420_), .B(new_n7400_), .ZN(new_n7428_));
  AOI21_X1   g06426(.A1(new_n7396_), .A2(new_n7397_), .B(new_n7392_), .ZN(new_n7429_));
  NOR2_X1    g06427(.A1(new_n7429_), .A2(new_n7393_), .ZN(new_n7430_));
  NOR3_X1    g06428(.A1(new_n7387_), .A2(new_n7390_), .A3(new_n7392_), .ZN(new_n7431_));
  AOI22_X1   g06429(.A1(new_n7396_), .A2(new_n7397_), .B1(new_n5708_), .B2(new_n5726_), .ZN(new_n7432_));
  OAI22_X1   g06430(.A1(new_n7430_), .A2(new_n5728_), .B1(new_n7431_), .B2(new_n7432_), .ZN(new_n7433_));
  NOR3_X1    g06431(.A1(new_n7409_), .A2(new_n7408_), .A3(new_n7410_), .ZN(new_n7434_));
  AOI21_X1   g06432(.A1(new_n7403_), .A2(new_n7406_), .B(new_n5698_), .ZN(new_n7435_));
  OAI22_X1   g06433(.A1(new_n7418_), .A2(new_n7415_), .B1(new_n7434_), .B2(new_n7435_), .ZN(new_n7436_));
  NOR2_X1    g06434(.A1(new_n7436_), .A2(new_n7422_), .ZN(new_n7437_));
  NAND3_X1   g06435(.A1(new_n7413_), .A2(new_n5699_), .A3(new_n5736_), .ZN(new_n7438_));
  NOR2_X1    g06436(.A1(new_n7426_), .A2(new_n7438_), .ZN(new_n7439_));
  OAI21_X1   g06437(.A1(new_n7439_), .A2(new_n7437_), .B(new_n7433_), .ZN(new_n7440_));
  NAND2_X1   g06438(.A1(new_n7440_), .A2(new_n7428_), .ZN(new_n7441_));
  NOR2_X1    g06439(.A1(new_n5655_), .A2(new_n5639_), .ZN(new_n7442_));
  NOR2_X1    g06440(.A1(new_n5653_), .A2(new_n5643_), .ZN(new_n7443_));
  OAI21_X1   g06441(.A1(new_n7443_), .A2(new_n7442_), .B(new_n5656_), .ZN(new_n7444_));
  NOR2_X1    g06442(.A1(new_n5639_), .A2(new_n5643_), .ZN(new_n7445_));
  INV_X1     g06443(.I(new_n7445_), .ZN(new_n7446_));
  NAND2_X1   g06444(.A1(new_n7444_), .A2(new_n7446_), .ZN(new_n7447_));
  NAND2_X1   g06445(.A1(new_n5653_), .A2(new_n5643_), .ZN(new_n7448_));
  NAND2_X1   g06446(.A1(new_n5655_), .A2(new_n5639_), .ZN(new_n7449_));
  NAND3_X1   g06447(.A1(new_n7448_), .A2(new_n7449_), .A3(new_n5656_), .ZN(new_n7450_));
  OAI21_X1   g06448(.A1(new_n7443_), .A2(new_n7442_), .B(new_n5644_), .ZN(new_n7451_));
  AOI22_X1   g06449(.A1(new_n7447_), .A2(new_n5650_), .B1(new_n7450_), .B2(new_n7451_), .ZN(new_n7452_));
  NAND2_X1   g06450(.A1(new_n5573_), .A2(new_n5574_), .ZN(new_n7453_));
  INV_X1     g06451(.I(new_n5602_), .ZN(new_n7454_));
  AOI21_X1   g06452(.A1(new_n7453_), .A2(\A[291] ), .B(new_n7454_), .ZN(new_n7455_));
  NAND2_X1   g06453(.A1(new_n5600_), .A2(new_n7455_), .ZN(new_n7456_));
  AOI21_X1   g06454(.A1(new_n5593_), .A2(\A[294] ), .B(new_n5598_), .ZN(new_n7457_));
  NAND2_X1   g06455(.A1(new_n5603_), .A2(new_n7457_), .ZN(new_n7458_));
  NAND3_X1   g06456(.A1(new_n7456_), .A2(new_n7458_), .A3(new_n5604_), .ZN(new_n7459_));
  NOR2_X1    g06457(.A1(new_n5603_), .A2(new_n7457_), .ZN(new_n7460_));
  NOR2_X1    g06458(.A1(new_n5600_), .A2(new_n7455_), .ZN(new_n7461_));
  NOR3_X1    g06459(.A1(new_n5583_), .A2(new_n5584_), .A3(new_n5580_), .ZN(new_n7462_));
  NAND2_X1   g06460(.A1(new_n5579_), .A2(\A[292] ), .ZN(new_n7463_));
  AOI21_X1   g06461(.A1(new_n5578_), .A2(new_n7463_), .B(\A[294] ), .ZN(new_n7464_));
  OAI22_X1   g06462(.A1(new_n7462_), .A2(new_n7464_), .B1(new_n5575_), .B2(new_n5572_), .ZN(new_n7465_));
  OAI21_X1   g06463(.A1(new_n7461_), .A2(new_n7460_), .B(new_n7465_), .ZN(new_n7466_));
  NAND2_X1   g06464(.A1(new_n7466_), .A2(new_n7459_), .ZN(new_n7467_));
  AOI22_X1   g06465(.A1(new_n5649_), .A2(new_n5648_), .B1(new_n5587_), .B2(new_n5595_), .ZN(new_n7468_));
  NAND3_X1   g06466(.A1(new_n7467_), .A2(new_n5605_), .A3(new_n7468_), .ZN(new_n7469_));
  NOR2_X1    g06467(.A1(new_n5592_), .A2(new_n5594_), .ZN(new_n7470_));
  NOR2_X1    g06468(.A1(new_n5586_), .A2(new_n5576_), .ZN(new_n7471_));
  NOR2_X1    g06469(.A1(new_n7471_), .A2(new_n7470_), .ZN(new_n7472_));
  AOI21_X1   g06470(.A1(new_n7456_), .A2(new_n7458_), .B(new_n7465_), .ZN(new_n7473_));
  NOR2_X1    g06471(.A1(new_n7455_), .A2(new_n7457_), .ZN(new_n7474_));
  NOR2_X1    g06472(.A1(new_n7473_), .A2(new_n7474_), .ZN(new_n7475_));
  OAI21_X1   g06473(.A1(new_n7475_), .A2(new_n7472_), .B(new_n5657_), .ZN(new_n7476_));
  NOR2_X1    g06474(.A1(new_n7469_), .A2(new_n7476_), .ZN(new_n7477_));
  NOR3_X1    g06475(.A1(new_n7465_), .A2(new_n7457_), .A3(new_n7455_), .ZN(new_n7478_));
  OAI22_X1   g06476(.A1(new_n5627_), .A2(new_n5635_), .B1(new_n7471_), .B2(new_n7470_), .ZN(new_n7479_));
  NOR3_X1    g06477(.A1(new_n7479_), .A2(new_n7478_), .A3(new_n5645_), .ZN(new_n7480_));
  NOR3_X1    g06478(.A1(new_n7461_), .A2(new_n7460_), .A3(new_n7465_), .ZN(new_n7481_));
  AOI21_X1   g06479(.A1(new_n7456_), .A2(new_n7458_), .B(new_n5604_), .ZN(new_n7482_));
  NOR2_X1    g06480(.A1(new_n7481_), .A2(new_n7482_), .ZN(new_n7483_));
  OAI21_X1   g06481(.A1(new_n7461_), .A2(new_n7460_), .B(new_n5604_), .ZN(new_n7484_));
  INV_X1     g06482(.I(new_n7474_), .ZN(new_n7485_));
  AOI21_X1   g06483(.A1(new_n7484_), .A2(new_n7485_), .B(new_n7472_), .ZN(new_n7486_));
  NOR2_X1    g06484(.A1(new_n7486_), .A2(new_n7483_), .ZN(new_n7487_));
  NOR2_X1    g06485(.A1(new_n7487_), .A2(new_n7480_), .ZN(new_n7488_));
  OAI21_X1   g06486(.A1(new_n7488_), .A2(new_n7477_), .B(new_n7452_), .ZN(new_n7489_));
  NAND2_X1   g06487(.A1(new_n7448_), .A2(new_n7449_), .ZN(new_n7490_));
  AOI21_X1   g06488(.A1(new_n7490_), .A2(new_n5656_), .B(new_n7445_), .ZN(new_n7491_));
  NOR3_X1    g06489(.A1(new_n7443_), .A2(new_n7442_), .A3(new_n5644_), .ZN(new_n7492_));
  AOI21_X1   g06490(.A1(new_n7448_), .A2(new_n7449_), .B(new_n5656_), .ZN(new_n7493_));
  OAI22_X1   g06491(.A1(new_n7491_), .A2(new_n5636_), .B1(new_n7492_), .B2(new_n7493_), .ZN(new_n7494_));
  NAND3_X1   g06492(.A1(new_n7468_), .A2(new_n5605_), .A3(new_n5657_), .ZN(new_n7495_));
  NOR2_X1    g06493(.A1(new_n7487_), .A2(new_n7495_), .ZN(new_n7496_));
  NOR3_X1    g06494(.A1(new_n7480_), .A2(new_n7483_), .A3(new_n7486_), .ZN(new_n7497_));
  OAI21_X1   g06495(.A1(new_n7496_), .A2(new_n7497_), .B(new_n7494_), .ZN(new_n7498_));
  AOI22_X1   g06496(.A1(new_n5739_), .A2(new_n5744_), .B1(new_n5659_), .B2(new_n5647_), .ZN(new_n7499_));
  NAND3_X1   g06497(.A1(new_n7489_), .A2(new_n7498_), .A3(new_n7499_), .ZN(new_n7500_));
  NOR3_X1    g06498(.A1(new_n7483_), .A2(new_n7478_), .A3(new_n7479_), .ZN(new_n7501_));
  NAND2_X1   g06499(.A1(new_n7484_), .A2(new_n7485_), .ZN(new_n7502_));
  AOI21_X1   g06500(.A1(new_n7502_), .A2(new_n5596_), .B(new_n5645_), .ZN(new_n7503_));
  NAND2_X1   g06501(.A1(new_n7501_), .A2(new_n7503_), .ZN(new_n7504_));
  OAI21_X1   g06502(.A1(new_n7483_), .A2(new_n7486_), .B(new_n7495_), .ZN(new_n7505_));
  AOI21_X1   g06503(.A1(new_n7504_), .A2(new_n7505_), .B(new_n7494_), .ZN(new_n7506_));
  OAI21_X1   g06504(.A1(new_n7483_), .A2(new_n7486_), .B(new_n7480_), .ZN(new_n7507_));
  OAI21_X1   g06505(.A1(new_n7473_), .A2(new_n7474_), .B(new_n5596_), .ZN(new_n7508_));
  NAND3_X1   g06506(.A1(new_n7495_), .A2(new_n7467_), .A3(new_n7508_), .ZN(new_n7509_));
  AOI21_X1   g06507(.A1(new_n7507_), .A2(new_n7509_), .B(new_n7452_), .ZN(new_n7510_));
  NAND2_X1   g06508(.A1(new_n5745_), .A2(new_n5747_), .ZN(new_n7511_));
  OAI21_X1   g06509(.A1(new_n7506_), .A2(new_n7510_), .B(new_n7511_), .ZN(new_n7512_));
  AOI21_X1   g06510(.A1(new_n7512_), .A2(new_n7500_), .B(new_n7441_), .ZN(new_n7513_));
  NOR2_X1    g06511(.A1(new_n7434_), .A2(new_n7435_), .ZN(new_n7514_));
  NOR4_X1    g06512(.A1(new_n7514_), .A2(new_n7425_), .A3(new_n7415_), .A4(new_n5728_), .ZN(new_n7515_));
  AOI21_X1   g06513(.A1(new_n7425_), .A2(new_n5689_), .B(new_n5737_), .ZN(new_n7516_));
  NAND2_X1   g06514(.A1(new_n7515_), .A2(new_n7516_), .ZN(new_n7517_));
  NAND2_X1   g06515(.A1(new_n7436_), .A2(new_n7438_), .ZN(new_n7518_));
  AOI21_X1   g06516(.A1(new_n7517_), .A2(new_n7518_), .B(new_n7433_), .ZN(new_n7519_));
  NAND2_X1   g06517(.A1(new_n7426_), .A2(new_n7438_), .ZN(new_n7520_));
  NAND2_X1   g06518(.A1(new_n7436_), .A2(new_n7422_), .ZN(new_n7521_));
  AOI21_X1   g06519(.A1(new_n7520_), .A2(new_n7521_), .B(new_n7400_), .ZN(new_n7522_));
  NOR2_X1    g06520(.A1(new_n7519_), .A2(new_n7522_), .ZN(new_n7523_));
  NAND3_X1   g06521(.A1(new_n7489_), .A2(new_n7498_), .A3(new_n7511_), .ZN(new_n7524_));
  OAI21_X1   g06522(.A1(new_n7506_), .A2(new_n7510_), .B(new_n7499_), .ZN(new_n7525_));
  AOI21_X1   g06523(.A1(new_n7524_), .A2(new_n7525_), .B(new_n7523_), .ZN(new_n7526_));
  NOR2_X1    g06524(.A1(new_n7526_), .A2(new_n7513_), .ZN(new_n7527_));
  NOR2_X1    g06525(.A1(new_n5521_), .A2(new_n5523_), .ZN(new_n7528_));
  INV_X1     g06526(.I(new_n5540_), .ZN(new_n7529_));
  OAI21_X1   g06527(.A1(new_n7528_), .A2(new_n5519_), .B(new_n7529_), .ZN(new_n7530_));
  NAND2_X1   g06528(.A1(new_n7530_), .A2(new_n5544_), .ZN(new_n7531_));
  NOR2_X1    g06529(.A1(new_n5515_), .A2(new_n5516_), .ZN(new_n7532_));
  INV_X1     g06530(.I(new_n5543_), .ZN(new_n7533_));
  OAI21_X1   g06531(.A1(new_n7532_), .A2(new_n5512_), .B(new_n7533_), .ZN(new_n7534_));
  NAND2_X1   g06532(.A1(new_n7534_), .A2(new_n5541_), .ZN(new_n7535_));
  NAND2_X1   g06533(.A1(new_n7531_), .A2(new_n7535_), .ZN(new_n7536_));
  AOI22_X1   g06534(.A1(new_n5514_), .A2(new_n5517_), .B1(new_n5535_), .B2(new_n5534_), .ZN(new_n7537_));
  NOR2_X1    g06535(.A1(new_n5544_), .A2(new_n5541_), .ZN(new_n7538_));
  AOI21_X1   g06536(.A1(new_n7536_), .A2(new_n7537_), .B(new_n7538_), .ZN(new_n7539_));
  NAND3_X1   g06537(.A1(new_n7531_), .A2(new_n7535_), .A3(new_n7537_), .ZN(new_n7540_));
  NOR2_X1    g06538(.A1(new_n7534_), .A2(new_n5541_), .ZN(new_n7541_));
  NOR2_X1    g06539(.A1(new_n7530_), .A2(new_n5544_), .ZN(new_n7542_));
  OAI21_X1   g06540(.A1(new_n7541_), .A2(new_n7542_), .B(new_n5545_), .ZN(new_n7543_));
  NAND2_X1   g06541(.A1(new_n7543_), .A2(new_n7540_), .ZN(new_n7544_));
  OAI21_X1   g06542(.A1(new_n5538_), .A2(new_n7539_), .B(new_n7544_), .ZN(new_n7545_));
  NOR2_X1    g06543(.A1(new_n5505_), .A2(new_n5553_), .ZN(new_n7546_));
  NOR2_X1    g06544(.A1(new_n5501_), .A2(new_n5555_), .ZN(new_n7547_));
  NOR3_X1    g06545(.A1(new_n7546_), .A2(new_n7547_), .A3(new_n5556_), .ZN(new_n7548_));
  NAND2_X1   g06546(.A1(new_n5501_), .A2(new_n5555_), .ZN(new_n7549_));
  NAND2_X1   g06547(.A1(new_n5505_), .A2(new_n5553_), .ZN(new_n7550_));
  AOI21_X1   g06548(.A1(new_n7549_), .A2(new_n7550_), .B(new_n5506_), .ZN(new_n7551_));
  NOR2_X1    g06549(.A1(new_n7551_), .A2(new_n7548_), .ZN(new_n7552_));
  OAI22_X1   g06550(.A1(new_n5529_), .A2(new_n5537_), .B1(new_n5549_), .B2(new_n5550_), .ZN(new_n7553_));
  NOR3_X1    g06551(.A1(new_n7552_), .A2(new_n5557_), .A3(new_n7553_), .ZN(new_n7554_));
  OAI21_X1   g06552(.A1(new_n7546_), .A2(new_n7547_), .B(new_n5506_), .ZN(new_n7555_));
  NOR2_X1    g06553(.A1(new_n5553_), .A2(new_n5555_), .ZN(new_n7556_));
  INV_X1     g06554(.I(new_n7556_), .ZN(new_n7557_));
  NAND2_X1   g06555(.A1(new_n7555_), .A2(new_n7557_), .ZN(new_n7558_));
  AOI21_X1   g06556(.A1(new_n7558_), .A2(new_n5497_), .B(new_n5546_), .ZN(new_n7559_));
  NAND2_X1   g06557(.A1(new_n7554_), .A2(new_n7559_), .ZN(new_n7560_));
  NAND4_X1   g06558(.A1(new_n5560_), .A2(new_n5559_), .A3(new_n5497_), .A4(new_n5507_), .ZN(new_n7561_));
  NAND3_X1   g06559(.A1(new_n7549_), .A2(new_n7550_), .A3(new_n5506_), .ZN(new_n7562_));
  OAI21_X1   g06560(.A1(new_n7546_), .A2(new_n7547_), .B(new_n5556_), .ZN(new_n7563_));
  NAND2_X1   g06561(.A1(new_n7563_), .A2(new_n7562_), .ZN(new_n7564_));
  AOI21_X1   g06562(.A1(new_n7550_), .A2(new_n7549_), .B(new_n5556_), .ZN(new_n7565_));
  OAI21_X1   g06563(.A1(new_n7565_), .A2(new_n7556_), .B(new_n5497_), .ZN(new_n7566_));
  NAND2_X1   g06564(.A1(new_n7566_), .A2(new_n7564_), .ZN(new_n7567_));
  NAND2_X1   g06565(.A1(new_n7567_), .A2(new_n7561_), .ZN(new_n7568_));
  AOI21_X1   g06566(.A1(new_n7560_), .A2(new_n7568_), .B(new_n7545_), .ZN(new_n7569_));
  OAI21_X1   g06567(.A1(new_n7542_), .A2(new_n7541_), .B(new_n7537_), .ZN(new_n7570_));
  INV_X1     g06568(.I(new_n7538_), .ZN(new_n7571_));
  NAND2_X1   g06569(.A1(new_n7570_), .A2(new_n7571_), .ZN(new_n7572_));
  NOR3_X1    g06570(.A1(new_n7541_), .A2(new_n7542_), .A3(new_n5545_), .ZN(new_n7573_));
  AOI21_X1   g06571(.A1(new_n7531_), .A2(new_n7535_), .B(new_n7537_), .ZN(new_n7574_));
  NOR2_X1    g06572(.A1(new_n7574_), .A2(new_n7573_), .ZN(new_n7575_));
  AOI21_X1   g06573(.A1(new_n5559_), .A2(new_n7572_), .B(new_n7575_), .ZN(new_n7576_));
  NAND3_X1   g06574(.A1(new_n7561_), .A2(new_n7566_), .A3(new_n7564_), .ZN(new_n7577_));
  NOR3_X1    g06575(.A1(new_n7553_), .A2(new_n5557_), .A3(new_n5546_), .ZN(new_n7578_));
  NAND2_X1   g06576(.A1(new_n7567_), .A2(new_n7578_), .ZN(new_n7579_));
  AOI21_X1   g06577(.A1(new_n7579_), .A2(new_n7577_), .B(new_n7576_), .ZN(new_n7580_));
  NOR2_X1    g06578(.A1(new_n7569_), .A2(new_n7580_), .ZN(new_n7581_));
  AOI22_X1   g06579(.A1(new_n5562_), .A2(new_n5548_), .B1(new_n5439_), .B2(new_n5467_), .ZN(new_n7582_));
  NAND2_X1   g06580(.A1(new_n5460_), .A2(new_n5436_), .ZN(new_n7583_));
  NAND2_X1   g06581(.A1(new_n5463_), .A2(new_n5434_), .ZN(new_n7584_));
  NAND2_X1   g06582(.A1(new_n7583_), .A2(new_n7584_), .ZN(new_n7585_));
  NOR2_X1    g06583(.A1(new_n5436_), .A2(new_n5434_), .ZN(new_n7586_));
  AOI21_X1   g06584(.A1(new_n7585_), .A2(new_n5464_), .B(new_n7586_), .ZN(new_n7587_));
  NOR2_X1    g06585(.A1(new_n5463_), .A2(new_n5434_), .ZN(new_n7588_));
  NOR2_X1    g06586(.A1(new_n5460_), .A2(new_n5436_), .ZN(new_n7589_));
  NOR4_X1    g06587(.A1(new_n7589_), .A2(new_n7588_), .A3(new_n5432_), .A4(new_n5428_), .ZN(new_n7590_));
  AOI21_X1   g06588(.A1(new_n7583_), .A2(new_n7584_), .B(new_n5464_), .ZN(new_n7591_));
  OAI22_X1   g06589(.A1(new_n7587_), .A2(new_n5429_), .B1(new_n7590_), .B2(new_n7591_), .ZN(new_n7592_));
  NOR2_X1    g06590(.A1(new_n5408_), .A2(new_n5444_), .ZN(new_n7593_));
  NOR2_X1    g06591(.A1(new_n5404_), .A2(new_n5446_), .ZN(new_n7594_));
  NOR3_X1    g06592(.A1(new_n7593_), .A2(new_n7594_), .A3(new_n5447_), .ZN(new_n7595_));
  NAND2_X1   g06593(.A1(new_n5404_), .A2(new_n5446_), .ZN(new_n7596_));
  NAND2_X1   g06594(.A1(new_n5408_), .A2(new_n5444_), .ZN(new_n7597_));
  AOI21_X1   g06595(.A1(new_n7597_), .A2(new_n7596_), .B(new_n5409_), .ZN(new_n7598_));
  NOR2_X1    g06596(.A1(new_n7598_), .A2(new_n7595_), .ZN(new_n7599_));
  OAI21_X1   g06597(.A1(new_n7593_), .A2(new_n7594_), .B(new_n5409_), .ZN(new_n7600_));
  NOR2_X1    g06598(.A1(new_n5444_), .A2(new_n5446_), .ZN(new_n7601_));
  INV_X1     g06599(.I(new_n7601_), .ZN(new_n7602_));
  NAND2_X1   g06600(.A1(new_n7600_), .A2(new_n7602_), .ZN(new_n7603_));
  NOR4_X1    g06601(.A1(new_n7599_), .A2(new_n7603_), .A3(new_n5442_), .A4(new_n5429_), .ZN(new_n7604_));
  AOI21_X1   g06602(.A1(new_n7603_), .A2(new_n5400_), .B(new_n5437_), .ZN(new_n7605_));
  NAND2_X1   g06603(.A1(new_n7604_), .A2(new_n7605_), .ZN(new_n7606_));
  NAND4_X1   g06604(.A1(new_n5400_), .A2(new_n5457_), .A3(new_n5410_), .A4(new_n5465_), .ZN(new_n7607_));
  NAND3_X1   g06605(.A1(new_n7597_), .A2(new_n7596_), .A3(new_n5409_), .ZN(new_n7608_));
  OAI21_X1   g06606(.A1(new_n7593_), .A2(new_n7594_), .B(new_n5447_), .ZN(new_n7609_));
  NAND2_X1   g06607(.A1(new_n7609_), .A2(new_n7608_), .ZN(new_n7610_));
  AOI21_X1   g06608(.A1(new_n7597_), .A2(new_n7596_), .B(new_n5447_), .ZN(new_n7611_));
  OAI21_X1   g06609(.A1(new_n7611_), .A2(new_n7601_), .B(new_n5400_), .ZN(new_n7612_));
  NAND2_X1   g06610(.A1(new_n7612_), .A2(new_n7610_), .ZN(new_n7613_));
  NAND2_X1   g06611(.A1(new_n7613_), .A2(new_n7607_), .ZN(new_n7614_));
  AOI21_X1   g06612(.A1(new_n7606_), .A2(new_n7614_), .B(new_n7592_), .ZN(new_n7615_));
  OAI21_X1   g06613(.A1(new_n7589_), .A2(new_n7588_), .B(new_n5464_), .ZN(new_n7616_));
  INV_X1     g06614(.I(new_n7586_), .ZN(new_n7617_));
  NAND2_X1   g06615(.A1(new_n7616_), .A2(new_n7617_), .ZN(new_n7618_));
  NAND3_X1   g06616(.A1(new_n7583_), .A2(new_n7584_), .A3(new_n5464_), .ZN(new_n7619_));
  OAI22_X1   g06617(.A1(new_n7589_), .A2(new_n7588_), .B1(new_n5432_), .B2(new_n5428_), .ZN(new_n7620_));
  AOI22_X1   g06618(.A1(new_n7618_), .A2(new_n5457_), .B1(new_n7619_), .B2(new_n7620_), .ZN(new_n7621_));
  NOR4_X1    g06619(.A1(new_n5429_), .A2(new_n5442_), .A3(new_n5448_), .A4(new_n5437_), .ZN(new_n7622_));
  NAND2_X1   g06620(.A1(new_n7613_), .A2(new_n7622_), .ZN(new_n7623_));
  NAND3_X1   g06621(.A1(new_n7612_), .A2(new_n7607_), .A3(new_n7610_), .ZN(new_n7624_));
  AOI21_X1   g06622(.A1(new_n7623_), .A2(new_n7624_), .B(new_n7621_), .ZN(new_n7625_));
  OAI21_X1   g06623(.A1(new_n7615_), .A2(new_n7625_), .B(new_n7582_), .ZN(new_n7626_));
  NAND2_X1   g06624(.A1(new_n5563_), .A2(new_n5565_), .ZN(new_n7627_));
  NAND4_X1   g06625(.A1(new_n7610_), .A2(new_n5400_), .A3(new_n5410_), .A4(new_n5457_), .ZN(new_n7628_));
  NOR2_X1    g06626(.A1(new_n7611_), .A2(new_n7601_), .ZN(new_n7629_));
  OAI21_X1   g06627(.A1(new_n7629_), .A2(new_n5442_), .B(new_n5465_), .ZN(new_n7630_));
  NOR2_X1    g06628(.A1(new_n7628_), .A2(new_n7630_), .ZN(new_n7631_));
  AOI21_X1   g06629(.A1(new_n7610_), .A2(new_n7612_), .B(new_n7622_), .ZN(new_n7632_));
  OAI21_X1   g06630(.A1(new_n7631_), .A2(new_n7632_), .B(new_n7621_), .ZN(new_n7633_));
  AOI21_X1   g06631(.A1(new_n7610_), .A2(new_n7612_), .B(new_n7607_), .ZN(new_n7634_));
  AOI21_X1   g06632(.A1(new_n7600_), .A2(new_n7602_), .B(new_n5442_), .ZN(new_n7635_));
  NOR3_X1    g06633(.A1(new_n7622_), .A2(new_n7635_), .A3(new_n7599_), .ZN(new_n7636_));
  OAI21_X1   g06634(.A1(new_n7636_), .A2(new_n7634_), .B(new_n7592_), .ZN(new_n7637_));
  NAND3_X1   g06635(.A1(new_n7633_), .A2(new_n7627_), .A3(new_n7637_), .ZN(new_n7638_));
  AOI21_X1   g06636(.A1(new_n7626_), .A2(new_n7638_), .B(new_n7581_), .ZN(new_n7639_));
  NAND4_X1   g06637(.A1(new_n7564_), .A2(new_n5497_), .A3(new_n5507_), .A4(new_n5559_), .ZN(new_n7640_));
  AOI21_X1   g06638(.A1(new_n7555_), .A2(new_n7557_), .B(new_n5551_), .ZN(new_n7641_));
  NOR3_X1    g06639(.A1(new_n7640_), .A2(new_n5546_), .A3(new_n7641_), .ZN(new_n7642_));
  NOR2_X1    g06640(.A1(new_n7641_), .A2(new_n7552_), .ZN(new_n7643_));
  NOR2_X1    g06641(.A1(new_n7643_), .A2(new_n7578_), .ZN(new_n7644_));
  OAI21_X1   g06642(.A1(new_n7642_), .A2(new_n7644_), .B(new_n7576_), .ZN(new_n7645_));
  NOR2_X1    g06643(.A1(new_n7567_), .A2(new_n7578_), .ZN(new_n7646_));
  NOR2_X1    g06644(.A1(new_n7643_), .A2(new_n7561_), .ZN(new_n7647_));
  OAI21_X1   g06645(.A1(new_n7647_), .A2(new_n7646_), .B(new_n7545_), .ZN(new_n7648_));
  NAND2_X1   g06646(.A1(new_n7645_), .A2(new_n7648_), .ZN(new_n7649_));
  OAI21_X1   g06647(.A1(new_n7615_), .A2(new_n7625_), .B(new_n7627_), .ZN(new_n7650_));
  NAND3_X1   g06648(.A1(new_n7633_), .A2(new_n7637_), .A3(new_n7582_), .ZN(new_n7651_));
  AOI21_X1   g06649(.A1(new_n7650_), .A2(new_n7651_), .B(new_n7649_), .ZN(new_n7652_));
  AOI22_X1   g06650(.A1(new_n5564_), .A2(new_n5566_), .B1(new_n5746_), .B2(new_n5748_), .ZN(new_n7653_));
  INV_X1     g06651(.I(new_n7653_), .ZN(new_n7654_));
  NOR3_X1    g06652(.A1(new_n7652_), .A2(new_n7639_), .A3(new_n7654_), .ZN(new_n7655_));
  AOI21_X1   g06653(.A1(new_n7633_), .A2(new_n7637_), .B(new_n7627_), .ZN(new_n7656_));
  NOR3_X1    g06654(.A1(new_n7615_), .A2(new_n7625_), .A3(new_n7582_), .ZN(new_n7657_));
  OAI21_X1   g06655(.A1(new_n7657_), .A2(new_n7656_), .B(new_n7649_), .ZN(new_n7658_));
  AOI21_X1   g06656(.A1(new_n7633_), .A2(new_n7637_), .B(new_n7582_), .ZN(new_n7659_));
  NOR3_X1    g06657(.A1(new_n7615_), .A2(new_n7625_), .A3(new_n7627_), .ZN(new_n7660_));
  OAI21_X1   g06658(.A1(new_n7660_), .A2(new_n7659_), .B(new_n7581_), .ZN(new_n7661_));
  AOI21_X1   g06659(.A1(new_n7658_), .A2(new_n7661_), .B(new_n7653_), .ZN(new_n7662_));
  OAI21_X1   g06660(.A1(new_n7655_), .A2(new_n7662_), .B(new_n7527_), .ZN(new_n7663_));
  NOR3_X1    g06661(.A1(new_n7506_), .A2(new_n7511_), .A3(new_n7510_), .ZN(new_n7664_));
  AOI21_X1   g06662(.A1(new_n7489_), .A2(new_n7498_), .B(new_n7499_), .ZN(new_n7665_));
  OAI21_X1   g06663(.A1(new_n7664_), .A2(new_n7665_), .B(new_n7523_), .ZN(new_n7666_));
  NOR3_X1    g06664(.A1(new_n7506_), .A2(new_n7510_), .A3(new_n7499_), .ZN(new_n7667_));
  AOI21_X1   g06665(.A1(new_n7489_), .A2(new_n7498_), .B(new_n7511_), .ZN(new_n7668_));
  OAI21_X1   g06666(.A1(new_n7667_), .A2(new_n7668_), .B(new_n7441_), .ZN(new_n7669_));
  NAND2_X1   g06667(.A1(new_n7666_), .A2(new_n7669_), .ZN(new_n7670_));
  NAND3_X1   g06668(.A1(new_n7658_), .A2(new_n7661_), .A3(new_n7654_), .ZN(new_n7671_));
  OAI21_X1   g06669(.A1(new_n7652_), .A2(new_n7639_), .B(new_n7653_), .ZN(new_n7672_));
  NAND2_X1   g06670(.A1(new_n7672_), .A2(new_n7671_), .ZN(new_n7673_));
  NAND2_X1   g06671(.A1(new_n7673_), .A2(new_n7670_), .ZN(new_n7674_));
  NAND2_X1   g06672(.A1(new_n7674_), .A2(new_n7663_), .ZN(new_n7675_));
  INV_X1     g06673(.I(new_n7675_), .ZN(new_n7676_));
  NAND2_X1   g06674(.A1(new_n5359_), .A2(new_n5340_), .ZN(new_n7677_));
  NAND2_X1   g06675(.A1(new_n5362_), .A2(new_n5337_), .ZN(new_n7678_));
  AOI21_X1   g06676(.A1(new_n7677_), .A2(new_n7678_), .B(new_n5345_), .ZN(new_n7679_));
  NOR2_X1    g06677(.A1(new_n5340_), .A2(new_n5337_), .ZN(new_n7680_));
  NOR2_X1    g06678(.A1(new_n7679_), .A2(new_n7680_), .ZN(new_n7681_));
  NOR2_X1    g06679(.A1(new_n5362_), .A2(new_n5337_), .ZN(new_n7682_));
  NOR2_X1    g06680(.A1(new_n5359_), .A2(new_n5340_), .ZN(new_n7683_));
  NOR3_X1    g06681(.A1(new_n7683_), .A2(new_n7682_), .A3(new_n5345_), .ZN(new_n7684_));
  AOI22_X1   g06682(.A1(new_n7677_), .A2(new_n7678_), .B1(new_n5354_), .B2(new_n5333_), .ZN(new_n7685_));
  OAI22_X1   g06683(.A1(new_n7681_), .A2(new_n5334_), .B1(new_n7684_), .B2(new_n7685_), .ZN(new_n7686_));
  NOR2_X1    g06684(.A1(new_n5279_), .A2(new_n5281_), .ZN(new_n7687_));
  INV_X1     g06685(.I(new_n5310_), .ZN(new_n7688_));
  OAI21_X1   g06686(.A1(new_n7687_), .A2(new_n5277_), .B(new_n7688_), .ZN(new_n7689_));
  NOR2_X1    g06687(.A1(new_n7689_), .A2(new_n5308_), .ZN(new_n7690_));
  NOR2_X1    g06688(.A1(new_n5293_), .A2(new_n5294_), .ZN(new_n7691_));
  INV_X1     g06689(.I(new_n5307_), .ZN(new_n7692_));
  OAI21_X1   g06690(.A1(new_n7691_), .A2(new_n5292_), .B(new_n7692_), .ZN(new_n7693_));
  NOR2_X1    g06691(.A1(new_n7693_), .A2(new_n5311_), .ZN(new_n7694_));
  NOR3_X1    g06692(.A1(new_n7690_), .A2(new_n7694_), .A3(new_n5312_), .ZN(new_n7695_));
  NAND2_X1   g06693(.A1(new_n7693_), .A2(new_n5311_), .ZN(new_n7696_));
  NAND2_X1   g06694(.A1(new_n7689_), .A2(new_n5308_), .ZN(new_n7697_));
  AOI22_X1   g06695(.A1(new_n5298_), .A2(new_n5299_), .B1(new_n5295_), .B2(new_n5291_), .ZN(new_n7698_));
  AOI21_X1   g06696(.A1(new_n7696_), .A2(new_n7697_), .B(new_n7698_), .ZN(new_n7699_));
  NOR2_X1    g06697(.A1(new_n7699_), .A2(new_n7695_), .ZN(new_n7700_));
  NOR4_X1    g06698(.A1(new_n7700_), .A2(new_n5351_), .A3(new_n5313_), .A4(new_n5334_), .ZN(new_n7701_));
  OAI21_X1   g06699(.A1(new_n7690_), .A2(new_n7694_), .B(new_n7698_), .ZN(new_n7702_));
  NOR2_X1    g06700(.A1(new_n5308_), .A2(new_n5311_), .ZN(new_n7703_));
  INV_X1     g06701(.I(new_n7703_), .ZN(new_n7704_));
  AOI22_X1   g06702(.A1(new_n7702_), .A2(new_n7704_), .B1(new_n5297_), .B2(new_n5304_), .ZN(new_n7705_));
  NOR2_X1    g06703(.A1(new_n7705_), .A2(new_n5346_), .ZN(new_n7706_));
  NAND2_X1   g06704(.A1(new_n7701_), .A2(new_n7706_), .ZN(new_n7707_));
  AOI22_X1   g06705(.A1(new_n5353_), .A2(new_n5356_), .B1(new_n5304_), .B2(new_n5297_), .ZN(new_n7708_));
  NAND3_X1   g06706(.A1(new_n7708_), .A2(new_n5314_), .A3(new_n5363_), .ZN(new_n7709_));
  AOI21_X1   g06707(.A1(new_n7696_), .A2(new_n7697_), .B(new_n5312_), .ZN(new_n7710_));
  NOR2_X1    g06708(.A1(new_n7710_), .A2(new_n7703_), .ZN(new_n7711_));
  OAI22_X1   g06709(.A1(new_n7711_), .A2(new_n5351_), .B1(new_n7695_), .B2(new_n7699_), .ZN(new_n7712_));
  NAND2_X1   g06710(.A1(new_n7712_), .A2(new_n7709_), .ZN(new_n7713_));
  AOI21_X1   g06711(.A1(new_n7707_), .A2(new_n7713_), .B(new_n7686_), .ZN(new_n7714_));
  NOR2_X1    g06712(.A1(new_n7683_), .A2(new_n7682_), .ZN(new_n7715_));
  INV_X1     g06713(.I(new_n7680_), .ZN(new_n7716_));
  OAI21_X1   g06714(.A1(new_n7715_), .A2(new_n5345_), .B(new_n7716_), .ZN(new_n7717_));
  NAND4_X1   g06715(.A1(new_n7677_), .A2(new_n7678_), .A3(new_n5354_), .A4(new_n5333_), .ZN(new_n7718_));
  OAI21_X1   g06716(.A1(new_n7683_), .A2(new_n7682_), .B(new_n5345_), .ZN(new_n7719_));
  AOI22_X1   g06717(.A1(new_n7717_), .A2(new_n5357_), .B1(new_n7718_), .B2(new_n7719_), .ZN(new_n7720_));
  NOR2_X1    g06718(.A1(new_n7705_), .A2(new_n7700_), .ZN(new_n7721_));
  NAND2_X1   g06719(.A1(new_n7721_), .A2(new_n7709_), .ZN(new_n7722_));
  NOR4_X1    g06720(.A1(new_n5334_), .A2(new_n5351_), .A3(new_n5313_), .A4(new_n5346_), .ZN(new_n7723_));
  NAND2_X1   g06721(.A1(new_n7712_), .A2(new_n7723_), .ZN(new_n7724_));
  AOI21_X1   g06722(.A1(new_n7722_), .A2(new_n7724_), .B(new_n7720_), .ZN(new_n7725_));
  NOR2_X1    g06723(.A1(new_n7714_), .A2(new_n7725_), .ZN(new_n7726_));
  NOR2_X1    g06724(.A1(new_n5229_), .A2(new_n5231_), .ZN(new_n7727_));
  OAI21_X1   g06725(.A1(new_n7727_), .A2(new_n5227_), .B(new_n5249_), .ZN(new_n7728_));
  NAND2_X1   g06726(.A1(new_n7728_), .A2(new_n5253_), .ZN(new_n7729_));
  NOR2_X1    g06727(.A1(new_n5223_), .A2(new_n5224_), .ZN(new_n7730_));
  INV_X1     g06728(.I(new_n5252_), .ZN(new_n7731_));
  OAI21_X1   g06729(.A1(new_n7730_), .A2(new_n5222_), .B(new_n7731_), .ZN(new_n7732_));
  NAND2_X1   g06730(.A1(new_n7732_), .A2(new_n5251_), .ZN(new_n7733_));
  NAND2_X1   g06731(.A1(new_n7733_), .A2(new_n7729_), .ZN(new_n7734_));
  AOI22_X1   g06732(.A1(new_n5239_), .A2(new_n5240_), .B1(new_n5232_), .B2(new_n5235_), .ZN(new_n7735_));
  NOR2_X1    g06733(.A1(new_n5251_), .A2(new_n5253_), .ZN(new_n7736_));
  AOI21_X1   g06734(.A1(new_n7734_), .A2(new_n7735_), .B(new_n7736_), .ZN(new_n7737_));
  NOR2_X1    g06735(.A1(new_n7732_), .A2(new_n5251_), .ZN(new_n7738_));
  NOR2_X1    g06736(.A1(new_n7728_), .A2(new_n5253_), .ZN(new_n7739_));
  NOR3_X1    g06737(.A1(new_n7738_), .A2(new_n7739_), .A3(new_n5254_), .ZN(new_n7740_));
  AOI21_X1   g06738(.A1(new_n7733_), .A2(new_n7729_), .B(new_n7735_), .ZN(new_n7741_));
  OAI22_X1   g06739(.A1(new_n7737_), .A2(new_n5273_), .B1(new_n7740_), .B2(new_n7741_), .ZN(new_n7742_));
  NOR2_X1    g06740(.A1(new_n5264_), .A2(new_n5213_), .ZN(new_n7743_));
  NOR2_X1    g06741(.A1(new_n5266_), .A2(new_n5209_), .ZN(new_n7744_));
  NOR3_X1    g06742(.A1(new_n7743_), .A2(new_n7744_), .A3(new_n5214_), .ZN(new_n7745_));
  NAND2_X1   g06743(.A1(new_n5266_), .A2(new_n5209_), .ZN(new_n7746_));
  NAND2_X1   g06744(.A1(new_n5264_), .A2(new_n5213_), .ZN(new_n7747_));
  AOI21_X1   g06745(.A1(new_n7747_), .A2(new_n7746_), .B(new_n5268_), .ZN(new_n7748_));
  NOR2_X1    g06746(.A1(new_n7748_), .A2(new_n7745_), .ZN(new_n7749_));
  NOR2_X1    g06747(.A1(new_n5209_), .A2(new_n5213_), .ZN(new_n7750_));
  INV_X1     g06748(.I(new_n7750_), .ZN(new_n7751_));
  OAI21_X1   g06749(.A1(new_n7743_), .A2(new_n7744_), .B(new_n5268_), .ZN(new_n7752_));
  NAND2_X1   g06750(.A1(new_n7752_), .A2(new_n7751_), .ZN(new_n7753_));
  NOR4_X1    g06751(.A1(new_n7749_), .A2(new_n7753_), .A3(new_n5206_), .A4(new_n5273_), .ZN(new_n7754_));
  AOI21_X1   g06752(.A1(new_n7753_), .A2(new_n5261_), .B(new_n5255_), .ZN(new_n7755_));
  NAND2_X1   g06753(.A1(new_n7754_), .A2(new_n7755_), .ZN(new_n7756_));
  AOI22_X1   g06754(.A1(new_n5246_), .A2(new_n5237_), .B1(new_n5260_), .B2(new_n5259_), .ZN(new_n7757_));
  NAND3_X1   g06755(.A1(new_n7757_), .A2(new_n5256_), .A3(new_n5269_), .ZN(new_n7758_));
  NAND3_X1   g06756(.A1(new_n7746_), .A2(new_n7747_), .A3(new_n5268_), .ZN(new_n7759_));
  OAI21_X1   g06757(.A1(new_n7743_), .A2(new_n7744_), .B(new_n5214_), .ZN(new_n7760_));
  NAND2_X1   g06758(.A1(new_n7760_), .A2(new_n7759_), .ZN(new_n7761_));
  AOI21_X1   g06759(.A1(new_n7747_), .A2(new_n7746_), .B(new_n5214_), .ZN(new_n7762_));
  OAI21_X1   g06760(.A1(new_n7750_), .A2(new_n7762_), .B(new_n5261_), .ZN(new_n7763_));
  NAND2_X1   g06761(.A1(new_n7763_), .A2(new_n7761_), .ZN(new_n7764_));
  NAND2_X1   g06762(.A1(new_n7764_), .A2(new_n7758_), .ZN(new_n7765_));
  AOI21_X1   g06763(.A1(new_n7756_), .A2(new_n7765_), .B(new_n7742_), .ZN(new_n7766_));
  OAI21_X1   g06764(.A1(new_n7738_), .A2(new_n7739_), .B(new_n7735_), .ZN(new_n7767_));
  INV_X1     g06765(.I(new_n7736_), .ZN(new_n7768_));
  NAND2_X1   g06766(.A1(new_n7767_), .A2(new_n7768_), .ZN(new_n7769_));
  NAND3_X1   g06767(.A1(new_n7729_), .A2(new_n7733_), .A3(new_n7735_), .ZN(new_n7770_));
  OAI21_X1   g06768(.A1(new_n7738_), .A2(new_n7739_), .B(new_n5254_), .ZN(new_n7771_));
  AOI22_X1   g06769(.A1(new_n7769_), .A2(new_n5247_), .B1(new_n7770_), .B2(new_n7771_), .ZN(new_n7772_));
  NAND3_X1   g06770(.A1(new_n7758_), .A2(new_n7761_), .A3(new_n7763_), .ZN(new_n7773_));
  NOR4_X1    g06771(.A1(new_n5273_), .A2(new_n5206_), .A3(new_n5215_), .A4(new_n5255_), .ZN(new_n7774_));
  NAND2_X1   g06772(.A1(new_n7764_), .A2(new_n7774_), .ZN(new_n7775_));
  AOI21_X1   g06773(.A1(new_n7775_), .A2(new_n7773_), .B(new_n7772_), .ZN(new_n7776_));
  NAND2_X1   g06774(.A1(new_n5367_), .A2(new_n5276_), .ZN(new_n7777_));
  NOR3_X1    g06775(.A1(new_n7766_), .A2(new_n7777_), .A3(new_n7776_), .ZN(new_n7778_));
  NAND3_X1   g06776(.A1(new_n7761_), .A2(new_n5269_), .A3(new_n7757_), .ZN(new_n7779_));
  NOR2_X1    g06777(.A1(new_n7762_), .A2(new_n7750_), .ZN(new_n7780_));
  OAI21_X1   g06778(.A1(new_n7780_), .A2(new_n5206_), .B(new_n5256_), .ZN(new_n7781_));
  NOR2_X1    g06779(.A1(new_n7779_), .A2(new_n7781_), .ZN(new_n7782_));
  AOI21_X1   g06780(.A1(new_n7751_), .A2(new_n7752_), .B(new_n5206_), .ZN(new_n7783_));
  NOR2_X1    g06781(.A1(new_n7783_), .A2(new_n7749_), .ZN(new_n7784_));
  NOR2_X1    g06782(.A1(new_n7784_), .A2(new_n7774_), .ZN(new_n7785_));
  OAI21_X1   g06783(.A1(new_n7785_), .A2(new_n7782_), .B(new_n7772_), .ZN(new_n7786_));
  NOR2_X1    g06784(.A1(new_n7764_), .A2(new_n7774_), .ZN(new_n7787_));
  NOR2_X1    g06785(.A1(new_n7784_), .A2(new_n7758_), .ZN(new_n7788_));
  OAI21_X1   g06786(.A1(new_n7788_), .A2(new_n7787_), .B(new_n7742_), .ZN(new_n7789_));
  AOI22_X1   g06787(.A1(new_n5348_), .A2(new_n5365_), .B1(new_n5258_), .B2(new_n5275_), .ZN(new_n7790_));
  AOI21_X1   g06788(.A1(new_n7789_), .A2(new_n7786_), .B(new_n7790_), .ZN(new_n7791_));
  OAI21_X1   g06789(.A1(new_n7778_), .A2(new_n7791_), .B(new_n7726_), .ZN(new_n7792_));
  NAND3_X1   g06790(.A1(new_n7696_), .A2(new_n7698_), .A3(new_n7697_), .ZN(new_n7793_));
  OAI21_X1   g06791(.A1(new_n7690_), .A2(new_n7694_), .B(new_n5312_), .ZN(new_n7794_));
  NAND2_X1   g06792(.A1(new_n7793_), .A2(new_n7794_), .ZN(new_n7795_));
  NAND3_X1   g06793(.A1(new_n7795_), .A2(new_n7708_), .A3(new_n5314_), .ZN(new_n7796_));
  OAI21_X1   g06794(.A1(new_n7711_), .A2(new_n5351_), .B(new_n5363_), .ZN(new_n7797_));
  NOR2_X1    g06795(.A1(new_n7796_), .A2(new_n7797_), .ZN(new_n7798_));
  NOR2_X1    g06796(.A1(new_n7721_), .A2(new_n7723_), .ZN(new_n7799_));
  OAI21_X1   g06797(.A1(new_n7799_), .A2(new_n7798_), .B(new_n7720_), .ZN(new_n7800_));
  NOR2_X1    g06798(.A1(new_n7712_), .A2(new_n7723_), .ZN(new_n7801_));
  NOR2_X1    g06799(.A1(new_n7721_), .A2(new_n7709_), .ZN(new_n7802_));
  OAI21_X1   g06800(.A1(new_n7802_), .A2(new_n7801_), .B(new_n7686_), .ZN(new_n7803_));
  NAND2_X1   g06801(.A1(new_n7803_), .A2(new_n7800_), .ZN(new_n7804_));
  NOR3_X1    g06802(.A1(new_n7766_), .A2(new_n7776_), .A3(new_n7790_), .ZN(new_n7805_));
  AOI21_X1   g06803(.A1(new_n7789_), .A2(new_n7786_), .B(new_n7777_), .ZN(new_n7806_));
  OAI21_X1   g06804(.A1(new_n7805_), .A2(new_n7806_), .B(new_n7804_), .ZN(new_n7807_));
  NAND2_X1   g06805(.A1(new_n7792_), .A2(new_n7807_), .ZN(new_n7808_));
  XOR2_X1    g06806(.A1(\A[346] ), .A2(\A[347] ), .Z(new_n7809_));
  AOI21_X1   g06807(.A1(new_n7809_), .A2(\A[348] ), .B(new_n5120_), .ZN(new_n7810_));
  NOR2_X1    g06808(.A1(new_n5129_), .A2(new_n7810_), .ZN(new_n7811_));
  INV_X1     g06809(.I(new_n5127_), .ZN(new_n7812_));
  AOI21_X1   g06810(.A1(new_n5145_), .A2(\A[345] ), .B(new_n7812_), .ZN(new_n7813_));
  NOR2_X1    g06811(.A1(new_n5125_), .A2(new_n7813_), .ZN(new_n7814_));
  NOR2_X1    g06812(.A1(new_n7814_), .A2(new_n7811_), .ZN(new_n7815_));
  NOR2_X1    g06813(.A1(new_n5128_), .A2(\A[345] ), .ZN(new_n7816_));
  OAI22_X1   g06814(.A1(new_n7816_), .A2(new_n5146_), .B1(new_n5141_), .B2(new_n5142_), .ZN(new_n7817_));
  NOR2_X1    g06815(.A1(new_n7810_), .A2(new_n7813_), .ZN(new_n7818_));
  INV_X1     g06816(.I(new_n7818_), .ZN(new_n7819_));
  OAI21_X1   g06817(.A1(new_n7815_), .A2(new_n7817_), .B(new_n7819_), .ZN(new_n7820_));
  NAND2_X1   g06818(.A1(new_n5125_), .A2(new_n7813_), .ZN(new_n7821_));
  NAND2_X1   g06819(.A1(new_n5129_), .A2(new_n7810_), .ZN(new_n7822_));
  NAND4_X1   g06820(.A1(new_n7821_), .A2(new_n7822_), .A3(new_n5134_), .A4(new_n5136_), .ZN(new_n7823_));
  OAI21_X1   g06821(.A1(new_n7811_), .A2(new_n7814_), .B(new_n7817_), .ZN(new_n7824_));
  AOI22_X1   g06822(.A1(new_n7820_), .A2(new_n5165_), .B1(new_n7823_), .B2(new_n7824_), .ZN(new_n7825_));
  NAND2_X1   g06823(.A1(new_n5093_), .A2(new_n5152_), .ZN(new_n7826_));
  NAND2_X1   g06824(.A1(new_n5084_), .A2(new_n5153_), .ZN(new_n7827_));
  NAND3_X1   g06825(.A1(new_n7826_), .A2(new_n7827_), .A3(new_n5103_), .ZN(new_n7828_));
  NOR2_X1    g06826(.A1(new_n5084_), .A2(new_n5153_), .ZN(new_n7829_));
  NOR2_X1    g06827(.A1(new_n5093_), .A2(new_n5152_), .ZN(new_n7830_));
  OAI21_X1   g06828(.A1(new_n7829_), .A2(new_n7830_), .B(new_n5157_), .ZN(new_n7831_));
  NAND2_X1   g06829(.A1(new_n7831_), .A2(new_n7828_), .ZN(new_n7832_));
  AOI22_X1   g06830(.A1(new_n5163_), .A2(new_n5164_), .B1(new_n5109_), .B2(new_n5114_), .ZN(new_n7833_));
  NAND3_X1   g06831(.A1(new_n7833_), .A2(new_n5104_), .A3(new_n5137_), .ZN(new_n7834_));
  NOR2_X1    g06832(.A1(new_n5152_), .A2(new_n5153_), .ZN(new_n7835_));
  AOI21_X1   g06833(.A1(new_n7826_), .A2(new_n7827_), .B(new_n5157_), .ZN(new_n7836_));
  OAI21_X1   g06834(.A1(new_n7835_), .A2(new_n7836_), .B(new_n5115_), .ZN(new_n7837_));
  NAND3_X1   g06835(.A1(new_n7834_), .A2(new_n7837_), .A3(new_n7832_), .ZN(new_n7838_));
  NOR3_X1    g06836(.A1(new_n7829_), .A2(new_n7830_), .A3(new_n5157_), .ZN(new_n7839_));
  AOI21_X1   g06837(.A1(new_n7826_), .A2(new_n7827_), .B(new_n5103_), .ZN(new_n7840_));
  NOR2_X1    g06838(.A1(new_n7840_), .A2(new_n7839_), .ZN(new_n7841_));
  OAI22_X1   g06839(.A1(new_n5144_), .A2(new_n5148_), .B1(new_n5160_), .B2(new_n5159_), .ZN(new_n7842_));
  NOR3_X1    g06840(.A1(new_n7842_), .A2(new_n5158_), .A3(new_n5138_), .ZN(new_n7843_));
  INV_X1     g06841(.I(new_n7835_), .ZN(new_n7844_));
  OAI21_X1   g06842(.A1(new_n7829_), .A2(new_n7830_), .B(new_n5103_), .ZN(new_n7845_));
  AOI21_X1   g06843(.A1(new_n7844_), .A2(new_n7845_), .B(new_n5161_), .ZN(new_n7846_));
  OAI21_X1   g06844(.A1(new_n7841_), .A2(new_n7846_), .B(new_n7843_), .ZN(new_n7847_));
  AOI21_X1   g06845(.A1(new_n7847_), .A2(new_n7838_), .B(new_n7825_), .ZN(new_n7848_));
  AOI21_X1   g06846(.A1(new_n7821_), .A2(new_n7822_), .B(new_n7817_), .ZN(new_n7849_));
  NOR2_X1    g06847(.A1(new_n7849_), .A2(new_n7818_), .ZN(new_n7850_));
  NOR3_X1    g06848(.A1(new_n7814_), .A2(new_n7817_), .A3(new_n7811_), .ZN(new_n7851_));
  AOI22_X1   g06849(.A1(new_n7821_), .A2(new_n7822_), .B1(new_n5134_), .B2(new_n5136_), .ZN(new_n7852_));
  OAI22_X1   g06850(.A1(new_n7850_), .A2(new_n5149_), .B1(new_n7851_), .B2(new_n7852_), .ZN(new_n7853_));
  NOR3_X1    g06851(.A1(new_n7841_), .A2(new_n5158_), .A3(new_n7842_), .ZN(new_n7854_));
  NAND2_X1   g06852(.A1(new_n7845_), .A2(new_n7844_), .ZN(new_n7855_));
  AOI21_X1   g06853(.A1(new_n7855_), .A2(new_n5115_), .B(new_n5138_), .ZN(new_n7856_));
  NAND2_X1   g06854(.A1(new_n7854_), .A2(new_n7856_), .ZN(new_n7857_));
  OAI21_X1   g06855(.A1(new_n7846_), .A2(new_n7841_), .B(new_n7834_), .ZN(new_n7858_));
  AOI21_X1   g06856(.A1(new_n7857_), .A2(new_n7858_), .B(new_n7853_), .ZN(new_n7859_));
  NOR2_X1    g06857(.A1(new_n7859_), .A2(new_n7848_), .ZN(new_n7860_));
  NOR2_X1    g06858(.A1(new_n5068_), .A2(new_n5015_), .ZN(new_n7861_));
  NOR2_X1    g06859(.A1(new_n5067_), .A2(new_n5019_), .ZN(new_n7862_));
  NOR2_X1    g06860(.A1(new_n7862_), .A2(new_n7861_), .ZN(new_n7863_));
  NOR2_X1    g06861(.A1(new_n5015_), .A2(new_n5019_), .ZN(new_n7864_));
  INV_X1     g06862(.I(new_n7864_), .ZN(new_n7865_));
  OAI21_X1   g06863(.A1(new_n7863_), .A2(new_n5038_), .B(new_n7865_), .ZN(new_n7866_));
  NOR3_X1    g06864(.A1(new_n7862_), .A2(new_n7861_), .A3(new_n5038_), .ZN(new_n7867_));
  NAND2_X1   g06865(.A1(new_n5067_), .A2(new_n5019_), .ZN(new_n7868_));
  NAND2_X1   g06866(.A1(new_n5068_), .A2(new_n5015_), .ZN(new_n7869_));
  AOI22_X1   g06867(.A1(new_n7868_), .A2(new_n7869_), .B1(new_n5042_), .B2(new_n5049_), .ZN(new_n7870_));
  NOR2_X1    g06868(.A1(new_n7870_), .A2(new_n7867_), .ZN(new_n7871_));
  AOI21_X1   g06869(.A1(new_n7866_), .A2(new_n5072_), .B(new_n7871_), .ZN(new_n7872_));
  NAND2_X1   g06870(.A1(new_n4981_), .A2(new_n5055_), .ZN(new_n7873_));
  NAND2_X1   g06871(.A1(new_n4977_), .A2(new_n5058_), .ZN(new_n7874_));
  NAND3_X1   g06872(.A1(new_n7873_), .A2(new_n7874_), .A3(new_n4998_), .ZN(new_n7875_));
  NOR2_X1    g06873(.A1(new_n4977_), .A2(new_n5058_), .ZN(new_n7876_));
  NOR2_X1    g06874(.A1(new_n4981_), .A2(new_n5055_), .ZN(new_n7877_));
  OAI21_X1   g06875(.A1(new_n7876_), .A2(new_n7877_), .B(new_n5061_), .ZN(new_n7878_));
  NAND2_X1   g06876(.A1(new_n7878_), .A2(new_n7875_), .ZN(new_n7879_));
  NAND4_X1   g06877(.A1(new_n7879_), .A2(new_n4999_), .A3(new_n5010_), .A4(new_n5072_), .ZN(new_n7880_));
  NOR2_X1    g06878(.A1(new_n5055_), .A2(new_n5058_), .ZN(new_n7881_));
  AOI21_X1   g06879(.A1(new_n7873_), .A2(new_n7874_), .B(new_n5061_), .ZN(new_n7882_));
  NOR2_X1    g06880(.A1(new_n7882_), .A2(new_n7881_), .ZN(new_n7883_));
  OAI21_X1   g06881(.A1(new_n7883_), .A2(new_n5065_), .B(new_n5069_), .ZN(new_n7884_));
  NOR2_X1    g06882(.A1(new_n7880_), .A2(new_n7884_), .ZN(new_n7885_));
  OAI21_X1   g06883(.A1(new_n7881_), .A2(new_n7882_), .B(new_n5010_), .ZN(new_n7886_));
  NOR4_X1    g06884(.A1(new_n5051_), .A2(new_n5065_), .A3(new_n5062_), .A4(new_n5039_), .ZN(new_n7887_));
  AOI21_X1   g06885(.A1(new_n7879_), .A2(new_n7886_), .B(new_n7887_), .ZN(new_n7888_));
  OAI21_X1   g06886(.A1(new_n7885_), .A2(new_n7888_), .B(new_n7872_), .ZN(new_n7889_));
  AOI21_X1   g06887(.A1(new_n7868_), .A2(new_n7869_), .B(new_n5038_), .ZN(new_n7890_));
  NOR2_X1    g06888(.A1(new_n7890_), .A2(new_n7864_), .ZN(new_n7891_));
  OAI22_X1   g06889(.A1(new_n7891_), .A2(new_n5051_), .B1(new_n7867_), .B2(new_n7870_), .ZN(new_n7892_));
  NOR3_X1    g06890(.A1(new_n7876_), .A2(new_n7877_), .A3(new_n5061_), .ZN(new_n7893_));
  AOI21_X1   g06891(.A1(new_n7873_), .A2(new_n7874_), .B(new_n4998_), .ZN(new_n7894_));
  NOR2_X1    g06892(.A1(new_n7893_), .A2(new_n7894_), .ZN(new_n7895_));
  INV_X1     g06893(.I(new_n7881_), .ZN(new_n7896_));
  OAI21_X1   g06894(.A1(new_n7876_), .A2(new_n7877_), .B(new_n4998_), .ZN(new_n7897_));
  AOI21_X1   g06895(.A1(new_n7896_), .A2(new_n7897_), .B(new_n5065_), .ZN(new_n7898_));
  NOR3_X1    g06896(.A1(new_n7887_), .A2(new_n7898_), .A3(new_n7895_), .ZN(new_n7899_));
  NAND4_X1   g06897(.A1(new_n5072_), .A2(new_n5010_), .A3(new_n4999_), .A4(new_n5069_), .ZN(new_n7900_));
  AOI21_X1   g06898(.A1(new_n7879_), .A2(new_n7886_), .B(new_n7900_), .ZN(new_n7901_));
  OAI21_X1   g06899(.A1(new_n7901_), .A2(new_n7899_), .B(new_n7892_), .ZN(new_n7902_));
  OAI22_X1   g06900(.A1(new_n5173_), .A2(new_n5174_), .B1(new_n5074_), .B2(new_n5053_), .ZN(new_n7903_));
  NAND3_X1   g06901(.A1(new_n7889_), .A2(new_n7902_), .A3(new_n7903_), .ZN(new_n7904_));
  NOR2_X1    g06902(.A1(new_n5051_), .A2(new_n5065_), .ZN(new_n7905_));
  NAND2_X1   g06903(.A1(new_n7897_), .A2(new_n7896_), .ZN(new_n7906_));
  AOI21_X1   g06904(.A1(new_n7906_), .A2(new_n5010_), .B(new_n5039_), .ZN(new_n7907_));
  NAND4_X1   g06905(.A1(new_n7907_), .A2(new_n7883_), .A3(new_n7879_), .A4(new_n7905_), .ZN(new_n7908_));
  OAI21_X1   g06906(.A1(new_n7895_), .A2(new_n7898_), .B(new_n7900_), .ZN(new_n7909_));
  AOI21_X1   g06907(.A1(new_n7908_), .A2(new_n7909_), .B(new_n7892_), .ZN(new_n7910_));
  NAND3_X1   g06908(.A1(new_n7900_), .A2(new_n7886_), .A3(new_n7879_), .ZN(new_n7911_));
  NAND2_X1   g06909(.A1(new_n7886_), .A2(new_n7879_), .ZN(new_n7912_));
  NAND2_X1   g06910(.A1(new_n7912_), .A2(new_n7887_), .ZN(new_n7913_));
  AOI21_X1   g06911(.A1(new_n7913_), .A2(new_n7911_), .B(new_n7872_), .ZN(new_n7914_));
  AOI22_X1   g06912(.A1(new_n5151_), .A2(new_n5167_), .B1(new_n5170_), .B2(new_n5171_), .ZN(new_n7915_));
  OAI21_X1   g06913(.A1(new_n7910_), .A2(new_n7914_), .B(new_n7915_), .ZN(new_n7916_));
  AOI21_X1   g06914(.A1(new_n7916_), .A2(new_n7904_), .B(new_n7860_), .ZN(new_n7917_));
  NOR3_X1    g06915(.A1(new_n7843_), .A2(new_n7841_), .A3(new_n7846_), .ZN(new_n7918_));
  NOR2_X1    g06916(.A1(new_n7846_), .A2(new_n7841_), .ZN(new_n7919_));
  NOR2_X1    g06917(.A1(new_n7919_), .A2(new_n7834_), .ZN(new_n7920_));
  OAI21_X1   g06918(.A1(new_n7920_), .A2(new_n7918_), .B(new_n7853_), .ZN(new_n7921_));
  NAND3_X1   g06919(.A1(new_n7832_), .A2(new_n5104_), .A3(new_n7833_), .ZN(new_n7922_));
  NOR2_X1    g06920(.A1(new_n7836_), .A2(new_n7835_), .ZN(new_n7923_));
  OAI21_X1   g06921(.A1(new_n7923_), .A2(new_n5161_), .B(new_n5137_), .ZN(new_n7924_));
  NOR2_X1    g06922(.A1(new_n7922_), .A2(new_n7924_), .ZN(new_n7925_));
  NOR2_X1    g06923(.A1(new_n7919_), .A2(new_n7843_), .ZN(new_n7926_));
  OAI21_X1   g06924(.A1(new_n7926_), .A2(new_n7925_), .B(new_n7825_), .ZN(new_n7927_));
  NAND2_X1   g06925(.A1(new_n7927_), .A2(new_n7921_), .ZN(new_n7928_));
  NAND3_X1   g06926(.A1(new_n7889_), .A2(new_n7902_), .A3(new_n7915_), .ZN(new_n7929_));
  OAI21_X1   g06927(.A1(new_n7910_), .A2(new_n7914_), .B(new_n7903_), .ZN(new_n7930_));
  AOI21_X1   g06928(.A1(new_n7930_), .A2(new_n7929_), .B(new_n7928_), .ZN(new_n7931_));
  AOI21_X1   g06929(.A1(new_n5366_), .A2(new_n5368_), .B(new_n5177_), .ZN(new_n7932_));
  NOR3_X1    g06930(.A1(new_n7931_), .A2(new_n7917_), .A3(new_n7932_), .ZN(new_n7933_));
  NOR3_X1    g06931(.A1(new_n7910_), .A2(new_n7914_), .A3(new_n7915_), .ZN(new_n7934_));
  AOI21_X1   g06932(.A1(new_n7889_), .A2(new_n7902_), .B(new_n7903_), .ZN(new_n7935_));
  OAI21_X1   g06933(.A1(new_n7934_), .A2(new_n7935_), .B(new_n7928_), .ZN(new_n7936_));
  NOR3_X1    g06934(.A1(new_n7910_), .A2(new_n7914_), .A3(new_n7903_), .ZN(new_n7937_));
  AOI21_X1   g06935(.A1(new_n7889_), .A2(new_n7902_), .B(new_n7915_), .ZN(new_n7938_));
  OAI21_X1   g06936(.A1(new_n7937_), .A2(new_n7938_), .B(new_n7860_), .ZN(new_n7939_));
  NAND2_X1   g06937(.A1(new_n5175_), .A2(new_n5172_), .ZN(new_n7940_));
  NAND2_X1   g06938(.A1(new_n5168_), .A2(new_n5075_), .ZN(new_n7941_));
  NAND2_X1   g06939(.A1(new_n7941_), .A2(new_n7940_), .ZN(new_n7942_));
  NAND2_X1   g06940(.A1(new_n5369_), .A2(new_n7942_), .ZN(new_n7943_));
  AOI21_X1   g06941(.A1(new_n7936_), .A2(new_n7939_), .B(new_n7943_), .ZN(new_n7944_));
  OAI21_X1   g06942(.A1(new_n7933_), .A2(new_n7944_), .B(new_n7808_), .ZN(new_n7945_));
  INV_X1     g06943(.I(new_n7945_), .ZN(new_n7946_));
  NAND3_X1   g06944(.A1(new_n7789_), .A2(new_n7786_), .A3(new_n7790_), .ZN(new_n7947_));
  OAI21_X1   g06945(.A1(new_n7766_), .A2(new_n7776_), .B(new_n7777_), .ZN(new_n7948_));
  AOI21_X1   g06946(.A1(new_n7948_), .A2(new_n7947_), .B(new_n7804_), .ZN(new_n7949_));
  NAND3_X1   g06947(.A1(new_n7786_), .A2(new_n7789_), .A3(new_n7777_), .ZN(new_n7950_));
  OAI21_X1   g06948(.A1(new_n7766_), .A2(new_n7776_), .B(new_n7790_), .ZN(new_n7951_));
  AOI21_X1   g06949(.A1(new_n7950_), .A2(new_n7951_), .B(new_n7726_), .ZN(new_n7952_));
  NOR2_X1    g06950(.A1(new_n7952_), .A2(new_n7949_), .ZN(new_n7953_));
  NOR3_X1    g06951(.A1(new_n7931_), .A2(new_n7917_), .A3(new_n7943_), .ZN(new_n7954_));
  AOI21_X1   g06952(.A1(new_n7936_), .A2(new_n7939_), .B(new_n7932_), .ZN(new_n7955_));
  OAI21_X1   g06953(.A1(new_n7954_), .A2(new_n7955_), .B(new_n7953_), .ZN(new_n7956_));
  INV_X1     g06954(.I(new_n7956_), .ZN(new_n7957_));
  INV_X1     g06955(.I(new_n5370_), .ZN(new_n7958_));
  NAND2_X1   g06956(.A1(new_n7958_), .A2(new_n5750_), .ZN(new_n7959_));
  NOR3_X1    g06957(.A1(new_n7957_), .A2(new_n7946_), .A3(new_n7959_), .ZN(new_n7960_));
  INV_X1     g06958(.I(new_n7959_), .ZN(new_n7961_));
  AOI21_X1   g06959(.A1(new_n7945_), .A2(new_n7956_), .B(new_n7961_), .ZN(new_n7962_));
  OAI21_X1   g06960(.A1(new_n7962_), .A2(new_n7960_), .B(new_n7676_), .ZN(new_n7963_));
  NAND3_X1   g06961(.A1(new_n7956_), .A2(new_n7945_), .A3(new_n7959_), .ZN(new_n7964_));
  NAND2_X1   g06962(.A1(new_n7956_), .A2(new_n7945_), .ZN(new_n7965_));
  NAND2_X1   g06963(.A1(new_n7965_), .A2(new_n7961_), .ZN(new_n7966_));
  NAND2_X1   g06964(.A1(new_n7966_), .A2(new_n7964_), .ZN(new_n7967_));
  NAND2_X1   g06965(.A1(new_n7967_), .A2(new_n7675_), .ZN(new_n7968_));
  NAND2_X1   g06966(.A1(new_n7968_), .A2(new_n7963_), .ZN(new_n7969_));
  INV_X1     g06967(.I(new_n7969_), .ZN(new_n7970_));
  NOR2_X1    g06968(.A1(new_n4540_), .A2(new_n4548_), .ZN(new_n7971_));
  NOR2_X1    g06969(.A1(new_n4536_), .A2(new_n4550_), .ZN(new_n7972_));
  OAI21_X1   g06970(.A1(new_n7972_), .A2(new_n7971_), .B(new_n4541_), .ZN(new_n7973_));
  NOR2_X1    g06971(.A1(new_n4550_), .A2(new_n4548_), .ZN(new_n7974_));
  INV_X1     g06972(.I(new_n7974_), .ZN(new_n7975_));
  NAND2_X1   g06973(.A1(new_n7973_), .A2(new_n7975_), .ZN(new_n7976_));
  NAND2_X1   g06974(.A1(new_n4536_), .A2(new_n4550_), .ZN(new_n7977_));
  NAND2_X1   g06975(.A1(new_n4540_), .A2(new_n4548_), .ZN(new_n7978_));
  NAND3_X1   g06976(.A1(new_n7977_), .A2(new_n7978_), .A3(new_n4541_), .ZN(new_n7979_));
  OAI21_X1   g06977(.A1(new_n7972_), .A2(new_n7971_), .B(new_n4554_), .ZN(new_n7980_));
  AOI22_X1   g06978(.A1(new_n7976_), .A2(new_n4532_), .B1(new_n7979_), .B2(new_n7980_), .ZN(new_n7981_));
  NAND2_X1   g06979(.A1(new_n4489_), .A2(new_n4492_), .ZN(new_n7982_));
  NAND2_X1   g06980(.A1(new_n4484_), .A2(new_n4474_), .ZN(new_n7983_));
  NAND2_X1   g06981(.A1(new_n7983_), .A2(new_n7982_), .ZN(new_n7984_));
  NOR2_X1    g06982(.A1(new_n4477_), .A2(new_n4479_), .ZN(new_n7985_));
  INV_X1     g06983(.I(new_n4496_), .ZN(new_n7986_));
  OAI21_X1   g06984(.A1(new_n7985_), .A2(new_n4475_), .B(new_n7986_), .ZN(new_n7987_));
  NAND2_X1   g06985(.A1(new_n7987_), .A2(new_n4500_), .ZN(new_n7988_));
  NOR2_X1    g06986(.A1(new_n4471_), .A2(new_n4472_), .ZN(new_n7989_));
  INV_X1     g06987(.I(new_n4499_), .ZN(new_n7990_));
  OAI21_X1   g06988(.A1(new_n7989_), .A2(new_n4468_), .B(new_n7990_), .ZN(new_n7991_));
  NAND2_X1   g06989(.A1(new_n7991_), .A2(new_n4497_), .ZN(new_n7992_));
  AOI22_X1   g06990(.A1(new_n4470_), .A2(new_n4473_), .B1(new_n4491_), .B2(new_n4490_), .ZN(new_n7993_));
  NAND3_X1   g06991(.A1(new_n7988_), .A2(new_n7992_), .A3(new_n7993_), .ZN(new_n7994_));
  NOR2_X1    g06992(.A1(new_n7991_), .A2(new_n4497_), .ZN(new_n7995_));
  NOR2_X1    g06993(.A1(new_n7987_), .A2(new_n4500_), .ZN(new_n7996_));
  OAI21_X1   g06994(.A1(new_n7995_), .A2(new_n7996_), .B(new_n4501_), .ZN(new_n7997_));
  NAND2_X1   g06995(.A1(new_n7997_), .A2(new_n7994_), .ZN(new_n7998_));
  NAND3_X1   g06996(.A1(new_n7993_), .A2(new_n7987_), .A3(new_n7991_), .ZN(new_n7999_));
  NAND4_X1   g06997(.A1(new_n7998_), .A2(new_n7984_), .A3(new_n7999_), .A4(new_n4532_), .ZN(new_n8000_));
  AOI21_X1   g06998(.A1(new_n7988_), .A2(new_n7992_), .B(new_n4501_), .ZN(new_n8001_));
  NOR2_X1    g06999(.A1(new_n4497_), .A2(new_n4500_), .ZN(new_n8002_));
  OAI21_X1   g07000(.A1(new_n8001_), .A2(new_n8002_), .B(new_n7984_), .ZN(new_n8003_));
  NAND2_X1   g07001(.A1(new_n8003_), .A2(new_n4542_), .ZN(new_n8004_));
  NOR2_X1    g07002(.A1(new_n8000_), .A2(new_n8004_), .ZN(new_n8005_));
  NOR4_X1    g07003(.A1(new_n4494_), .A2(new_n4547_), .A3(new_n4502_), .A4(new_n4555_), .ZN(new_n8006_));
  AOI21_X1   g07004(.A1(new_n7998_), .A2(new_n8003_), .B(new_n8006_), .ZN(new_n8007_));
  OAI21_X1   g07005(.A1(new_n8005_), .A2(new_n8007_), .B(new_n7981_), .ZN(new_n8008_));
  NAND2_X1   g07006(.A1(new_n7977_), .A2(new_n7978_), .ZN(new_n8009_));
  AOI21_X1   g07007(.A1(new_n8009_), .A2(new_n4541_), .B(new_n7974_), .ZN(new_n8010_));
  NAND2_X1   g07008(.A1(new_n7980_), .A2(new_n7979_), .ZN(new_n8011_));
  OAI21_X1   g07009(.A1(new_n4547_), .A2(new_n8010_), .B(new_n8011_), .ZN(new_n8012_));
  NAND4_X1   g07010(.A1(new_n7984_), .A2(new_n4532_), .A3(new_n7999_), .A4(new_n4542_), .ZN(new_n8013_));
  NAND3_X1   g07011(.A1(new_n8003_), .A2(new_n8013_), .A3(new_n7998_), .ZN(new_n8014_));
  INV_X1     g07012(.I(new_n8014_), .ZN(new_n8015_));
  AOI21_X1   g07013(.A1(new_n8003_), .A2(new_n7998_), .B(new_n8013_), .ZN(new_n8016_));
  OAI21_X1   g07014(.A1(new_n8015_), .A2(new_n8016_), .B(new_n8012_), .ZN(new_n8017_));
  NAND2_X1   g07015(.A1(new_n8008_), .A2(new_n8017_), .ZN(new_n8018_));
  NOR2_X1    g07016(.A1(new_n4429_), .A2(new_n4430_), .ZN(new_n8019_));
  INV_X1     g07017(.I(new_n4439_), .ZN(new_n8020_));
  OAI21_X1   g07018(.A1(new_n8019_), .A2(new_n4410_), .B(new_n8020_), .ZN(new_n8021_));
  NOR2_X1    g07019(.A1(new_n8021_), .A2(new_n4438_), .ZN(new_n8022_));
  NOR2_X1    g07020(.A1(new_n4423_), .A2(new_n4424_), .ZN(new_n8023_));
  INV_X1     g07021(.I(new_n4437_), .ZN(new_n8024_));
  OAI21_X1   g07022(.A1(new_n8023_), .A2(new_n4420_), .B(new_n8024_), .ZN(new_n8025_));
  NOR2_X1    g07023(.A1(new_n8025_), .A2(new_n4440_), .ZN(new_n8026_));
  AOI22_X1   g07024(.A1(new_n4428_), .A2(new_n4431_), .B1(new_n4422_), .B2(new_n4425_), .ZN(new_n8027_));
  OAI21_X1   g07025(.A1(new_n8022_), .A2(new_n8026_), .B(new_n8027_), .ZN(new_n8028_));
  NOR2_X1    g07026(.A1(new_n4438_), .A2(new_n4440_), .ZN(new_n8029_));
  INV_X1     g07027(.I(new_n8029_), .ZN(new_n8030_));
  NAND2_X1   g07028(.A1(new_n8028_), .A2(new_n8030_), .ZN(new_n8031_));
  NAND2_X1   g07029(.A1(new_n8025_), .A2(new_n4440_), .ZN(new_n8032_));
  NAND2_X1   g07030(.A1(new_n8021_), .A2(new_n4438_), .ZN(new_n8033_));
  NAND3_X1   g07031(.A1(new_n8032_), .A2(new_n8033_), .A3(new_n8027_), .ZN(new_n8034_));
  OAI22_X1   g07032(.A1(new_n8022_), .A2(new_n8026_), .B1(new_n4416_), .B2(new_n4434_), .ZN(new_n8035_));
  AOI22_X1   g07033(.A1(new_n8031_), .A2(new_n4436_), .B1(new_n8034_), .B2(new_n8035_), .ZN(new_n8036_));
  NAND2_X1   g07034(.A1(new_n4453_), .A2(new_n4398_), .ZN(new_n8037_));
  NAND2_X1   g07035(.A1(new_n4455_), .A2(new_n4394_), .ZN(new_n8038_));
  NAND3_X1   g07036(.A1(new_n8037_), .A2(new_n8038_), .A3(new_n4456_), .ZN(new_n8039_));
  NOR2_X1    g07037(.A1(new_n4455_), .A2(new_n4394_), .ZN(new_n8040_));
  NOR2_X1    g07038(.A1(new_n4453_), .A2(new_n4398_), .ZN(new_n8041_));
  OAI21_X1   g07039(.A1(new_n8040_), .A2(new_n8041_), .B(new_n4407_), .ZN(new_n8042_));
  NAND2_X1   g07040(.A1(new_n8042_), .A2(new_n8039_), .ZN(new_n8043_));
  NAND4_X1   g07041(.A1(new_n8043_), .A2(new_n4451_), .A3(new_n4457_), .A4(new_n4436_), .ZN(new_n8044_));
  AOI21_X1   g07042(.A1(new_n8037_), .A2(new_n8038_), .B(new_n4407_), .ZN(new_n8045_));
  NOR2_X1    g07043(.A1(new_n4394_), .A2(new_n4398_), .ZN(new_n8046_));
  OAI21_X1   g07044(.A1(new_n8045_), .A2(new_n8046_), .B(new_n4451_), .ZN(new_n8047_));
  NAND2_X1   g07045(.A1(new_n8047_), .A2(new_n4442_), .ZN(new_n8048_));
  NOR2_X1    g07046(.A1(new_n8044_), .A2(new_n8048_), .ZN(new_n8049_));
  NOR4_X1    g07047(.A1(new_n4391_), .A2(new_n4461_), .A3(new_n4408_), .A4(new_n4441_), .ZN(new_n8050_));
  AOI21_X1   g07048(.A1(new_n8043_), .A2(new_n8047_), .B(new_n8050_), .ZN(new_n8051_));
  OAI21_X1   g07049(.A1(new_n8049_), .A2(new_n8051_), .B(new_n8036_), .ZN(new_n8052_));
  NAND2_X1   g07050(.A1(new_n8032_), .A2(new_n8033_), .ZN(new_n8053_));
  AOI21_X1   g07051(.A1(new_n8053_), .A2(new_n8027_), .B(new_n8029_), .ZN(new_n8054_));
  NOR4_X1    g07052(.A1(new_n8022_), .A2(new_n8026_), .A3(new_n4416_), .A4(new_n4434_), .ZN(new_n8055_));
  AOI21_X1   g07053(.A1(new_n8032_), .A2(new_n8033_), .B(new_n8027_), .ZN(new_n8056_));
  OAI22_X1   g07054(.A1(new_n8054_), .A2(new_n4461_), .B1(new_n8055_), .B2(new_n8056_), .ZN(new_n8057_));
  NAND4_X1   g07055(.A1(new_n4451_), .A2(new_n4436_), .A3(new_n4442_), .A4(new_n4457_), .ZN(new_n8058_));
  AOI21_X1   g07056(.A1(new_n8043_), .A2(new_n8047_), .B(new_n8058_), .ZN(new_n8059_));
  NOR3_X1    g07057(.A1(new_n8040_), .A2(new_n8041_), .A3(new_n4407_), .ZN(new_n8060_));
  AOI21_X1   g07058(.A1(new_n8037_), .A2(new_n8038_), .B(new_n4456_), .ZN(new_n8061_));
  NOR2_X1    g07059(.A1(new_n8061_), .A2(new_n8060_), .ZN(new_n8062_));
  OAI21_X1   g07060(.A1(new_n8040_), .A2(new_n8041_), .B(new_n4456_), .ZN(new_n8063_));
  INV_X1     g07061(.I(new_n8046_), .ZN(new_n8064_));
  AOI21_X1   g07062(.A1(new_n8063_), .A2(new_n8064_), .B(new_n4391_), .ZN(new_n8065_));
  NOR3_X1    g07063(.A1(new_n8065_), .A2(new_n8050_), .A3(new_n8062_), .ZN(new_n8066_));
  OAI21_X1   g07064(.A1(new_n8066_), .A2(new_n8059_), .B(new_n8057_), .ZN(new_n8067_));
  NOR2_X1    g07065(.A1(new_n4464_), .A2(new_n4559_), .ZN(new_n8068_));
  NAND3_X1   g07066(.A1(new_n8052_), .A2(new_n8068_), .A3(new_n8067_), .ZN(new_n8069_));
  NAND2_X1   g07067(.A1(new_n8063_), .A2(new_n8064_), .ZN(new_n8070_));
  NOR4_X1    g07068(.A1(new_n8062_), .A2(new_n8070_), .A3(new_n4391_), .A4(new_n4461_), .ZN(new_n8071_));
  AOI21_X1   g07069(.A1(new_n8070_), .A2(new_n4451_), .B(new_n4441_), .ZN(new_n8072_));
  NAND2_X1   g07070(.A1(new_n8071_), .A2(new_n8072_), .ZN(new_n8073_));
  NAND2_X1   g07071(.A1(new_n8047_), .A2(new_n8043_), .ZN(new_n8074_));
  NAND2_X1   g07072(.A1(new_n8074_), .A2(new_n8058_), .ZN(new_n8075_));
  AOI21_X1   g07073(.A1(new_n8073_), .A2(new_n8075_), .B(new_n8057_), .ZN(new_n8076_));
  NAND2_X1   g07074(.A1(new_n8074_), .A2(new_n8050_), .ZN(new_n8077_));
  NAND3_X1   g07075(.A1(new_n8058_), .A2(new_n8047_), .A3(new_n8043_), .ZN(new_n8078_));
  AOI21_X1   g07076(.A1(new_n8077_), .A2(new_n8078_), .B(new_n8036_), .ZN(new_n8079_));
  OAI22_X1   g07077(.A1(new_n4444_), .A2(new_n4463_), .B1(new_n4557_), .B2(new_n4544_), .ZN(new_n8080_));
  OAI21_X1   g07078(.A1(new_n8076_), .A2(new_n8079_), .B(new_n8080_), .ZN(new_n8081_));
  AOI21_X1   g07079(.A1(new_n8081_), .A2(new_n8069_), .B(new_n8018_), .ZN(new_n8082_));
  OAI21_X1   g07080(.A1(new_n7995_), .A2(new_n7996_), .B(new_n7993_), .ZN(new_n8083_));
  INV_X1     g07081(.I(new_n8002_), .ZN(new_n8084_));
  NAND2_X1   g07082(.A1(new_n8083_), .A2(new_n8084_), .ZN(new_n8085_));
  NOR3_X1    g07083(.A1(new_n7995_), .A2(new_n7996_), .A3(new_n4501_), .ZN(new_n8086_));
  AOI21_X1   g07084(.A1(new_n7988_), .A2(new_n7992_), .B(new_n7993_), .ZN(new_n8087_));
  NOR2_X1    g07085(.A1(new_n8087_), .A2(new_n8086_), .ZN(new_n8088_));
  NOR4_X1    g07086(.A1(new_n8088_), .A2(new_n8085_), .A3(new_n4494_), .A4(new_n4547_), .ZN(new_n8089_));
  AOI21_X1   g07087(.A1(new_n8083_), .A2(new_n8084_), .B(new_n4494_), .ZN(new_n8090_));
  NOR2_X1    g07088(.A1(new_n8090_), .A2(new_n4555_), .ZN(new_n8091_));
  NAND2_X1   g07089(.A1(new_n8089_), .A2(new_n8091_), .ZN(new_n8092_));
  NAND2_X1   g07090(.A1(new_n8003_), .A2(new_n7998_), .ZN(new_n8093_));
  NAND2_X1   g07091(.A1(new_n8093_), .A2(new_n8013_), .ZN(new_n8094_));
  AOI21_X1   g07092(.A1(new_n8092_), .A2(new_n8094_), .B(new_n8012_), .ZN(new_n8095_));
  INV_X1     g07093(.I(new_n8016_), .ZN(new_n8096_));
  AOI21_X1   g07094(.A1(new_n8096_), .A2(new_n8014_), .B(new_n7981_), .ZN(new_n8097_));
  NOR2_X1    g07095(.A1(new_n8095_), .A2(new_n8097_), .ZN(new_n8098_));
  NAND3_X1   g07096(.A1(new_n8052_), .A2(new_n8067_), .A3(new_n8080_), .ZN(new_n8099_));
  OAI21_X1   g07097(.A1(new_n8076_), .A2(new_n8079_), .B(new_n8068_), .ZN(new_n8100_));
  AOI21_X1   g07098(.A1(new_n8099_), .A2(new_n8100_), .B(new_n8098_), .ZN(new_n8101_));
  NOR2_X1    g07099(.A1(new_n8101_), .A2(new_n8082_), .ZN(new_n8102_));
  AOI22_X1   g07100(.A1(new_n4558_), .A2(new_n4560_), .B1(new_n4372_), .B2(new_n4358_), .ZN(new_n8103_));
  NAND2_X1   g07101(.A1(new_n4339_), .A2(new_n4336_), .ZN(new_n8104_));
  NAND2_X1   g07102(.A1(new_n4324_), .A2(new_n4334_), .ZN(new_n8105_));
  NAND2_X1   g07103(.A1(new_n8105_), .A2(new_n8104_), .ZN(new_n8106_));
  NOR2_X1    g07104(.A1(new_n4347_), .A2(new_n4350_), .ZN(new_n8107_));
  INV_X1     g07105(.I(new_n4345_), .ZN(new_n8108_));
  OAI21_X1   g07106(.A1(new_n8107_), .A2(new_n4316_), .B(new_n8108_), .ZN(new_n8109_));
  NOR2_X1    g07107(.A1(new_n8109_), .A2(new_n4344_), .ZN(new_n8110_));
  NOR2_X1    g07108(.A1(new_n4331_), .A2(new_n4332_), .ZN(new_n8111_));
  INV_X1     g07109(.I(new_n4343_), .ZN(new_n8112_));
  OAI21_X1   g07110(.A1(new_n8111_), .A2(new_n4330_), .B(new_n8112_), .ZN(new_n8113_));
  NOR2_X1    g07111(.A1(new_n8113_), .A2(new_n4346_), .ZN(new_n8114_));
  AOI22_X1   g07112(.A1(new_n4318_), .A2(new_n4323_), .B1(new_n4337_), .B2(new_n4338_), .ZN(new_n8115_));
  OAI21_X1   g07113(.A1(new_n8110_), .A2(new_n8114_), .B(new_n8115_), .ZN(new_n8116_));
  NOR2_X1    g07114(.A1(new_n4344_), .A2(new_n4346_), .ZN(new_n8117_));
  INV_X1     g07115(.I(new_n8117_), .ZN(new_n8118_));
  NAND2_X1   g07116(.A1(new_n8116_), .A2(new_n8118_), .ZN(new_n8119_));
  NAND2_X1   g07117(.A1(new_n8113_), .A2(new_n4346_), .ZN(new_n8120_));
  NAND2_X1   g07118(.A1(new_n8109_), .A2(new_n4344_), .ZN(new_n8121_));
  NAND3_X1   g07119(.A1(new_n8121_), .A2(new_n8120_), .A3(new_n8115_), .ZN(new_n8122_));
  OAI21_X1   g07120(.A1(new_n8110_), .A2(new_n8114_), .B(new_n4352_), .ZN(new_n8123_));
  AOI22_X1   g07121(.A1(new_n8119_), .A2(new_n8106_), .B1(new_n8122_), .B2(new_n8123_), .ZN(new_n8124_));
  NOR2_X1    g07122(.A1(new_n4290_), .A2(new_n4363_), .ZN(new_n8125_));
  NOR2_X1    g07123(.A1(new_n4281_), .A2(new_n4364_), .ZN(new_n8126_));
  OAI21_X1   g07124(.A1(new_n8125_), .A2(new_n8126_), .B(new_n4365_), .ZN(new_n8127_));
  NAND2_X1   g07125(.A1(new_n4281_), .A2(new_n4364_), .ZN(new_n8128_));
  NAND2_X1   g07126(.A1(new_n4290_), .A2(new_n4363_), .ZN(new_n8129_));
  NAND3_X1   g07127(.A1(new_n8128_), .A2(new_n8129_), .A3(new_n4300_), .ZN(new_n8130_));
  NAND2_X1   g07128(.A1(new_n8127_), .A2(new_n8130_), .ZN(new_n8131_));
  NAND3_X1   g07129(.A1(new_n8115_), .A2(new_n8113_), .A3(new_n8109_), .ZN(new_n8132_));
  AOI22_X1   g07130(.A1(new_n8105_), .A2(new_n8104_), .B1(new_n4313_), .B2(new_n4307_), .ZN(new_n8133_));
  NAND3_X1   g07131(.A1(new_n8133_), .A2(new_n4301_), .A3(new_n8132_), .ZN(new_n8134_));
  NOR2_X1    g07132(.A1(new_n4363_), .A2(new_n4364_), .ZN(new_n8135_));
  AOI21_X1   g07133(.A1(new_n8128_), .A2(new_n8129_), .B(new_n4365_), .ZN(new_n8136_));
  OAI21_X1   g07134(.A1(new_n8135_), .A2(new_n8136_), .B(new_n4314_), .ZN(new_n8137_));
  NAND3_X1   g07135(.A1(new_n8134_), .A2(new_n8137_), .A3(new_n8131_), .ZN(new_n8138_));
  NOR4_X1    g07136(.A1(new_n4341_), .A2(new_n4369_), .A3(new_n4353_), .A4(new_n4366_), .ZN(new_n8139_));
  NAND2_X1   g07137(.A1(new_n8137_), .A2(new_n8131_), .ZN(new_n8140_));
  NAND2_X1   g07138(.A1(new_n8140_), .A2(new_n8139_), .ZN(new_n8141_));
  AOI21_X1   g07139(.A1(new_n8141_), .A2(new_n8138_), .B(new_n8124_), .ZN(new_n8142_));
  NAND2_X1   g07140(.A1(new_n8121_), .A2(new_n8120_), .ZN(new_n8143_));
  AOI21_X1   g07141(.A1(new_n8143_), .A2(new_n8115_), .B(new_n8117_), .ZN(new_n8144_));
  NOR3_X1    g07142(.A1(new_n8110_), .A2(new_n8114_), .A3(new_n4352_), .ZN(new_n8145_));
  AOI21_X1   g07143(.A1(new_n8121_), .A2(new_n8120_), .B(new_n8115_), .ZN(new_n8146_));
  OAI22_X1   g07144(.A1(new_n8144_), .A2(new_n4341_), .B1(new_n8145_), .B2(new_n8146_), .ZN(new_n8147_));
  INV_X1     g07145(.I(new_n8135_), .ZN(new_n8148_));
  OAI21_X1   g07146(.A1(new_n8125_), .A2(new_n8126_), .B(new_n4300_), .ZN(new_n8149_));
  NAND2_X1   g07147(.A1(new_n8149_), .A2(new_n8148_), .ZN(new_n8150_));
  AOI21_X1   g07148(.A1(new_n8128_), .A2(new_n8129_), .B(new_n4300_), .ZN(new_n8151_));
  NOR3_X1    g07149(.A1(new_n8125_), .A2(new_n8126_), .A3(new_n4365_), .ZN(new_n8152_));
  NOR2_X1    g07150(.A1(new_n8151_), .A2(new_n8152_), .ZN(new_n8153_));
  NOR4_X1    g07151(.A1(new_n8153_), .A2(new_n8150_), .A3(new_n4369_), .A4(new_n4341_), .ZN(new_n8154_));
  AOI21_X1   g07152(.A1(new_n8150_), .A2(new_n4314_), .B(new_n4353_), .ZN(new_n8155_));
  NAND2_X1   g07153(.A1(new_n8154_), .A2(new_n8155_), .ZN(new_n8156_));
  NAND2_X1   g07154(.A1(new_n8140_), .A2(new_n8134_), .ZN(new_n8157_));
  AOI21_X1   g07155(.A1(new_n8156_), .A2(new_n8157_), .B(new_n8147_), .ZN(new_n8158_));
  NOR2_X1    g07156(.A1(new_n8158_), .A2(new_n8142_), .ZN(new_n8159_));
  NAND2_X1   g07157(.A1(new_n4266_), .A2(new_n4242_), .ZN(new_n8160_));
  NAND2_X1   g07158(.A1(new_n4268_), .A2(new_n4238_), .ZN(new_n8161_));
  AOI21_X1   g07159(.A1(new_n8160_), .A2(new_n8161_), .B(new_n4246_), .ZN(new_n8162_));
  NOR2_X1    g07160(.A1(new_n4242_), .A2(new_n4238_), .ZN(new_n8163_));
  NOR2_X1    g07161(.A1(new_n8162_), .A2(new_n8163_), .ZN(new_n8164_));
  NOR2_X1    g07162(.A1(new_n4268_), .A2(new_n4238_), .ZN(new_n8165_));
  NOR2_X1    g07163(.A1(new_n4266_), .A2(new_n4242_), .ZN(new_n8166_));
  NOR3_X1    g07164(.A1(new_n8166_), .A2(new_n8165_), .A3(new_n4246_), .ZN(new_n8167_));
  AOI22_X1   g07165(.A1(new_n8160_), .A2(new_n8161_), .B1(new_n4216_), .B2(new_n4234_), .ZN(new_n8168_));
  OAI22_X1   g07166(.A1(new_n8164_), .A2(new_n4236_), .B1(new_n8167_), .B2(new_n8168_), .ZN(new_n8169_));
  NAND2_X1   g07167(.A1(new_n4175_), .A2(new_n4255_), .ZN(new_n8170_));
  NAND2_X1   g07168(.A1(new_n4179_), .A2(new_n4252_), .ZN(new_n8171_));
  AOI21_X1   g07169(.A1(new_n8170_), .A2(new_n8171_), .B(new_n4196_), .ZN(new_n8172_));
  NOR2_X1    g07170(.A1(new_n4179_), .A2(new_n4252_), .ZN(new_n8173_));
  NOR2_X1    g07171(.A1(new_n4175_), .A2(new_n4255_), .ZN(new_n8174_));
  NOR3_X1    g07172(.A1(new_n8173_), .A2(new_n8174_), .A3(new_n4256_), .ZN(new_n8175_));
  NOR2_X1    g07173(.A1(new_n8172_), .A2(new_n8175_), .ZN(new_n8176_));
  OAI22_X1   g07174(.A1(new_n4258_), .A2(new_n4259_), .B1(new_n4235_), .B2(new_n4224_), .ZN(new_n8177_));
  NOR3_X1    g07175(.A1(new_n8176_), .A2(new_n4257_), .A3(new_n8177_), .ZN(new_n8178_));
  NOR2_X1    g07176(.A1(new_n4252_), .A2(new_n4255_), .ZN(new_n8179_));
  INV_X1     g07177(.I(new_n8179_), .ZN(new_n8180_));
  OAI21_X1   g07178(.A1(new_n8173_), .A2(new_n8174_), .B(new_n4196_), .ZN(new_n8181_));
  NAND2_X1   g07179(.A1(new_n8181_), .A2(new_n8180_), .ZN(new_n8182_));
  AOI21_X1   g07180(.A1(new_n8182_), .A2(new_n4209_), .B(new_n4247_), .ZN(new_n8183_));
  NAND2_X1   g07181(.A1(new_n8178_), .A2(new_n8183_), .ZN(new_n8184_));
  AOI21_X1   g07182(.A1(new_n8180_), .A2(new_n8181_), .B(new_n4260_), .ZN(new_n8185_));
  NAND4_X1   g07183(.A1(new_n4209_), .A2(new_n4264_), .A3(new_n4197_), .A4(new_n4269_), .ZN(new_n8186_));
  OAI21_X1   g07184(.A1(new_n8185_), .A2(new_n8176_), .B(new_n8186_), .ZN(new_n8187_));
  AOI21_X1   g07185(.A1(new_n8184_), .A2(new_n8187_), .B(new_n8169_), .ZN(new_n8188_));
  NOR2_X1    g07186(.A1(new_n8166_), .A2(new_n8165_), .ZN(new_n8189_));
  INV_X1     g07187(.I(new_n8163_), .ZN(new_n8190_));
  OAI21_X1   g07188(.A1(new_n8189_), .A2(new_n4246_), .B(new_n8190_), .ZN(new_n8191_));
  NOR2_X1    g07189(.A1(new_n8168_), .A2(new_n8167_), .ZN(new_n8192_));
  AOI21_X1   g07190(.A1(new_n4264_), .A2(new_n8191_), .B(new_n8192_), .ZN(new_n8193_));
  OAI21_X1   g07191(.A1(new_n8173_), .A2(new_n8174_), .B(new_n4256_), .ZN(new_n8194_));
  NAND3_X1   g07192(.A1(new_n8170_), .A2(new_n8171_), .A3(new_n4196_), .ZN(new_n8195_));
  NAND2_X1   g07193(.A1(new_n8194_), .A2(new_n8195_), .ZN(new_n8196_));
  AOI21_X1   g07194(.A1(new_n8170_), .A2(new_n8171_), .B(new_n4256_), .ZN(new_n8197_));
  OAI21_X1   g07195(.A1(new_n8179_), .A2(new_n8197_), .B(new_n4209_), .ZN(new_n8198_));
  NAND3_X1   g07196(.A1(new_n8198_), .A2(new_n8186_), .A3(new_n8196_), .ZN(new_n8199_));
  NOR4_X1    g07197(.A1(new_n4260_), .A2(new_n4236_), .A3(new_n4257_), .A4(new_n4247_), .ZN(new_n8200_));
  NAND2_X1   g07198(.A1(new_n8198_), .A2(new_n8196_), .ZN(new_n8201_));
  NAND2_X1   g07199(.A1(new_n8201_), .A2(new_n8200_), .ZN(new_n8202_));
  AOI21_X1   g07200(.A1(new_n8202_), .A2(new_n8199_), .B(new_n8193_), .ZN(new_n8203_));
  OAI22_X1   g07201(.A1(new_n4355_), .A2(new_n4371_), .B1(new_n4360_), .B2(new_n4359_), .ZN(new_n8204_));
  NOR3_X1    g07202(.A1(new_n8203_), .A2(new_n8188_), .A3(new_n8204_), .ZN(new_n8205_));
  NAND4_X1   g07203(.A1(new_n8196_), .A2(new_n4197_), .A3(new_n4209_), .A4(new_n4264_), .ZN(new_n8206_));
  NOR2_X1    g07204(.A1(new_n8197_), .A2(new_n8179_), .ZN(new_n8207_));
  OAI21_X1   g07205(.A1(new_n8207_), .A2(new_n4260_), .B(new_n4269_), .ZN(new_n8208_));
  NOR2_X1    g07206(.A1(new_n8206_), .A2(new_n8208_), .ZN(new_n8209_));
  AOI21_X1   g07207(.A1(new_n8196_), .A2(new_n8198_), .B(new_n8200_), .ZN(new_n8210_));
  OAI21_X1   g07208(.A1(new_n8209_), .A2(new_n8210_), .B(new_n8193_), .ZN(new_n8211_));
  NOR3_X1    g07209(.A1(new_n8185_), .A2(new_n8200_), .A3(new_n8176_), .ZN(new_n8212_));
  AOI21_X1   g07210(.A1(new_n8196_), .A2(new_n8198_), .B(new_n8186_), .ZN(new_n8213_));
  OAI21_X1   g07211(.A1(new_n8213_), .A2(new_n8212_), .B(new_n8169_), .ZN(new_n8214_));
  AOI22_X1   g07212(.A1(new_n4356_), .A2(new_n4357_), .B1(new_n4249_), .B2(new_n4271_), .ZN(new_n8215_));
  AOI21_X1   g07213(.A1(new_n8211_), .A2(new_n8214_), .B(new_n8215_), .ZN(new_n8216_));
  OAI21_X1   g07214(.A1(new_n8205_), .A2(new_n8216_), .B(new_n8159_), .ZN(new_n8217_));
  AOI21_X1   g07215(.A1(new_n8148_), .A2(new_n8149_), .B(new_n4369_), .ZN(new_n8218_));
  NOR3_X1    g07216(.A1(new_n8139_), .A2(new_n8218_), .A3(new_n8153_), .ZN(new_n8219_));
  AOI21_X1   g07217(.A1(new_n8131_), .A2(new_n8137_), .B(new_n8134_), .ZN(new_n8220_));
  OAI21_X1   g07218(.A1(new_n8220_), .A2(new_n8219_), .B(new_n8147_), .ZN(new_n8221_));
  NAND3_X1   g07219(.A1(new_n8131_), .A2(new_n4301_), .A3(new_n8133_), .ZN(new_n8222_));
  NOR2_X1    g07220(.A1(new_n8136_), .A2(new_n8135_), .ZN(new_n8223_));
  OAI21_X1   g07221(.A1(new_n8223_), .A2(new_n4369_), .B(new_n8132_), .ZN(new_n8224_));
  NOR2_X1    g07222(.A1(new_n8222_), .A2(new_n8224_), .ZN(new_n8225_));
  AOI21_X1   g07223(.A1(new_n8131_), .A2(new_n8137_), .B(new_n8139_), .ZN(new_n8226_));
  OAI21_X1   g07224(.A1(new_n8225_), .A2(new_n8226_), .B(new_n8124_), .ZN(new_n8227_));
  NAND2_X1   g07225(.A1(new_n8227_), .A2(new_n8221_), .ZN(new_n8228_));
  NOR3_X1    g07226(.A1(new_n8203_), .A2(new_n8188_), .A3(new_n8215_), .ZN(new_n8229_));
  AOI21_X1   g07227(.A1(new_n8211_), .A2(new_n8214_), .B(new_n8204_), .ZN(new_n8230_));
  OAI21_X1   g07228(.A1(new_n8229_), .A2(new_n8230_), .B(new_n8228_), .ZN(new_n8231_));
  AOI21_X1   g07229(.A1(new_n8217_), .A2(new_n8231_), .B(new_n8103_), .ZN(new_n8232_));
  NAND2_X1   g07230(.A1(new_n4561_), .A2(new_n4373_), .ZN(new_n8233_));
  NAND3_X1   g07231(.A1(new_n8211_), .A2(new_n8215_), .A3(new_n8214_), .ZN(new_n8234_));
  OAI21_X1   g07232(.A1(new_n8203_), .A2(new_n8188_), .B(new_n8204_), .ZN(new_n8235_));
  AOI21_X1   g07233(.A1(new_n8235_), .A2(new_n8234_), .B(new_n8228_), .ZN(new_n8236_));
  NAND3_X1   g07234(.A1(new_n8211_), .A2(new_n8214_), .A3(new_n8204_), .ZN(new_n8237_));
  OAI21_X1   g07235(.A1(new_n8203_), .A2(new_n8188_), .B(new_n8215_), .ZN(new_n8238_));
  AOI21_X1   g07236(.A1(new_n8238_), .A2(new_n8237_), .B(new_n8159_), .ZN(new_n8239_));
  NOR3_X1    g07237(.A1(new_n8239_), .A2(new_n8236_), .A3(new_n8233_), .ZN(new_n8240_));
  OAI21_X1   g07238(.A1(new_n8232_), .A2(new_n8240_), .B(new_n8102_), .ZN(new_n8241_));
  NOR3_X1    g07239(.A1(new_n8076_), .A2(new_n8079_), .A3(new_n8080_), .ZN(new_n8242_));
  AOI21_X1   g07240(.A1(new_n8052_), .A2(new_n8067_), .B(new_n8068_), .ZN(new_n8243_));
  OAI21_X1   g07241(.A1(new_n8242_), .A2(new_n8243_), .B(new_n8098_), .ZN(new_n8244_));
  NOR3_X1    g07242(.A1(new_n8076_), .A2(new_n8079_), .A3(new_n8068_), .ZN(new_n8245_));
  AOI21_X1   g07243(.A1(new_n8052_), .A2(new_n8067_), .B(new_n8080_), .ZN(new_n8246_));
  OAI21_X1   g07244(.A1(new_n8245_), .A2(new_n8246_), .B(new_n8018_), .ZN(new_n8247_));
  NAND2_X1   g07245(.A1(new_n8244_), .A2(new_n8247_), .ZN(new_n8248_));
  AOI21_X1   g07246(.A1(new_n8217_), .A2(new_n8231_), .B(new_n8233_), .ZN(new_n8249_));
  NOR3_X1    g07247(.A1(new_n8239_), .A2(new_n8236_), .A3(new_n8103_), .ZN(new_n8250_));
  OAI21_X1   g07248(.A1(new_n8249_), .A2(new_n8250_), .B(new_n8248_), .ZN(new_n8251_));
  NAND2_X1   g07249(.A1(new_n8241_), .A2(new_n8251_), .ZN(new_n8252_));
  INV_X1     g07250(.I(new_n8252_), .ZN(new_n8253_));
  NAND2_X1   g07251(.A1(new_n4935_), .A2(new_n4958_), .ZN(new_n8254_));
  NAND2_X1   g07252(.A1(new_n4939_), .A2(new_n4957_), .ZN(new_n8255_));
  NAND2_X1   g07253(.A1(new_n8254_), .A2(new_n8255_), .ZN(new_n8256_));
  NOR2_X1    g07254(.A1(new_n4958_), .A2(new_n4957_), .ZN(new_n8257_));
  AOI21_X1   g07255(.A1(new_n8256_), .A2(new_n4940_), .B(new_n8257_), .ZN(new_n8258_));
  NOR2_X1    g07256(.A1(new_n4939_), .A2(new_n4957_), .ZN(new_n8259_));
  NOR2_X1    g07257(.A1(new_n4935_), .A2(new_n4958_), .ZN(new_n8260_));
  NOR4_X1    g07258(.A1(new_n8260_), .A2(new_n8259_), .A3(new_n4911_), .A4(new_n4929_), .ZN(new_n8261_));
  AOI21_X1   g07259(.A1(new_n8254_), .A2(new_n8255_), .B(new_n4940_), .ZN(new_n8262_));
  OAI22_X1   g07260(.A1(new_n8258_), .A2(new_n4956_), .B1(new_n8261_), .B2(new_n8262_), .ZN(new_n8263_));
  NOR2_X1    g07261(.A1(new_n4952_), .A2(new_n4896_), .ZN(new_n8264_));
  NOR2_X1    g07262(.A1(new_n4949_), .A2(new_n4899_), .ZN(new_n8265_));
  NOR3_X1    g07263(.A1(new_n8264_), .A2(new_n8265_), .A3(new_n4900_), .ZN(new_n8266_));
  NAND2_X1   g07264(.A1(new_n4949_), .A2(new_n4899_), .ZN(new_n8267_));
  NAND2_X1   g07265(.A1(new_n4952_), .A2(new_n4896_), .ZN(new_n8268_));
  AOI21_X1   g07266(.A1(new_n8267_), .A2(new_n8268_), .B(new_n4953_), .ZN(new_n8269_));
  NOR2_X1    g07267(.A1(new_n8269_), .A2(new_n8266_), .ZN(new_n8270_));
  NOR4_X1    g07268(.A1(new_n8270_), .A2(new_n4893_), .A3(new_n4901_), .A4(new_n4956_), .ZN(new_n8271_));
  OAI21_X1   g07269(.A1(new_n8264_), .A2(new_n8265_), .B(new_n4953_), .ZN(new_n8272_));
  NOR2_X1    g07270(.A1(new_n4896_), .A2(new_n4899_), .ZN(new_n8273_));
  INV_X1     g07271(.I(new_n8273_), .ZN(new_n8274_));
  AOI21_X1   g07272(.A1(new_n8272_), .A2(new_n8274_), .B(new_n4893_), .ZN(new_n8275_));
  NOR2_X1    g07273(.A1(new_n8275_), .A2(new_n4959_), .ZN(new_n8276_));
  NAND2_X1   g07274(.A1(new_n8276_), .A2(new_n8271_), .ZN(new_n8277_));
  NAND4_X1   g07275(.A1(new_n4946_), .A2(new_n4931_), .A3(new_n4954_), .A4(new_n4941_), .ZN(new_n8278_));
  NAND3_X1   g07276(.A1(new_n8267_), .A2(new_n8268_), .A3(new_n4953_), .ZN(new_n8279_));
  OAI21_X1   g07277(.A1(new_n8264_), .A2(new_n8265_), .B(new_n4900_), .ZN(new_n8280_));
  NAND2_X1   g07278(.A1(new_n8279_), .A2(new_n8280_), .ZN(new_n8281_));
  AOI21_X1   g07279(.A1(new_n8268_), .A2(new_n8267_), .B(new_n4900_), .ZN(new_n8282_));
  OAI22_X1   g07280(.A1(new_n8282_), .A2(new_n8273_), .B1(new_n4884_), .B2(new_n4892_), .ZN(new_n8283_));
  NAND2_X1   g07281(.A1(new_n8283_), .A2(new_n8281_), .ZN(new_n8284_));
  NAND2_X1   g07282(.A1(new_n8284_), .A2(new_n8278_), .ZN(new_n8285_));
  AOI21_X1   g07283(.A1(new_n8277_), .A2(new_n8285_), .B(new_n8263_), .ZN(new_n8286_));
  OAI21_X1   g07284(.A1(new_n8260_), .A2(new_n8259_), .B(new_n4940_), .ZN(new_n8287_));
  INV_X1     g07285(.I(new_n8257_), .ZN(new_n8288_));
  NAND2_X1   g07286(.A1(new_n8287_), .A2(new_n8288_), .ZN(new_n8289_));
  NAND3_X1   g07287(.A1(new_n8254_), .A2(new_n8255_), .A3(new_n4940_), .ZN(new_n8290_));
  OAI22_X1   g07288(.A1(new_n8260_), .A2(new_n8259_), .B1(new_n4911_), .B2(new_n4929_), .ZN(new_n8291_));
  AOI22_X1   g07289(.A1(new_n8289_), .A2(new_n4931_), .B1(new_n8290_), .B2(new_n8291_), .ZN(new_n8292_));
  NOR2_X1    g07290(.A1(new_n8275_), .A2(new_n8270_), .ZN(new_n8293_));
  NAND2_X1   g07291(.A1(new_n8293_), .A2(new_n8278_), .ZN(new_n8294_));
  NOR4_X1    g07292(.A1(new_n4956_), .A2(new_n4893_), .A3(new_n4901_), .A4(new_n4959_), .ZN(new_n8295_));
  NAND2_X1   g07293(.A1(new_n8284_), .A2(new_n8295_), .ZN(new_n8296_));
  AOI21_X1   g07294(.A1(new_n8294_), .A2(new_n8296_), .B(new_n8292_), .ZN(new_n8297_));
  NOR2_X1    g07295(.A1(new_n8286_), .A2(new_n8297_), .ZN(new_n8298_));
  NOR2_X1    g07296(.A1(new_n4823_), .A2(new_n4825_), .ZN(new_n8299_));
  INV_X1     g07297(.I(new_n4839_), .ZN(new_n8300_));
  OAI21_X1   g07298(.A1(new_n8299_), .A2(new_n4821_), .B(new_n8300_), .ZN(new_n8301_));
  NAND2_X1   g07299(.A1(new_n8301_), .A2(new_n4842_), .ZN(new_n8302_));
  INV_X1     g07300(.I(new_n4841_), .ZN(new_n8303_));
  OAI21_X1   g07301(.A1(new_n4833_), .A2(new_n4813_), .B(new_n8303_), .ZN(new_n8304_));
  NAND2_X1   g07302(.A1(new_n8304_), .A2(new_n4840_), .ZN(new_n8305_));
  NAND2_X1   g07303(.A1(new_n8302_), .A2(new_n8305_), .ZN(new_n8306_));
  NAND2_X1   g07304(.A1(new_n4814_), .A2(new_n4813_), .ZN(new_n8307_));
  NAND2_X1   g07305(.A1(new_n4815_), .A2(\A[427] ), .ZN(new_n8308_));
  NAND2_X1   g07306(.A1(new_n4817_), .A2(\A[428] ), .ZN(new_n8309_));
  NAND3_X1   g07307(.A1(new_n8308_), .A2(new_n8309_), .A3(\A[429] ), .ZN(new_n8310_));
  AOI22_X1   g07308(.A1(new_n8307_), .A2(new_n8310_), .B1(new_n4826_), .B2(new_n4829_), .ZN(new_n8311_));
  NOR2_X1    g07309(.A1(new_n4840_), .A2(new_n4842_), .ZN(new_n8312_));
  AOI21_X1   g07310(.A1(new_n8306_), .A2(new_n8311_), .B(new_n8312_), .ZN(new_n8313_));
  NOR2_X1    g07311(.A1(new_n8304_), .A2(new_n4840_), .ZN(new_n8314_));
  NOR2_X1    g07312(.A1(new_n8301_), .A2(new_n4842_), .ZN(new_n8315_));
  NOR4_X1    g07313(.A1(new_n8315_), .A2(new_n8314_), .A3(new_n4820_), .A4(new_n4836_), .ZN(new_n8316_));
  AOI21_X1   g07314(.A1(new_n8302_), .A2(new_n8305_), .B(new_n8311_), .ZN(new_n8317_));
  OAI22_X1   g07315(.A1(new_n8313_), .A2(new_n4860_), .B1(new_n8316_), .B2(new_n8317_), .ZN(new_n8318_));
  NAND2_X1   g07316(.A1(new_n4854_), .A2(new_n4802_), .ZN(new_n8319_));
  NAND2_X1   g07317(.A1(new_n4852_), .A2(new_n4806_), .ZN(new_n8320_));
  NAND3_X1   g07318(.A1(new_n8320_), .A2(new_n8319_), .A3(new_n4855_), .ZN(new_n8321_));
  NOR2_X1    g07319(.A1(new_n4852_), .A2(new_n4806_), .ZN(new_n8322_));
  NOR2_X1    g07320(.A1(new_n4854_), .A2(new_n4802_), .ZN(new_n8323_));
  OAI21_X1   g07321(.A1(new_n8322_), .A2(new_n8323_), .B(new_n4810_), .ZN(new_n8324_));
  NAND2_X1   g07322(.A1(new_n8324_), .A2(new_n8321_), .ZN(new_n8325_));
  NAND2_X1   g07323(.A1(new_n8320_), .A2(new_n8319_), .ZN(new_n8326_));
  NOR2_X1    g07324(.A1(new_n4802_), .A2(new_n4806_), .ZN(new_n8327_));
  AOI21_X1   g07325(.A1(new_n8326_), .A2(new_n4855_), .B(new_n8327_), .ZN(new_n8328_));
  NOR2_X1    g07326(.A1(new_n4860_), .A2(new_n4800_), .ZN(new_n8329_));
  INV_X1     g07327(.I(new_n8327_), .ZN(new_n8330_));
  OAI21_X1   g07328(.A1(new_n8322_), .A2(new_n8323_), .B(new_n4855_), .ZN(new_n8331_));
  NAND2_X1   g07329(.A1(new_n8331_), .A2(new_n8330_), .ZN(new_n8332_));
  AOI21_X1   g07330(.A1(new_n8332_), .A2(new_n4849_), .B(new_n4843_), .ZN(new_n8333_));
  NAND4_X1   g07331(.A1(new_n8333_), .A2(new_n8325_), .A3(new_n8328_), .A4(new_n8329_), .ZN(new_n8334_));
  NAND4_X1   g07332(.A1(new_n4844_), .A2(new_n4838_), .A3(new_n4849_), .A4(new_n4856_), .ZN(new_n8335_));
  OAI21_X1   g07333(.A1(new_n4800_), .A2(new_n8328_), .B(new_n8325_), .ZN(new_n8336_));
  NAND2_X1   g07334(.A1(new_n8336_), .A2(new_n8335_), .ZN(new_n8337_));
  AOI21_X1   g07335(.A1(new_n8337_), .A2(new_n8334_), .B(new_n8318_), .ZN(new_n8338_));
  OAI21_X1   g07336(.A1(new_n8315_), .A2(new_n8314_), .B(new_n8311_), .ZN(new_n8339_));
  INV_X1     g07337(.I(new_n8312_), .ZN(new_n8340_));
  NAND2_X1   g07338(.A1(new_n8339_), .A2(new_n8340_), .ZN(new_n8341_));
  NAND3_X1   g07339(.A1(new_n8302_), .A2(new_n8305_), .A3(new_n8311_), .ZN(new_n8342_));
  OAI22_X1   g07340(.A1(new_n8315_), .A2(new_n8314_), .B1(new_n4820_), .B2(new_n4836_), .ZN(new_n8343_));
  AOI22_X1   g07341(.A1(new_n8341_), .A2(new_n4838_), .B1(new_n8342_), .B2(new_n8343_), .ZN(new_n8344_));
  AOI22_X1   g07342(.A1(new_n8332_), .A2(new_n4849_), .B1(new_n8321_), .B2(new_n8324_), .ZN(new_n8345_));
  NAND2_X1   g07343(.A1(new_n8345_), .A2(new_n8335_), .ZN(new_n8346_));
  NOR4_X1    g07344(.A1(new_n4860_), .A2(new_n4800_), .A3(new_n4811_), .A4(new_n4843_), .ZN(new_n8347_));
  NAND2_X1   g07345(.A1(new_n8336_), .A2(new_n8347_), .ZN(new_n8348_));
  AOI21_X1   g07346(.A1(new_n8348_), .A2(new_n8346_), .B(new_n8344_), .ZN(new_n8349_));
  NAND2_X1   g07347(.A1(new_n4969_), .A2(new_n4863_), .ZN(new_n8350_));
  NOR3_X1    g07348(.A1(new_n8338_), .A2(new_n8349_), .A3(new_n8350_), .ZN(new_n8351_));
  NAND4_X1   g07349(.A1(new_n8325_), .A2(new_n4849_), .A3(new_n4856_), .A4(new_n4838_), .ZN(new_n8352_));
  OAI21_X1   g07350(.A1(new_n8328_), .A2(new_n4800_), .B(new_n4844_), .ZN(new_n8353_));
  NOR2_X1    g07351(.A1(new_n8352_), .A2(new_n8353_), .ZN(new_n8354_));
  NOR2_X1    g07352(.A1(new_n8345_), .A2(new_n8347_), .ZN(new_n8355_));
  OAI21_X1   g07353(.A1(new_n8354_), .A2(new_n8355_), .B(new_n8344_), .ZN(new_n8356_));
  NOR3_X1    g07354(.A1(new_n8322_), .A2(new_n8323_), .A3(new_n4810_), .ZN(new_n8357_));
  AOI21_X1   g07355(.A1(new_n8320_), .A2(new_n8319_), .B(new_n4855_), .ZN(new_n8358_));
  NOR2_X1    g07356(.A1(new_n8357_), .A2(new_n8358_), .ZN(new_n8359_));
  NOR2_X1    g07357(.A1(new_n8328_), .A2(new_n4800_), .ZN(new_n8360_));
  NOR3_X1    g07358(.A1(new_n8360_), .A2(new_n8359_), .A3(new_n8347_), .ZN(new_n8361_));
  NOR2_X1    g07359(.A1(new_n8345_), .A2(new_n8335_), .ZN(new_n8362_));
  OAI21_X1   g07360(.A1(new_n8362_), .A2(new_n8361_), .B(new_n8318_), .ZN(new_n8363_));
  NOR2_X1    g07361(.A1(new_n4962_), .A2(new_n4966_), .ZN(new_n8364_));
  AOI21_X1   g07362(.A1(new_n8356_), .A2(new_n8363_), .B(new_n8364_), .ZN(new_n8365_));
  OAI21_X1   g07363(.A1(new_n8351_), .A2(new_n8365_), .B(new_n8298_), .ZN(new_n8366_));
  NOR2_X1    g07364(.A1(new_n8282_), .A2(new_n8273_), .ZN(new_n8367_));
  NAND4_X1   g07365(.A1(new_n8281_), .A2(new_n8367_), .A3(new_n4946_), .A4(new_n4931_), .ZN(new_n8368_));
  NAND2_X1   g07366(.A1(new_n8283_), .A2(new_n4941_), .ZN(new_n8369_));
  NOR2_X1    g07367(.A1(new_n8368_), .A2(new_n8369_), .ZN(new_n8370_));
  NOR2_X1    g07368(.A1(new_n8293_), .A2(new_n8295_), .ZN(new_n8371_));
  OAI21_X1   g07369(.A1(new_n8371_), .A2(new_n8370_), .B(new_n8292_), .ZN(new_n8372_));
  NOR2_X1    g07370(.A1(new_n8284_), .A2(new_n8295_), .ZN(new_n8373_));
  NOR2_X1    g07371(.A1(new_n8293_), .A2(new_n8278_), .ZN(new_n8374_));
  OAI21_X1   g07372(.A1(new_n8374_), .A2(new_n8373_), .B(new_n8263_), .ZN(new_n8375_));
  NAND2_X1   g07373(.A1(new_n8372_), .A2(new_n8375_), .ZN(new_n8376_));
  NOR3_X1    g07374(.A1(new_n8338_), .A2(new_n8349_), .A3(new_n8364_), .ZN(new_n8377_));
  AOI21_X1   g07375(.A1(new_n8356_), .A2(new_n8363_), .B(new_n8350_), .ZN(new_n8378_));
  OAI21_X1   g07376(.A1(new_n8377_), .A2(new_n8378_), .B(new_n8376_), .ZN(new_n8379_));
  NAND2_X1   g07377(.A1(new_n8379_), .A2(new_n8366_), .ZN(new_n8380_));
  NOR2_X1    g07378(.A1(new_n4724_), .A2(new_n4761_), .ZN(new_n8381_));
  NOR2_X1    g07379(.A1(new_n4715_), .A2(new_n4762_), .ZN(new_n8382_));
  OAI21_X1   g07380(.A1(new_n8381_), .A2(new_n8382_), .B(new_n4734_), .ZN(new_n8383_));
  NOR2_X1    g07381(.A1(new_n4761_), .A2(new_n4762_), .ZN(new_n8384_));
  INV_X1     g07382(.I(new_n8384_), .ZN(new_n8385_));
  NAND2_X1   g07383(.A1(new_n8383_), .A2(new_n8385_), .ZN(new_n8386_));
  NAND2_X1   g07384(.A1(new_n4715_), .A2(new_n4762_), .ZN(new_n8387_));
  NAND2_X1   g07385(.A1(new_n4724_), .A2(new_n4761_), .ZN(new_n8388_));
  NAND3_X1   g07386(.A1(new_n8387_), .A2(new_n8388_), .A3(new_n4734_), .ZN(new_n8389_));
  OAI22_X1   g07387(.A1(new_n8381_), .A2(new_n8382_), .B1(new_n4737_), .B2(new_n4743_), .ZN(new_n8390_));
  AOI22_X1   g07388(.A1(new_n8386_), .A2(new_n4745_), .B1(new_n8389_), .B2(new_n8390_), .ZN(new_n8391_));
  NAND2_X1   g07389(.A1(new_n4753_), .A2(new_n4673_), .ZN(new_n8392_));
  NAND2_X1   g07390(.A1(new_n4750_), .A2(new_n4678_), .ZN(new_n8393_));
  NAND3_X1   g07391(.A1(new_n8392_), .A2(new_n8393_), .A3(new_n4755_), .ZN(new_n8394_));
  NOR2_X1    g07392(.A1(new_n4750_), .A2(new_n4678_), .ZN(new_n8395_));
  NOR2_X1    g07393(.A1(new_n4753_), .A2(new_n4673_), .ZN(new_n8396_));
  OAI21_X1   g07394(.A1(new_n8395_), .A2(new_n8396_), .B(new_n4692_), .ZN(new_n8397_));
  NAND2_X1   g07395(.A1(new_n8397_), .A2(new_n8394_), .ZN(new_n8398_));
  AOI22_X1   g07396(.A1(new_n4744_), .A2(new_n4739_), .B1(new_n4757_), .B2(new_n4758_), .ZN(new_n8399_));
  NAND3_X1   g07397(.A1(new_n8399_), .A2(new_n4756_), .A3(new_n4735_), .ZN(new_n8400_));
  NOR2_X1    g07398(.A1(new_n4673_), .A2(new_n4678_), .ZN(new_n8401_));
  AOI21_X1   g07399(.A1(new_n8392_), .A2(new_n8393_), .B(new_n4692_), .ZN(new_n8402_));
  OAI21_X1   g07400(.A1(new_n8401_), .A2(new_n8402_), .B(new_n4759_), .ZN(new_n8403_));
  NAND3_X1   g07401(.A1(new_n8400_), .A2(new_n8403_), .A3(new_n8398_), .ZN(new_n8404_));
  OAI22_X1   g07402(.A1(new_n4764_), .A2(new_n4765_), .B1(new_n4704_), .B2(new_n4698_), .ZN(new_n8405_));
  NOR3_X1    g07403(.A1(new_n8405_), .A2(new_n4693_), .A3(new_n4763_), .ZN(new_n8406_));
  NAND2_X1   g07404(.A1(new_n8403_), .A2(new_n8398_), .ZN(new_n8407_));
  NAND2_X1   g07405(.A1(new_n8407_), .A2(new_n8406_), .ZN(new_n8408_));
  AOI21_X1   g07406(.A1(new_n8408_), .A2(new_n8404_), .B(new_n8391_), .ZN(new_n8409_));
  NAND2_X1   g07407(.A1(new_n8387_), .A2(new_n8388_), .ZN(new_n8410_));
  AOI21_X1   g07408(.A1(new_n8410_), .A2(new_n4734_), .B(new_n8384_), .ZN(new_n8411_));
  NOR4_X1    g07409(.A1(new_n8381_), .A2(new_n8382_), .A3(new_n4737_), .A4(new_n4743_), .ZN(new_n8412_));
  AOI21_X1   g07410(.A1(new_n8387_), .A2(new_n8388_), .B(new_n4734_), .ZN(new_n8413_));
  OAI22_X1   g07411(.A1(new_n8411_), .A2(new_n4766_), .B1(new_n8412_), .B2(new_n8413_), .ZN(new_n8414_));
  NOR3_X1    g07412(.A1(new_n8395_), .A2(new_n8396_), .A3(new_n4692_), .ZN(new_n8415_));
  AOI21_X1   g07413(.A1(new_n8392_), .A2(new_n8393_), .B(new_n4755_), .ZN(new_n8416_));
  NOR2_X1    g07414(.A1(new_n8416_), .A2(new_n8415_), .ZN(new_n8417_));
  NOR3_X1    g07415(.A1(new_n8417_), .A2(new_n4693_), .A3(new_n8405_), .ZN(new_n8418_));
  INV_X1     g07416(.I(new_n8401_), .ZN(new_n8419_));
  OAI21_X1   g07417(.A1(new_n8395_), .A2(new_n8396_), .B(new_n4755_), .ZN(new_n8420_));
  NAND2_X1   g07418(.A1(new_n8420_), .A2(new_n8419_), .ZN(new_n8421_));
  AOI21_X1   g07419(.A1(new_n8421_), .A2(new_n4759_), .B(new_n4763_), .ZN(new_n8422_));
  NAND2_X1   g07420(.A1(new_n8418_), .A2(new_n8422_), .ZN(new_n8423_));
  NAND2_X1   g07421(.A1(new_n8407_), .A2(new_n8400_), .ZN(new_n8424_));
  AOI21_X1   g07422(.A1(new_n8423_), .A2(new_n8424_), .B(new_n8414_), .ZN(new_n8425_));
  NOR2_X1    g07423(.A1(new_n8425_), .A2(new_n8409_), .ZN(new_n8426_));
  NOR2_X1    g07424(.A1(new_n4660_), .A2(new_n4603_), .ZN(new_n8427_));
  NOR2_X1    g07425(.A1(new_n4658_), .A2(new_n4607_), .ZN(new_n8428_));
  OAI21_X1   g07426(.A1(new_n8427_), .A2(new_n8428_), .B(new_n4661_), .ZN(new_n8429_));
  NOR2_X1    g07427(.A1(new_n4603_), .A2(new_n4607_), .ZN(new_n8430_));
  INV_X1     g07428(.I(new_n8430_), .ZN(new_n8431_));
  NAND2_X1   g07429(.A1(new_n8429_), .A2(new_n8431_), .ZN(new_n8432_));
  NAND2_X1   g07430(.A1(new_n4658_), .A2(new_n4607_), .ZN(new_n8433_));
  NAND2_X1   g07431(.A1(new_n4660_), .A2(new_n4603_), .ZN(new_n8434_));
  NAND3_X1   g07432(.A1(new_n8433_), .A2(new_n8434_), .A3(new_n4661_), .ZN(new_n8435_));
  OAI21_X1   g07433(.A1(new_n8427_), .A2(new_n8428_), .B(new_n4625_), .ZN(new_n8436_));
  AOI22_X1   g07434(.A1(new_n8432_), .A2(new_n4665_), .B1(new_n8435_), .B2(new_n8436_), .ZN(new_n8437_));
  NAND2_X1   g07435(.A1(new_n4574_), .A2(new_n4645_), .ZN(new_n8438_));
  NAND2_X1   g07436(.A1(new_n4570_), .A2(new_n4647_), .ZN(new_n8439_));
  NAND3_X1   g07437(.A1(new_n8439_), .A2(new_n8438_), .A3(new_n4587_), .ZN(new_n8440_));
  NOR2_X1    g07438(.A1(new_n4570_), .A2(new_n4647_), .ZN(new_n8441_));
  NOR2_X1    g07439(.A1(new_n4574_), .A2(new_n4645_), .ZN(new_n8442_));
  OAI21_X1   g07440(.A1(new_n8441_), .A2(new_n8442_), .B(new_n4651_), .ZN(new_n8443_));
  NAND2_X1   g07441(.A1(new_n8443_), .A2(new_n8440_), .ZN(new_n8444_));
  NAND4_X1   g07442(.A1(new_n8444_), .A2(new_n4588_), .A3(new_n4598_), .A4(new_n4665_), .ZN(new_n8445_));
  NOR2_X1    g07443(.A1(new_n4645_), .A2(new_n4647_), .ZN(new_n8446_));
  AOI21_X1   g07444(.A1(new_n8439_), .A2(new_n8438_), .B(new_n4651_), .ZN(new_n8447_));
  NOR2_X1    g07445(.A1(new_n8447_), .A2(new_n8446_), .ZN(new_n8448_));
  OAI21_X1   g07446(.A1(new_n8448_), .A2(new_n4655_), .B(new_n4662_), .ZN(new_n8449_));
  NOR2_X1    g07447(.A1(new_n8445_), .A2(new_n8449_), .ZN(new_n8450_));
  OAI21_X1   g07448(.A1(new_n8446_), .A2(new_n8447_), .B(new_n4598_), .ZN(new_n8451_));
  OAI22_X1   g07449(.A1(new_n4653_), .A2(new_n4654_), .B1(new_n4632_), .B2(new_n4639_), .ZN(new_n8452_));
  NOR3_X1    g07450(.A1(new_n8452_), .A2(new_n4652_), .A3(new_n4626_), .ZN(new_n8453_));
  AOI21_X1   g07451(.A1(new_n8444_), .A2(new_n8451_), .B(new_n8453_), .ZN(new_n8454_));
  OAI21_X1   g07452(.A1(new_n8450_), .A2(new_n8454_), .B(new_n8437_), .ZN(new_n8455_));
  NAND2_X1   g07453(.A1(new_n8436_), .A2(new_n8435_), .ZN(new_n8456_));
  AOI21_X1   g07454(.A1(new_n8433_), .A2(new_n8434_), .B(new_n4625_), .ZN(new_n8457_));
  OAI22_X1   g07455(.A1(new_n8457_), .A2(new_n8430_), .B1(new_n4632_), .B2(new_n4639_), .ZN(new_n8458_));
  NAND2_X1   g07456(.A1(new_n8458_), .A2(new_n8456_), .ZN(new_n8459_));
  NOR3_X1    g07457(.A1(new_n8441_), .A2(new_n8442_), .A3(new_n4651_), .ZN(new_n8460_));
  AOI21_X1   g07458(.A1(new_n8439_), .A2(new_n8438_), .B(new_n4587_), .ZN(new_n8461_));
  NOR2_X1    g07459(.A1(new_n8460_), .A2(new_n8461_), .ZN(new_n8462_));
  INV_X1     g07460(.I(new_n8446_), .ZN(new_n8463_));
  OAI21_X1   g07461(.A1(new_n8441_), .A2(new_n8442_), .B(new_n4587_), .ZN(new_n8464_));
  AOI22_X1   g07462(.A1(new_n8464_), .A2(new_n8463_), .B1(new_n4593_), .B2(new_n4597_), .ZN(new_n8465_));
  NOR3_X1    g07463(.A1(new_n8453_), .A2(new_n8465_), .A3(new_n8462_), .ZN(new_n8466_));
  NAND4_X1   g07464(.A1(new_n4598_), .A2(new_n4665_), .A3(new_n4588_), .A4(new_n4662_), .ZN(new_n8467_));
  AOI21_X1   g07465(.A1(new_n8444_), .A2(new_n8451_), .B(new_n8467_), .ZN(new_n8468_));
  OAI21_X1   g07466(.A1(new_n8466_), .A2(new_n8468_), .B(new_n8459_), .ZN(new_n8469_));
  OAI22_X1   g07467(.A1(new_n4747_), .A2(new_n4768_), .B1(new_n4642_), .B2(new_n4667_), .ZN(new_n8470_));
  NAND3_X1   g07468(.A1(new_n8455_), .A2(new_n8469_), .A3(new_n8470_), .ZN(new_n8471_));
  NOR3_X1    g07469(.A1(new_n8462_), .A2(new_n4652_), .A3(new_n8452_), .ZN(new_n8472_));
  NAND2_X1   g07470(.A1(new_n8464_), .A2(new_n8463_), .ZN(new_n8473_));
  AOI21_X1   g07471(.A1(new_n8473_), .A2(new_n4598_), .B(new_n4626_), .ZN(new_n8474_));
  NAND2_X1   g07472(.A1(new_n8472_), .A2(new_n8474_), .ZN(new_n8475_));
  NAND2_X1   g07473(.A1(new_n8451_), .A2(new_n8444_), .ZN(new_n8476_));
  NAND2_X1   g07474(.A1(new_n8476_), .A2(new_n8467_), .ZN(new_n8477_));
  AOI21_X1   g07475(.A1(new_n8477_), .A2(new_n8475_), .B(new_n8459_), .ZN(new_n8478_));
  NAND3_X1   g07476(.A1(new_n8451_), .A2(new_n8467_), .A3(new_n8444_), .ZN(new_n8479_));
  NAND2_X1   g07477(.A1(new_n8476_), .A2(new_n8453_), .ZN(new_n8480_));
  AOI21_X1   g07478(.A1(new_n8480_), .A2(new_n8479_), .B(new_n8437_), .ZN(new_n8481_));
  NOR2_X1    g07479(.A1(new_n4770_), .A2(new_n4668_), .ZN(new_n8482_));
  OAI21_X1   g07480(.A1(new_n8478_), .A2(new_n8481_), .B(new_n8482_), .ZN(new_n8483_));
  AOI21_X1   g07481(.A1(new_n8483_), .A2(new_n8471_), .B(new_n8426_), .ZN(new_n8484_));
  AOI21_X1   g07482(.A1(new_n8419_), .A2(new_n8420_), .B(new_n4705_), .ZN(new_n8485_));
  NOR3_X1    g07483(.A1(new_n8406_), .A2(new_n8417_), .A3(new_n8485_), .ZN(new_n8486_));
  AOI21_X1   g07484(.A1(new_n8398_), .A2(new_n8403_), .B(new_n8400_), .ZN(new_n8487_));
  OAI21_X1   g07485(.A1(new_n8487_), .A2(new_n8486_), .B(new_n8414_), .ZN(new_n8488_));
  NAND3_X1   g07486(.A1(new_n8398_), .A2(new_n4756_), .A3(new_n8399_), .ZN(new_n8489_));
  NOR2_X1    g07487(.A1(new_n8402_), .A2(new_n8401_), .ZN(new_n8490_));
  OAI21_X1   g07488(.A1(new_n8490_), .A2(new_n4705_), .B(new_n4735_), .ZN(new_n8491_));
  NOR2_X1    g07489(.A1(new_n8489_), .A2(new_n8491_), .ZN(new_n8492_));
  AOI21_X1   g07490(.A1(new_n8398_), .A2(new_n8403_), .B(new_n8406_), .ZN(new_n8493_));
  OAI21_X1   g07491(.A1(new_n8492_), .A2(new_n8493_), .B(new_n8391_), .ZN(new_n8494_));
  NAND2_X1   g07492(.A1(new_n8494_), .A2(new_n8488_), .ZN(new_n8495_));
  NAND3_X1   g07493(.A1(new_n8455_), .A2(new_n8482_), .A3(new_n8469_), .ZN(new_n8496_));
  OAI21_X1   g07494(.A1(new_n8478_), .A2(new_n8481_), .B(new_n8470_), .ZN(new_n8497_));
  AOI21_X1   g07495(.A1(new_n8497_), .A2(new_n8496_), .B(new_n8495_), .ZN(new_n8498_));
  AOI21_X1   g07496(.A1(new_n4963_), .A2(new_n4970_), .B(new_n4772_), .ZN(new_n8499_));
  NOR3_X1    g07497(.A1(new_n8484_), .A2(new_n8498_), .A3(new_n8499_), .ZN(new_n8500_));
  NOR3_X1    g07498(.A1(new_n8478_), .A2(new_n8481_), .A3(new_n8482_), .ZN(new_n8501_));
  AOI21_X1   g07499(.A1(new_n8455_), .A2(new_n8469_), .B(new_n8470_), .ZN(new_n8502_));
  OAI21_X1   g07500(.A1(new_n8501_), .A2(new_n8502_), .B(new_n8495_), .ZN(new_n8503_));
  NOR3_X1    g07501(.A1(new_n8478_), .A2(new_n8481_), .A3(new_n8470_), .ZN(new_n8504_));
  AOI21_X1   g07502(.A1(new_n8455_), .A2(new_n8469_), .B(new_n8482_), .ZN(new_n8505_));
  OAI21_X1   g07503(.A1(new_n8505_), .A2(new_n8504_), .B(new_n8426_), .ZN(new_n8506_));
  OAI21_X1   g07504(.A1(new_n4769_), .A2(new_n4771_), .B(new_n4971_), .ZN(new_n8507_));
  AOI21_X1   g07505(.A1(new_n8506_), .A2(new_n8503_), .B(new_n8507_), .ZN(new_n8508_));
  OAI21_X1   g07506(.A1(new_n8500_), .A2(new_n8508_), .B(new_n8380_), .ZN(new_n8509_));
  NAND3_X1   g07507(.A1(new_n8356_), .A2(new_n8364_), .A3(new_n8363_), .ZN(new_n8510_));
  OAI21_X1   g07508(.A1(new_n8338_), .A2(new_n8349_), .B(new_n8350_), .ZN(new_n8511_));
  AOI21_X1   g07509(.A1(new_n8511_), .A2(new_n8510_), .B(new_n8376_), .ZN(new_n8512_));
  NAND3_X1   g07510(.A1(new_n8356_), .A2(new_n8363_), .A3(new_n8350_), .ZN(new_n8513_));
  OAI21_X1   g07511(.A1(new_n8338_), .A2(new_n8349_), .B(new_n8364_), .ZN(new_n8514_));
  AOI21_X1   g07512(.A1(new_n8513_), .A2(new_n8514_), .B(new_n8298_), .ZN(new_n8515_));
  NOR2_X1    g07513(.A1(new_n8512_), .A2(new_n8515_), .ZN(new_n8516_));
  NOR3_X1    g07514(.A1(new_n8484_), .A2(new_n8498_), .A3(new_n8507_), .ZN(new_n8517_));
  AOI21_X1   g07515(.A1(new_n8506_), .A2(new_n8503_), .B(new_n8499_), .ZN(new_n8518_));
  OAI21_X1   g07516(.A1(new_n8517_), .A2(new_n8518_), .B(new_n8516_), .ZN(new_n8519_));
  NAND2_X1   g07517(.A1(new_n4562_), .A2(new_n4972_), .ZN(new_n8520_));
  NAND3_X1   g07518(.A1(new_n8519_), .A2(new_n8509_), .A3(new_n8520_), .ZN(new_n8521_));
  INV_X1     g07519(.I(new_n8520_), .ZN(new_n8522_));
  NAND2_X1   g07520(.A1(new_n8519_), .A2(new_n8509_), .ZN(new_n8523_));
  NAND2_X1   g07521(.A1(new_n8523_), .A2(new_n8522_), .ZN(new_n8524_));
  AOI21_X1   g07522(.A1(new_n8524_), .A2(new_n8521_), .B(new_n8253_), .ZN(new_n8525_));
  INV_X1     g07523(.I(new_n8525_), .ZN(new_n8526_));
  NAND3_X1   g07524(.A1(new_n8522_), .A2(new_n8519_), .A3(new_n8509_), .ZN(new_n8527_));
  NAND2_X1   g07525(.A1(new_n8523_), .A2(new_n8520_), .ZN(new_n8528_));
  NAND2_X1   g07526(.A1(new_n8528_), .A2(new_n8527_), .ZN(new_n8529_));
  NAND2_X1   g07527(.A1(new_n8529_), .A2(new_n8253_), .ZN(new_n8530_));
  NOR2_X1    g07528(.A1(new_n4973_), .A2(new_n5751_), .ZN(new_n8531_));
  NAND3_X1   g07529(.A1(new_n8526_), .A2(new_n8530_), .A3(new_n8531_), .ZN(new_n8532_));
  AOI21_X1   g07530(.A1(new_n8528_), .A2(new_n8527_), .B(new_n8252_), .ZN(new_n8533_));
  INV_X1     g07531(.I(new_n8531_), .ZN(new_n8534_));
  OAI21_X1   g07532(.A1(new_n8525_), .A2(new_n8533_), .B(new_n8534_), .ZN(new_n8535_));
  NAND2_X1   g07533(.A1(new_n8532_), .A2(new_n8535_), .ZN(new_n8536_));
  NAND2_X1   g07534(.A1(new_n8536_), .A2(new_n7970_), .ZN(new_n8537_));
  NOR3_X1    g07535(.A1(new_n8525_), .A2(new_n8533_), .A3(new_n8531_), .ZN(new_n8538_));
  AOI21_X1   g07536(.A1(new_n8526_), .A2(new_n8530_), .B(new_n8534_), .ZN(new_n8539_));
  OAI21_X1   g07537(.A1(new_n8539_), .A2(new_n8538_), .B(new_n7969_), .ZN(new_n8540_));
  NAND2_X1   g07538(.A1(new_n8537_), .A2(new_n8540_), .ZN(new_n8541_));
  NAND2_X1   g07539(.A1(new_n8541_), .A2(new_n7384_), .ZN(new_n8542_));
  NOR2_X1    g07540(.A1(new_n7371_), .A2(new_n7350_), .ZN(new_n8543_));
  NOR2_X1    g07541(.A1(new_n7369_), .A2(new_n7354_), .ZN(new_n8544_));
  OAI21_X1   g07542(.A1(new_n8544_), .A2(new_n8543_), .B(new_n7372_), .ZN(new_n8545_));
  NOR2_X1    g07543(.A1(new_n7350_), .A2(new_n7354_), .ZN(new_n8546_));
  INV_X1     g07544(.I(new_n8546_), .ZN(new_n8547_));
  NAND2_X1   g07545(.A1(new_n8545_), .A2(new_n8547_), .ZN(new_n8548_));
  NAND2_X1   g07546(.A1(new_n7369_), .A2(new_n7354_), .ZN(new_n8549_));
  NAND2_X1   g07547(.A1(new_n7371_), .A2(new_n7350_), .ZN(new_n8550_));
  NAND3_X1   g07548(.A1(new_n8549_), .A2(new_n8550_), .A3(new_n7372_), .ZN(new_n8551_));
  OAI21_X1   g07549(.A1(new_n8544_), .A2(new_n8543_), .B(new_n7355_), .ZN(new_n8552_));
  AOI22_X1   g07550(.A1(new_n8548_), .A2(new_n7366_), .B1(new_n8551_), .B2(new_n8552_), .ZN(new_n8553_));
  NAND2_X1   g07551(.A1(new_n7284_), .A2(new_n7285_), .ZN(new_n8554_));
  AOI21_X1   g07552(.A1(new_n8554_), .A2(\A[87] ), .B(new_n7312_), .ZN(new_n8555_));
  NAND2_X1   g07553(.A1(new_n7310_), .A2(new_n8555_), .ZN(new_n8556_));
  XOR2_X1    g07554(.A1(\A[88] ), .A2(\A[89] ), .Z(new_n8557_));
  AOI21_X1   g07555(.A1(new_n8557_), .A2(\A[90] ), .B(new_n7308_), .ZN(new_n8558_));
  NAND2_X1   g07556(.A1(new_n7314_), .A2(new_n8558_), .ZN(new_n8559_));
  NAND3_X1   g07557(.A1(new_n8556_), .A2(new_n8559_), .A3(new_n7315_), .ZN(new_n8560_));
  NOR2_X1    g07558(.A1(new_n7314_), .A2(new_n8558_), .ZN(new_n8561_));
  NOR2_X1    g07559(.A1(new_n7310_), .A2(new_n8555_), .ZN(new_n8562_));
  OAI22_X1   g07560(.A1(new_n7283_), .A2(new_n7286_), .B1(new_n7303_), .B2(new_n7302_), .ZN(new_n8563_));
  OAI21_X1   g07561(.A1(new_n8562_), .A2(new_n8561_), .B(new_n8563_), .ZN(new_n8564_));
  NAND2_X1   g07562(.A1(new_n8564_), .A2(new_n8560_), .ZN(new_n8565_));
  AOI22_X1   g07563(.A1(new_n7298_), .A2(new_n7305_), .B1(new_n7365_), .B2(new_n7364_), .ZN(new_n8566_));
  NAND3_X1   g07564(.A1(new_n8565_), .A2(new_n7316_), .A3(new_n8566_), .ZN(new_n8567_));
  AOI21_X1   g07565(.A1(new_n8556_), .A2(new_n8559_), .B(new_n8563_), .ZN(new_n8568_));
  NOR2_X1    g07566(.A1(new_n8555_), .A2(new_n8558_), .ZN(new_n8569_));
  NOR2_X1    g07567(.A1(new_n8568_), .A2(new_n8569_), .ZN(new_n8570_));
  OAI21_X1   g07568(.A1(new_n8570_), .A2(new_n7361_), .B(new_n7373_), .ZN(new_n8571_));
  NOR2_X1    g07569(.A1(new_n8567_), .A2(new_n8571_), .ZN(new_n8572_));
  NOR4_X1    g07570(.A1(new_n7362_), .A2(new_n7361_), .A3(new_n7347_), .A4(new_n7356_), .ZN(new_n8573_));
  OAI21_X1   g07571(.A1(new_n8562_), .A2(new_n8561_), .B(new_n7315_), .ZN(new_n8574_));
  INV_X1     g07572(.I(new_n8569_), .ZN(new_n8575_));
  NAND2_X1   g07573(.A1(new_n8574_), .A2(new_n8575_), .ZN(new_n8576_));
  NOR3_X1    g07574(.A1(new_n8562_), .A2(new_n8561_), .A3(new_n8563_), .ZN(new_n8577_));
  AOI21_X1   g07575(.A1(new_n8556_), .A2(new_n8559_), .B(new_n7315_), .ZN(new_n8578_));
  NOR2_X1    g07576(.A1(new_n8578_), .A2(new_n8577_), .ZN(new_n8579_));
  AOI21_X1   g07577(.A1(new_n7306_), .A2(new_n8576_), .B(new_n8579_), .ZN(new_n8580_));
  NOR2_X1    g07578(.A1(new_n8580_), .A2(new_n8573_), .ZN(new_n8581_));
  OAI21_X1   g07579(.A1(new_n8581_), .A2(new_n8572_), .B(new_n8553_), .ZN(new_n8582_));
  NAND2_X1   g07580(.A1(new_n8549_), .A2(new_n8550_), .ZN(new_n8583_));
  AOI21_X1   g07581(.A1(new_n8583_), .A2(new_n7372_), .B(new_n8546_), .ZN(new_n8584_));
  NAND2_X1   g07582(.A1(new_n8552_), .A2(new_n8551_), .ZN(new_n8585_));
  OAI21_X1   g07583(.A1(new_n7347_), .A2(new_n8584_), .B(new_n8585_), .ZN(new_n8586_));
  OAI21_X1   g07584(.A1(new_n8568_), .A2(new_n8569_), .B(new_n7306_), .ZN(new_n8587_));
  NAND2_X1   g07585(.A1(new_n8587_), .A2(new_n8565_), .ZN(new_n8588_));
  NOR2_X1    g07586(.A1(new_n8588_), .A2(new_n8573_), .ZN(new_n8589_));
  NAND3_X1   g07587(.A1(new_n8566_), .A2(new_n7316_), .A3(new_n7373_), .ZN(new_n8590_));
  NOR2_X1    g07588(.A1(new_n8580_), .A2(new_n8590_), .ZN(new_n8591_));
  OAI21_X1   g07589(.A1(new_n8591_), .A2(new_n8589_), .B(new_n8586_), .ZN(new_n8592_));
  NAND2_X1   g07590(.A1(new_n8582_), .A2(new_n8592_), .ZN(new_n8593_));
  NAND2_X1   g07591(.A1(new_n7271_), .A2(new_n7245_), .ZN(new_n8594_));
  NAND2_X1   g07592(.A1(new_n7273_), .A2(new_n7242_), .ZN(new_n8595_));
  NAND2_X1   g07593(.A1(new_n8594_), .A2(new_n8595_), .ZN(new_n8596_));
  NOR2_X1    g07594(.A1(new_n7242_), .A2(new_n7245_), .ZN(new_n8597_));
  AOI21_X1   g07595(.A1(new_n8596_), .A2(new_n7274_), .B(new_n8597_), .ZN(new_n8598_));
  NOR2_X1    g07596(.A1(new_n7273_), .A2(new_n7242_), .ZN(new_n8599_));
  NOR2_X1    g07597(.A1(new_n7271_), .A2(new_n7245_), .ZN(new_n8600_));
  NOR3_X1    g07598(.A1(new_n8599_), .A2(new_n8600_), .A3(new_n7251_), .ZN(new_n8601_));
  AOI21_X1   g07599(.A1(new_n8594_), .A2(new_n8595_), .B(new_n7274_), .ZN(new_n8602_));
  OAI22_X1   g07600(.A1(new_n8598_), .A2(new_n7239_), .B1(new_n8601_), .B2(new_n8602_), .ZN(new_n8603_));
  NAND2_X1   g07601(.A1(new_n7205_), .A2(new_n7261_), .ZN(new_n8604_));
  NAND2_X1   g07602(.A1(new_n7208_), .A2(new_n7258_), .ZN(new_n8605_));
  AOI21_X1   g07603(.A1(new_n8604_), .A2(new_n8605_), .B(new_n7264_), .ZN(new_n8606_));
  NOR2_X1    g07604(.A1(new_n7258_), .A2(new_n7261_), .ZN(new_n8607_));
  NOR2_X1    g07605(.A1(new_n8606_), .A2(new_n8607_), .ZN(new_n8608_));
  NAND3_X1   g07606(.A1(new_n8604_), .A2(new_n8605_), .A3(new_n7209_), .ZN(new_n8609_));
  NOR2_X1    g07607(.A1(new_n7208_), .A2(new_n7258_), .ZN(new_n8610_));
  NOR2_X1    g07608(.A1(new_n7205_), .A2(new_n7261_), .ZN(new_n8611_));
  OAI21_X1   g07609(.A1(new_n8611_), .A2(new_n8610_), .B(new_n7264_), .ZN(new_n8612_));
  NAND2_X1   g07610(.A1(new_n8612_), .A2(new_n8609_), .ZN(new_n8613_));
  AOI22_X1   g07611(.A1(new_n7193_), .A2(new_n7200_), .B1(new_n7268_), .B2(new_n7267_), .ZN(new_n8614_));
  OAI21_X1   g07612(.A1(new_n8611_), .A2(new_n8610_), .B(new_n7209_), .ZN(new_n8615_));
  INV_X1     g07613(.I(new_n8607_), .ZN(new_n8616_));
  NAND2_X1   g07614(.A1(new_n8615_), .A2(new_n8616_), .ZN(new_n8617_));
  AOI21_X1   g07615(.A1(new_n8617_), .A2(new_n7201_), .B(new_n7252_), .ZN(new_n8618_));
  NAND4_X1   g07616(.A1(new_n8618_), .A2(new_n8608_), .A3(new_n8613_), .A4(new_n8614_), .ZN(new_n8619_));
  NOR3_X1    g07617(.A1(new_n8611_), .A2(new_n8610_), .A3(new_n7264_), .ZN(new_n8620_));
  AOI21_X1   g07618(.A1(new_n8604_), .A2(new_n8605_), .B(new_n7209_), .ZN(new_n8621_));
  NOR2_X1    g07619(.A1(new_n8620_), .A2(new_n8621_), .ZN(new_n8622_));
  AOI21_X1   g07620(.A1(new_n8615_), .A2(new_n8616_), .B(new_n7257_), .ZN(new_n8623_));
  NAND3_X1   g07621(.A1(new_n8614_), .A2(new_n7210_), .A3(new_n7275_), .ZN(new_n8624_));
  OAI21_X1   g07622(.A1(new_n8622_), .A2(new_n8623_), .B(new_n8624_), .ZN(new_n8625_));
  AOI21_X1   g07623(.A1(new_n8619_), .A2(new_n8625_), .B(new_n8603_), .ZN(new_n8626_));
  OAI21_X1   g07624(.A1(new_n8599_), .A2(new_n8600_), .B(new_n7274_), .ZN(new_n8627_));
  INV_X1     g07625(.I(new_n8597_), .ZN(new_n8628_));
  NAND2_X1   g07626(.A1(new_n8627_), .A2(new_n8628_), .ZN(new_n8629_));
  NAND3_X1   g07627(.A1(new_n8594_), .A2(new_n8595_), .A3(new_n7274_), .ZN(new_n8630_));
  OAI21_X1   g07628(.A1(new_n8599_), .A2(new_n8600_), .B(new_n7251_), .ZN(new_n8631_));
  AOI22_X1   g07629(.A1(new_n8629_), .A2(new_n7269_), .B1(new_n8630_), .B2(new_n8631_), .ZN(new_n8632_));
  NOR4_X1    g07630(.A1(new_n7257_), .A2(new_n7239_), .A3(new_n7265_), .A4(new_n7252_), .ZN(new_n8633_));
  OAI21_X1   g07631(.A1(new_n8622_), .A2(new_n8623_), .B(new_n8633_), .ZN(new_n8634_));
  OAI21_X1   g07632(.A1(new_n8606_), .A2(new_n8607_), .B(new_n7201_), .ZN(new_n8635_));
  NAND3_X1   g07633(.A1(new_n8624_), .A2(new_n8613_), .A3(new_n8635_), .ZN(new_n8636_));
  AOI21_X1   g07634(.A1(new_n8634_), .A2(new_n8636_), .B(new_n8632_), .ZN(new_n8637_));
  NAND2_X1   g07635(.A1(new_n7376_), .A2(new_n7378_), .ZN(new_n8638_));
  NOR3_X1    g07636(.A1(new_n8626_), .A2(new_n8638_), .A3(new_n8637_), .ZN(new_n8639_));
  NAND3_X1   g07637(.A1(new_n8613_), .A2(new_n7210_), .A3(new_n8614_), .ZN(new_n8640_));
  OAI21_X1   g07638(.A1(new_n8608_), .A2(new_n7257_), .B(new_n7275_), .ZN(new_n8641_));
  NOR2_X1    g07639(.A1(new_n8640_), .A2(new_n8641_), .ZN(new_n8642_));
  AOI21_X1   g07640(.A1(new_n8613_), .A2(new_n8635_), .B(new_n8633_), .ZN(new_n8643_));
  OAI21_X1   g07641(.A1(new_n8642_), .A2(new_n8643_), .B(new_n8632_), .ZN(new_n8644_));
  AOI21_X1   g07642(.A1(new_n8613_), .A2(new_n8635_), .B(new_n8624_), .ZN(new_n8645_));
  NOR3_X1    g07643(.A1(new_n8633_), .A2(new_n8623_), .A3(new_n8622_), .ZN(new_n8646_));
  OAI21_X1   g07644(.A1(new_n8645_), .A2(new_n8646_), .B(new_n8603_), .ZN(new_n8647_));
  AOI22_X1   g07645(.A1(new_n7375_), .A2(new_n7358_), .B1(new_n7254_), .B2(new_n7277_), .ZN(new_n8648_));
  AOI21_X1   g07646(.A1(new_n8644_), .A2(new_n8647_), .B(new_n8648_), .ZN(new_n8649_));
  NOR2_X1    g07647(.A1(new_n8639_), .A2(new_n8649_), .ZN(new_n8650_));
  NOR2_X1    g07648(.A1(new_n8650_), .A2(new_n8593_), .ZN(new_n8651_));
  NOR4_X1    g07649(.A1(new_n8579_), .A2(new_n8576_), .A3(new_n7361_), .A4(new_n7347_), .ZN(new_n8652_));
  AOI21_X1   g07650(.A1(new_n8576_), .A2(new_n7306_), .B(new_n7356_), .ZN(new_n8653_));
  NAND2_X1   g07651(.A1(new_n8652_), .A2(new_n8653_), .ZN(new_n8654_));
  NAND2_X1   g07652(.A1(new_n8588_), .A2(new_n8590_), .ZN(new_n8655_));
  AOI21_X1   g07653(.A1(new_n8654_), .A2(new_n8655_), .B(new_n8586_), .ZN(new_n8656_));
  NAND3_X1   g07654(.A1(new_n8590_), .A2(new_n8587_), .A3(new_n8565_), .ZN(new_n8657_));
  NAND2_X1   g07655(.A1(new_n8588_), .A2(new_n8573_), .ZN(new_n8658_));
  AOI21_X1   g07656(.A1(new_n8658_), .A2(new_n8657_), .B(new_n8553_), .ZN(new_n8659_));
  NOR2_X1    g07657(.A1(new_n8656_), .A2(new_n8659_), .ZN(new_n8660_));
  NAND3_X1   g07658(.A1(new_n8644_), .A2(new_n8638_), .A3(new_n8647_), .ZN(new_n8661_));
  OAI21_X1   g07659(.A1(new_n8626_), .A2(new_n8637_), .B(new_n8648_), .ZN(new_n8662_));
  AOI21_X1   g07660(.A1(new_n8661_), .A2(new_n8662_), .B(new_n8660_), .ZN(new_n8663_));
  NOR2_X1    g07661(.A1(new_n8651_), .A2(new_n8663_), .ZN(new_n8664_));
  NAND2_X1   g07662(.A1(new_n7161_), .A2(new_n7151_), .ZN(new_n8665_));
  NAND2_X1   g07663(.A1(new_n7163_), .A2(new_n7147_), .ZN(new_n8666_));
  NAND2_X1   g07664(.A1(new_n8665_), .A2(new_n8666_), .ZN(new_n8667_));
  NOR2_X1    g07665(.A1(new_n7151_), .A2(new_n7147_), .ZN(new_n8668_));
  AOI21_X1   g07666(.A1(new_n8667_), .A2(new_n7164_), .B(new_n8668_), .ZN(new_n8669_));
  NOR2_X1    g07667(.A1(new_n7163_), .A2(new_n7147_), .ZN(new_n8670_));
  NOR2_X1    g07668(.A1(new_n7161_), .A2(new_n7151_), .ZN(new_n8671_));
  NOR3_X1    g07669(.A1(new_n8671_), .A2(new_n8670_), .A3(new_n7152_), .ZN(new_n8672_));
  AOI21_X1   g07670(.A1(new_n8665_), .A2(new_n8666_), .B(new_n7164_), .ZN(new_n8673_));
  OAI22_X1   g07671(.A1(new_n8669_), .A2(new_n7145_), .B1(new_n8672_), .B2(new_n8673_), .ZN(new_n8674_));
  NAND2_X1   g07672(.A1(new_n7082_), .A2(new_n7084_), .ZN(new_n8675_));
  AOI21_X1   g07673(.A1(new_n8675_), .A2(\A[114] ), .B(new_n7104_), .ZN(new_n8676_));
  NOR2_X1    g07674(.A1(new_n7110_), .A2(new_n8676_), .ZN(new_n8677_));
  AOI21_X1   g07675(.A1(new_n7079_), .A2(\A[111] ), .B(new_n7108_), .ZN(new_n8678_));
  NOR2_X1    g07676(.A1(new_n7106_), .A2(new_n8678_), .ZN(new_n8679_));
  NOR3_X1    g07677(.A1(new_n7093_), .A2(new_n7094_), .A3(new_n7074_), .ZN(new_n8680_));
  NAND2_X1   g07678(.A1(new_n7077_), .A2(\A[109] ), .ZN(new_n8681_));
  AOI21_X1   g07679(.A1(new_n7076_), .A2(new_n8681_), .B(\A[111] ), .ZN(new_n8682_));
  OAI22_X1   g07680(.A1(new_n8680_), .A2(new_n8682_), .B1(new_n7099_), .B2(new_n7098_), .ZN(new_n8683_));
  NOR3_X1    g07681(.A1(new_n8677_), .A2(new_n8679_), .A3(new_n8683_), .ZN(new_n8684_));
  NAND2_X1   g07682(.A1(new_n7106_), .A2(new_n8678_), .ZN(new_n8685_));
  NAND2_X1   g07683(.A1(new_n7110_), .A2(new_n8676_), .ZN(new_n8686_));
  AOI21_X1   g07684(.A1(new_n8686_), .A2(new_n8685_), .B(new_n7111_), .ZN(new_n8687_));
  NOR2_X1    g07685(.A1(new_n8687_), .A2(new_n8684_), .ZN(new_n8688_));
  NOR3_X1    g07686(.A1(new_n8683_), .A2(new_n8676_), .A3(new_n8678_), .ZN(new_n8689_));
  NOR2_X1    g07687(.A1(new_n7096_), .A2(new_n7100_), .ZN(new_n8690_));
  NOR2_X1    g07688(.A1(new_n7090_), .A2(new_n7080_), .ZN(new_n8691_));
  OAI22_X1   g07689(.A1(new_n7144_), .A2(new_n7134_), .B1(new_n8690_), .B2(new_n8691_), .ZN(new_n8692_));
  NOR3_X1    g07690(.A1(new_n8688_), .A2(new_n8689_), .A3(new_n8692_), .ZN(new_n8693_));
  OAI21_X1   g07691(.A1(new_n8677_), .A2(new_n8679_), .B(new_n7111_), .ZN(new_n8694_));
  NOR2_X1    g07692(.A1(new_n8676_), .A2(new_n8678_), .ZN(new_n8695_));
  INV_X1     g07693(.I(new_n8695_), .ZN(new_n8696_));
  NAND2_X1   g07694(.A1(new_n8694_), .A2(new_n8696_), .ZN(new_n8697_));
  AOI21_X1   g07695(.A1(new_n8697_), .A2(new_n7102_), .B(new_n7153_), .ZN(new_n8698_));
  NAND2_X1   g07696(.A1(new_n8693_), .A2(new_n8698_), .ZN(new_n8699_));
  NOR2_X1    g07697(.A1(new_n8690_), .A2(new_n8691_), .ZN(new_n8700_));
  AOI21_X1   g07698(.A1(new_n8694_), .A2(new_n8696_), .B(new_n8700_), .ZN(new_n8701_));
  NAND4_X1   g07699(.A1(new_n7158_), .A2(new_n7102_), .A3(new_n7165_), .A4(new_n7112_), .ZN(new_n8702_));
  OAI21_X1   g07700(.A1(new_n8688_), .A2(new_n8701_), .B(new_n8702_), .ZN(new_n8703_));
  AOI21_X1   g07701(.A1(new_n8699_), .A2(new_n8703_), .B(new_n8674_), .ZN(new_n8704_));
  OAI21_X1   g07702(.A1(new_n8671_), .A2(new_n8670_), .B(new_n7164_), .ZN(new_n8705_));
  INV_X1     g07703(.I(new_n8668_), .ZN(new_n8706_));
  NAND2_X1   g07704(.A1(new_n8705_), .A2(new_n8706_), .ZN(new_n8707_));
  NOR2_X1    g07705(.A1(new_n8673_), .A2(new_n8672_), .ZN(new_n8708_));
  AOI21_X1   g07706(.A1(new_n7158_), .A2(new_n8707_), .B(new_n8708_), .ZN(new_n8709_));
  NAND3_X1   g07707(.A1(new_n8686_), .A2(new_n8685_), .A3(new_n7111_), .ZN(new_n8710_));
  OAI21_X1   g07708(.A1(new_n8677_), .A2(new_n8679_), .B(new_n8683_), .ZN(new_n8711_));
  NAND2_X1   g07709(.A1(new_n8711_), .A2(new_n8710_), .ZN(new_n8712_));
  AOI21_X1   g07710(.A1(new_n8686_), .A2(new_n8685_), .B(new_n8683_), .ZN(new_n8713_));
  OAI21_X1   g07711(.A1(new_n8713_), .A2(new_n8695_), .B(new_n7102_), .ZN(new_n8714_));
  NAND3_X1   g07712(.A1(new_n8702_), .A2(new_n8714_), .A3(new_n8712_), .ZN(new_n8715_));
  NOR3_X1    g07713(.A1(new_n8692_), .A2(new_n8689_), .A3(new_n7153_), .ZN(new_n8716_));
  NAND2_X1   g07714(.A1(new_n8714_), .A2(new_n8712_), .ZN(new_n8717_));
  NAND2_X1   g07715(.A1(new_n8717_), .A2(new_n8716_), .ZN(new_n8718_));
  AOI21_X1   g07716(.A1(new_n8718_), .A2(new_n8715_), .B(new_n8709_), .ZN(new_n8719_));
  NOR2_X1    g07717(.A1(new_n8704_), .A2(new_n8719_), .ZN(new_n8720_));
  AOI22_X1   g07718(.A1(new_n7167_), .A2(new_n7155_), .B1(new_n7060_), .B2(new_n7073_), .ZN(new_n8721_));
  NAND2_X1   g07719(.A1(new_n7066_), .A2(new_n7053_), .ZN(new_n8722_));
  NAND2_X1   g07720(.A1(new_n7069_), .A2(new_n7051_), .ZN(new_n8723_));
  NAND2_X1   g07721(.A1(new_n8723_), .A2(new_n8722_), .ZN(new_n8724_));
  NOR2_X1    g07722(.A1(new_n7051_), .A2(new_n7053_), .ZN(new_n8725_));
  AOI21_X1   g07723(.A1(new_n8724_), .A2(new_n7070_), .B(new_n8725_), .ZN(new_n8726_));
  NAND3_X1   g07724(.A1(new_n8723_), .A2(new_n8722_), .A3(new_n7070_), .ZN(new_n8727_));
  NOR2_X1    g07725(.A1(new_n7069_), .A2(new_n7051_), .ZN(new_n8728_));
  NOR2_X1    g07726(.A1(new_n7066_), .A2(new_n7053_), .ZN(new_n8729_));
  OAI21_X1   g07727(.A1(new_n8728_), .A2(new_n8729_), .B(new_n7057_), .ZN(new_n8730_));
  NAND2_X1   g07728(.A1(new_n8730_), .A2(new_n8727_), .ZN(new_n8731_));
  OAI21_X1   g07729(.A1(new_n7048_), .A2(new_n8726_), .B(new_n8731_), .ZN(new_n8732_));
  NOR2_X1    g07730(.A1(new_n7006_), .A2(new_n7008_), .ZN(new_n8733_));
  NOR2_X1    g07731(.A1(new_n7000_), .A2(new_n6990_), .ZN(new_n8734_));
  NOR2_X1    g07732(.A1(new_n8733_), .A2(new_n8734_), .ZN(new_n8735_));
  INV_X1     g07733(.I(new_n7012_), .ZN(new_n8736_));
  AOI21_X1   g07734(.A1(new_n7007_), .A2(\A[126] ), .B(new_n8736_), .ZN(new_n8737_));
  NOR2_X1    g07735(.A1(new_n7016_), .A2(new_n8737_), .ZN(new_n8738_));
  INV_X1     g07736(.I(new_n7015_), .ZN(new_n8739_));
  AOI21_X1   g07737(.A1(new_n6989_), .A2(\A[123] ), .B(new_n8739_), .ZN(new_n8740_));
  NOR2_X1    g07738(.A1(new_n7013_), .A2(new_n8740_), .ZN(new_n8741_));
  OAI21_X1   g07739(.A1(new_n8738_), .A2(new_n8741_), .B(new_n7017_), .ZN(new_n8742_));
  NOR2_X1    g07740(.A1(new_n8737_), .A2(new_n8740_), .ZN(new_n8743_));
  INV_X1     g07741(.I(new_n8743_), .ZN(new_n8744_));
  NAND2_X1   g07742(.A1(new_n8742_), .A2(new_n8744_), .ZN(new_n8745_));
  NOR3_X1    g07743(.A1(new_n7003_), .A2(new_n7004_), .A3(new_n6984_), .ZN(new_n8746_));
  NAND2_X1   g07744(.A1(new_n6987_), .A2(\A[121] ), .ZN(new_n8747_));
  AOI21_X1   g07745(.A1(new_n6986_), .A2(new_n8747_), .B(\A[123] ), .ZN(new_n8748_));
  NOR3_X1    g07746(.A1(new_n6997_), .A2(new_n6998_), .A3(new_n6994_), .ZN(new_n8749_));
  NAND2_X1   g07747(.A1(new_n6993_), .A2(\A[124] ), .ZN(new_n8750_));
  AOI21_X1   g07748(.A1(new_n6992_), .A2(new_n8750_), .B(\A[126] ), .ZN(new_n8751_));
  OAI22_X1   g07749(.A1(new_n8746_), .A2(new_n8748_), .B1(new_n8751_), .B2(new_n8749_), .ZN(new_n8752_));
  NOR3_X1    g07750(.A1(new_n8738_), .A2(new_n8741_), .A3(new_n8752_), .ZN(new_n8753_));
  NAND2_X1   g07751(.A1(new_n7013_), .A2(new_n8740_), .ZN(new_n8754_));
  NAND2_X1   g07752(.A1(new_n7016_), .A2(new_n8737_), .ZN(new_n8755_));
  AOI21_X1   g07753(.A1(new_n8754_), .A2(new_n8755_), .B(new_n7017_), .ZN(new_n8756_));
  NOR2_X1    g07754(.A1(new_n8756_), .A2(new_n8753_), .ZN(new_n8757_));
  NOR4_X1    g07755(.A1(new_n8757_), .A2(new_n8745_), .A3(new_n8735_), .A4(new_n7048_), .ZN(new_n8758_));
  AOI21_X1   g07756(.A1(new_n8745_), .A2(new_n7010_), .B(new_n7058_), .ZN(new_n8759_));
  NAND2_X1   g07757(.A1(new_n8758_), .A2(new_n8759_), .ZN(new_n8760_));
  AOI21_X1   g07758(.A1(new_n8742_), .A2(new_n8744_), .B(new_n8735_), .ZN(new_n8761_));
  AOI22_X1   g07759(.A1(new_n7001_), .A2(new_n7009_), .B1(new_n7062_), .B2(new_n7061_), .ZN(new_n8762_));
  NAND3_X1   g07760(.A1(new_n8762_), .A2(new_n7018_), .A3(new_n7071_), .ZN(new_n8763_));
  OAI21_X1   g07761(.A1(new_n8757_), .A2(new_n8761_), .B(new_n8763_), .ZN(new_n8764_));
  AOI21_X1   g07762(.A1(new_n8760_), .A2(new_n8764_), .B(new_n8732_), .ZN(new_n8765_));
  OAI21_X1   g07763(.A1(new_n8728_), .A2(new_n8729_), .B(new_n7070_), .ZN(new_n8766_));
  INV_X1     g07764(.I(new_n8725_), .ZN(new_n8767_));
  NAND2_X1   g07765(.A1(new_n8766_), .A2(new_n8767_), .ZN(new_n8768_));
  AOI22_X1   g07766(.A1(new_n8768_), .A2(new_n7063_), .B1(new_n8727_), .B2(new_n8730_), .ZN(new_n8769_));
  NOR3_X1    g07767(.A1(new_n8752_), .A2(new_n8737_), .A3(new_n8740_), .ZN(new_n8770_));
  NOR4_X1    g07768(.A1(new_n8735_), .A2(new_n7048_), .A3(new_n8770_), .A4(new_n7058_), .ZN(new_n8771_));
  OAI21_X1   g07769(.A1(new_n8757_), .A2(new_n8761_), .B(new_n8771_), .ZN(new_n8772_));
  NAND3_X1   g07770(.A1(new_n8754_), .A2(new_n8755_), .A3(new_n7017_), .ZN(new_n8773_));
  OAI21_X1   g07771(.A1(new_n8738_), .A2(new_n8741_), .B(new_n8752_), .ZN(new_n8774_));
  NAND2_X1   g07772(.A1(new_n8774_), .A2(new_n8773_), .ZN(new_n8775_));
  AOI21_X1   g07773(.A1(new_n8754_), .A2(new_n8755_), .B(new_n8752_), .ZN(new_n8776_));
  OAI21_X1   g07774(.A1(new_n8776_), .A2(new_n8743_), .B(new_n7010_), .ZN(new_n8777_));
  NAND3_X1   g07775(.A1(new_n8763_), .A2(new_n8777_), .A3(new_n8775_), .ZN(new_n8778_));
  AOI21_X1   g07776(.A1(new_n8772_), .A2(new_n8778_), .B(new_n8769_), .ZN(new_n8779_));
  OAI21_X1   g07777(.A1(new_n8765_), .A2(new_n8779_), .B(new_n8721_), .ZN(new_n8780_));
  NAND2_X1   g07778(.A1(new_n7168_), .A2(new_n7170_), .ZN(new_n8781_));
  NAND3_X1   g07779(.A1(new_n8775_), .A2(new_n7018_), .A3(new_n8762_), .ZN(new_n8782_));
  NOR2_X1    g07780(.A1(new_n8776_), .A2(new_n8743_), .ZN(new_n8783_));
  OAI21_X1   g07781(.A1(new_n8783_), .A2(new_n8735_), .B(new_n7071_), .ZN(new_n8784_));
  NOR2_X1    g07782(.A1(new_n8782_), .A2(new_n8784_), .ZN(new_n8785_));
  AOI21_X1   g07783(.A1(new_n8775_), .A2(new_n8777_), .B(new_n8771_), .ZN(new_n8786_));
  OAI21_X1   g07784(.A1(new_n8785_), .A2(new_n8786_), .B(new_n8769_), .ZN(new_n8787_));
  AOI21_X1   g07785(.A1(new_n8775_), .A2(new_n8777_), .B(new_n8763_), .ZN(new_n8788_));
  NOR3_X1    g07786(.A1(new_n8771_), .A2(new_n8761_), .A3(new_n8757_), .ZN(new_n8789_));
  OAI21_X1   g07787(.A1(new_n8788_), .A2(new_n8789_), .B(new_n8732_), .ZN(new_n8790_));
  NAND3_X1   g07788(.A1(new_n8787_), .A2(new_n8790_), .A3(new_n8781_), .ZN(new_n8791_));
  AOI21_X1   g07789(.A1(new_n8780_), .A2(new_n8791_), .B(new_n8720_), .ZN(new_n8792_));
  NAND4_X1   g07790(.A1(new_n8712_), .A2(new_n7102_), .A3(new_n7112_), .A4(new_n7158_), .ZN(new_n8793_));
  NAND2_X1   g07791(.A1(new_n8714_), .A2(new_n7165_), .ZN(new_n8794_));
  NOR2_X1    g07792(.A1(new_n8793_), .A2(new_n8794_), .ZN(new_n8795_));
  NOR2_X1    g07793(.A1(new_n8701_), .A2(new_n8688_), .ZN(new_n8796_));
  NOR2_X1    g07794(.A1(new_n8796_), .A2(new_n8716_), .ZN(new_n8797_));
  OAI21_X1   g07795(.A1(new_n8795_), .A2(new_n8797_), .B(new_n8709_), .ZN(new_n8798_));
  NOR2_X1    g07796(.A1(new_n8717_), .A2(new_n8716_), .ZN(new_n8799_));
  NOR2_X1    g07797(.A1(new_n8796_), .A2(new_n8702_), .ZN(new_n8800_));
  OAI21_X1   g07798(.A1(new_n8800_), .A2(new_n8799_), .B(new_n8674_), .ZN(new_n8801_));
  NAND2_X1   g07799(.A1(new_n8798_), .A2(new_n8801_), .ZN(new_n8802_));
  OAI21_X1   g07800(.A1(new_n8765_), .A2(new_n8779_), .B(new_n8781_), .ZN(new_n8803_));
  NAND3_X1   g07801(.A1(new_n8787_), .A2(new_n8790_), .A3(new_n8721_), .ZN(new_n8804_));
  AOI21_X1   g07802(.A1(new_n8803_), .A2(new_n8804_), .B(new_n8802_), .ZN(new_n8805_));
  AOI22_X1   g07803(.A1(new_n7377_), .A2(new_n7379_), .B1(new_n7169_), .B2(new_n7171_), .ZN(new_n8806_));
  INV_X1     g07804(.I(new_n8806_), .ZN(new_n8807_));
  NOR3_X1    g07805(.A1(new_n8805_), .A2(new_n8792_), .A3(new_n8807_), .ZN(new_n8808_));
  AOI21_X1   g07806(.A1(new_n8787_), .A2(new_n8790_), .B(new_n8781_), .ZN(new_n8809_));
  NOR3_X1    g07807(.A1(new_n8765_), .A2(new_n8721_), .A3(new_n8779_), .ZN(new_n8810_));
  OAI21_X1   g07808(.A1(new_n8810_), .A2(new_n8809_), .B(new_n8802_), .ZN(new_n8811_));
  AOI21_X1   g07809(.A1(new_n8787_), .A2(new_n8790_), .B(new_n8721_), .ZN(new_n8812_));
  NOR3_X1    g07810(.A1(new_n8765_), .A2(new_n8781_), .A3(new_n8779_), .ZN(new_n8813_));
  OAI21_X1   g07811(.A1(new_n8813_), .A2(new_n8812_), .B(new_n8720_), .ZN(new_n8814_));
  AOI21_X1   g07812(.A1(new_n8811_), .A2(new_n8814_), .B(new_n8806_), .ZN(new_n8815_));
  OAI21_X1   g07813(.A1(new_n8808_), .A2(new_n8815_), .B(new_n8664_), .ZN(new_n8816_));
  OAI21_X1   g07814(.A1(new_n8639_), .A2(new_n8649_), .B(new_n8660_), .ZN(new_n8817_));
  NOR3_X1    g07815(.A1(new_n8626_), .A2(new_n8637_), .A3(new_n8648_), .ZN(new_n8818_));
  AOI21_X1   g07816(.A1(new_n8644_), .A2(new_n8647_), .B(new_n8638_), .ZN(new_n8819_));
  OAI21_X1   g07817(.A1(new_n8818_), .A2(new_n8819_), .B(new_n8593_), .ZN(new_n8820_));
  NAND2_X1   g07818(.A1(new_n8820_), .A2(new_n8817_), .ZN(new_n8821_));
  NOR3_X1    g07819(.A1(new_n8805_), .A2(new_n8792_), .A3(new_n8806_), .ZN(new_n8822_));
  AOI21_X1   g07820(.A1(new_n8811_), .A2(new_n8814_), .B(new_n8807_), .ZN(new_n8823_));
  OAI21_X1   g07821(.A1(new_n8822_), .A2(new_n8823_), .B(new_n8821_), .ZN(new_n8824_));
  NAND2_X1   g07822(.A1(new_n8816_), .A2(new_n8824_), .ZN(new_n8825_));
  NAND2_X1   g07823(.A1(new_n6966_), .A2(new_n6952_), .ZN(new_n8826_));
  NAND2_X1   g07824(.A1(new_n6969_), .A2(new_n6949_), .ZN(new_n8827_));
  AOI21_X1   g07825(.A1(new_n8826_), .A2(new_n8827_), .B(new_n6953_), .ZN(new_n8828_));
  NOR2_X1    g07826(.A1(new_n6949_), .A2(new_n6952_), .ZN(new_n8829_));
  NOR2_X1    g07827(.A1(new_n8828_), .A2(new_n8829_), .ZN(new_n8830_));
  NOR2_X1    g07828(.A1(new_n6969_), .A2(new_n6949_), .ZN(new_n8831_));
  NOR2_X1    g07829(.A1(new_n6966_), .A2(new_n6952_), .ZN(new_n8832_));
  NOR3_X1    g07830(.A1(new_n8831_), .A2(new_n8832_), .A3(new_n6953_), .ZN(new_n8833_));
  AOI22_X1   g07831(.A1(new_n8826_), .A2(new_n8827_), .B1(new_n6925_), .B2(new_n6944_), .ZN(new_n8834_));
  OAI22_X1   g07832(.A1(new_n8830_), .A2(new_n6946_), .B1(new_n8833_), .B2(new_n8834_), .ZN(new_n8835_));
  NAND2_X1   g07833(.A1(new_n6888_), .A2(new_n6890_), .ZN(new_n8836_));
  AOI21_X1   g07834(.A1(new_n8836_), .A2(\A[138] ), .B(new_n6909_), .ZN(new_n8837_));
  NOR2_X1    g07835(.A1(new_n6915_), .A2(new_n8837_), .ZN(new_n8838_));
  NAND2_X1   g07836(.A1(new_n6880_), .A2(new_n6882_), .ZN(new_n8839_));
  AOI21_X1   g07837(.A1(new_n8839_), .A2(\A[135] ), .B(new_n6913_), .ZN(new_n8840_));
  NOR2_X1    g07838(.A1(new_n6911_), .A2(new_n8840_), .ZN(new_n8841_));
  OAI21_X1   g07839(.A1(new_n8841_), .A2(new_n8838_), .B(new_n6916_), .ZN(new_n8842_));
  NOR2_X1    g07840(.A1(new_n8840_), .A2(new_n8837_), .ZN(new_n8843_));
  INV_X1     g07841(.I(new_n8843_), .ZN(new_n8844_));
  NAND2_X1   g07842(.A1(new_n8842_), .A2(new_n8844_), .ZN(new_n8845_));
  OAI22_X1   g07843(.A1(new_n6884_), .A2(new_n6885_), .B1(new_n6904_), .B2(new_n6903_), .ZN(new_n8846_));
  NOR3_X1    g07844(.A1(new_n8841_), .A2(new_n8838_), .A3(new_n8846_), .ZN(new_n8847_));
  NAND2_X1   g07845(.A1(new_n6911_), .A2(new_n8840_), .ZN(new_n8848_));
  NAND2_X1   g07846(.A1(new_n6915_), .A2(new_n8837_), .ZN(new_n8849_));
  AOI21_X1   g07847(.A1(new_n8848_), .A2(new_n8849_), .B(new_n6916_), .ZN(new_n8850_));
  NOR2_X1    g07848(.A1(new_n8847_), .A2(new_n8850_), .ZN(new_n8851_));
  NOR4_X1    g07849(.A1(new_n8851_), .A2(new_n8845_), .A3(new_n6959_), .A4(new_n6946_), .ZN(new_n8852_));
  AOI21_X1   g07850(.A1(new_n8845_), .A2(new_n6907_), .B(new_n6954_), .ZN(new_n8853_));
  NAND2_X1   g07851(.A1(new_n8852_), .A2(new_n8853_), .ZN(new_n8854_));
  AOI22_X1   g07852(.A1(new_n6897_), .A2(new_n6906_), .B1(new_n6963_), .B2(new_n6962_), .ZN(new_n8855_));
  NAND3_X1   g07853(.A1(new_n8855_), .A2(new_n6917_), .A3(new_n6970_), .ZN(new_n8856_));
  AOI21_X1   g07854(.A1(new_n8848_), .A2(new_n8849_), .B(new_n8846_), .ZN(new_n8857_));
  NOR2_X1    g07855(.A1(new_n8857_), .A2(new_n8843_), .ZN(new_n8858_));
  OAI22_X1   g07856(.A1(new_n8858_), .A2(new_n6959_), .B1(new_n8847_), .B2(new_n8850_), .ZN(new_n8859_));
  NAND2_X1   g07857(.A1(new_n8859_), .A2(new_n8856_), .ZN(new_n8860_));
  AOI21_X1   g07858(.A1(new_n8854_), .A2(new_n8860_), .B(new_n8835_), .ZN(new_n8861_));
  NOR2_X1    g07859(.A1(new_n8831_), .A2(new_n8832_), .ZN(new_n8862_));
  INV_X1     g07860(.I(new_n8829_), .ZN(new_n8863_));
  OAI21_X1   g07861(.A1(new_n8862_), .A2(new_n6953_), .B(new_n8863_), .ZN(new_n8864_));
  NAND4_X1   g07862(.A1(new_n8826_), .A2(new_n8827_), .A3(new_n6925_), .A4(new_n6944_), .ZN(new_n8865_));
  OAI21_X1   g07863(.A1(new_n8831_), .A2(new_n8832_), .B(new_n6953_), .ZN(new_n8866_));
  AOI22_X1   g07864(.A1(new_n8864_), .A2(new_n6964_), .B1(new_n8865_), .B2(new_n8866_), .ZN(new_n8867_));
  NAND3_X1   g07865(.A1(new_n8848_), .A2(new_n8849_), .A3(new_n6916_), .ZN(new_n8868_));
  OAI21_X1   g07866(.A1(new_n8838_), .A2(new_n8841_), .B(new_n8846_), .ZN(new_n8869_));
  AOI22_X1   g07867(.A1(new_n8845_), .A2(new_n6907_), .B1(new_n8868_), .B2(new_n8869_), .ZN(new_n8870_));
  NAND2_X1   g07868(.A1(new_n8870_), .A2(new_n8856_), .ZN(new_n8871_));
  NOR4_X1    g07869(.A1(new_n6959_), .A2(new_n6960_), .A3(new_n6946_), .A4(new_n6954_), .ZN(new_n8872_));
  NAND2_X1   g07870(.A1(new_n8859_), .A2(new_n8872_), .ZN(new_n8873_));
  AOI21_X1   g07871(.A1(new_n8873_), .A2(new_n8871_), .B(new_n8867_), .ZN(new_n8874_));
  NOR2_X1    g07872(.A1(new_n8861_), .A2(new_n8874_), .ZN(new_n8875_));
  NAND2_X1   g07873(.A1(new_n6844_), .A2(new_n6870_), .ZN(new_n8876_));
  NAND2_X1   g07874(.A1(new_n6848_), .A2(new_n6869_), .ZN(new_n8877_));
  NAND2_X1   g07875(.A1(new_n8877_), .A2(new_n8876_), .ZN(new_n8878_));
  NOR2_X1    g07876(.A1(new_n6869_), .A2(new_n6870_), .ZN(new_n8879_));
  AOI21_X1   g07877(.A1(new_n8878_), .A2(new_n6849_), .B(new_n8879_), .ZN(new_n8880_));
  NOR2_X1    g07878(.A1(new_n6848_), .A2(new_n6869_), .ZN(new_n8881_));
  NOR2_X1    g07879(.A1(new_n6844_), .A2(new_n6870_), .ZN(new_n8882_));
  NOR3_X1    g07880(.A1(new_n8881_), .A2(new_n8882_), .A3(new_n6874_), .ZN(new_n8883_));
  AOI21_X1   g07881(.A1(new_n8877_), .A2(new_n8876_), .B(new_n6849_), .ZN(new_n8884_));
  OAI22_X1   g07882(.A1(new_n8880_), .A2(new_n6866_), .B1(new_n8883_), .B2(new_n8884_), .ZN(new_n8885_));
  NOR2_X1    g07883(.A1(new_n6860_), .A2(new_n6803_), .ZN(new_n8886_));
  NOR2_X1    g07884(.A1(new_n6858_), .A2(new_n6807_), .ZN(new_n8887_));
  NOR3_X1    g07885(.A1(new_n8887_), .A2(new_n8886_), .A3(new_n6811_), .ZN(new_n8888_));
  NAND2_X1   g07886(.A1(new_n6858_), .A2(new_n6807_), .ZN(new_n8889_));
  NAND2_X1   g07887(.A1(new_n6860_), .A2(new_n6803_), .ZN(new_n8890_));
  AOI21_X1   g07888(.A1(new_n8889_), .A2(new_n8890_), .B(new_n6861_), .ZN(new_n8891_));
  NOR2_X1    g07889(.A1(new_n8888_), .A2(new_n8891_), .ZN(new_n8892_));
  OAI22_X1   g07890(.A1(new_n6864_), .A2(new_n6865_), .B1(new_n6800_), .B2(new_n6791_), .ZN(new_n8893_));
  NOR2_X1    g07891(.A1(new_n8892_), .A2(new_n8893_), .ZN(new_n8894_));
  AOI21_X1   g07892(.A1(new_n8889_), .A2(new_n8890_), .B(new_n6811_), .ZN(new_n8895_));
  NOR2_X1    g07893(.A1(new_n6807_), .A2(new_n6803_), .ZN(new_n8896_));
  OAI21_X1   g07894(.A1(new_n8895_), .A2(new_n8896_), .B(new_n6855_), .ZN(new_n8897_));
  NAND4_X1   g07895(.A1(new_n8894_), .A2(new_n6862_), .A3(new_n6850_), .A4(new_n8897_), .ZN(new_n8898_));
  AOI22_X1   g07896(.A1(new_n6831_), .A2(new_n6840_), .B1(new_n6853_), .B2(new_n6854_), .ZN(new_n8899_));
  NAND3_X1   g07897(.A1(new_n8899_), .A2(new_n6862_), .A3(new_n6850_), .ZN(new_n8900_));
  NAND3_X1   g07898(.A1(new_n8889_), .A2(new_n8890_), .A3(new_n6861_), .ZN(new_n8901_));
  OAI21_X1   g07899(.A1(new_n8887_), .A2(new_n8886_), .B(new_n6811_), .ZN(new_n8902_));
  NAND2_X1   g07900(.A1(new_n8902_), .A2(new_n8901_), .ZN(new_n8903_));
  NAND2_X1   g07901(.A1(new_n8897_), .A2(new_n8903_), .ZN(new_n8904_));
  NAND2_X1   g07902(.A1(new_n8904_), .A2(new_n8900_), .ZN(new_n8905_));
  AOI21_X1   g07903(.A1(new_n8898_), .A2(new_n8905_), .B(new_n8885_), .ZN(new_n8906_));
  OAI21_X1   g07904(.A1(new_n8881_), .A2(new_n8882_), .B(new_n6849_), .ZN(new_n8907_));
  INV_X1     g07905(.I(new_n8879_), .ZN(new_n8908_));
  NAND2_X1   g07906(.A1(new_n8907_), .A2(new_n8908_), .ZN(new_n8909_));
  NAND3_X1   g07907(.A1(new_n8877_), .A2(new_n8876_), .A3(new_n6849_), .ZN(new_n8910_));
  OAI21_X1   g07908(.A1(new_n8881_), .A2(new_n8882_), .B(new_n6874_), .ZN(new_n8911_));
  AOI22_X1   g07909(.A1(new_n8909_), .A2(new_n6841_), .B1(new_n8910_), .B2(new_n8911_), .ZN(new_n8912_));
  NOR3_X1    g07910(.A1(new_n8893_), .A2(new_n6812_), .A3(new_n6875_), .ZN(new_n8913_));
  NAND2_X1   g07911(.A1(new_n8904_), .A2(new_n8913_), .ZN(new_n8914_));
  NAND3_X1   g07912(.A1(new_n8900_), .A2(new_n8903_), .A3(new_n8897_), .ZN(new_n8915_));
  AOI21_X1   g07913(.A1(new_n8914_), .A2(new_n8915_), .B(new_n8912_), .ZN(new_n8916_));
  NAND2_X1   g07914(.A1(new_n6973_), .A2(new_n6977_), .ZN(new_n8917_));
  NOR3_X1    g07915(.A1(new_n8906_), .A2(new_n8916_), .A3(new_n8917_), .ZN(new_n8918_));
  NAND3_X1   g07916(.A1(new_n8903_), .A2(new_n6862_), .A3(new_n8899_), .ZN(new_n8919_));
  NOR2_X1    g07917(.A1(new_n8895_), .A2(new_n8896_), .ZN(new_n8920_));
  OAI21_X1   g07918(.A1(new_n8920_), .A2(new_n6801_), .B(new_n6850_), .ZN(new_n8921_));
  NOR2_X1    g07919(.A1(new_n8919_), .A2(new_n8921_), .ZN(new_n8922_));
  AOI21_X1   g07920(.A1(new_n8903_), .A2(new_n8897_), .B(new_n8913_), .ZN(new_n8923_));
  OAI21_X1   g07921(.A1(new_n8923_), .A2(new_n8922_), .B(new_n8912_), .ZN(new_n8924_));
  AOI21_X1   g07922(.A1(new_n8903_), .A2(new_n8897_), .B(new_n8900_), .ZN(new_n8925_));
  OAI21_X1   g07923(.A1(new_n8887_), .A2(new_n8886_), .B(new_n6861_), .ZN(new_n8926_));
  INV_X1     g07924(.I(new_n8896_), .ZN(new_n8927_));
  AOI21_X1   g07925(.A1(new_n8926_), .A2(new_n8927_), .B(new_n6801_), .ZN(new_n8928_));
  NOR3_X1    g07926(.A1(new_n8913_), .A2(new_n8892_), .A3(new_n8928_), .ZN(new_n8929_));
  OAI21_X1   g07927(.A1(new_n8925_), .A2(new_n8929_), .B(new_n8885_), .ZN(new_n8930_));
  NOR2_X1    g07928(.A1(new_n6980_), .A2(new_n6878_), .ZN(new_n8931_));
  AOI21_X1   g07929(.A1(new_n8924_), .A2(new_n8930_), .B(new_n8931_), .ZN(new_n8932_));
  OAI21_X1   g07930(.A1(new_n8918_), .A2(new_n8932_), .B(new_n8875_), .ZN(new_n8933_));
  NAND2_X1   g07931(.A1(new_n8869_), .A2(new_n8868_), .ZN(new_n8934_));
  NAND3_X1   g07932(.A1(new_n8934_), .A2(new_n6917_), .A3(new_n8855_), .ZN(new_n8935_));
  OAI21_X1   g07933(.A1(new_n8858_), .A2(new_n6959_), .B(new_n6970_), .ZN(new_n8936_));
  NOR2_X1    g07934(.A1(new_n8936_), .A2(new_n8935_), .ZN(new_n8937_));
  NOR2_X1    g07935(.A1(new_n8870_), .A2(new_n8872_), .ZN(new_n8938_));
  OAI21_X1   g07936(.A1(new_n8937_), .A2(new_n8938_), .B(new_n8867_), .ZN(new_n8939_));
  NOR2_X1    g07937(.A1(new_n8858_), .A2(new_n6959_), .ZN(new_n8940_));
  NOR3_X1    g07938(.A1(new_n8940_), .A2(new_n8872_), .A3(new_n8851_), .ZN(new_n8941_));
  NOR2_X1    g07939(.A1(new_n8870_), .A2(new_n8856_), .ZN(new_n8942_));
  OAI21_X1   g07940(.A1(new_n8942_), .A2(new_n8941_), .B(new_n8835_), .ZN(new_n8943_));
  NAND2_X1   g07941(.A1(new_n8939_), .A2(new_n8943_), .ZN(new_n8944_));
  NOR3_X1    g07942(.A1(new_n8906_), .A2(new_n8916_), .A3(new_n8931_), .ZN(new_n8945_));
  AOI21_X1   g07943(.A1(new_n8924_), .A2(new_n8930_), .B(new_n8917_), .ZN(new_n8946_));
  OAI21_X1   g07944(.A1(new_n8945_), .A2(new_n8946_), .B(new_n8944_), .ZN(new_n8947_));
  NAND2_X1   g07945(.A1(new_n8933_), .A2(new_n8947_), .ZN(new_n8948_));
  NAND2_X1   g07946(.A1(new_n6763_), .A2(new_n6753_), .ZN(new_n8949_));
  NAND2_X1   g07947(.A1(new_n6765_), .A2(new_n6750_), .ZN(new_n8950_));
  AOI21_X1   g07948(.A1(new_n8949_), .A2(new_n8950_), .B(new_n6754_), .ZN(new_n8951_));
  NOR2_X1    g07949(.A1(new_n6753_), .A2(new_n6750_), .ZN(new_n8952_));
  NOR2_X1    g07950(.A1(new_n8951_), .A2(new_n8952_), .ZN(new_n8953_));
  NOR2_X1    g07951(.A1(new_n6765_), .A2(new_n6750_), .ZN(new_n8954_));
  NOR2_X1    g07952(.A1(new_n6763_), .A2(new_n6753_), .ZN(new_n8955_));
  NOR3_X1    g07953(.A1(new_n8955_), .A2(new_n8954_), .A3(new_n6754_), .ZN(new_n8956_));
  AOI22_X1   g07954(.A1(new_n8949_), .A2(new_n8950_), .B1(new_n6725_), .B2(new_n6745_), .ZN(new_n8957_));
  OAI22_X1   g07955(.A1(new_n8953_), .A2(new_n6747_), .B1(new_n8956_), .B2(new_n8957_), .ZN(new_n8958_));
  NAND2_X1   g07956(.A1(new_n6687_), .A2(new_n6689_), .ZN(new_n8959_));
  AOI21_X1   g07957(.A1(new_n8959_), .A2(\A[162] ), .B(new_n6708_), .ZN(new_n8960_));
  NOR2_X1    g07958(.A1(new_n6714_), .A2(new_n8960_), .ZN(new_n8961_));
  AOI21_X1   g07959(.A1(new_n6699_), .A2(\A[159] ), .B(new_n6712_), .ZN(new_n8962_));
  NOR2_X1    g07960(.A1(new_n6710_), .A2(new_n8962_), .ZN(new_n8963_));
  OAI22_X1   g07961(.A1(new_n6681_), .A2(new_n6684_), .B1(new_n6703_), .B2(new_n6702_), .ZN(new_n8964_));
  NOR3_X1    g07962(.A1(new_n8961_), .A2(new_n8963_), .A3(new_n8964_), .ZN(new_n8965_));
  NAND2_X1   g07963(.A1(new_n6710_), .A2(new_n8962_), .ZN(new_n8966_));
  NAND2_X1   g07964(.A1(new_n6714_), .A2(new_n8960_), .ZN(new_n8967_));
  AOI21_X1   g07965(.A1(new_n8967_), .A2(new_n8966_), .B(new_n6715_), .ZN(new_n8968_));
  NOR2_X1    g07966(.A1(new_n8968_), .A2(new_n8965_), .ZN(new_n8969_));
  NOR3_X1    g07967(.A1(new_n8964_), .A2(new_n8960_), .A3(new_n8962_), .ZN(new_n8970_));
  NOR2_X1    g07968(.A1(new_n6701_), .A2(new_n6704_), .ZN(new_n8971_));
  NOR2_X1    g07969(.A1(new_n6685_), .A2(new_n6695_), .ZN(new_n8972_));
  OAI22_X1   g07970(.A1(new_n6736_), .A2(new_n6746_), .B1(new_n8971_), .B2(new_n8972_), .ZN(new_n8973_));
  NOR3_X1    g07971(.A1(new_n8969_), .A2(new_n8970_), .A3(new_n8973_), .ZN(new_n8974_));
  OAI21_X1   g07972(.A1(new_n8961_), .A2(new_n8963_), .B(new_n6715_), .ZN(new_n8975_));
  NOR2_X1    g07973(.A1(new_n8960_), .A2(new_n8962_), .ZN(new_n8976_));
  INV_X1     g07974(.I(new_n8976_), .ZN(new_n8977_));
  NAND2_X1   g07975(.A1(new_n8975_), .A2(new_n8977_), .ZN(new_n8978_));
  AOI21_X1   g07976(.A1(new_n8978_), .A2(new_n6706_), .B(new_n6755_), .ZN(new_n8979_));
  NAND2_X1   g07977(.A1(new_n8974_), .A2(new_n8979_), .ZN(new_n8980_));
  NOR2_X1    g07978(.A1(new_n8971_), .A2(new_n8972_), .ZN(new_n8981_));
  AOI21_X1   g07979(.A1(new_n8975_), .A2(new_n8977_), .B(new_n8981_), .ZN(new_n8982_));
  NAND4_X1   g07980(.A1(new_n6761_), .A2(new_n6706_), .A3(new_n6716_), .A4(new_n6766_), .ZN(new_n8983_));
  OAI21_X1   g07981(.A1(new_n8969_), .A2(new_n8982_), .B(new_n8983_), .ZN(new_n8984_));
  AOI21_X1   g07982(.A1(new_n8980_), .A2(new_n8984_), .B(new_n8958_), .ZN(new_n8985_));
  NOR2_X1    g07983(.A1(new_n8955_), .A2(new_n8954_), .ZN(new_n8986_));
  INV_X1     g07984(.I(new_n8952_), .ZN(new_n8987_));
  OAI21_X1   g07985(.A1(new_n8986_), .A2(new_n6754_), .B(new_n8987_), .ZN(new_n8988_));
  NOR2_X1    g07986(.A1(new_n8957_), .A2(new_n8956_), .ZN(new_n8989_));
  AOI21_X1   g07987(.A1(new_n6761_), .A2(new_n8988_), .B(new_n8989_), .ZN(new_n8990_));
  NAND3_X1   g07988(.A1(new_n8967_), .A2(new_n8966_), .A3(new_n6715_), .ZN(new_n8991_));
  OAI21_X1   g07989(.A1(new_n8961_), .A2(new_n8963_), .B(new_n8964_), .ZN(new_n8992_));
  NAND2_X1   g07990(.A1(new_n8992_), .A2(new_n8991_), .ZN(new_n8993_));
  AOI21_X1   g07991(.A1(new_n8967_), .A2(new_n8966_), .B(new_n8964_), .ZN(new_n8994_));
  OAI21_X1   g07992(.A1(new_n8994_), .A2(new_n8976_), .B(new_n6706_), .ZN(new_n8995_));
  NAND3_X1   g07993(.A1(new_n8983_), .A2(new_n8995_), .A3(new_n8993_), .ZN(new_n8996_));
  NOR4_X1    g07994(.A1(new_n6747_), .A2(new_n8981_), .A3(new_n8970_), .A4(new_n6755_), .ZN(new_n8997_));
  OAI21_X1   g07995(.A1(new_n8969_), .A2(new_n8982_), .B(new_n8997_), .ZN(new_n8998_));
  AOI21_X1   g07996(.A1(new_n8998_), .A2(new_n8996_), .B(new_n8990_), .ZN(new_n8999_));
  NOR2_X1    g07997(.A1(new_n8985_), .A2(new_n8999_), .ZN(new_n9000_));
  AOI22_X1   g07998(.A1(new_n6768_), .A2(new_n6757_), .B1(new_n6652_), .B2(new_n6675_), .ZN(new_n9001_));
  NAND2_X1   g07999(.A1(new_n6668_), .A2(new_n6645_), .ZN(new_n9002_));
  NAND2_X1   g08000(.A1(new_n6671_), .A2(new_n6643_), .ZN(new_n9003_));
  NAND2_X1   g08001(.A1(new_n9003_), .A2(new_n9002_), .ZN(new_n9004_));
  NOR2_X1    g08002(.A1(new_n6643_), .A2(new_n6645_), .ZN(new_n9005_));
  AOI21_X1   g08003(.A1(new_n9004_), .A2(new_n6672_), .B(new_n9005_), .ZN(new_n9006_));
  NAND3_X1   g08004(.A1(new_n9003_), .A2(new_n9002_), .A3(new_n6672_), .ZN(new_n9007_));
  NOR2_X1    g08005(.A1(new_n6671_), .A2(new_n6643_), .ZN(new_n9008_));
  NOR2_X1    g08006(.A1(new_n6668_), .A2(new_n6645_), .ZN(new_n9009_));
  OAI21_X1   g08007(.A1(new_n9008_), .A2(new_n9009_), .B(new_n6649_), .ZN(new_n9010_));
  NAND2_X1   g08008(.A1(new_n9010_), .A2(new_n9007_), .ZN(new_n9011_));
  OAI21_X1   g08009(.A1(new_n6640_), .A2(new_n9006_), .B(new_n9011_), .ZN(new_n9012_));
  NAND2_X1   g08010(.A1(new_n6604_), .A2(new_n6656_), .ZN(new_n9013_));
  NAND2_X1   g08011(.A1(new_n6608_), .A2(new_n6654_), .ZN(new_n9014_));
  AOI21_X1   g08012(.A1(new_n9013_), .A2(new_n9014_), .B(new_n6660_), .ZN(new_n9015_));
  NOR2_X1    g08013(.A1(new_n6654_), .A2(new_n6656_), .ZN(new_n9016_));
  NOR2_X1    g08014(.A1(new_n9015_), .A2(new_n9016_), .ZN(new_n9017_));
  NAND3_X1   g08015(.A1(new_n9013_), .A2(new_n9014_), .A3(new_n6609_), .ZN(new_n9018_));
  NOR2_X1    g08016(.A1(new_n6608_), .A2(new_n6654_), .ZN(new_n9019_));
  NOR2_X1    g08017(.A1(new_n6604_), .A2(new_n6656_), .ZN(new_n9020_));
  OAI21_X1   g08018(.A1(new_n9019_), .A2(new_n9020_), .B(new_n6660_), .ZN(new_n9021_));
  NAND2_X1   g08019(.A1(new_n9021_), .A2(new_n9018_), .ZN(new_n9022_));
  NOR2_X1    g08020(.A1(new_n6653_), .A2(new_n6640_), .ZN(new_n9023_));
  OAI21_X1   g08021(.A1(new_n9019_), .A2(new_n9020_), .B(new_n6609_), .ZN(new_n9024_));
  INV_X1     g08022(.I(new_n9016_), .ZN(new_n9025_));
  NAND2_X1   g08023(.A1(new_n9024_), .A2(new_n9025_), .ZN(new_n9026_));
  AOI21_X1   g08024(.A1(new_n9026_), .A2(new_n6600_), .B(new_n6650_), .ZN(new_n9027_));
  NAND4_X1   g08025(.A1(new_n9027_), .A2(new_n9017_), .A3(new_n9022_), .A4(new_n9023_), .ZN(new_n9028_));
  NAND4_X1   g08026(.A1(new_n6665_), .A2(new_n6600_), .A3(new_n6610_), .A4(new_n6673_), .ZN(new_n9029_));
  OAI21_X1   g08027(.A1(new_n9015_), .A2(new_n9016_), .B(new_n6600_), .ZN(new_n9030_));
  NAND2_X1   g08028(.A1(new_n9030_), .A2(new_n9022_), .ZN(new_n9031_));
  NAND2_X1   g08029(.A1(new_n9031_), .A2(new_n9029_), .ZN(new_n9032_));
  AOI21_X1   g08030(.A1(new_n9028_), .A2(new_n9032_), .B(new_n9012_), .ZN(new_n9033_));
  OAI21_X1   g08031(.A1(new_n9008_), .A2(new_n9009_), .B(new_n6672_), .ZN(new_n9034_));
  INV_X1     g08032(.I(new_n9005_), .ZN(new_n9035_));
  NAND2_X1   g08033(.A1(new_n9034_), .A2(new_n9035_), .ZN(new_n9036_));
  AOI22_X1   g08034(.A1(new_n9036_), .A2(new_n6665_), .B1(new_n9007_), .B2(new_n9010_), .ZN(new_n9037_));
  NOR4_X1    g08035(.A1(new_n6653_), .A2(new_n6640_), .A3(new_n6661_), .A4(new_n6650_), .ZN(new_n9038_));
  NAND2_X1   g08036(.A1(new_n9031_), .A2(new_n9038_), .ZN(new_n9039_));
  NAND3_X1   g08037(.A1(new_n9029_), .A2(new_n9030_), .A3(new_n9022_), .ZN(new_n9040_));
  AOI21_X1   g08038(.A1(new_n9039_), .A2(new_n9040_), .B(new_n9037_), .ZN(new_n9041_));
  OAI21_X1   g08039(.A1(new_n9033_), .A2(new_n9041_), .B(new_n9001_), .ZN(new_n9042_));
  NOR2_X1    g08040(.A1(new_n6662_), .A2(new_n6674_), .ZN(new_n9043_));
  NOR2_X1    g08041(.A1(new_n6651_), .A2(new_n6611_), .ZN(new_n9044_));
  NOR2_X1    g08042(.A1(new_n6758_), .A2(new_n6767_), .ZN(new_n9045_));
  NOR2_X1    g08043(.A1(new_n6756_), .A2(new_n6717_), .ZN(new_n9046_));
  OAI22_X1   g08044(.A1(new_n9045_), .A2(new_n9046_), .B1(new_n9043_), .B2(new_n9044_), .ZN(new_n9047_));
  NAND4_X1   g08045(.A1(new_n9022_), .A2(new_n6600_), .A3(new_n6610_), .A4(new_n6665_), .ZN(new_n9048_));
  OAI21_X1   g08046(.A1(new_n9017_), .A2(new_n6653_), .B(new_n6673_), .ZN(new_n9049_));
  NOR2_X1    g08047(.A1(new_n9048_), .A2(new_n9049_), .ZN(new_n9050_));
  AOI21_X1   g08048(.A1(new_n9022_), .A2(new_n9030_), .B(new_n9038_), .ZN(new_n9051_));
  OAI21_X1   g08049(.A1(new_n9050_), .A2(new_n9051_), .B(new_n9037_), .ZN(new_n9052_));
  AOI21_X1   g08050(.A1(new_n9022_), .A2(new_n9030_), .B(new_n9029_), .ZN(new_n9053_));
  NOR3_X1    g08051(.A1(new_n9019_), .A2(new_n9020_), .A3(new_n6660_), .ZN(new_n9054_));
  AOI21_X1   g08052(.A1(new_n9013_), .A2(new_n9014_), .B(new_n6609_), .ZN(new_n9055_));
  NOR2_X1    g08053(.A1(new_n9055_), .A2(new_n9054_), .ZN(new_n9056_));
  AOI21_X1   g08054(.A1(new_n9024_), .A2(new_n9025_), .B(new_n6653_), .ZN(new_n9057_));
  NOR3_X1    g08055(.A1(new_n9057_), .A2(new_n9038_), .A3(new_n9056_), .ZN(new_n9058_));
  OAI21_X1   g08056(.A1(new_n9058_), .A2(new_n9053_), .B(new_n9012_), .ZN(new_n9059_));
  NAND3_X1   g08057(.A1(new_n9052_), .A2(new_n9059_), .A3(new_n9047_), .ZN(new_n9060_));
  AOI21_X1   g08058(.A1(new_n9042_), .A2(new_n9060_), .B(new_n9000_), .ZN(new_n9061_));
  NAND4_X1   g08059(.A1(new_n8993_), .A2(new_n6706_), .A3(new_n6716_), .A4(new_n6761_), .ZN(new_n9062_));
  NOR3_X1    g08060(.A1(new_n9062_), .A2(new_n6755_), .A3(new_n8982_), .ZN(new_n9063_));
  AOI21_X1   g08061(.A1(new_n8993_), .A2(new_n8995_), .B(new_n8997_), .ZN(new_n9064_));
  OAI21_X1   g08062(.A1(new_n9063_), .A2(new_n9064_), .B(new_n8990_), .ZN(new_n9065_));
  NOR3_X1    g08063(.A1(new_n8997_), .A2(new_n8982_), .A3(new_n8969_), .ZN(new_n9066_));
  AOI21_X1   g08064(.A1(new_n8993_), .A2(new_n8995_), .B(new_n8983_), .ZN(new_n9067_));
  OAI21_X1   g08065(.A1(new_n9067_), .A2(new_n9066_), .B(new_n8958_), .ZN(new_n9068_));
  NAND2_X1   g08066(.A1(new_n9065_), .A2(new_n9068_), .ZN(new_n9069_));
  OAI21_X1   g08067(.A1(new_n9033_), .A2(new_n9041_), .B(new_n9047_), .ZN(new_n9070_));
  NAND3_X1   g08068(.A1(new_n9052_), .A2(new_n9059_), .A3(new_n9001_), .ZN(new_n9071_));
  AOI21_X1   g08069(.A1(new_n9070_), .A2(new_n9071_), .B(new_n9069_), .ZN(new_n9072_));
  AOI22_X1   g08070(.A1(new_n6770_), .A2(new_n6772_), .B1(new_n6974_), .B2(new_n6981_), .ZN(new_n9073_));
  NOR3_X1    g08071(.A1(new_n9072_), .A2(new_n9061_), .A3(new_n9073_), .ZN(new_n9074_));
  AOI21_X1   g08072(.A1(new_n9052_), .A2(new_n9059_), .B(new_n9047_), .ZN(new_n9075_));
  NOR3_X1    g08073(.A1(new_n9033_), .A2(new_n9041_), .A3(new_n9001_), .ZN(new_n9076_));
  OAI21_X1   g08074(.A1(new_n9076_), .A2(new_n9075_), .B(new_n9069_), .ZN(new_n9077_));
  AOI21_X1   g08075(.A1(new_n9052_), .A2(new_n9059_), .B(new_n9001_), .ZN(new_n9078_));
  NOR3_X1    g08076(.A1(new_n9033_), .A2(new_n9041_), .A3(new_n9047_), .ZN(new_n9079_));
  OAI21_X1   g08077(.A1(new_n9079_), .A2(new_n9078_), .B(new_n9000_), .ZN(new_n9080_));
  INV_X1     g08078(.I(new_n9073_), .ZN(new_n9081_));
  AOI21_X1   g08079(.A1(new_n9077_), .A2(new_n9080_), .B(new_n9081_), .ZN(new_n9082_));
  OAI21_X1   g08080(.A1(new_n9082_), .A2(new_n9074_), .B(new_n8948_), .ZN(new_n9083_));
  NAND2_X1   g08081(.A1(new_n6983_), .A2(new_n7381_), .ZN(new_n9084_));
  NAND3_X1   g08082(.A1(new_n8924_), .A2(new_n8931_), .A3(new_n8930_), .ZN(new_n9085_));
  OAI21_X1   g08083(.A1(new_n8906_), .A2(new_n8916_), .B(new_n8917_), .ZN(new_n9086_));
  AOI21_X1   g08084(.A1(new_n9086_), .A2(new_n9085_), .B(new_n8944_), .ZN(new_n9087_));
  NAND3_X1   g08085(.A1(new_n8924_), .A2(new_n8930_), .A3(new_n8917_), .ZN(new_n9088_));
  OAI21_X1   g08086(.A1(new_n8906_), .A2(new_n8916_), .B(new_n8931_), .ZN(new_n9089_));
  AOI21_X1   g08087(.A1(new_n9088_), .A2(new_n9089_), .B(new_n8875_), .ZN(new_n9090_));
  NOR2_X1    g08088(.A1(new_n9090_), .A2(new_n9087_), .ZN(new_n9091_));
  NOR3_X1    g08089(.A1(new_n9072_), .A2(new_n9061_), .A3(new_n9081_), .ZN(new_n9092_));
  AOI21_X1   g08090(.A1(new_n9077_), .A2(new_n9080_), .B(new_n9073_), .ZN(new_n9093_));
  OAI21_X1   g08091(.A1(new_n9092_), .A2(new_n9093_), .B(new_n9091_), .ZN(new_n9094_));
  INV_X1     g08092(.I(new_n9094_), .ZN(new_n9095_));
  NOR2_X1    g08093(.A1(new_n9095_), .A2(new_n9084_), .ZN(new_n9096_));
  NAND2_X1   g08094(.A1(new_n9094_), .A2(new_n9083_), .ZN(new_n9097_));
  AOI22_X1   g08095(.A1(new_n9096_), .A2(new_n9083_), .B1(new_n9084_), .B2(new_n9097_), .ZN(new_n9098_));
  NAND3_X1   g08096(.A1(new_n9094_), .A2(new_n9083_), .A3(new_n9084_), .ZN(new_n9099_));
  INV_X1     g08097(.I(new_n9084_), .ZN(new_n9100_));
  NAND2_X1   g08098(.A1(new_n9097_), .A2(new_n9100_), .ZN(new_n9101_));
  NAND2_X1   g08099(.A1(new_n9101_), .A2(new_n9099_), .ZN(new_n9102_));
  NAND2_X1   g08100(.A1(new_n9102_), .A2(new_n8825_), .ZN(new_n9103_));
  OAI21_X1   g08101(.A1(new_n8825_), .A2(new_n9098_), .B(new_n9103_), .ZN(new_n9104_));
  NOR2_X1    g08102(.A1(new_n6571_), .A2(new_n7382_), .ZN(new_n9105_));
  INV_X1     g08103(.I(new_n9105_), .ZN(new_n9106_));
  NOR2_X1    g08104(.A1(new_n6125_), .A2(new_n6127_), .ZN(new_n9107_));
  INV_X1     g08105(.I(new_n6144_), .ZN(new_n9108_));
  OAI21_X1   g08106(.A1(new_n9107_), .A2(new_n6123_), .B(new_n9108_), .ZN(new_n9109_));
  NAND2_X1   g08107(.A1(new_n9109_), .A2(new_n6148_), .ZN(new_n9110_));
  NOR2_X1    g08108(.A1(new_n6119_), .A2(new_n6120_), .ZN(new_n9111_));
  INV_X1     g08109(.I(new_n6147_), .ZN(new_n9112_));
  OAI21_X1   g08110(.A1(new_n9111_), .A2(new_n6116_), .B(new_n9112_), .ZN(new_n9113_));
  NAND2_X1   g08111(.A1(new_n9113_), .A2(new_n6145_), .ZN(new_n9114_));
  NAND2_X1   g08112(.A1(new_n9110_), .A2(new_n9114_), .ZN(new_n9115_));
  AOI22_X1   g08113(.A1(new_n6118_), .A2(new_n6121_), .B1(new_n6139_), .B2(new_n6138_), .ZN(new_n9116_));
  NOR2_X1    g08114(.A1(new_n6148_), .A2(new_n6145_), .ZN(new_n9117_));
  AOI21_X1   g08115(.A1(new_n9115_), .A2(new_n9116_), .B(new_n9117_), .ZN(new_n9118_));
  NAND3_X1   g08116(.A1(new_n9110_), .A2(new_n9114_), .A3(new_n9116_), .ZN(new_n9119_));
  NOR2_X1    g08117(.A1(new_n9113_), .A2(new_n6145_), .ZN(new_n9120_));
  NOR2_X1    g08118(.A1(new_n9109_), .A2(new_n6148_), .ZN(new_n9121_));
  OAI21_X1   g08119(.A1(new_n9120_), .A2(new_n9121_), .B(new_n6149_), .ZN(new_n9122_));
  NAND2_X1   g08120(.A1(new_n9122_), .A2(new_n9119_), .ZN(new_n9123_));
  OAI21_X1   g08121(.A1(new_n6142_), .A2(new_n9118_), .B(new_n9123_), .ZN(new_n9124_));
  NOR2_X1    g08122(.A1(new_n6109_), .A2(new_n6157_), .ZN(new_n9125_));
  NOR2_X1    g08123(.A1(new_n6105_), .A2(new_n6159_), .ZN(new_n9126_));
  OAI21_X1   g08124(.A1(new_n9125_), .A2(new_n9126_), .B(new_n6110_), .ZN(new_n9127_));
  NOR2_X1    g08125(.A1(new_n6157_), .A2(new_n6159_), .ZN(new_n9128_));
  INV_X1     g08126(.I(new_n9128_), .ZN(new_n9129_));
  NAND2_X1   g08127(.A1(new_n9127_), .A2(new_n9129_), .ZN(new_n9130_));
  NOR3_X1    g08128(.A1(new_n9125_), .A2(new_n9126_), .A3(new_n6160_), .ZN(new_n9131_));
  NAND2_X1   g08129(.A1(new_n6105_), .A2(new_n6159_), .ZN(new_n9132_));
  NAND2_X1   g08130(.A1(new_n6109_), .A2(new_n6157_), .ZN(new_n9133_));
  AOI21_X1   g08131(.A1(new_n9132_), .A2(new_n9133_), .B(new_n6110_), .ZN(new_n9134_));
  NOR2_X1    g08132(.A1(new_n9134_), .A2(new_n9131_), .ZN(new_n9135_));
  NOR4_X1    g08133(.A1(new_n9135_), .A2(new_n9130_), .A3(new_n6155_), .A4(new_n6142_), .ZN(new_n9136_));
  AOI21_X1   g08134(.A1(new_n9130_), .A2(new_n6101_), .B(new_n6150_), .ZN(new_n9137_));
  NAND2_X1   g08135(.A1(new_n9136_), .A2(new_n9137_), .ZN(new_n9138_));
  INV_X1     g08136(.I(new_n6150_), .ZN(new_n9139_));
  NAND2_X1   g08137(.A1(new_n6137_), .A2(new_n6140_), .ZN(new_n9140_));
  NAND2_X1   g08138(.A1(new_n6132_), .A2(new_n6122_), .ZN(new_n9141_));
  AOI22_X1   g08139(.A1(new_n9140_), .A2(new_n9141_), .B1(new_n6100_), .B2(new_n6092_), .ZN(new_n9142_));
  NAND3_X1   g08140(.A1(new_n9142_), .A2(new_n9139_), .A3(new_n6111_), .ZN(new_n9143_));
  NAND3_X1   g08141(.A1(new_n9132_), .A2(new_n9133_), .A3(new_n6110_), .ZN(new_n9144_));
  OAI21_X1   g08142(.A1(new_n9125_), .A2(new_n9126_), .B(new_n6160_), .ZN(new_n9145_));
  NAND2_X1   g08143(.A1(new_n9145_), .A2(new_n9144_), .ZN(new_n9146_));
  AOI21_X1   g08144(.A1(new_n9132_), .A2(new_n9133_), .B(new_n6160_), .ZN(new_n9147_));
  OAI21_X1   g08145(.A1(new_n9147_), .A2(new_n9128_), .B(new_n6101_), .ZN(new_n9148_));
  NAND2_X1   g08146(.A1(new_n9148_), .A2(new_n9146_), .ZN(new_n9149_));
  NAND2_X1   g08147(.A1(new_n9149_), .A2(new_n9143_), .ZN(new_n9150_));
  AOI21_X1   g08148(.A1(new_n9138_), .A2(new_n9150_), .B(new_n9124_), .ZN(new_n9151_));
  INV_X1     g08149(.I(new_n6142_), .ZN(new_n9152_));
  OAI21_X1   g08150(.A1(new_n9121_), .A2(new_n9120_), .B(new_n9116_), .ZN(new_n9153_));
  INV_X1     g08151(.I(new_n9117_), .ZN(new_n9154_));
  NAND2_X1   g08152(.A1(new_n9153_), .A2(new_n9154_), .ZN(new_n9155_));
  AOI22_X1   g08153(.A1(new_n9155_), .A2(new_n9152_), .B1(new_n9119_), .B2(new_n9122_), .ZN(new_n9156_));
  NAND3_X1   g08154(.A1(new_n9143_), .A2(new_n9148_), .A3(new_n9146_), .ZN(new_n9157_));
  NOR4_X1    g08155(.A1(new_n6142_), .A2(new_n6155_), .A3(new_n6161_), .A4(new_n6150_), .ZN(new_n9158_));
  NAND2_X1   g08156(.A1(new_n9149_), .A2(new_n9158_), .ZN(new_n9159_));
  AOI21_X1   g08157(.A1(new_n9159_), .A2(new_n9157_), .B(new_n9156_), .ZN(new_n9160_));
  NOR2_X1    g08158(.A1(new_n9151_), .A2(new_n9160_), .ZN(new_n9161_));
  NAND2_X1   g08159(.A1(new_n6064_), .A2(new_n6039_), .ZN(new_n9162_));
  NAND2_X1   g08160(.A1(new_n6067_), .A2(new_n6036_), .ZN(new_n9163_));
  NAND2_X1   g08161(.A1(new_n9162_), .A2(new_n9163_), .ZN(new_n9164_));
  NOR2_X1    g08162(.A1(new_n6036_), .A2(new_n6039_), .ZN(new_n9165_));
  AOI21_X1   g08163(.A1(new_n9164_), .A2(new_n6068_), .B(new_n9165_), .ZN(new_n9166_));
  NOR2_X1    g08164(.A1(new_n6067_), .A2(new_n6036_), .ZN(new_n9167_));
  NOR2_X1    g08165(.A1(new_n6064_), .A2(new_n6039_), .ZN(new_n9168_));
  NOR3_X1    g08166(.A1(new_n9167_), .A2(new_n9168_), .A3(new_n6040_), .ZN(new_n9169_));
  AOI21_X1   g08167(.A1(new_n9162_), .A2(new_n9163_), .B(new_n6068_), .ZN(new_n9170_));
  OAI22_X1   g08168(.A1(new_n9166_), .A2(new_n6033_), .B1(new_n9169_), .B2(new_n9170_), .ZN(new_n9171_));
  NAND2_X1   g08169(.A1(new_n5997_), .A2(new_n6049_), .ZN(new_n9172_));
  NAND2_X1   g08170(.A1(new_n6000_), .A2(new_n6047_), .ZN(new_n9173_));
  AOI21_X1   g08171(.A1(new_n9172_), .A2(new_n9173_), .B(new_n6056_), .ZN(new_n9174_));
  NOR2_X1    g08172(.A1(new_n6047_), .A2(new_n6049_), .ZN(new_n9175_));
  NOR2_X1    g08173(.A1(new_n9174_), .A2(new_n9175_), .ZN(new_n9176_));
  NAND3_X1   g08174(.A1(new_n9172_), .A2(new_n9173_), .A3(new_n6001_), .ZN(new_n9177_));
  NOR2_X1    g08175(.A1(new_n6000_), .A2(new_n6047_), .ZN(new_n9178_));
  NOR2_X1    g08176(.A1(new_n5997_), .A2(new_n6049_), .ZN(new_n9179_));
  OAI21_X1   g08177(.A1(new_n9179_), .A2(new_n9178_), .B(new_n6056_), .ZN(new_n9180_));
  NAND2_X1   g08178(.A1(new_n9180_), .A2(new_n9177_), .ZN(new_n9181_));
  AOI22_X1   g08179(.A1(new_n6059_), .A2(new_n6060_), .B1(new_n5984_), .B2(new_n5992_), .ZN(new_n9182_));
  OAI21_X1   g08180(.A1(new_n9179_), .A2(new_n9178_), .B(new_n6001_), .ZN(new_n9183_));
  INV_X1     g08181(.I(new_n9175_), .ZN(new_n9184_));
  NAND2_X1   g08182(.A1(new_n9183_), .A2(new_n9184_), .ZN(new_n9185_));
  AOI21_X1   g08183(.A1(new_n9185_), .A2(new_n5993_), .B(new_n6041_), .ZN(new_n9186_));
  NAND4_X1   g08184(.A1(new_n9186_), .A2(new_n9176_), .A3(new_n9181_), .A4(new_n9182_), .ZN(new_n9187_));
  NAND3_X1   g08185(.A1(new_n9182_), .A2(new_n6002_), .A3(new_n6069_), .ZN(new_n9188_));
  OAI21_X1   g08186(.A1(new_n9174_), .A2(new_n9175_), .B(new_n5993_), .ZN(new_n9189_));
  NAND2_X1   g08187(.A1(new_n9189_), .A2(new_n9181_), .ZN(new_n9190_));
  NAND2_X1   g08188(.A1(new_n9190_), .A2(new_n9188_), .ZN(new_n9191_));
  AOI21_X1   g08189(.A1(new_n9187_), .A2(new_n9191_), .B(new_n9171_), .ZN(new_n9192_));
  OAI21_X1   g08190(.A1(new_n9167_), .A2(new_n9168_), .B(new_n6068_), .ZN(new_n9193_));
  INV_X1     g08191(.I(new_n9165_), .ZN(new_n9194_));
  NAND2_X1   g08192(.A1(new_n9193_), .A2(new_n9194_), .ZN(new_n9195_));
  NAND3_X1   g08193(.A1(new_n9162_), .A2(new_n9163_), .A3(new_n6068_), .ZN(new_n9196_));
  OAI21_X1   g08194(.A1(new_n9167_), .A2(new_n9168_), .B(new_n6040_), .ZN(new_n9197_));
  AOI22_X1   g08195(.A1(new_n9195_), .A2(new_n6061_), .B1(new_n9196_), .B2(new_n9197_), .ZN(new_n9198_));
  NOR4_X1    g08196(.A1(new_n6033_), .A2(new_n6046_), .A3(new_n6057_), .A4(new_n6041_), .ZN(new_n9199_));
  NAND2_X1   g08197(.A1(new_n9190_), .A2(new_n9199_), .ZN(new_n9200_));
  NAND3_X1   g08198(.A1(new_n9188_), .A2(new_n9189_), .A3(new_n9181_), .ZN(new_n9201_));
  AOI21_X1   g08199(.A1(new_n9200_), .A2(new_n9201_), .B(new_n9198_), .ZN(new_n9202_));
  NOR2_X1    g08200(.A1(new_n6070_), .A2(new_n6058_), .ZN(new_n9203_));
  NOR2_X1    g08201(.A1(new_n6042_), .A2(new_n6003_), .ZN(new_n9204_));
  NOR2_X1    g08202(.A1(new_n6163_), .A2(new_n6162_), .ZN(new_n9205_));
  NOR2_X1    g08203(.A1(new_n6151_), .A2(new_n6112_), .ZN(new_n9206_));
  OAI22_X1   g08204(.A1(new_n9205_), .A2(new_n9206_), .B1(new_n9203_), .B2(new_n9204_), .ZN(new_n9207_));
  NOR3_X1    g08205(.A1(new_n9192_), .A2(new_n9202_), .A3(new_n9207_), .ZN(new_n9208_));
  NAND3_X1   g08206(.A1(new_n9181_), .A2(new_n6002_), .A3(new_n9182_), .ZN(new_n9209_));
  OAI21_X1   g08207(.A1(new_n9176_), .A2(new_n6046_), .B(new_n6069_), .ZN(new_n9210_));
  NOR2_X1    g08208(.A1(new_n9209_), .A2(new_n9210_), .ZN(new_n9211_));
  AOI21_X1   g08209(.A1(new_n9181_), .A2(new_n9189_), .B(new_n9199_), .ZN(new_n9212_));
  OAI21_X1   g08210(.A1(new_n9211_), .A2(new_n9212_), .B(new_n9198_), .ZN(new_n9213_));
  AOI21_X1   g08211(.A1(new_n9181_), .A2(new_n9189_), .B(new_n9188_), .ZN(new_n9214_));
  NOR3_X1    g08212(.A1(new_n9179_), .A2(new_n9178_), .A3(new_n6056_), .ZN(new_n9215_));
  AOI21_X1   g08213(.A1(new_n9172_), .A2(new_n9173_), .B(new_n6001_), .ZN(new_n9216_));
  NOR2_X1    g08214(.A1(new_n9216_), .A2(new_n9215_), .ZN(new_n9217_));
  AOI21_X1   g08215(.A1(new_n9183_), .A2(new_n9184_), .B(new_n6046_), .ZN(new_n9218_));
  NOR3_X1    g08216(.A1(new_n9199_), .A2(new_n9218_), .A3(new_n9217_), .ZN(new_n9219_));
  OAI21_X1   g08217(.A1(new_n9214_), .A2(new_n9219_), .B(new_n9171_), .ZN(new_n9220_));
  AOI22_X1   g08218(.A1(new_n6164_), .A2(new_n6152_), .B1(new_n6043_), .B2(new_n6071_), .ZN(new_n9221_));
  AOI21_X1   g08219(.A1(new_n9213_), .A2(new_n9220_), .B(new_n9221_), .ZN(new_n9222_));
  OAI21_X1   g08220(.A1(new_n9208_), .A2(new_n9222_), .B(new_n9161_), .ZN(new_n9223_));
  NAND3_X1   g08221(.A1(new_n9146_), .A2(new_n6111_), .A3(new_n9142_), .ZN(new_n9224_));
  NOR2_X1    g08222(.A1(new_n9147_), .A2(new_n9128_), .ZN(new_n9225_));
  OAI21_X1   g08223(.A1(new_n9225_), .A2(new_n6155_), .B(new_n9139_), .ZN(new_n9226_));
  NOR2_X1    g08224(.A1(new_n9224_), .A2(new_n9226_), .ZN(new_n9227_));
  AOI21_X1   g08225(.A1(new_n9146_), .A2(new_n9148_), .B(new_n9158_), .ZN(new_n9228_));
  OAI21_X1   g08226(.A1(new_n9227_), .A2(new_n9228_), .B(new_n9156_), .ZN(new_n9229_));
  AOI21_X1   g08227(.A1(new_n9127_), .A2(new_n9129_), .B(new_n6155_), .ZN(new_n9230_));
  NOR3_X1    g08228(.A1(new_n9158_), .A2(new_n9230_), .A3(new_n9135_), .ZN(new_n9231_));
  AOI21_X1   g08229(.A1(new_n9146_), .A2(new_n9148_), .B(new_n9143_), .ZN(new_n9232_));
  OAI21_X1   g08230(.A1(new_n9232_), .A2(new_n9231_), .B(new_n9124_), .ZN(new_n9233_));
  NAND2_X1   g08231(.A1(new_n9229_), .A2(new_n9233_), .ZN(new_n9234_));
  NOR3_X1    g08232(.A1(new_n9192_), .A2(new_n9202_), .A3(new_n9221_), .ZN(new_n9235_));
  AOI21_X1   g08233(.A1(new_n9213_), .A2(new_n9220_), .B(new_n9207_), .ZN(new_n9236_));
  OAI21_X1   g08234(.A1(new_n9235_), .A2(new_n9236_), .B(new_n9234_), .ZN(new_n9237_));
  NAND2_X1   g08235(.A1(new_n9223_), .A2(new_n9237_), .ZN(new_n9238_));
  NAND2_X1   g08236(.A1(new_n6169_), .A2(new_n5966_), .ZN(new_n9239_));
  NOR2_X1    g08237(.A1(new_n5936_), .A2(new_n5957_), .ZN(new_n9240_));
  NOR2_X1    g08238(.A1(new_n5932_), .A2(new_n5958_), .ZN(new_n9241_));
  OAI21_X1   g08239(.A1(new_n9240_), .A2(new_n9241_), .B(new_n5937_), .ZN(new_n9242_));
  NOR2_X1    g08240(.A1(new_n5957_), .A2(new_n5958_), .ZN(new_n9243_));
  INV_X1     g08241(.I(new_n9243_), .ZN(new_n9244_));
  NAND2_X1   g08242(.A1(new_n9242_), .A2(new_n9244_), .ZN(new_n9245_));
  NAND2_X1   g08243(.A1(new_n5932_), .A2(new_n5958_), .ZN(new_n9246_));
  NAND2_X1   g08244(.A1(new_n5936_), .A2(new_n5957_), .ZN(new_n9247_));
  NAND3_X1   g08245(.A1(new_n9246_), .A2(new_n9247_), .A3(new_n5937_), .ZN(new_n9248_));
  OAI21_X1   g08246(.A1(new_n9240_), .A2(new_n9241_), .B(new_n5959_), .ZN(new_n9249_));
  AOI22_X1   g08247(.A1(new_n9245_), .A2(new_n5928_), .B1(new_n9248_), .B2(new_n9249_), .ZN(new_n9250_));
  NOR2_X1    g08248(.A1(new_n5946_), .A2(new_n5864_), .ZN(new_n9251_));
  NOR2_X1    g08249(.A1(new_n5943_), .A2(new_n5869_), .ZN(new_n9252_));
  OAI21_X1   g08250(.A1(new_n9251_), .A2(new_n9252_), .B(new_n5883_), .ZN(new_n9253_));
  NAND2_X1   g08251(.A1(new_n5943_), .A2(new_n5869_), .ZN(new_n9254_));
  NAND2_X1   g08252(.A1(new_n5946_), .A2(new_n5864_), .ZN(new_n9255_));
  NAND3_X1   g08253(.A1(new_n9254_), .A2(new_n9255_), .A3(new_n5949_), .ZN(new_n9256_));
  NAND2_X1   g08254(.A1(new_n9253_), .A2(new_n9256_), .ZN(new_n9257_));
  AOI22_X1   g08255(.A1(new_n5927_), .A2(new_n5918_), .B1(new_n5952_), .B2(new_n5951_), .ZN(new_n9258_));
  NAND3_X1   g08256(.A1(new_n9258_), .A2(new_n5950_), .A3(new_n5938_), .ZN(new_n9259_));
  NOR2_X1    g08257(.A1(new_n5864_), .A2(new_n5869_), .ZN(new_n9260_));
  AOI21_X1   g08258(.A1(new_n9254_), .A2(new_n9255_), .B(new_n5883_), .ZN(new_n9261_));
  OAI21_X1   g08259(.A1(new_n9260_), .A2(new_n9261_), .B(new_n5953_), .ZN(new_n9262_));
  NAND3_X1   g08260(.A1(new_n9259_), .A2(new_n9262_), .A3(new_n9257_), .ZN(new_n9263_));
  NOR4_X1    g08261(.A1(new_n5955_), .A2(new_n5896_), .A3(new_n5884_), .A4(new_n5960_), .ZN(new_n9264_));
  NAND2_X1   g08262(.A1(new_n9262_), .A2(new_n9257_), .ZN(new_n9265_));
  NAND2_X1   g08263(.A1(new_n9265_), .A2(new_n9264_), .ZN(new_n9266_));
  AOI21_X1   g08264(.A1(new_n9266_), .A2(new_n9263_), .B(new_n9250_), .ZN(new_n9267_));
  NAND2_X1   g08265(.A1(new_n9246_), .A2(new_n9247_), .ZN(new_n9268_));
  AOI21_X1   g08266(.A1(new_n9268_), .A2(new_n5937_), .B(new_n9243_), .ZN(new_n9269_));
  NOR3_X1    g08267(.A1(new_n9240_), .A2(new_n9241_), .A3(new_n5959_), .ZN(new_n9270_));
  AOI21_X1   g08268(.A1(new_n9246_), .A2(new_n9247_), .B(new_n5937_), .ZN(new_n9271_));
  OAI22_X1   g08269(.A1(new_n9269_), .A2(new_n5955_), .B1(new_n9270_), .B2(new_n9271_), .ZN(new_n9272_));
  INV_X1     g08270(.I(new_n9260_), .ZN(new_n9273_));
  OAI21_X1   g08271(.A1(new_n9251_), .A2(new_n9252_), .B(new_n5949_), .ZN(new_n9274_));
  NAND2_X1   g08272(.A1(new_n9274_), .A2(new_n9273_), .ZN(new_n9275_));
  AOI21_X1   g08273(.A1(new_n9254_), .A2(new_n9255_), .B(new_n5949_), .ZN(new_n9276_));
  NOR3_X1    g08274(.A1(new_n9251_), .A2(new_n9252_), .A3(new_n5883_), .ZN(new_n9277_));
  NOR2_X1    g08275(.A1(new_n9276_), .A2(new_n9277_), .ZN(new_n9278_));
  NOR4_X1    g08276(.A1(new_n9278_), .A2(new_n9275_), .A3(new_n5896_), .A4(new_n5955_), .ZN(new_n9279_));
  AOI21_X1   g08277(.A1(new_n9275_), .A2(new_n5953_), .B(new_n5960_), .ZN(new_n9280_));
  NAND2_X1   g08278(.A1(new_n9279_), .A2(new_n9280_), .ZN(new_n9281_));
  NAND2_X1   g08279(.A1(new_n9265_), .A2(new_n9259_), .ZN(new_n9282_));
  AOI21_X1   g08280(.A1(new_n9281_), .A2(new_n9282_), .B(new_n9272_), .ZN(new_n9283_));
  NOR2_X1    g08281(.A1(new_n9283_), .A2(new_n9267_), .ZN(new_n9284_));
  NAND2_X1   g08282(.A1(new_n5851_), .A2(new_n5830_), .ZN(new_n9285_));
  NAND2_X1   g08283(.A1(new_n5854_), .A2(new_n5827_), .ZN(new_n9286_));
  NAND2_X1   g08284(.A1(new_n9286_), .A2(new_n9285_), .ZN(new_n9287_));
  NOR2_X1    g08285(.A1(new_n5827_), .A2(new_n5830_), .ZN(new_n9288_));
  AOI21_X1   g08286(.A1(new_n9287_), .A2(new_n5855_), .B(new_n9288_), .ZN(new_n9289_));
  NOR2_X1    g08287(.A1(new_n5854_), .A2(new_n5827_), .ZN(new_n9290_));
  NOR2_X1    g08288(.A1(new_n5851_), .A2(new_n5830_), .ZN(new_n9291_));
  NOR3_X1    g08289(.A1(new_n9290_), .A2(new_n9291_), .A3(new_n5831_), .ZN(new_n9292_));
  AOI21_X1   g08290(.A1(new_n9286_), .A2(new_n9285_), .B(new_n5855_), .ZN(new_n9293_));
  OAI22_X1   g08291(.A1(new_n9289_), .A2(new_n5823_), .B1(new_n9292_), .B2(new_n9293_), .ZN(new_n9294_));
  NAND2_X1   g08292(.A1(new_n5756_), .A2(new_n5840_), .ZN(new_n9295_));
  NAND2_X1   g08293(.A1(new_n5760_), .A2(new_n5837_), .ZN(new_n9296_));
  AOI21_X1   g08294(.A1(new_n9295_), .A2(new_n9296_), .B(new_n5777_), .ZN(new_n9297_));
  NOR2_X1    g08295(.A1(new_n5760_), .A2(new_n5837_), .ZN(new_n9298_));
  NOR2_X1    g08296(.A1(new_n5756_), .A2(new_n5840_), .ZN(new_n9299_));
  NOR3_X1    g08297(.A1(new_n9298_), .A2(new_n9299_), .A3(new_n5841_), .ZN(new_n9300_));
  NOR2_X1    g08298(.A1(new_n9297_), .A2(new_n9300_), .ZN(new_n9301_));
  OAI22_X1   g08299(.A1(new_n5843_), .A2(new_n5844_), .B1(new_n5812_), .B2(new_n5822_), .ZN(new_n9302_));
  NOR2_X1    g08300(.A1(new_n9301_), .A2(new_n9302_), .ZN(new_n9303_));
  NOR2_X1    g08301(.A1(new_n5837_), .A2(new_n5840_), .ZN(new_n9304_));
  AOI21_X1   g08302(.A1(new_n9295_), .A2(new_n9296_), .B(new_n5841_), .ZN(new_n9305_));
  OAI21_X1   g08303(.A1(new_n9304_), .A2(new_n9305_), .B(new_n5791_), .ZN(new_n9306_));
  NAND4_X1   g08304(.A1(new_n9303_), .A2(new_n5778_), .A3(new_n5856_), .A4(new_n9306_), .ZN(new_n9307_));
  INV_X1     g08305(.I(new_n9304_), .ZN(new_n9308_));
  OAI21_X1   g08306(.A1(new_n9298_), .A2(new_n9299_), .B(new_n5777_), .ZN(new_n9309_));
  AOI21_X1   g08307(.A1(new_n9308_), .A2(new_n9309_), .B(new_n5845_), .ZN(new_n9310_));
  NAND4_X1   g08308(.A1(new_n5791_), .A2(new_n5849_), .A3(new_n5778_), .A4(new_n5856_), .ZN(new_n9311_));
  OAI21_X1   g08309(.A1(new_n9301_), .A2(new_n9310_), .B(new_n9311_), .ZN(new_n9312_));
  AOI21_X1   g08310(.A1(new_n9307_), .A2(new_n9312_), .B(new_n9294_), .ZN(new_n9313_));
  OAI21_X1   g08311(.A1(new_n9290_), .A2(new_n9291_), .B(new_n5855_), .ZN(new_n9314_));
  INV_X1     g08312(.I(new_n9288_), .ZN(new_n9315_));
  NAND2_X1   g08313(.A1(new_n9314_), .A2(new_n9315_), .ZN(new_n9316_));
  NOR2_X1    g08314(.A1(new_n9292_), .A2(new_n9293_), .ZN(new_n9317_));
  AOI21_X1   g08315(.A1(new_n5849_), .A2(new_n9316_), .B(new_n9317_), .ZN(new_n9318_));
  OAI21_X1   g08316(.A1(new_n9298_), .A2(new_n9299_), .B(new_n5841_), .ZN(new_n9319_));
  NAND3_X1   g08317(.A1(new_n9295_), .A2(new_n9296_), .A3(new_n5777_), .ZN(new_n9320_));
  NAND2_X1   g08318(.A1(new_n9319_), .A2(new_n9320_), .ZN(new_n9321_));
  NAND3_X1   g08319(.A1(new_n9311_), .A2(new_n9306_), .A3(new_n9321_), .ZN(new_n9322_));
  NOR4_X1    g08320(.A1(new_n5845_), .A2(new_n5823_), .A3(new_n5842_), .A4(new_n5832_), .ZN(new_n9323_));
  OAI21_X1   g08321(.A1(new_n9301_), .A2(new_n9310_), .B(new_n9323_), .ZN(new_n9324_));
  AOI21_X1   g08322(.A1(new_n9324_), .A2(new_n9322_), .B(new_n9318_), .ZN(new_n9325_));
  NOR2_X1    g08323(.A1(new_n5846_), .A2(new_n5857_), .ZN(new_n9326_));
  NOR2_X1    g08324(.A1(new_n5833_), .A2(new_n5792_), .ZN(new_n9327_));
  NOR2_X1    g08325(.A1(new_n5961_), .A2(new_n5954_), .ZN(new_n9328_));
  NOR2_X1    g08326(.A1(new_n5939_), .A2(new_n5897_), .ZN(new_n9329_));
  OAI22_X1   g08327(.A1(new_n9328_), .A2(new_n9329_), .B1(new_n9326_), .B2(new_n9327_), .ZN(new_n9330_));
  NOR3_X1    g08328(.A1(new_n9313_), .A2(new_n9325_), .A3(new_n9330_), .ZN(new_n9331_));
  NAND4_X1   g08329(.A1(new_n9321_), .A2(new_n5778_), .A3(new_n5791_), .A4(new_n5849_), .ZN(new_n9332_));
  NOR2_X1    g08330(.A1(new_n9305_), .A2(new_n9304_), .ZN(new_n9333_));
  OAI21_X1   g08331(.A1(new_n9333_), .A2(new_n5845_), .B(new_n5856_), .ZN(new_n9334_));
  NOR2_X1    g08332(.A1(new_n9332_), .A2(new_n9334_), .ZN(new_n9335_));
  AOI21_X1   g08333(.A1(new_n9321_), .A2(new_n9306_), .B(new_n9323_), .ZN(new_n9336_));
  OAI21_X1   g08334(.A1(new_n9335_), .A2(new_n9336_), .B(new_n9318_), .ZN(new_n9337_));
  NOR3_X1    g08335(.A1(new_n9323_), .A2(new_n9310_), .A3(new_n9301_), .ZN(new_n9338_));
  AOI21_X1   g08336(.A1(new_n9321_), .A2(new_n9306_), .B(new_n9311_), .ZN(new_n9339_));
  OAI21_X1   g08337(.A1(new_n9339_), .A2(new_n9338_), .B(new_n9294_), .ZN(new_n9340_));
  AOI22_X1   g08338(.A1(new_n5962_), .A2(new_n5940_), .B1(new_n5834_), .B2(new_n5858_), .ZN(new_n9341_));
  AOI21_X1   g08339(.A1(new_n9337_), .A2(new_n9340_), .B(new_n9341_), .ZN(new_n9342_));
  OAI21_X1   g08340(.A1(new_n9331_), .A2(new_n9342_), .B(new_n9284_), .ZN(new_n9343_));
  AOI21_X1   g08341(.A1(new_n9273_), .A2(new_n9274_), .B(new_n5896_), .ZN(new_n9344_));
  NOR3_X1    g08342(.A1(new_n9264_), .A2(new_n9344_), .A3(new_n9278_), .ZN(new_n9345_));
  AOI21_X1   g08343(.A1(new_n9257_), .A2(new_n9262_), .B(new_n9259_), .ZN(new_n9346_));
  OAI21_X1   g08344(.A1(new_n9346_), .A2(new_n9345_), .B(new_n9272_), .ZN(new_n9347_));
  NAND3_X1   g08345(.A1(new_n9257_), .A2(new_n5950_), .A3(new_n9258_), .ZN(new_n9348_));
  NOR2_X1    g08346(.A1(new_n9261_), .A2(new_n9260_), .ZN(new_n9349_));
  OAI21_X1   g08347(.A1(new_n9349_), .A2(new_n5896_), .B(new_n5938_), .ZN(new_n9350_));
  NOR2_X1    g08348(.A1(new_n9348_), .A2(new_n9350_), .ZN(new_n9351_));
  AOI21_X1   g08349(.A1(new_n9257_), .A2(new_n9262_), .B(new_n9264_), .ZN(new_n9352_));
  OAI21_X1   g08350(.A1(new_n9351_), .A2(new_n9352_), .B(new_n9250_), .ZN(new_n9353_));
  NAND2_X1   g08351(.A1(new_n9353_), .A2(new_n9347_), .ZN(new_n9354_));
  NOR3_X1    g08352(.A1(new_n9313_), .A2(new_n9325_), .A3(new_n9341_), .ZN(new_n9355_));
  AOI21_X1   g08353(.A1(new_n9337_), .A2(new_n9340_), .B(new_n9330_), .ZN(new_n9356_));
  OAI21_X1   g08354(.A1(new_n9355_), .A2(new_n9356_), .B(new_n9354_), .ZN(new_n9357_));
  NAND2_X1   g08355(.A1(new_n9343_), .A2(new_n9357_), .ZN(new_n9358_));
  NAND2_X1   g08356(.A1(new_n9358_), .A2(new_n9239_), .ZN(new_n9359_));
  AOI22_X1   g08357(.A1(new_n6166_), .A2(new_n6168_), .B1(new_n5963_), .B2(new_n5965_), .ZN(new_n9360_));
  NAND3_X1   g08358(.A1(new_n9343_), .A2(new_n9357_), .A3(new_n9360_), .ZN(new_n9361_));
  AOI21_X1   g08359(.A1(new_n9359_), .A2(new_n9361_), .B(new_n9238_), .ZN(new_n9362_));
  NAND3_X1   g08360(.A1(new_n9213_), .A2(new_n9220_), .A3(new_n9221_), .ZN(new_n9363_));
  OAI21_X1   g08361(.A1(new_n9192_), .A2(new_n9202_), .B(new_n9207_), .ZN(new_n9364_));
  AOI21_X1   g08362(.A1(new_n9364_), .A2(new_n9363_), .B(new_n9234_), .ZN(new_n9365_));
  NAND3_X1   g08363(.A1(new_n9213_), .A2(new_n9220_), .A3(new_n9207_), .ZN(new_n9366_));
  OAI21_X1   g08364(.A1(new_n9192_), .A2(new_n9202_), .B(new_n9221_), .ZN(new_n9367_));
  AOI21_X1   g08365(.A1(new_n9366_), .A2(new_n9367_), .B(new_n9161_), .ZN(new_n9368_));
  NOR2_X1    g08366(.A1(new_n9368_), .A2(new_n9365_), .ZN(new_n9369_));
  NAND3_X1   g08367(.A1(new_n9337_), .A2(new_n9340_), .A3(new_n9341_), .ZN(new_n9370_));
  OAI21_X1   g08368(.A1(new_n9313_), .A2(new_n9325_), .B(new_n9330_), .ZN(new_n9371_));
  AOI21_X1   g08369(.A1(new_n9371_), .A2(new_n9370_), .B(new_n9354_), .ZN(new_n9372_));
  NAND3_X1   g08370(.A1(new_n9337_), .A2(new_n9340_), .A3(new_n9330_), .ZN(new_n9373_));
  OAI21_X1   g08371(.A1(new_n9313_), .A2(new_n9325_), .B(new_n9341_), .ZN(new_n9374_));
  AOI21_X1   g08372(.A1(new_n9373_), .A2(new_n9374_), .B(new_n9284_), .ZN(new_n9375_));
  OAI21_X1   g08373(.A1(new_n9375_), .A2(new_n9372_), .B(new_n9360_), .ZN(new_n9376_));
  NAND3_X1   g08374(.A1(new_n9343_), .A2(new_n9357_), .A3(new_n9239_), .ZN(new_n9377_));
  AOI21_X1   g08375(.A1(new_n9376_), .A2(new_n9377_), .B(new_n9369_), .ZN(new_n9378_));
  NOR2_X1    g08376(.A1(new_n9362_), .A2(new_n9378_), .ZN(new_n9379_));
  INV_X1     g08377(.I(new_n9379_), .ZN(new_n9380_));
  NOR2_X1    g08378(.A1(new_n6537_), .A2(new_n6555_), .ZN(new_n9381_));
  NOR2_X1    g08379(.A1(new_n6533_), .A2(new_n6556_), .ZN(new_n9382_));
  OAI21_X1   g08380(.A1(new_n9381_), .A2(new_n9382_), .B(new_n6538_), .ZN(new_n9383_));
  NOR2_X1    g08381(.A1(new_n6555_), .A2(new_n6556_), .ZN(new_n9384_));
  INV_X1     g08382(.I(new_n9384_), .ZN(new_n9385_));
  NAND2_X1   g08383(.A1(new_n9383_), .A2(new_n9385_), .ZN(new_n9386_));
  NOR4_X1    g08384(.A1(new_n9381_), .A2(new_n9382_), .A3(new_n6508_), .A4(new_n6527_), .ZN(new_n9387_));
  NAND2_X1   g08385(.A1(new_n6533_), .A2(new_n6556_), .ZN(new_n9388_));
  NAND2_X1   g08386(.A1(new_n6537_), .A2(new_n6555_), .ZN(new_n9389_));
  AOI21_X1   g08387(.A1(new_n9388_), .A2(new_n9389_), .B(new_n6538_), .ZN(new_n9390_));
  NOR2_X1    g08388(.A1(new_n9387_), .A2(new_n9390_), .ZN(new_n9391_));
  AOI21_X1   g08389(.A1(new_n6529_), .A2(new_n9386_), .B(new_n9391_), .ZN(new_n9392_));
  NAND2_X1   g08390(.A1(new_n6545_), .A2(new_n6497_), .ZN(new_n9393_));
  NAND2_X1   g08391(.A1(new_n6548_), .A2(new_n6494_), .ZN(new_n9394_));
  NAND3_X1   g08392(.A1(new_n9393_), .A2(new_n9394_), .A3(new_n6549_), .ZN(new_n9395_));
  NOR2_X1    g08393(.A1(new_n6548_), .A2(new_n6494_), .ZN(new_n9396_));
  NOR2_X1    g08394(.A1(new_n6545_), .A2(new_n6497_), .ZN(new_n9397_));
  OAI21_X1   g08395(.A1(new_n9396_), .A2(new_n9397_), .B(new_n6498_), .ZN(new_n9398_));
  NAND2_X1   g08396(.A1(new_n9398_), .A2(new_n9395_), .ZN(new_n9399_));
  NAND4_X1   g08397(.A1(new_n9399_), .A2(new_n6542_), .A3(new_n6550_), .A4(new_n6529_), .ZN(new_n9400_));
  AOI21_X1   g08398(.A1(new_n9393_), .A2(new_n9394_), .B(new_n6498_), .ZN(new_n9401_));
  NOR2_X1    g08399(.A1(new_n6494_), .A2(new_n6497_), .ZN(new_n9402_));
  OAI21_X1   g08400(.A1(new_n9401_), .A2(new_n9402_), .B(new_n6542_), .ZN(new_n9403_));
  NAND2_X1   g08401(.A1(new_n9403_), .A2(new_n6539_), .ZN(new_n9404_));
  NOR2_X1    g08402(.A1(new_n9404_), .A2(new_n9400_), .ZN(new_n9405_));
  NOR4_X1    g08403(.A1(new_n6491_), .A2(new_n6554_), .A3(new_n6499_), .A4(new_n6557_), .ZN(new_n9406_));
  AOI21_X1   g08404(.A1(new_n9399_), .A2(new_n9403_), .B(new_n9406_), .ZN(new_n9407_));
  OAI21_X1   g08405(.A1(new_n9405_), .A2(new_n9407_), .B(new_n9392_), .ZN(new_n9408_));
  NAND2_X1   g08406(.A1(new_n9388_), .A2(new_n9389_), .ZN(new_n9409_));
  AOI21_X1   g08407(.A1(new_n9409_), .A2(new_n6538_), .B(new_n9384_), .ZN(new_n9410_));
  NAND3_X1   g08408(.A1(new_n9388_), .A2(new_n9389_), .A3(new_n6538_), .ZN(new_n9411_));
  OAI22_X1   g08409(.A1(new_n9381_), .A2(new_n9382_), .B1(new_n6508_), .B2(new_n6527_), .ZN(new_n9412_));
  NAND2_X1   g08410(.A1(new_n9412_), .A2(new_n9411_), .ZN(new_n9413_));
  OAI21_X1   g08411(.A1(new_n6554_), .A2(new_n9410_), .B(new_n9413_), .ZN(new_n9414_));
  NOR3_X1    g08412(.A1(new_n9396_), .A2(new_n6498_), .A3(new_n9397_), .ZN(new_n9415_));
  AOI21_X1   g08413(.A1(new_n9393_), .A2(new_n9394_), .B(new_n6549_), .ZN(new_n9416_));
  NOR2_X1    g08414(.A1(new_n9415_), .A2(new_n9416_), .ZN(new_n9417_));
  OAI21_X1   g08415(.A1(new_n9396_), .A2(new_n9397_), .B(new_n6549_), .ZN(new_n9418_));
  INV_X1     g08416(.I(new_n9402_), .ZN(new_n9419_));
  AOI21_X1   g08417(.A1(new_n9418_), .A2(new_n9419_), .B(new_n6491_), .ZN(new_n9420_));
  NOR3_X1    g08418(.A1(new_n9420_), .A2(new_n9406_), .A3(new_n9417_), .ZN(new_n9421_));
  NAND4_X1   g08419(.A1(new_n6542_), .A2(new_n6529_), .A3(new_n6550_), .A4(new_n6539_), .ZN(new_n9422_));
  AOI21_X1   g08420(.A1(new_n9403_), .A2(new_n9399_), .B(new_n9422_), .ZN(new_n9423_));
  OAI21_X1   g08421(.A1(new_n9423_), .A2(new_n9421_), .B(new_n9414_), .ZN(new_n9424_));
  NAND2_X1   g08422(.A1(new_n9408_), .A2(new_n9424_), .ZN(new_n9425_));
  NOR2_X1    g08423(.A1(new_n6425_), .A2(new_n6453_), .ZN(new_n9426_));
  NOR2_X1    g08424(.A1(new_n6419_), .A2(new_n6454_), .ZN(new_n9427_));
  OAI21_X1   g08425(.A1(new_n9426_), .A2(new_n9427_), .B(new_n6431_), .ZN(new_n9428_));
  NOR2_X1    g08426(.A1(new_n6453_), .A2(new_n6454_), .ZN(new_n9429_));
  INV_X1     g08427(.I(new_n9429_), .ZN(new_n9430_));
  NAND2_X1   g08428(.A1(new_n9428_), .A2(new_n9430_), .ZN(new_n9431_));
  NAND2_X1   g08429(.A1(new_n6419_), .A2(new_n6454_), .ZN(new_n9432_));
  NAND2_X1   g08430(.A1(new_n6425_), .A2(new_n6453_), .ZN(new_n9433_));
  NAND3_X1   g08431(.A1(new_n9432_), .A2(new_n9433_), .A3(new_n6431_), .ZN(new_n9434_));
  OAI21_X1   g08432(.A1(new_n9426_), .A2(new_n9427_), .B(new_n6458_), .ZN(new_n9435_));
  AOI22_X1   g08433(.A1(new_n9431_), .A2(new_n6413_), .B1(new_n9434_), .B2(new_n9435_), .ZN(new_n9436_));
  NAND2_X1   g08434(.A1(new_n6444_), .A2(new_n6391_), .ZN(new_n9437_));
  NAND2_X1   g08435(.A1(new_n6440_), .A2(new_n6393_), .ZN(new_n9438_));
  NAND3_X1   g08436(.A1(new_n9437_), .A2(new_n9438_), .A3(new_n6445_), .ZN(new_n9439_));
  NOR2_X1    g08437(.A1(new_n6440_), .A2(new_n6393_), .ZN(new_n9440_));
  NOR2_X1    g08438(.A1(new_n6444_), .A2(new_n6391_), .ZN(new_n9441_));
  OAI21_X1   g08439(.A1(new_n9440_), .A2(new_n9441_), .B(new_n6394_), .ZN(new_n9442_));
  NAND2_X1   g08440(.A1(new_n9442_), .A2(new_n9439_), .ZN(new_n9443_));
  NAND4_X1   g08441(.A1(new_n9443_), .A2(new_n6437_), .A3(new_n6446_), .A4(new_n6413_), .ZN(new_n9444_));
  NOR2_X1    g08442(.A1(new_n6391_), .A2(new_n6393_), .ZN(new_n9445_));
  AOI21_X1   g08443(.A1(new_n9437_), .A2(new_n9438_), .B(new_n6394_), .ZN(new_n9446_));
  OAI21_X1   g08444(.A1(new_n9445_), .A2(new_n9446_), .B(new_n6437_), .ZN(new_n9447_));
  NAND2_X1   g08445(.A1(new_n9447_), .A2(new_n6432_), .ZN(new_n9448_));
  NOR2_X1    g08446(.A1(new_n9444_), .A2(new_n9448_), .ZN(new_n9449_));
  OAI22_X1   g08447(.A1(new_n6378_), .A2(new_n6387_), .B1(new_n6449_), .B2(new_n6451_), .ZN(new_n9450_));
  NOR3_X1    g08448(.A1(new_n9450_), .A2(new_n6395_), .A3(new_n6459_), .ZN(new_n9451_));
  AOI21_X1   g08449(.A1(new_n9443_), .A2(new_n9447_), .B(new_n9451_), .ZN(new_n9452_));
  OAI21_X1   g08450(.A1(new_n9449_), .A2(new_n9452_), .B(new_n9436_), .ZN(new_n9453_));
  NAND2_X1   g08451(.A1(new_n6567_), .A2(new_n6462_), .ZN(new_n9454_));
  NAND4_X1   g08452(.A1(new_n6413_), .A2(new_n6437_), .A3(new_n6446_), .A4(new_n6432_), .ZN(new_n9455_));
  NOR3_X1    g08453(.A1(new_n9440_), .A2(new_n9441_), .A3(new_n6394_), .ZN(new_n9456_));
  AOI21_X1   g08454(.A1(new_n9437_), .A2(new_n9438_), .B(new_n6445_), .ZN(new_n9457_));
  NOR2_X1    g08455(.A1(new_n9457_), .A2(new_n9456_), .ZN(new_n9458_));
  INV_X1     g08456(.I(new_n9445_), .ZN(new_n9459_));
  OAI21_X1   g08457(.A1(new_n9440_), .A2(new_n9441_), .B(new_n6445_), .ZN(new_n9460_));
  AOI21_X1   g08458(.A1(new_n9459_), .A2(new_n9460_), .B(new_n6388_), .ZN(new_n9461_));
  NOR2_X1    g08459(.A1(new_n9461_), .A2(new_n9458_), .ZN(new_n9462_));
  NAND2_X1   g08460(.A1(new_n9462_), .A2(new_n9455_), .ZN(new_n9463_));
  NAND2_X1   g08461(.A1(new_n9447_), .A2(new_n9443_), .ZN(new_n9464_));
  NAND2_X1   g08462(.A1(new_n9464_), .A2(new_n9451_), .ZN(new_n9465_));
  AOI21_X1   g08463(.A1(new_n9463_), .A2(new_n9465_), .B(new_n9436_), .ZN(new_n9466_));
  NOR2_X1    g08464(.A1(new_n9466_), .A2(new_n9454_), .ZN(new_n9467_));
  NAND2_X1   g08465(.A1(new_n9432_), .A2(new_n9433_), .ZN(new_n9468_));
  AOI21_X1   g08466(.A1(new_n9468_), .A2(new_n6431_), .B(new_n9429_), .ZN(new_n9469_));
  NOR3_X1    g08467(.A1(new_n9426_), .A2(new_n9427_), .A3(new_n6458_), .ZN(new_n9470_));
  AOI21_X1   g08468(.A1(new_n9432_), .A2(new_n9433_), .B(new_n6431_), .ZN(new_n9471_));
  OAI22_X1   g08469(.A1(new_n9469_), .A2(new_n6452_), .B1(new_n9470_), .B2(new_n9471_), .ZN(new_n9472_));
  NOR2_X1    g08470(.A1(new_n9464_), .A2(new_n9451_), .ZN(new_n9473_));
  AOI21_X1   g08471(.A1(new_n9443_), .A2(new_n9447_), .B(new_n9455_), .ZN(new_n9474_));
  OAI21_X1   g08472(.A1(new_n9473_), .A2(new_n9474_), .B(new_n9472_), .ZN(new_n9475_));
  NAND2_X1   g08473(.A1(new_n9453_), .A2(new_n9475_), .ZN(new_n9476_));
  AOI22_X1   g08474(.A1(new_n9453_), .A2(new_n9467_), .B1(new_n9476_), .B2(new_n9454_), .ZN(new_n9477_));
  NOR2_X1    g08475(.A1(new_n9458_), .A2(new_n9450_), .ZN(new_n9478_));
  NAND4_X1   g08476(.A1(new_n9478_), .A2(new_n6446_), .A3(new_n6432_), .A4(new_n9447_), .ZN(new_n9479_));
  NAND2_X1   g08477(.A1(new_n9464_), .A2(new_n9455_), .ZN(new_n9480_));
  AOI21_X1   g08478(.A1(new_n9479_), .A2(new_n9480_), .B(new_n9472_), .ZN(new_n9481_));
  NOR2_X1    g08479(.A1(new_n6560_), .A2(new_n6564_), .ZN(new_n9482_));
  NOR3_X1    g08480(.A1(new_n9481_), .A2(new_n9466_), .A3(new_n9482_), .ZN(new_n9483_));
  AOI21_X1   g08481(.A1(new_n9453_), .A2(new_n9475_), .B(new_n9454_), .ZN(new_n9484_));
  OAI21_X1   g08482(.A1(new_n9483_), .A2(new_n9484_), .B(new_n9425_), .ZN(new_n9485_));
  OAI21_X1   g08483(.A1(new_n9425_), .A2(new_n9477_), .B(new_n9485_), .ZN(new_n9486_));
  XOR2_X1    g08484(.A1(\A[250] ), .A2(\A[251] ), .Z(new_n9487_));
  AOI21_X1   g08485(.A1(new_n9487_), .A2(\A[252] ), .B(new_n6303_), .ZN(new_n9488_));
  NOR2_X1    g08486(.A1(new_n6317_), .A2(new_n9488_), .ZN(new_n9489_));
  NAND2_X1   g08487(.A1(new_n6318_), .A2(new_n6325_), .ZN(new_n9490_));
  AOI21_X1   g08488(.A1(new_n9490_), .A2(\A[249] ), .B(new_n6312_), .ZN(new_n9491_));
  NOR2_X1    g08489(.A1(new_n6308_), .A2(new_n9491_), .ZN(new_n9492_));
  NOR2_X1    g08490(.A1(new_n9492_), .A2(new_n9489_), .ZN(new_n9493_));
  OAI22_X1   g08491(.A1(new_n6326_), .A2(new_n6327_), .B1(new_n6331_), .B2(new_n6332_), .ZN(new_n9494_));
  NOR2_X1    g08492(.A1(new_n9491_), .A2(new_n9488_), .ZN(new_n9495_));
  INV_X1     g08493(.I(new_n9495_), .ZN(new_n9496_));
  OAI21_X1   g08494(.A1(new_n9493_), .A2(new_n9494_), .B(new_n9496_), .ZN(new_n9497_));
  NAND2_X1   g08495(.A1(new_n6308_), .A2(new_n9491_), .ZN(new_n9498_));
  NAND2_X1   g08496(.A1(new_n6317_), .A2(new_n9488_), .ZN(new_n9499_));
  NAND4_X1   g08497(.A1(new_n9498_), .A2(new_n9499_), .A3(new_n6320_), .A4(new_n6323_), .ZN(new_n9500_));
  OAI21_X1   g08498(.A1(new_n9492_), .A2(new_n9489_), .B(new_n9494_), .ZN(new_n9501_));
  AOI22_X1   g08499(.A1(new_n9497_), .A2(new_n6335_), .B1(new_n9500_), .B2(new_n9501_), .ZN(new_n9502_));
  NAND2_X1   g08500(.A1(new_n6277_), .A2(new_n6338_), .ZN(new_n9503_));
  NAND2_X1   g08501(.A1(new_n6268_), .A2(new_n6340_), .ZN(new_n9504_));
  NAND3_X1   g08502(.A1(new_n9504_), .A2(new_n9503_), .A3(new_n6286_), .ZN(new_n9505_));
  NOR2_X1    g08503(.A1(new_n6268_), .A2(new_n6340_), .ZN(new_n9506_));
  NOR2_X1    g08504(.A1(new_n6277_), .A2(new_n6338_), .ZN(new_n9507_));
  OAI21_X1   g08505(.A1(new_n9506_), .A2(new_n9507_), .B(new_n6341_), .ZN(new_n9508_));
  NAND2_X1   g08506(.A1(new_n9508_), .A2(new_n9505_), .ZN(new_n9509_));
  AOI22_X1   g08507(.A1(new_n6329_), .A2(new_n6334_), .B1(new_n6292_), .B2(new_n6297_), .ZN(new_n9510_));
  NAND3_X1   g08508(.A1(new_n9510_), .A2(new_n6287_), .A3(new_n6324_), .ZN(new_n9511_));
  NOR2_X1    g08509(.A1(new_n6340_), .A2(new_n6338_), .ZN(new_n9512_));
  AOI21_X1   g08510(.A1(new_n9504_), .A2(new_n9503_), .B(new_n6341_), .ZN(new_n9513_));
  OAI21_X1   g08511(.A1(new_n9512_), .A2(new_n9513_), .B(new_n6298_), .ZN(new_n9514_));
  NAND3_X1   g08512(.A1(new_n9511_), .A2(new_n9514_), .A3(new_n9509_), .ZN(new_n9515_));
  NOR3_X1    g08513(.A1(new_n9494_), .A2(new_n9488_), .A3(new_n9491_), .ZN(new_n9516_));
  NOR2_X1    g08514(.A1(new_n6320_), .A2(new_n6333_), .ZN(new_n9517_));
  NOR2_X1    g08515(.A1(new_n6323_), .A2(new_n6328_), .ZN(new_n9518_));
  NOR2_X1    g08516(.A1(new_n9518_), .A2(new_n9517_), .ZN(new_n9519_));
  NOR4_X1    g08517(.A1(new_n9519_), .A2(new_n6345_), .A3(new_n6342_), .A4(new_n9516_), .ZN(new_n9520_));
  NAND2_X1   g08518(.A1(new_n9514_), .A2(new_n9509_), .ZN(new_n9521_));
  NAND2_X1   g08519(.A1(new_n9521_), .A2(new_n9520_), .ZN(new_n9522_));
  AOI21_X1   g08520(.A1(new_n9522_), .A2(new_n9515_), .B(new_n9502_), .ZN(new_n9523_));
  AOI21_X1   g08521(.A1(new_n9498_), .A2(new_n9499_), .B(new_n9494_), .ZN(new_n9524_));
  NOR2_X1    g08522(.A1(new_n9524_), .A2(new_n9495_), .ZN(new_n9525_));
  NOR3_X1    g08523(.A1(new_n9492_), .A2(new_n9489_), .A3(new_n9494_), .ZN(new_n9526_));
  AOI22_X1   g08524(.A1(new_n9498_), .A2(new_n9499_), .B1(new_n6320_), .B2(new_n6323_), .ZN(new_n9527_));
  OAI22_X1   g08525(.A1(new_n9525_), .A2(new_n9519_), .B1(new_n9526_), .B2(new_n9527_), .ZN(new_n9528_));
  INV_X1     g08526(.I(new_n9512_), .ZN(new_n9529_));
  OAI21_X1   g08527(.A1(new_n9506_), .A2(new_n9507_), .B(new_n6286_), .ZN(new_n9530_));
  NAND2_X1   g08528(.A1(new_n9530_), .A2(new_n9529_), .ZN(new_n9531_));
  NOR3_X1    g08529(.A1(new_n9506_), .A2(new_n9507_), .A3(new_n6341_), .ZN(new_n9532_));
  AOI21_X1   g08530(.A1(new_n9504_), .A2(new_n9503_), .B(new_n6286_), .ZN(new_n9533_));
  NOR2_X1    g08531(.A1(new_n9533_), .A2(new_n9532_), .ZN(new_n9534_));
  NOR4_X1    g08532(.A1(new_n9534_), .A2(new_n9531_), .A3(new_n6345_), .A4(new_n9519_), .ZN(new_n9535_));
  AOI21_X1   g08533(.A1(new_n9531_), .A2(new_n6298_), .B(new_n9516_), .ZN(new_n9536_));
  NAND2_X1   g08534(.A1(new_n9535_), .A2(new_n9536_), .ZN(new_n9537_));
  NAND2_X1   g08535(.A1(new_n9521_), .A2(new_n9511_), .ZN(new_n9538_));
  AOI21_X1   g08536(.A1(new_n9537_), .A2(new_n9538_), .B(new_n9528_), .ZN(new_n9539_));
  NOR2_X1    g08537(.A1(new_n9539_), .A2(new_n9523_), .ZN(new_n9540_));
  INV_X1     g08538(.I(new_n6212_), .ZN(new_n9541_));
  AOI21_X1   g08539(.A1(new_n6232_), .A2(\A[264] ), .B(new_n9541_), .ZN(new_n9542_));
  NOR2_X1    g08540(.A1(new_n6218_), .A2(new_n9542_), .ZN(new_n9543_));
  INV_X1     g08541(.I(new_n6216_), .ZN(new_n9544_));
  XOR2_X1    g08542(.A1(\A[259] ), .A2(\A[260] ), .Z(new_n9545_));
  AOI21_X1   g08543(.A1(new_n9545_), .A2(\A[261] ), .B(new_n9544_), .ZN(new_n9546_));
  NOR2_X1    g08544(.A1(new_n6214_), .A2(new_n9546_), .ZN(new_n9547_));
  NOR2_X1    g08545(.A1(new_n9543_), .A2(new_n9547_), .ZN(new_n9548_));
  NAND2_X1   g08546(.A1(new_n6224_), .A2(\A[262] ), .ZN(new_n9549_));
  AOI21_X1   g08547(.A1(new_n9549_), .A2(new_n6231_), .B(\A[264] ), .ZN(new_n9550_));
  NOR2_X1    g08548(.A1(new_n6226_), .A2(\A[263] ), .ZN(new_n9551_));
  NOR3_X1    g08549(.A1(new_n9551_), .A2(new_n6225_), .A3(new_n6211_), .ZN(new_n9552_));
  OAI22_X1   g08550(.A1(new_n9550_), .A2(new_n9552_), .B1(new_n6251_), .B2(new_n6252_), .ZN(new_n9553_));
  NOR2_X1    g08551(.A1(new_n9542_), .A2(new_n9546_), .ZN(new_n9554_));
  INV_X1     g08552(.I(new_n9554_), .ZN(new_n9555_));
  OAI21_X1   g08553(.A1(new_n9548_), .A2(new_n9553_), .B(new_n9555_), .ZN(new_n9556_));
  NAND2_X1   g08554(.A1(new_n6214_), .A2(new_n9546_), .ZN(new_n9557_));
  NAND2_X1   g08555(.A1(new_n6218_), .A2(new_n9542_), .ZN(new_n9558_));
  NAND4_X1   g08556(.A1(new_n9557_), .A2(new_n9558_), .A3(new_n6223_), .A4(new_n6228_), .ZN(new_n9559_));
  OAI21_X1   g08557(.A1(new_n9543_), .A2(new_n9547_), .B(new_n9553_), .ZN(new_n9560_));
  AOI22_X1   g08558(.A1(new_n9556_), .A2(new_n6256_), .B1(new_n9559_), .B2(new_n9560_), .ZN(new_n9561_));
  NAND2_X1   g08559(.A1(new_n6183_), .A2(new_n6239_), .ZN(new_n9562_));
  NAND2_X1   g08560(.A1(new_n6179_), .A2(new_n6242_), .ZN(new_n9563_));
  NAND3_X1   g08561(.A1(new_n9563_), .A2(new_n9562_), .A3(new_n6196_), .ZN(new_n9564_));
  NOR2_X1    g08562(.A1(new_n6179_), .A2(new_n6242_), .ZN(new_n9565_));
  NOR2_X1    g08563(.A1(new_n6183_), .A2(new_n6239_), .ZN(new_n9566_));
  OAI21_X1   g08564(.A1(new_n9565_), .A2(new_n9566_), .B(new_n6243_), .ZN(new_n9567_));
  NAND2_X1   g08565(.A1(new_n9567_), .A2(new_n9564_), .ZN(new_n9568_));
  NAND4_X1   g08566(.A1(new_n9568_), .A2(new_n6197_), .A3(new_n6209_), .A4(new_n6256_), .ZN(new_n9569_));
  NOR2_X1    g08567(.A1(new_n6239_), .A2(new_n6242_), .ZN(new_n9570_));
  AOI21_X1   g08568(.A1(new_n9563_), .A2(new_n9562_), .B(new_n6243_), .ZN(new_n9571_));
  NOR2_X1    g08569(.A1(new_n9571_), .A2(new_n9570_), .ZN(new_n9572_));
  OAI21_X1   g08570(.A1(new_n9572_), .A2(new_n6247_), .B(new_n6229_), .ZN(new_n9573_));
  NOR2_X1    g08571(.A1(new_n9569_), .A2(new_n9573_), .ZN(new_n9574_));
  OAI21_X1   g08572(.A1(new_n9570_), .A2(new_n9571_), .B(new_n6209_), .ZN(new_n9575_));
  NOR4_X1    g08573(.A1(new_n6235_), .A2(new_n6247_), .A3(new_n6230_), .A4(new_n6244_), .ZN(new_n9576_));
  AOI21_X1   g08574(.A1(new_n9568_), .A2(new_n9575_), .B(new_n9576_), .ZN(new_n9577_));
  OAI21_X1   g08575(.A1(new_n9574_), .A2(new_n9577_), .B(new_n9561_), .ZN(new_n9578_));
  AOI21_X1   g08576(.A1(new_n9557_), .A2(new_n9558_), .B(new_n9553_), .ZN(new_n9579_));
  NOR2_X1    g08577(.A1(new_n9579_), .A2(new_n9554_), .ZN(new_n9580_));
  NOR3_X1    g08578(.A1(new_n9543_), .A2(new_n9547_), .A3(new_n9553_), .ZN(new_n9581_));
  AOI22_X1   g08579(.A1(new_n9557_), .A2(new_n9558_), .B1(new_n6223_), .B2(new_n6228_), .ZN(new_n9582_));
  OAI22_X1   g08580(.A1(new_n9580_), .A2(new_n6235_), .B1(new_n9581_), .B2(new_n9582_), .ZN(new_n9583_));
  NOR3_X1    g08581(.A1(new_n9565_), .A2(new_n9566_), .A3(new_n6243_), .ZN(new_n9584_));
  AOI21_X1   g08582(.A1(new_n9563_), .A2(new_n9562_), .B(new_n6196_), .ZN(new_n9585_));
  NOR2_X1    g08583(.A1(new_n9584_), .A2(new_n9585_), .ZN(new_n9586_));
  INV_X1     g08584(.I(new_n9570_), .ZN(new_n9587_));
  OAI21_X1   g08585(.A1(new_n9565_), .A2(new_n9566_), .B(new_n6196_), .ZN(new_n9588_));
  AOI21_X1   g08586(.A1(new_n9587_), .A2(new_n9588_), .B(new_n6247_), .ZN(new_n9589_));
  NOR3_X1    g08587(.A1(new_n9576_), .A2(new_n9589_), .A3(new_n9586_), .ZN(new_n9590_));
  NAND4_X1   g08588(.A1(new_n6209_), .A2(new_n6256_), .A3(new_n6197_), .A4(new_n6229_), .ZN(new_n9591_));
  AOI21_X1   g08589(.A1(new_n9568_), .A2(new_n9575_), .B(new_n9591_), .ZN(new_n9592_));
  OAI21_X1   g08590(.A1(new_n9590_), .A2(new_n9592_), .B(new_n9583_), .ZN(new_n9593_));
  NAND2_X1   g08591(.A1(new_n6349_), .A2(new_n6353_), .ZN(new_n9594_));
  NAND3_X1   g08592(.A1(new_n9578_), .A2(new_n9594_), .A3(new_n9593_), .ZN(new_n9595_));
  NOR2_X1    g08593(.A1(new_n6247_), .A2(new_n6235_), .ZN(new_n9596_));
  NAND2_X1   g08594(.A1(new_n9588_), .A2(new_n9587_), .ZN(new_n9597_));
  AOI21_X1   g08595(.A1(new_n9597_), .A2(new_n6209_), .B(new_n6230_), .ZN(new_n9598_));
  NAND4_X1   g08596(.A1(new_n9598_), .A2(new_n9572_), .A3(new_n9568_), .A4(new_n9596_), .ZN(new_n9599_));
  NAND2_X1   g08597(.A1(new_n9575_), .A2(new_n9568_), .ZN(new_n9600_));
  NAND2_X1   g08598(.A1(new_n9600_), .A2(new_n9591_), .ZN(new_n9601_));
  AOI21_X1   g08599(.A1(new_n9599_), .A2(new_n9601_), .B(new_n9583_), .ZN(new_n9602_));
  NAND3_X1   g08600(.A1(new_n9575_), .A2(new_n9591_), .A3(new_n9568_), .ZN(new_n9603_));
  NAND2_X1   g08601(.A1(new_n9600_), .A2(new_n9576_), .ZN(new_n9604_));
  AOI21_X1   g08602(.A1(new_n9604_), .A2(new_n9603_), .B(new_n9561_), .ZN(new_n9605_));
  NOR2_X1    g08603(.A1(new_n6356_), .A2(new_n6259_), .ZN(new_n9606_));
  OAI21_X1   g08604(.A1(new_n9602_), .A2(new_n9605_), .B(new_n9606_), .ZN(new_n9607_));
  AOI21_X1   g08605(.A1(new_n9607_), .A2(new_n9595_), .B(new_n9540_), .ZN(new_n9608_));
  NOR2_X1    g08606(.A1(new_n9521_), .A2(new_n9520_), .ZN(new_n9609_));
  AOI21_X1   g08607(.A1(new_n9509_), .A2(new_n9514_), .B(new_n9511_), .ZN(new_n9610_));
  OAI21_X1   g08608(.A1(new_n9609_), .A2(new_n9610_), .B(new_n9528_), .ZN(new_n9611_));
  NAND3_X1   g08609(.A1(new_n9509_), .A2(new_n6287_), .A3(new_n9510_), .ZN(new_n9612_));
  NOR2_X1    g08610(.A1(new_n9513_), .A2(new_n9512_), .ZN(new_n9613_));
  OAI21_X1   g08611(.A1(new_n9613_), .A2(new_n6345_), .B(new_n6324_), .ZN(new_n9614_));
  NOR2_X1    g08612(.A1(new_n9612_), .A2(new_n9614_), .ZN(new_n9615_));
  AOI21_X1   g08613(.A1(new_n9509_), .A2(new_n9514_), .B(new_n9520_), .ZN(new_n9616_));
  OAI21_X1   g08614(.A1(new_n9615_), .A2(new_n9616_), .B(new_n9502_), .ZN(new_n9617_));
  NAND2_X1   g08615(.A1(new_n9611_), .A2(new_n9617_), .ZN(new_n9618_));
  NAND3_X1   g08616(.A1(new_n9578_), .A2(new_n9606_), .A3(new_n9593_), .ZN(new_n9619_));
  OAI21_X1   g08617(.A1(new_n9602_), .A2(new_n9605_), .B(new_n9594_), .ZN(new_n9620_));
  AOI21_X1   g08618(.A1(new_n9620_), .A2(new_n9619_), .B(new_n9618_), .ZN(new_n9621_));
  AOI21_X1   g08619(.A1(new_n6561_), .A2(new_n6568_), .B(new_n6358_), .ZN(new_n9622_));
  NOR3_X1    g08620(.A1(new_n9608_), .A2(new_n9621_), .A3(new_n9622_), .ZN(new_n9623_));
  NOR3_X1    g08621(.A1(new_n9602_), .A2(new_n9605_), .A3(new_n9606_), .ZN(new_n9624_));
  AOI21_X1   g08622(.A1(new_n9578_), .A2(new_n9593_), .B(new_n9594_), .ZN(new_n9625_));
  OAI21_X1   g08623(.A1(new_n9624_), .A2(new_n9625_), .B(new_n9618_), .ZN(new_n9626_));
  NOR3_X1    g08624(.A1(new_n9602_), .A2(new_n9605_), .A3(new_n9594_), .ZN(new_n9627_));
  AOI21_X1   g08625(.A1(new_n9578_), .A2(new_n9593_), .B(new_n9606_), .ZN(new_n9628_));
  OAI21_X1   g08626(.A1(new_n9628_), .A2(new_n9627_), .B(new_n9540_), .ZN(new_n9629_));
  OAI21_X1   g08627(.A1(new_n6350_), .A2(new_n6357_), .B(new_n6569_), .ZN(new_n9630_));
  AOI21_X1   g08628(.A1(new_n9629_), .A2(new_n9626_), .B(new_n9630_), .ZN(new_n9631_));
  OAI21_X1   g08629(.A1(new_n9631_), .A2(new_n9623_), .B(new_n9486_), .ZN(new_n9632_));
  NOR2_X1    g08630(.A1(new_n9477_), .A2(new_n9425_), .ZN(new_n9633_));
  INV_X1     g08631(.I(new_n9485_), .ZN(new_n9634_));
  NOR2_X1    g08632(.A1(new_n9633_), .A2(new_n9634_), .ZN(new_n9635_));
  NAND3_X1   g08633(.A1(new_n9629_), .A2(new_n9626_), .A3(new_n9622_), .ZN(new_n9636_));
  OAI21_X1   g08634(.A1(new_n9608_), .A2(new_n9621_), .B(new_n9630_), .ZN(new_n9637_));
  NAND2_X1   g08635(.A1(new_n9637_), .A2(new_n9636_), .ZN(new_n9638_));
  NAND2_X1   g08636(.A1(new_n9638_), .A2(new_n9635_), .ZN(new_n9639_));
  NAND2_X1   g08637(.A1(new_n6170_), .A2(new_n6570_), .ZN(new_n9640_));
  INV_X1     g08638(.I(new_n9640_), .ZN(new_n9641_));
  NAND3_X1   g08639(.A1(new_n9639_), .A2(new_n9632_), .A3(new_n9641_), .ZN(new_n9642_));
  NAND2_X1   g08640(.A1(new_n9639_), .A2(new_n9632_), .ZN(new_n9643_));
  NAND2_X1   g08641(.A1(new_n9643_), .A2(new_n9640_), .ZN(new_n9644_));
  AOI21_X1   g08642(.A1(new_n9644_), .A2(new_n9642_), .B(new_n9380_), .ZN(new_n9645_));
  NAND3_X1   g08643(.A1(new_n9639_), .A2(new_n9632_), .A3(new_n9640_), .ZN(new_n9646_));
  NAND3_X1   g08644(.A1(new_n9629_), .A2(new_n9626_), .A3(new_n9630_), .ZN(new_n9647_));
  OAI21_X1   g08645(.A1(new_n9608_), .A2(new_n9621_), .B(new_n9622_), .ZN(new_n9648_));
  AOI21_X1   g08646(.A1(new_n9647_), .A2(new_n9648_), .B(new_n9635_), .ZN(new_n9649_));
  AOI21_X1   g08647(.A1(new_n9637_), .A2(new_n9636_), .B(new_n9486_), .ZN(new_n9650_));
  OAI21_X1   g08648(.A1(new_n9649_), .A2(new_n9650_), .B(new_n9641_), .ZN(new_n9651_));
  AOI21_X1   g08649(.A1(new_n9651_), .A2(new_n9646_), .B(new_n9379_), .ZN(new_n9652_));
  OAI21_X1   g08650(.A1(new_n9645_), .A2(new_n9652_), .B(new_n9106_), .ZN(new_n9653_));
  NAND2_X1   g08651(.A1(new_n9644_), .A2(new_n9642_), .ZN(new_n9654_));
  NAND2_X1   g08652(.A1(new_n9654_), .A2(new_n9379_), .ZN(new_n9655_));
  INV_X1     g08653(.I(new_n9652_), .ZN(new_n9656_));
  NAND3_X1   g08654(.A1(new_n9655_), .A2(new_n9105_), .A3(new_n9656_), .ZN(new_n9657_));
  AOI21_X1   g08655(.A1(new_n9657_), .A2(new_n9653_), .B(new_n9104_), .ZN(new_n9658_));
  NOR2_X1    g08656(.A1(new_n9098_), .A2(new_n8825_), .ZN(new_n9659_));
  AOI21_X1   g08657(.A1(new_n8825_), .A2(new_n9102_), .B(new_n9659_), .ZN(new_n9660_));
  OAI21_X1   g08658(.A1(new_n9645_), .A2(new_n9652_), .B(new_n9105_), .ZN(new_n9661_));
  NOR3_X1    g08659(.A1(new_n9645_), .A2(new_n9105_), .A3(new_n9652_), .ZN(new_n9662_));
  INV_X1     g08660(.I(new_n9662_), .ZN(new_n9663_));
  AOI21_X1   g08661(.A1(new_n9663_), .A2(new_n9661_), .B(new_n9660_), .ZN(new_n9664_));
  NOR2_X1    g08662(.A1(new_n9664_), .A2(new_n9658_), .ZN(new_n9665_));
  INV_X1     g08663(.I(new_n7384_), .ZN(new_n9666_));
  NAND3_X1   g08664(.A1(new_n8537_), .A2(new_n9666_), .A3(new_n8540_), .ZN(new_n9667_));
  INV_X1     g08665(.I(new_n9667_), .ZN(new_n9668_));
  OAI21_X1   g08666(.A1(new_n9665_), .A2(new_n9668_), .B(new_n8542_), .ZN(new_n9669_));
  NAND2_X1   g08667(.A1(new_n9655_), .A2(new_n9656_), .ZN(new_n9670_));
  AOI22_X1   g08668(.A1(new_n9663_), .A2(new_n9104_), .B1(new_n9670_), .B2(new_n9105_), .ZN(new_n9671_));
  NAND2_X1   g08669(.A1(new_n8825_), .A2(new_n9099_), .ZN(new_n9672_));
  NAND2_X1   g08670(.A1(new_n9672_), .A2(new_n9101_), .ZN(new_n9673_));
  NAND3_X1   g08671(.A1(new_n8811_), .A2(new_n8814_), .A3(new_n8807_), .ZN(new_n9674_));
  AOI21_X1   g08672(.A1(new_n8821_), .A2(new_n9674_), .B(new_n8823_), .ZN(new_n9675_));
  OAI21_X1   g08673(.A1(new_n8660_), .A2(new_n8818_), .B(new_n8662_), .ZN(new_n9676_));
  OAI21_X1   g08674(.A1(new_n8579_), .A2(new_n7361_), .B(new_n8576_), .ZN(new_n9677_));
  AOI21_X1   g08675(.A1(new_n8585_), .A2(new_n7366_), .B(new_n8584_), .ZN(new_n9678_));
  NAND2_X1   g08676(.A1(new_n9677_), .A2(new_n9678_), .ZN(new_n9679_));
  AOI21_X1   g08677(.A1(new_n8565_), .A2(new_n7306_), .B(new_n8570_), .ZN(new_n9680_));
  NOR3_X1    g08678(.A1(new_n8544_), .A2(new_n8543_), .A3(new_n7355_), .ZN(new_n9681_));
  AOI21_X1   g08679(.A1(new_n8549_), .A2(new_n8550_), .B(new_n7372_), .ZN(new_n9682_));
  NOR2_X1    g08680(.A1(new_n9681_), .A2(new_n9682_), .ZN(new_n9683_));
  OAI21_X1   g08681(.A1(new_n9683_), .A2(new_n7347_), .B(new_n8548_), .ZN(new_n9684_));
  NAND2_X1   g08682(.A1(new_n9680_), .A2(new_n9684_), .ZN(new_n9685_));
  OAI21_X1   g08683(.A1(new_n8580_), .A2(new_n8573_), .B(new_n8553_), .ZN(new_n9686_));
  AOI22_X1   g08684(.A1(new_n9686_), .A2(new_n8654_), .B1(new_n9679_), .B2(new_n9685_), .ZN(new_n9687_));
  NOR2_X1    g08685(.A1(new_n9677_), .A2(new_n9678_), .ZN(new_n9688_));
  AOI21_X1   g08686(.A1(new_n8590_), .A2(new_n8588_), .B(new_n8586_), .ZN(new_n9689_));
  OAI22_X1   g08687(.A1(new_n9680_), .A2(new_n9684_), .B1(new_n8567_), .B2(new_n8571_), .ZN(new_n9690_));
  NOR3_X1    g08688(.A1(new_n9690_), .A2(new_n9689_), .A3(new_n9688_), .ZN(new_n9691_));
  NOR2_X1    g08689(.A1(new_n9687_), .A2(new_n9691_), .ZN(new_n9692_));
  AOI21_X1   g08690(.A1(new_n8613_), .A2(new_n7201_), .B(new_n8608_), .ZN(new_n9693_));
  NOR2_X1    g08691(.A1(new_n8601_), .A2(new_n8602_), .ZN(new_n9694_));
  OAI21_X1   g08692(.A1(new_n9694_), .A2(new_n7239_), .B(new_n8629_), .ZN(new_n9695_));
  NOR2_X1    g08693(.A1(new_n9693_), .A2(new_n9695_), .ZN(new_n9696_));
  OAI21_X1   g08694(.A1(new_n8622_), .A2(new_n7257_), .B(new_n8617_), .ZN(new_n9697_));
  NAND2_X1   g08695(.A1(new_n8631_), .A2(new_n8630_), .ZN(new_n9698_));
  AOI21_X1   g08696(.A1(new_n9698_), .A2(new_n7269_), .B(new_n8598_), .ZN(new_n9699_));
  NOR2_X1    g08697(.A1(new_n9699_), .A2(new_n9697_), .ZN(new_n9700_));
  NAND2_X1   g08698(.A1(new_n8635_), .A2(new_n8613_), .ZN(new_n9701_));
  AOI21_X1   g08699(.A1(new_n8624_), .A2(new_n9701_), .B(new_n8603_), .ZN(new_n9702_));
  OAI22_X1   g08700(.A1(new_n9702_), .A2(new_n8642_), .B1(new_n9696_), .B2(new_n9700_), .ZN(new_n9703_));
  NAND2_X1   g08701(.A1(new_n9699_), .A2(new_n9697_), .ZN(new_n9704_));
  NAND2_X1   g08702(.A1(new_n9693_), .A2(new_n9695_), .ZN(new_n9705_));
  NOR2_X1    g08703(.A1(new_n8623_), .A2(new_n8622_), .ZN(new_n9706_));
  OAI21_X1   g08704(.A1(new_n9706_), .A2(new_n8633_), .B(new_n8632_), .ZN(new_n9707_));
  NAND4_X1   g08705(.A1(new_n9707_), .A2(new_n9704_), .A3(new_n9705_), .A4(new_n8619_), .ZN(new_n9708_));
  NAND2_X1   g08706(.A1(new_n9703_), .A2(new_n9708_), .ZN(new_n9709_));
  NOR2_X1    g08707(.A1(new_n9692_), .A2(new_n9709_), .ZN(new_n9710_));
  NOR2_X1    g08708(.A1(new_n9680_), .A2(new_n9684_), .ZN(new_n9711_));
  OAI22_X1   g08709(.A1(new_n9689_), .A2(new_n8572_), .B1(new_n9711_), .B2(new_n9688_), .ZN(new_n9712_));
  NAND4_X1   g08710(.A1(new_n9686_), .A2(new_n8654_), .A3(new_n9679_), .A4(new_n9685_), .ZN(new_n9713_));
  NAND2_X1   g08711(.A1(new_n9712_), .A2(new_n9713_), .ZN(new_n9714_));
  AOI22_X1   g08712(.A1(new_n9707_), .A2(new_n8619_), .B1(new_n9704_), .B2(new_n9705_), .ZN(new_n9715_));
  OAI22_X1   g08713(.A1(new_n9693_), .A2(new_n9695_), .B1(new_n8640_), .B2(new_n8641_), .ZN(new_n9716_));
  NOR3_X1    g08714(.A1(new_n9716_), .A2(new_n9702_), .A3(new_n9700_), .ZN(new_n9717_));
  NOR2_X1    g08715(.A1(new_n9715_), .A2(new_n9717_), .ZN(new_n9718_));
  NOR2_X1    g08716(.A1(new_n9714_), .A2(new_n9718_), .ZN(new_n9719_));
  OAI21_X1   g08717(.A1(new_n9710_), .A2(new_n9719_), .B(new_n9676_), .ZN(new_n9720_));
  AOI21_X1   g08718(.A1(new_n8593_), .A2(new_n8661_), .B(new_n8819_), .ZN(new_n9721_));
  NAND2_X1   g08719(.A1(new_n9714_), .A2(new_n9718_), .ZN(new_n9722_));
  NAND2_X1   g08720(.A1(new_n9692_), .A2(new_n9709_), .ZN(new_n9723_));
  NAND3_X1   g08721(.A1(new_n9722_), .A2(new_n9723_), .A3(new_n9721_), .ZN(new_n9724_));
  NAND2_X1   g08722(.A1(new_n9720_), .A2(new_n9724_), .ZN(new_n9725_));
  AOI21_X1   g08723(.A1(new_n8802_), .A2(new_n8791_), .B(new_n8809_), .ZN(new_n9726_));
  AOI22_X1   g08724(.A1(new_n8712_), .A2(new_n7102_), .B1(new_n8694_), .B2(new_n8696_), .ZN(new_n9727_));
  OAI21_X1   g08725(.A1(new_n8708_), .A2(new_n7145_), .B(new_n8707_), .ZN(new_n9728_));
  NOR2_X1    g08726(.A1(new_n9727_), .A2(new_n9728_), .ZN(new_n9729_));
  OAI21_X1   g08727(.A1(new_n8688_), .A2(new_n8700_), .B(new_n8697_), .ZN(new_n9730_));
  NAND3_X1   g08728(.A1(new_n8665_), .A2(new_n8666_), .A3(new_n7164_), .ZN(new_n9731_));
  OAI21_X1   g08729(.A1(new_n8671_), .A2(new_n8670_), .B(new_n7152_), .ZN(new_n9732_));
  NAND2_X1   g08730(.A1(new_n9732_), .A2(new_n9731_), .ZN(new_n9733_));
  AOI21_X1   g08731(.A1(new_n9733_), .A2(new_n7158_), .B(new_n8669_), .ZN(new_n9734_));
  NOR2_X1    g08732(.A1(new_n9730_), .A2(new_n9734_), .ZN(new_n9735_));
  AOI21_X1   g08733(.A1(new_n8702_), .A2(new_n8717_), .B(new_n8674_), .ZN(new_n9736_));
  OAI22_X1   g08734(.A1(new_n9736_), .A2(new_n8795_), .B1(new_n9735_), .B2(new_n9729_), .ZN(new_n9737_));
  NAND2_X1   g08735(.A1(new_n9730_), .A2(new_n9734_), .ZN(new_n9738_));
  NAND2_X1   g08736(.A1(new_n9727_), .A2(new_n9728_), .ZN(new_n9739_));
  NAND2_X1   g08737(.A1(new_n8703_), .A2(new_n8709_), .ZN(new_n9740_));
  NAND4_X1   g08738(.A1(new_n9740_), .A2(new_n9738_), .A3(new_n9739_), .A4(new_n8699_), .ZN(new_n9741_));
  NAND2_X1   g08739(.A1(new_n9737_), .A2(new_n9741_), .ZN(new_n9742_));
  OAI21_X1   g08740(.A1(new_n8757_), .A2(new_n8735_), .B(new_n8745_), .ZN(new_n9743_));
  AOI21_X1   g08741(.A1(new_n8731_), .A2(new_n7063_), .B(new_n8726_), .ZN(new_n9744_));
  NAND2_X1   g08742(.A1(new_n9744_), .A2(new_n9743_), .ZN(new_n9745_));
  AOI21_X1   g08743(.A1(new_n8775_), .A2(new_n7010_), .B(new_n8783_), .ZN(new_n9746_));
  NOR3_X1    g08744(.A1(new_n8728_), .A2(new_n8729_), .A3(new_n7057_), .ZN(new_n9747_));
  AOI21_X1   g08745(.A1(new_n8723_), .A2(new_n8722_), .B(new_n7070_), .ZN(new_n9748_));
  NOR2_X1    g08746(.A1(new_n9748_), .A2(new_n9747_), .ZN(new_n9749_));
  OAI21_X1   g08747(.A1(new_n9749_), .A2(new_n7048_), .B(new_n8768_), .ZN(new_n9750_));
  NAND2_X1   g08748(.A1(new_n9750_), .A2(new_n9746_), .ZN(new_n9751_));
  NOR2_X1    g08749(.A1(new_n8761_), .A2(new_n8757_), .ZN(new_n9752_));
  OAI21_X1   g08750(.A1(new_n9752_), .A2(new_n8771_), .B(new_n8769_), .ZN(new_n9753_));
  AOI22_X1   g08751(.A1(new_n9753_), .A2(new_n8760_), .B1(new_n9751_), .B2(new_n9745_), .ZN(new_n9754_));
  NOR2_X1    g08752(.A1(new_n9750_), .A2(new_n9746_), .ZN(new_n9755_));
  NOR2_X1    g08753(.A1(new_n9744_), .A2(new_n9743_), .ZN(new_n9756_));
  NOR2_X1    g08754(.A1(new_n8786_), .A2(new_n8732_), .ZN(new_n9757_));
  NOR4_X1    g08755(.A1(new_n9757_), .A2(new_n9755_), .A3(new_n9756_), .A4(new_n8785_), .ZN(new_n9758_));
  NOR2_X1    g08756(.A1(new_n9754_), .A2(new_n9758_), .ZN(new_n9759_));
  NAND2_X1   g08757(.A1(new_n9759_), .A2(new_n9742_), .ZN(new_n9760_));
  AOI22_X1   g08758(.A1(new_n9740_), .A2(new_n8699_), .B1(new_n9738_), .B2(new_n9739_), .ZN(new_n9761_));
  NOR4_X1    g08759(.A1(new_n9736_), .A2(new_n9735_), .A3(new_n9729_), .A4(new_n8795_), .ZN(new_n9762_));
  NOR2_X1    g08760(.A1(new_n9761_), .A2(new_n9762_), .ZN(new_n9763_));
  OAI22_X1   g08761(.A1(new_n9757_), .A2(new_n8785_), .B1(new_n9755_), .B2(new_n9756_), .ZN(new_n9764_));
  NAND4_X1   g08762(.A1(new_n9753_), .A2(new_n9745_), .A3(new_n9751_), .A4(new_n8760_), .ZN(new_n9765_));
  NAND2_X1   g08763(.A1(new_n9764_), .A2(new_n9765_), .ZN(new_n9766_));
  NAND2_X1   g08764(.A1(new_n9763_), .A2(new_n9766_), .ZN(new_n9767_));
  AOI21_X1   g08765(.A1(new_n9767_), .A2(new_n9760_), .B(new_n9726_), .ZN(new_n9768_));
  OAI21_X1   g08766(.A1(new_n8720_), .A2(new_n8810_), .B(new_n8780_), .ZN(new_n9769_));
  NOR2_X1    g08767(.A1(new_n9763_), .A2(new_n9766_), .ZN(new_n9770_));
  NOR2_X1    g08768(.A1(new_n9759_), .A2(new_n9742_), .ZN(new_n9771_));
  NOR3_X1    g08769(.A1(new_n9770_), .A2(new_n9771_), .A3(new_n9769_), .ZN(new_n9772_));
  NOR2_X1    g08770(.A1(new_n9768_), .A2(new_n9772_), .ZN(new_n9773_));
  NAND2_X1   g08771(.A1(new_n9773_), .A2(new_n9725_), .ZN(new_n9774_));
  AOI21_X1   g08772(.A1(new_n9723_), .A2(new_n9722_), .B(new_n9721_), .ZN(new_n9775_));
  NOR3_X1    g08773(.A1(new_n9710_), .A2(new_n9719_), .A3(new_n9676_), .ZN(new_n9776_));
  NOR2_X1    g08774(.A1(new_n9775_), .A2(new_n9776_), .ZN(new_n9777_));
  OAI21_X1   g08775(.A1(new_n9770_), .A2(new_n9771_), .B(new_n9769_), .ZN(new_n9778_));
  NAND3_X1   g08776(.A1(new_n9767_), .A2(new_n9760_), .A3(new_n9726_), .ZN(new_n9779_));
  NAND2_X1   g08777(.A1(new_n9778_), .A2(new_n9779_), .ZN(new_n9780_));
  NAND2_X1   g08778(.A1(new_n9780_), .A2(new_n9777_), .ZN(new_n9781_));
  AOI21_X1   g08779(.A1(new_n9781_), .A2(new_n9774_), .B(new_n9675_), .ZN(new_n9782_));
  OAI21_X1   g08780(.A1(new_n8805_), .A2(new_n8792_), .B(new_n8806_), .ZN(new_n9783_));
  OAI21_X1   g08781(.A1(new_n8664_), .A2(new_n8822_), .B(new_n9783_), .ZN(new_n9784_));
  NOR2_X1    g08782(.A1(new_n9780_), .A2(new_n9777_), .ZN(new_n9785_));
  NOR2_X1    g08783(.A1(new_n9773_), .A2(new_n9725_), .ZN(new_n9786_));
  NOR3_X1    g08784(.A1(new_n9785_), .A2(new_n9786_), .A3(new_n9784_), .ZN(new_n9787_));
  NOR2_X1    g08785(.A1(new_n9782_), .A2(new_n9787_), .ZN(new_n9788_));
  OAI21_X1   g08786(.A1(new_n9072_), .A2(new_n9061_), .B(new_n9073_), .ZN(new_n9789_));
  OAI21_X1   g08787(.A1(new_n9091_), .A2(new_n9074_), .B(new_n9789_), .ZN(new_n9790_));
  AOI21_X1   g08788(.A1(new_n8944_), .A2(new_n9088_), .B(new_n8946_), .ZN(new_n9791_));
  AOI21_X1   g08789(.A1(new_n8934_), .A2(new_n6907_), .B(new_n8858_), .ZN(new_n9792_));
  NOR2_X1    g08790(.A1(new_n8834_), .A2(new_n8833_), .ZN(new_n9793_));
  OAI21_X1   g08791(.A1(new_n9793_), .A2(new_n6946_), .B(new_n8864_), .ZN(new_n9794_));
  NOR2_X1    g08792(.A1(new_n9792_), .A2(new_n9794_), .ZN(new_n9795_));
  OAI21_X1   g08793(.A1(new_n8851_), .A2(new_n6959_), .B(new_n8845_), .ZN(new_n9796_));
  NAND2_X1   g08794(.A1(new_n8865_), .A2(new_n8866_), .ZN(new_n9797_));
  AOI21_X1   g08795(.A1(new_n9797_), .A2(new_n6964_), .B(new_n8830_), .ZN(new_n9798_));
  NOR2_X1    g08796(.A1(new_n9796_), .A2(new_n9798_), .ZN(new_n9799_));
  AOI21_X1   g08797(.A1(new_n8859_), .A2(new_n8856_), .B(new_n8835_), .ZN(new_n9800_));
  OAI22_X1   g08798(.A1(new_n8937_), .A2(new_n9800_), .B1(new_n9799_), .B2(new_n9795_), .ZN(new_n9801_));
  NAND2_X1   g08799(.A1(new_n9796_), .A2(new_n9798_), .ZN(new_n9802_));
  NAND2_X1   g08800(.A1(new_n9792_), .A2(new_n9794_), .ZN(new_n9803_));
  OAI21_X1   g08801(.A1(new_n8870_), .A2(new_n8872_), .B(new_n8867_), .ZN(new_n9804_));
  NAND4_X1   g08802(.A1(new_n8854_), .A2(new_n9804_), .A3(new_n9802_), .A4(new_n9803_), .ZN(new_n9805_));
  NAND2_X1   g08803(.A1(new_n9801_), .A2(new_n9805_), .ZN(new_n9806_));
  NAND2_X1   g08804(.A1(new_n8926_), .A2(new_n8927_), .ZN(new_n9807_));
  OAI21_X1   g08805(.A1(new_n8892_), .A2(new_n6801_), .B(new_n9807_), .ZN(new_n9808_));
  NAND2_X1   g08806(.A1(new_n8911_), .A2(new_n8910_), .ZN(new_n9809_));
  AOI21_X1   g08807(.A1(new_n9809_), .A2(new_n6841_), .B(new_n8880_), .ZN(new_n9810_));
  NAND2_X1   g08808(.A1(new_n9810_), .A2(new_n9808_), .ZN(new_n9811_));
  AOI21_X1   g08809(.A1(new_n8903_), .A2(new_n6855_), .B(new_n8920_), .ZN(new_n9812_));
  NOR2_X1    g08810(.A1(new_n8884_), .A2(new_n8883_), .ZN(new_n9813_));
  OAI21_X1   g08811(.A1(new_n9813_), .A2(new_n6866_), .B(new_n8909_), .ZN(new_n9814_));
  NAND2_X1   g08812(.A1(new_n9814_), .A2(new_n9812_), .ZN(new_n9815_));
  NOR2_X1    g08813(.A1(new_n8928_), .A2(new_n8892_), .ZN(new_n9816_));
  OAI21_X1   g08814(.A1(new_n8913_), .A2(new_n9816_), .B(new_n8912_), .ZN(new_n9817_));
  AOI22_X1   g08815(.A1(new_n9817_), .A2(new_n8898_), .B1(new_n9815_), .B2(new_n9811_), .ZN(new_n9818_));
  NOR2_X1    g08816(.A1(new_n9814_), .A2(new_n9812_), .ZN(new_n9819_));
  NOR2_X1    g08817(.A1(new_n9810_), .A2(new_n9808_), .ZN(new_n9820_));
  AOI21_X1   g08818(.A1(new_n8900_), .A2(new_n8904_), .B(new_n8885_), .ZN(new_n9821_));
  NOR4_X1    g08819(.A1(new_n9821_), .A2(new_n9819_), .A3(new_n9820_), .A4(new_n8922_), .ZN(new_n9822_));
  NOR2_X1    g08820(.A1(new_n9818_), .A2(new_n9822_), .ZN(new_n9823_));
  NAND2_X1   g08821(.A1(new_n9806_), .A2(new_n9823_), .ZN(new_n9824_));
  AOI22_X1   g08822(.A1(new_n9804_), .A2(new_n8854_), .B1(new_n9802_), .B2(new_n9803_), .ZN(new_n9825_));
  NOR4_X1    g08823(.A1(new_n9800_), .A2(new_n9799_), .A3(new_n9795_), .A4(new_n8937_), .ZN(new_n9826_));
  NOR2_X1    g08824(.A1(new_n9825_), .A2(new_n9826_), .ZN(new_n9827_));
  OAI22_X1   g08825(.A1(new_n9821_), .A2(new_n8922_), .B1(new_n9819_), .B2(new_n9820_), .ZN(new_n9828_));
  NAND4_X1   g08826(.A1(new_n9817_), .A2(new_n9811_), .A3(new_n9815_), .A4(new_n8898_), .ZN(new_n9829_));
  NAND2_X1   g08827(.A1(new_n9828_), .A2(new_n9829_), .ZN(new_n9830_));
  NAND2_X1   g08828(.A1(new_n9827_), .A2(new_n9830_), .ZN(new_n9831_));
  AOI21_X1   g08829(.A1(new_n9824_), .A2(new_n9831_), .B(new_n9791_), .ZN(new_n9832_));
  OAI21_X1   g08830(.A1(new_n8875_), .A2(new_n8945_), .B(new_n9089_), .ZN(new_n9833_));
  NOR2_X1    g08831(.A1(new_n9827_), .A2(new_n9830_), .ZN(new_n9834_));
  NOR2_X1    g08832(.A1(new_n9806_), .A2(new_n9823_), .ZN(new_n9835_));
  NOR3_X1    g08833(.A1(new_n9835_), .A2(new_n9834_), .A3(new_n9833_), .ZN(new_n9836_));
  NOR2_X1    g08834(.A1(new_n9832_), .A2(new_n9836_), .ZN(new_n9837_));
  OAI21_X1   g08835(.A1(new_n9000_), .A2(new_n9076_), .B(new_n9042_), .ZN(new_n9838_));
  OAI21_X1   g08836(.A1(new_n8969_), .A2(new_n8981_), .B(new_n8978_), .ZN(new_n9839_));
  NAND4_X1   g08837(.A1(new_n8949_), .A2(new_n8950_), .A3(new_n6725_), .A4(new_n6745_), .ZN(new_n9840_));
  OAI21_X1   g08838(.A1(new_n8955_), .A2(new_n8954_), .B(new_n6754_), .ZN(new_n9841_));
  NAND2_X1   g08839(.A1(new_n9840_), .A2(new_n9841_), .ZN(new_n9842_));
  AOI21_X1   g08840(.A1(new_n9842_), .A2(new_n6761_), .B(new_n8953_), .ZN(new_n9843_));
  NAND2_X1   g08841(.A1(new_n9843_), .A2(new_n9839_), .ZN(new_n9844_));
  AOI22_X1   g08842(.A1(new_n8993_), .A2(new_n6706_), .B1(new_n8975_), .B2(new_n8977_), .ZN(new_n9845_));
  OAI21_X1   g08843(.A1(new_n8989_), .A2(new_n6747_), .B(new_n8988_), .ZN(new_n9846_));
  NAND2_X1   g08844(.A1(new_n9845_), .A2(new_n9846_), .ZN(new_n9847_));
  NAND2_X1   g08845(.A1(new_n8984_), .A2(new_n8990_), .ZN(new_n9848_));
  AOI22_X1   g08846(.A1(new_n9848_), .A2(new_n8980_), .B1(new_n9847_), .B2(new_n9844_), .ZN(new_n9849_));
  NOR2_X1    g08847(.A1(new_n9845_), .A2(new_n9846_), .ZN(new_n9850_));
  NOR2_X1    g08848(.A1(new_n9843_), .A2(new_n9839_), .ZN(new_n9851_));
  NOR2_X1    g08849(.A1(new_n9064_), .A2(new_n8958_), .ZN(new_n9852_));
  NOR4_X1    g08850(.A1(new_n9852_), .A2(new_n9851_), .A3(new_n9850_), .A4(new_n9063_), .ZN(new_n9853_));
  NOR2_X1    g08851(.A1(new_n9853_), .A2(new_n9849_), .ZN(new_n9854_));
  AOI21_X1   g08852(.A1(new_n9022_), .A2(new_n6600_), .B(new_n9017_), .ZN(new_n9855_));
  NOR3_X1    g08853(.A1(new_n9008_), .A2(new_n9009_), .A3(new_n6649_), .ZN(new_n9856_));
  AOI21_X1   g08854(.A1(new_n9003_), .A2(new_n9002_), .B(new_n6672_), .ZN(new_n9857_));
  NOR2_X1    g08855(.A1(new_n9856_), .A2(new_n9857_), .ZN(new_n9858_));
  OAI21_X1   g08856(.A1(new_n9858_), .A2(new_n6640_), .B(new_n9036_), .ZN(new_n9859_));
  NOR2_X1    g08857(.A1(new_n9855_), .A2(new_n9859_), .ZN(new_n9860_));
  OAI21_X1   g08858(.A1(new_n9056_), .A2(new_n6653_), .B(new_n9026_), .ZN(new_n9861_));
  AOI21_X1   g08859(.A1(new_n9011_), .A2(new_n6665_), .B(new_n9006_), .ZN(new_n9862_));
  NOR2_X1    g08860(.A1(new_n9862_), .A2(new_n9861_), .ZN(new_n9863_));
  AOI21_X1   g08861(.A1(new_n9029_), .A2(new_n9031_), .B(new_n9012_), .ZN(new_n9864_));
  OAI22_X1   g08862(.A1(new_n9864_), .A2(new_n9050_), .B1(new_n9860_), .B2(new_n9863_), .ZN(new_n9865_));
  NAND2_X1   g08863(.A1(new_n9862_), .A2(new_n9861_), .ZN(new_n9866_));
  NAND2_X1   g08864(.A1(new_n9855_), .A2(new_n9859_), .ZN(new_n9867_));
  NOR2_X1    g08865(.A1(new_n9057_), .A2(new_n9056_), .ZN(new_n9868_));
  OAI21_X1   g08866(.A1(new_n9868_), .A2(new_n9038_), .B(new_n9037_), .ZN(new_n9869_));
  NAND4_X1   g08867(.A1(new_n9869_), .A2(new_n9866_), .A3(new_n9867_), .A4(new_n9028_), .ZN(new_n9870_));
  NAND2_X1   g08868(.A1(new_n9865_), .A2(new_n9870_), .ZN(new_n9871_));
  NOR2_X1    g08869(.A1(new_n9854_), .A2(new_n9871_), .ZN(new_n9872_));
  OAI22_X1   g08870(.A1(new_n9852_), .A2(new_n9063_), .B1(new_n9850_), .B2(new_n9851_), .ZN(new_n9873_));
  NAND4_X1   g08871(.A1(new_n9848_), .A2(new_n9847_), .A3(new_n9844_), .A4(new_n8980_), .ZN(new_n9874_));
  NAND2_X1   g08872(.A1(new_n9873_), .A2(new_n9874_), .ZN(new_n9875_));
  AOI22_X1   g08873(.A1(new_n9869_), .A2(new_n9028_), .B1(new_n9866_), .B2(new_n9867_), .ZN(new_n9876_));
  NOR4_X1    g08874(.A1(new_n9864_), .A2(new_n9860_), .A3(new_n9863_), .A4(new_n9050_), .ZN(new_n9877_));
  NOR2_X1    g08875(.A1(new_n9877_), .A2(new_n9876_), .ZN(new_n9878_));
  NOR2_X1    g08876(.A1(new_n9878_), .A2(new_n9875_), .ZN(new_n9879_));
  OAI21_X1   g08877(.A1(new_n9879_), .A2(new_n9872_), .B(new_n9838_), .ZN(new_n9880_));
  AOI21_X1   g08878(.A1(new_n9069_), .A2(new_n9060_), .B(new_n9075_), .ZN(new_n9881_));
  NAND2_X1   g08879(.A1(new_n9878_), .A2(new_n9875_), .ZN(new_n9882_));
  NAND2_X1   g08880(.A1(new_n9854_), .A2(new_n9871_), .ZN(new_n9883_));
  NAND3_X1   g08881(.A1(new_n9882_), .A2(new_n9883_), .A3(new_n9881_), .ZN(new_n9884_));
  NAND2_X1   g08882(.A1(new_n9880_), .A2(new_n9884_), .ZN(new_n9885_));
  NOR2_X1    g08883(.A1(new_n9837_), .A2(new_n9885_), .ZN(new_n9886_));
  OAI21_X1   g08884(.A1(new_n9835_), .A2(new_n9834_), .B(new_n9833_), .ZN(new_n9887_));
  NAND3_X1   g08885(.A1(new_n9824_), .A2(new_n9831_), .A3(new_n9791_), .ZN(new_n9888_));
  NAND2_X1   g08886(.A1(new_n9887_), .A2(new_n9888_), .ZN(new_n9889_));
  AOI21_X1   g08887(.A1(new_n9882_), .A2(new_n9883_), .B(new_n9881_), .ZN(new_n9890_));
  NOR3_X1    g08888(.A1(new_n9879_), .A2(new_n9872_), .A3(new_n9838_), .ZN(new_n9891_));
  NOR2_X1    g08889(.A1(new_n9890_), .A2(new_n9891_), .ZN(new_n9892_));
  NOR2_X1    g08890(.A1(new_n9892_), .A2(new_n9889_), .ZN(new_n9893_));
  OAI21_X1   g08891(.A1(new_n9886_), .A2(new_n9893_), .B(new_n9790_), .ZN(new_n9894_));
  NAND3_X1   g08892(.A1(new_n9077_), .A2(new_n9080_), .A3(new_n9081_), .ZN(new_n9895_));
  AOI21_X1   g08893(.A1(new_n8948_), .A2(new_n9895_), .B(new_n9082_), .ZN(new_n9896_));
  NAND2_X1   g08894(.A1(new_n9892_), .A2(new_n9889_), .ZN(new_n9897_));
  NAND2_X1   g08895(.A1(new_n9837_), .A2(new_n9885_), .ZN(new_n9898_));
  NAND3_X1   g08896(.A1(new_n9898_), .A2(new_n9897_), .A3(new_n9896_), .ZN(new_n9899_));
  NAND2_X1   g08897(.A1(new_n9894_), .A2(new_n9899_), .ZN(new_n9900_));
  NOR2_X1    g08898(.A1(new_n9788_), .A2(new_n9900_), .ZN(new_n9901_));
  OAI21_X1   g08899(.A1(new_n9785_), .A2(new_n9786_), .B(new_n9784_), .ZN(new_n9902_));
  NAND3_X1   g08900(.A1(new_n9781_), .A2(new_n9774_), .A3(new_n9675_), .ZN(new_n9903_));
  NAND2_X1   g08901(.A1(new_n9902_), .A2(new_n9903_), .ZN(new_n9904_));
  AOI21_X1   g08902(.A1(new_n9898_), .A2(new_n9897_), .B(new_n9896_), .ZN(new_n9905_));
  NOR3_X1    g08903(.A1(new_n9886_), .A2(new_n9893_), .A3(new_n9790_), .ZN(new_n9906_));
  NOR2_X1    g08904(.A1(new_n9905_), .A2(new_n9906_), .ZN(new_n9907_));
  NOR2_X1    g08905(.A1(new_n9907_), .A2(new_n9904_), .ZN(new_n9908_));
  OAI21_X1   g08906(.A1(new_n9901_), .A2(new_n9908_), .B(new_n9673_), .ZN(new_n9909_));
  AOI22_X1   g08907(.A1(new_n8825_), .A2(new_n9099_), .B1(new_n9097_), .B2(new_n9100_), .ZN(new_n9910_));
  NAND2_X1   g08908(.A1(new_n9907_), .A2(new_n9904_), .ZN(new_n9911_));
  NAND2_X1   g08909(.A1(new_n9788_), .A2(new_n9900_), .ZN(new_n9912_));
  NAND3_X1   g08910(.A1(new_n9912_), .A2(new_n9911_), .A3(new_n9910_), .ZN(new_n9913_));
  NAND2_X1   g08911(.A1(new_n9909_), .A2(new_n9913_), .ZN(new_n9914_));
  AOI22_X1   g08912(.A1(new_n9380_), .A2(new_n9646_), .B1(new_n9641_), .B2(new_n9643_), .ZN(new_n9915_));
  NOR3_X1    g08913(.A1(new_n9375_), .A2(new_n9372_), .A3(new_n9360_), .ZN(new_n9916_));
  OAI21_X1   g08914(.A1(new_n9369_), .A2(new_n9916_), .B(new_n9376_), .ZN(new_n9917_));
  AOI21_X1   g08915(.A1(new_n9234_), .A2(new_n9366_), .B(new_n9236_), .ZN(new_n9918_));
  AOI21_X1   g08916(.A1(new_n9146_), .A2(new_n6101_), .B(new_n9225_), .ZN(new_n9919_));
  NOR3_X1    g08917(.A1(new_n9120_), .A2(new_n9121_), .A3(new_n6149_), .ZN(new_n9920_));
  AOI21_X1   g08918(.A1(new_n9110_), .A2(new_n9114_), .B(new_n9116_), .ZN(new_n9921_));
  NOR2_X1    g08919(.A1(new_n9921_), .A2(new_n9920_), .ZN(new_n9922_));
  OAI21_X1   g08920(.A1(new_n9922_), .A2(new_n6142_), .B(new_n9155_), .ZN(new_n9923_));
  NOR2_X1    g08921(.A1(new_n9919_), .A2(new_n9923_), .ZN(new_n9924_));
  OAI21_X1   g08922(.A1(new_n9135_), .A2(new_n6155_), .B(new_n9130_), .ZN(new_n9925_));
  AOI21_X1   g08923(.A1(new_n9123_), .A2(new_n9152_), .B(new_n9118_), .ZN(new_n9926_));
  NOR2_X1    g08924(.A1(new_n9926_), .A2(new_n9925_), .ZN(new_n9927_));
  NOR2_X1    g08925(.A1(new_n9228_), .A2(new_n9124_), .ZN(new_n9928_));
  OAI22_X1   g08926(.A1(new_n9928_), .A2(new_n9227_), .B1(new_n9924_), .B2(new_n9927_), .ZN(new_n9929_));
  NAND2_X1   g08927(.A1(new_n9926_), .A2(new_n9925_), .ZN(new_n9930_));
  NAND2_X1   g08928(.A1(new_n9919_), .A2(new_n9923_), .ZN(new_n9931_));
  NOR2_X1    g08929(.A1(new_n9230_), .A2(new_n9135_), .ZN(new_n9932_));
  OAI21_X1   g08930(.A1(new_n9932_), .A2(new_n9158_), .B(new_n9156_), .ZN(new_n9933_));
  NAND4_X1   g08931(.A1(new_n9933_), .A2(new_n9930_), .A3(new_n9931_), .A4(new_n9138_), .ZN(new_n9934_));
  NAND2_X1   g08932(.A1(new_n9929_), .A2(new_n9934_), .ZN(new_n9935_));
  OAI21_X1   g08933(.A1(new_n9217_), .A2(new_n6046_), .B(new_n9185_), .ZN(new_n9936_));
  NAND2_X1   g08934(.A1(new_n9197_), .A2(new_n9196_), .ZN(new_n9937_));
  AOI21_X1   g08935(.A1(new_n9937_), .A2(new_n6061_), .B(new_n9166_), .ZN(new_n9938_));
  NAND2_X1   g08936(.A1(new_n9938_), .A2(new_n9936_), .ZN(new_n9939_));
  AOI21_X1   g08937(.A1(new_n9181_), .A2(new_n5993_), .B(new_n9176_), .ZN(new_n9940_));
  NOR2_X1    g08938(.A1(new_n9170_), .A2(new_n9169_), .ZN(new_n9941_));
  OAI21_X1   g08939(.A1(new_n9941_), .A2(new_n6033_), .B(new_n9195_), .ZN(new_n9942_));
  NAND2_X1   g08940(.A1(new_n9942_), .A2(new_n9940_), .ZN(new_n9943_));
  NOR2_X1    g08941(.A1(new_n9218_), .A2(new_n9217_), .ZN(new_n9944_));
  OAI21_X1   g08942(.A1(new_n9944_), .A2(new_n9199_), .B(new_n9198_), .ZN(new_n9945_));
  AOI22_X1   g08943(.A1(new_n9945_), .A2(new_n9187_), .B1(new_n9943_), .B2(new_n9939_), .ZN(new_n9946_));
  NOR2_X1    g08944(.A1(new_n9942_), .A2(new_n9940_), .ZN(new_n9947_));
  NOR2_X1    g08945(.A1(new_n9938_), .A2(new_n9936_), .ZN(new_n9948_));
  NOR2_X1    g08946(.A1(new_n9212_), .A2(new_n9171_), .ZN(new_n9949_));
  NOR4_X1    g08947(.A1(new_n9949_), .A2(new_n9947_), .A3(new_n9948_), .A4(new_n9211_), .ZN(new_n9950_));
  NOR2_X1    g08948(.A1(new_n9946_), .A2(new_n9950_), .ZN(new_n9951_));
  NAND2_X1   g08949(.A1(new_n9935_), .A2(new_n9951_), .ZN(new_n9952_));
  AOI22_X1   g08950(.A1(new_n9933_), .A2(new_n9138_), .B1(new_n9930_), .B2(new_n9931_), .ZN(new_n9953_));
  NOR4_X1    g08951(.A1(new_n9928_), .A2(new_n9924_), .A3(new_n9927_), .A4(new_n9227_), .ZN(new_n9954_));
  NOR2_X1    g08952(.A1(new_n9953_), .A2(new_n9954_), .ZN(new_n9955_));
  OAI22_X1   g08953(.A1(new_n9949_), .A2(new_n9211_), .B1(new_n9947_), .B2(new_n9948_), .ZN(new_n9956_));
  NAND4_X1   g08954(.A1(new_n9945_), .A2(new_n9939_), .A3(new_n9943_), .A4(new_n9187_), .ZN(new_n9957_));
  NAND2_X1   g08955(.A1(new_n9956_), .A2(new_n9957_), .ZN(new_n9958_));
  NAND2_X1   g08956(.A1(new_n9955_), .A2(new_n9958_), .ZN(new_n9959_));
  AOI21_X1   g08957(.A1(new_n9952_), .A2(new_n9959_), .B(new_n9918_), .ZN(new_n9960_));
  OAI21_X1   g08958(.A1(new_n9161_), .A2(new_n9235_), .B(new_n9367_), .ZN(new_n9961_));
  NOR2_X1    g08959(.A1(new_n9955_), .A2(new_n9958_), .ZN(new_n9962_));
  NOR2_X1    g08960(.A1(new_n9935_), .A2(new_n9951_), .ZN(new_n9963_));
  NOR3_X1    g08961(.A1(new_n9963_), .A2(new_n9962_), .A3(new_n9961_), .ZN(new_n9964_));
  NOR2_X1    g08962(.A1(new_n9960_), .A2(new_n9964_), .ZN(new_n9965_));
  OAI21_X1   g08963(.A1(new_n9284_), .A2(new_n9355_), .B(new_n9374_), .ZN(new_n9966_));
  OAI21_X1   g08964(.A1(new_n9278_), .A2(new_n5896_), .B(new_n9275_), .ZN(new_n9967_));
  NAND2_X1   g08965(.A1(new_n9249_), .A2(new_n9248_), .ZN(new_n9968_));
  AOI21_X1   g08966(.A1(new_n9968_), .A2(new_n5928_), .B(new_n9269_), .ZN(new_n9969_));
  NAND2_X1   g08967(.A1(new_n9969_), .A2(new_n9967_), .ZN(new_n9970_));
  AOI21_X1   g08968(.A1(new_n9257_), .A2(new_n5953_), .B(new_n9349_), .ZN(new_n9971_));
  NOR2_X1    g08969(.A1(new_n9271_), .A2(new_n9270_), .ZN(new_n9972_));
  OAI21_X1   g08970(.A1(new_n9972_), .A2(new_n5955_), .B(new_n9245_), .ZN(new_n9973_));
  NAND2_X1   g08971(.A1(new_n9971_), .A2(new_n9973_), .ZN(new_n9974_));
  NOR2_X1    g08972(.A1(new_n9344_), .A2(new_n9278_), .ZN(new_n9975_));
  OAI21_X1   g08973(.A1(new_n9264_), .A2(new_n9975_), .B(new_n9250_), .ZN(new_n9976_));
  AOI22_X1   g08974(.A1(new_n9976_), .A2(new_n9281_), .B1(new_n9970_), .B2(new_n9974_), .ZN(new_n9977_));
  NOR2_X1    g08975(.A1(new_n9971_), .A2(new_n9973_), .ZN(new_n9978_));
  NOR2_X1    g08976(.A1(new_n9969_), .A2(new_n9967_), .ZN(new_n9979_));
  AOI21_X1   g08977(.A1(new_n9259_), .A2(new_n9265_), .B(new_n9272_), .ZN(new_n9980_));
  NOR4_X1    g08978(.A1(new_n9980_), .A2(new_n9979_), .A3(new_n9978_), .A4(new_n9351_), .ZN(new_n9981_));
  NOR2_X1    g08979(.A1(new_n9977_), .A2(new_n9981_), .ZN(new_n9982_));
  AOI21_X1   g08980(.A1(new_n9321_), .A2(new_n5791_), .B(new_n9333_), .ZN(new_n9983_));
  OAI21_X1   g08981(.A1(new_n9317_), .A2(new_n5823_), .B(new_n9316_), .ZN(new_n9984_));
  NOR2_X1    g08982(.A1(new_n9983_), .A2(new_n9984_), .ZN(new_n9985_));
  NAND2_X1   g08983(.A1(new_n9309_), .A2(new_n9308_), .ZN(new_n9986_));
  OAI21_X1   g08984(.A1(new_n9301_), .A2(new_n5845_), .B(new_n9986_), .ZN(new_n9987_));
  NAND3_X1   g08985(.A1(new_n9286_), .A2(new_n9285_), .A3(new_n5855_), .ZN(new_n9988_));
  OAI21_X1   g08986(.A1(new_n9290_), .A2(new_n9291_), .B(new_n5831_), .ZN(new_n9989_));
  NAND2_X1   g08987(.A1(new_n9989_), .A2(new_n9988_), .ZN(new_n9990_));
  AOI21_X1   g08988(.A1(new_n9990_), .A2(new_n5849_), .B(new_n9289_), .ZN(new_n9991_));
  NOR2_X1    g08989(.A1(new_n9991_), .A2(new_n9987_), .ZN(new_n9992_));
  NAND2_X1   g08990(.A1(new_n9306_), .A2(new_n9321_), .ZN(new_n9993_));
  AOI21_X1   g08991(.A1(new_n9993_), .A2(new_n9311_), .B(new_n9294_), .ZN(new_n9994_));
  OAI22_X1   g08992(.A1(new_n9994_), .A2(new_n9335_), .B1(new_n9985_), .B2(new_n9992_), .ZN(new_n9995_));
  NAND2_X1   g08993(.A1(new_n9991_), .A2(new_n9987_), .ZN(new_n9996_));
  NAND2_X1   g08994(.A1(new_n9983_), .A2(new_n9984_), .ZN(new_n9997_));
  NAND2_X1   g08995(.A1(new_n9312_), .A2(new_n9318_), .ZN(new_n9998_));
  NAND4_X1   g08996(.A1(new_n9998_), .A2(new_n9996_), .A3(new_n9997_), .A4(new_n9307_), .ZN(new_n9999_));
  NAND2_X1   g08997(.A1(new_n9995_), .A2(new_n9999_), .ZN(new_n10000_));
  NOR2_X1    g08998(.A1(new_n9982_), .A2(new_n10000_), .ZN(new_n10001_));
  OAI22_X1   g08999(.A1(new_n9980_), .A2(new_n9351_), .B1(new_n9979_), .B2(new_n9978_), .ZN(new_n10002_));
  NAND4_X1   g09000(.A1(new_n9976_), .A2(new_n9970_), .A3(new_n9974_), .A4(new_n9281_), .ZN(new_n10003_));
  NAND2_X1   g09001(.A1(new_n10002_), .A2(new_n10003_), .ZN(new_n10004_));
  AOI22_X1   g09002(.A1(new_n9998_), .A2(new_n9307_), .B1(new_n9996_), .B2(new_n9997_), .ZN(new_n10005_));
  NOR4_X1    g09003(.A1(new_n9994_), .A2(new_n9985_), .A3(new_n9992_), .A4(new_n9335_), .ZN(new_n10006_));
  NOR2_X1    g09004(.A1(new_n10005_), .A2(new_n10006_), .ZN(new_n10007_));
  NOR2_X1    g09005(.A1(new_n10004_), .A2(new_n10007_), .ZN(new_n10008_));
  OAI21_X1   g09006(.A1(new_n10008_), .A2(new_n10001_), .B(new_n9966_), .ZN(new_n10009_));
  AOI21_X1   g09007(.A1(new_n9354_), .A2(new_n9373_), .B(new_n9356_), .ZN(new_n10010_));
  NAND2_X1   g09008(.A1(new_n10004_), .A2(new_n10007_), .ZN(new_n10011_));
  NAND2_X1   g09009(.A1(new_n9982_), .A2(new_n10000_), .ZN(new_n10012_));
  NAND3_X1   g09010(.A1(new_n10011_), .A2(new_n10012_), .A3(new_n10010_), .ZN(new_n10013_));
  NAND2_X1   g09011(.A1(new_n10009_), .A2(new_n10013_), .ZN(new_n10014_));
  NOR2_X1    g09012(.A1(new_n9965_), .A2(new_n10014_), .ZN(new_n10015_));
  OAI21_X1   g09013(.A1(new_n9963_), .A2(new_n9962_), .B(new_n9961_), .ZN(new_n10016_));
  NAND3_X1   g09014(.A1(new_n9952_), .A2(new_n9959_), .A3(new_n9918_), .ZN(new_n10017_));
  NAND2_X1   g09015(.A1(new_n10016_), .A2(new_n10017_), .ZN(new_n10018_));
  AOI21_X1   g09016(.A1(new_n10011_), .A2(new_n10012_), .B(new_n10010_), .ZN(new_n10019_));
  NOR3_X1    g09017(.A1(new_n10008_), .A2(new_n10001_), .A3(new_n9966_), .ZN(new_n10020_));
  NOR2_X1    g09018(.A1(new_n10019_), .A2(new_n10020_), .ZN(new_n10021_));
  NOR2_X1    g09019(.A1(new_n10018_), .A2(new_n10021_), .ZN(new_n10022_));
  OAI21_X1   g09020(.A1(new_n10022_), .A2(new_n10015_), .B(new_n9917_), .ZN(new_n10023_));
  AOI22_X1   g09021(.A1(new_n9377_), .A2(new_n9238_), .B1(new_n9358_), .B2(new_n9360_), .ZN(new_n10024_));
  NAND2_X1   g09022(.A1(new_n10018_), .A2(new_n10021_), .ZN(new_n10025_));
  NAND2_X1   g09023(.A1(new_n9965_), .A2(new_n10014_), .ZN(new_n10026_));
  NAND3_X1   g09024(.A1(new_n10025_), .A2(new_n10026_), .A3(new_n10024_), .ZN(new_n10027_));
  NAND2_X1   g09025(.A1(new_n10023_), .A2(new_n10027_), .ZN(new_n10028_));
  AOI21_X1   g09026(.A1(new_n9486_), .A2(new_n9647_), .B(new_n9631_), .ZN(new_n10029_));
  NAND2_X1   g09027(.A1(new_n9418_), .A2(new_n9419_), .ZN(new_n10030_));
  NOR4_X1    g09028(.A1(new_n9417_), .A2(new_n10030_), .A3(new_n6491_), .A4(new_n6554_), .ZN(new_n10031_));
  AOI21_X1   g09029(.A1(new_n10030_), .A2(new_n6542_), .B(new_n6557_), .ZN(new_n10032_));
  NAND2_X1   g09030(.A1(new_n10031_), .A2(new_n10032_), .ZN(new_n10033_));
  OAI21_X1   g09031(.A1(new_n9420_), .A2(new_n9417_), .B(new_n9422_), .ZN(new_n10034_));
  AOI21_X1   g09032(.A1(new_n10033_), .A2(new_n10034_), .B(new_n9414_), .ZN(new_n10035_));
  INV_X1     g09033(.I(new_n9424_), .ZN(new_n10036_));
  NOR2_X1    g09034(.A1(new_n10036_), .A2(new_n10035_), .ZN(new_n10037_));
  OAI21_X1   g09035(.A1(new_n9481_), .A2(new_n9466_), .B(new_n9482_), .ZN(new_n10038_));
  OAI21_X1   g09036(.A1(new_n10037_), .A2(new_n9483_), .B(new_n10038_), .ZN(new_n10039_));
  AOI22_X1   g09037(.A1(new_n9399_), .A2(new_n6542_), .B1(new_n9418_), .B2(new_n9419_), .ZN(new_n10040_));
  OAI21_X1   g09038(.A1(new_n9391_), .A2(new_n6554_), .B(new_n9386_), .ZN(new_n10041_));
  NOR2_X1    g09039(.A1(new_n10040_), .A2(new_n10041_), .ZN(new_n10042_));
  OAI21_X1   g09040(.A1(new_n9417_), .A2(new_n6491_), .B(new_n10030_), .ZN(new_n10043_));
  AOI21_X1   g09041(.A1(new_n9413_), .A2(new_n6529_), .B(new_n9410_), .ZN(new_n10044_));
  NOR2_X1    g09042(.A1(new_n10044_), .A2(new_n10043_), .ZN(new_n10045_));
  NOR2_X1    g09043(.A1(new_n9407_), .A2(new_n9414_), .ZN(new_n10046_));
  OAI22_X1   g09044(.A1(new_n10046_), .A2(new_n9405_), .B1(new_n10042_), .B2(new_n10045_), .ZN(new_n10047_));
  NAND2_X1   g09045(.A1(new_n10044_), .A2(new_n10043_), .ZN(new_n10048_));
  NAND2_X1   g09046(.A1(new_n10040_), .A2(new_n10041_), .ZN(new_n10049_));
  NAND2_X1   g09047(.A1(new_n10034_), .A2(new_n9392_), .ZN(new_n10050_));
  NAND4_X1   g09048(.A1(new_n10050_), .A2(new_n10048_), .A3(new_n10049_), .A4(new_n10033_), .ZN(new_n10051_));
  AOI22_X1   g09049(.A1(new_n9443_), .A2(new_n6437_), .B1(new_n9459_), .B2(new_n9460_), .ZN(new_n10052_));
  NOR2_X1    g09050(.A1(new_n9470_), .A2(new_n9471_), .ZN(new_n10053_));
  OAI21_X1   g09051(.A1(new_n10053_), .A2(new_n6452_), .B(new_n9431_), .ZN(new_n10054_));
  NOR2_X1    g09052(.A1(new_n10052_), .A2(new_n10054_), .ZN(new_n10055_));
  NAND2_X1   g09053(.A1(new_n9460_), .A2(new_n9459_), .ZN(new_n10056_));
  OAI21_X1   g09054(.A1(new_n9458_), .A2(new_n6388_), .B(new_n10056_), .ZN(new_n10057_));
  NAND2_X1   g09055(.A1(new_n9435_), .A2(new_n9434_), .ZN(new_n10058_));
  AOI21_X1   g09056(.A1(new_n10058_), .A2(new_n6413_), .B(new_n9469_), .ZN(new_n10059_));
  NOR2_X1    g09057(.A1(new_n10059_), .A2(new_n10057_), .ZN(new_n10060_));
  AOI21_X1   g09058(.A1(new_n9455_), .A2(new_n9464_), .B(new_n9472_), .ZN(new_n10061_));
  OAI22_X1   g09059(.A1(new_n9449_), .A2(new_n10061_), .B1(new_n10055_), .B2(new_n10060_), .ZN(new_n10062_));
  NAND2_X1   g09060(.A1(new_n10059_), .A2(new_n10057_), .ZN(new_n10063_));
  NAND2_X1   g09061(.A1(new_n10052_), .A2(new_n10054_), .ZN(new_n10064_));
  OAI21_X1   g09062(.A1(new_n9462_), .A2(new_n9451_), .B(new_n9436_), .ZN(new_n10065_));
  NAND4_X1   g09063(.A1(new_n10065_), .A2(new_n10063_), .A3(new_n10064_), .A4(new_n9479_), .ZN(new_n10066_));
  NAND2_X1   g09064(.A1(new_n10062_), .A2(new_n10066_), .ZN(new_n10067_));
  AOI21_X1   g09065(.A1(new_n10047_), .A2(new_n10051_), .B(new_n10067_), .ZN(new_n10068_));
  NAND2_X1   g09066(.A1(new_n10047_), .A2(new_n10051_), .ZN(new_n10069_));
  AOI22_X1   g09067(.A1(new_n10065_), .A2(new_n9479_), .B1(new_n10063_), .B2(new_n10064_), .ZN(new_n10070_));
  NOR4_X1    g09068(.A1(new_n10061_), .A2(new_n10055_), .A3(new_n10060_), .A4(new_n9449_), .ZN(new_n10071_));
  NOR2_X1    g09069(.A1(new_n10070_), .A2(new_n10071_), .ZN(new_n10072_));
  NOR2_X1    g09070(.A1(new_n10072_), .A2(new_n10069_), .ZN(new_n10073_));
  OAI21_X1   g09071(.A1(new_n10068_), .A2(new_n10073_), .B(new_n10039_), .ZN(new_n10074_));
  NAND3_X1   g09072(.A1(new_n9453_), .A2(new_n9475_), .A3(new_n9454_), .ZN(new_n10075_));
  AOI21_X1   g09073(.A1(new_n9425_), .A2(new_n10075_), .B(new_n9484_), .ZN(new_n10076_));
  NAND2_X1   g09074(.A1(new_n10072_), .A2(new_n10069_), .ZN(new_n10077_));
  NAND3_X1   g09075(.A1(new_n10067_), .A2(new_n10047_), .A3(new_n10051_), .ZN(new_n10078_));
  NAND3_X1   g09076(.A1(new_n10077_), .A2(new_n10078_), .A3(new_n10076_), .ZN(new_n10079_));
  NAND2_X1   g09077(.A1(new_n10074_), .A2(new_n10079_), .ZN(new_n10080_));
  AOI21_X1   g09078(.A1(new_n9618_), .A2(new_n9595_), .B(new_n9625_), .ZN(new_n10081_));
  AOI21_X1   g09079(.A1(new_n9509_), .A2(new_n6298_), .B(new_n9613_), .ZN(new_n10082_));
  NOR2_X1    g09080(.A1(new_n9527_), .A2(new_n9526_), .ZN(new_n10083_));
  OAI21_X1   g09081(.A1(new_n10083_), .A2(new_n9519_), .B(new_n9497_), .ZN(new_n10084_));
  NOR2_X1    g09082(.A1(new_n10082_), .A2(new_n10084_), .ZN(new_n10085_));
  OAI21_X1   g09083(.A1(new_n9534_), .A2(new_n6345_), .B(new_n9531_), .ZN(new_n10086_));
  NAND2_X1   g09084(.A1(new_n9500_), .A2(new_n9501_), .ZN(new_n10087_));
  AOI21_X1   g09085(.A1(new_n10087_), .A2(new_n6335_), .B(new_n9525_), .ZN(new_n10088_));
  NOR2_X1    g09086(.A1(new_n10088_), .A2(new_n10086_), .ZN(new_n10089_));
  AOI21_X1   g09087(.A1(new_n9521_), .A2(new_n9511_), .B(new_n9528_), .ZN(new_n10090_));
  OAI22_X1   g09088(.A1(new_n10090_), .A2(new_n9615_), .B1(new_n10085_), .B2(new_n10089_), .ZN(new_n10091_));
  NAND2_X1   g09089(.A1(new_n10088_), .A2(new_n10086_), .ZN(new_n10092_));
  NAND2_X1   g09090(.A1(new_n10082_), .A2(new_n10084_), .ZN(new_n10093_));
  AOI21_X1   g09091(.A1(new_n9531_), .A2(new_n6298_), .B(new_n9534_), .ZN(new_n10094_));
  OAI21_X1   g09092(.A1(new_n10094_), .A2(new_n9520_), .B(new_n9502_), .ZN(new_n10095_));
  NAND4_X1   g09093(.A1(new_n10095_), .A2(new_n10092_), .A3(new_n10093_), .A4(new_n9537_), .ZN(new_n10096_));
  NAND2_X1   g09094(.A1(new_n10091_), .A2(new_n10096_), .ZN(new_n10097_));
  OAI21_X1   g09095(.A1(new_n9586_), .A2(new_n6247_), .B(new_n9597_), .ZN(new_n10098_));
  NAND2_X1   g09096(.A1(new_n9559_), .A2(new_n9560_), .ZN(new_n10099_));
  AOI21_X1   g09097(.A1(new_n10099_), .A2(new_n6256_), .B(new_n9580_), .ZN(new_n10100_));
  NAND2_X1   g09098(.A1(new_n10100_), .A2(new_n10098_), .ZN(new_n10101_));
  AOI21_X1   g09099(.A1(new_n9568_), .A2(new_n6209_), .B(new_n9572_), .ZN(new_n10102_));
  NOR2_X1    g09100(.A1(new_n9582_), .A2(new_n9581_), .ZN(new_n10103_));
  OAI21_X1   g09101(.A1(new_n10103_), .A2(new_n6235_), .B(new_n9556_), .ZN(new_n10104_));
  NAND2_X1   g09102(.A1(new_n10102_), .A2(new_n10104_), .ZN(new_n10105_));
  NOR2_X1    g09103(.A1(new_n9589_), .A2(new_n9586_), .ZN(new_n10106_));
  OAI21_X1   g09104(.A1(new_n10106_), .A2(new_n9576_), .B(new_n9561_), .ZN(new_n10107_));
  AOI22_X1   g09105(.A1(new_n10107_), .A2(new_n9599_), .B1(new_n10105_), .B2(new_n10101_), .ZN(new_n10108_));
  NOR2_X1    g09106(.A1(new_n10102_), .A2(new_n10104_), .ZN(new_n10109_));
  NOR2_X1    g09107(.A1(new_n10100_), .A2(new_n10098_), .ZN(new_n10110_));
  AOI21_X1   g09108(.A1(new_n9600_), .A2(new_n9591_), .B(new_n9583_), .ZN(new_n10111_));
  NOR4_X1    g09109(.A1(new_n10111_), .A2(new_n10109_), .A3(new_n10110_), .A4(new_n9574_), .ZN(new_n10112_));
  NOR2_X1    g09110(.A1(new_n10108_), .A2(new_n10112_), .ZN(new_n10113_));
  NAND2_X1   g09111(.A1(new_n10097_), .A2(new_n10113_), .ZN(new_n10114_));
  AOI22_X1   g09112(.A1(new_n10095_), .A2(new_n9537_), .B1(new_n10093_), .B2(new_n10092_), .ZN(new_n10115_));
  NOR4_X1    g09113(.A1(new_n10090_), .A2(new_n10085_), .A3(new_n10089_), .A4(new_n9615_), .ZN(new_n10116_));
  NOR2_X1    g09114(.A1(new_n10115_), .A2(new_n10116_), .ZN(new_n10117_));
  OAI22_X1   g09115(.A1(new_n10111_), .A2(new_n9574_), .B1(new_n10109_), .B2(new_n10110_), .ZN(new_n10118_));
  NAND4_X1   g09116(.A1(new_n10107_), .A2(new_n10101_), .A3(new_n10105_), .A4(new_n9599_), .ZN(new_n10119_));
  NAND2_X1   g09117(.A1(new_n10118_), .A2(new_n10119_), .ZN(new_n10120_));
  NAND2_X1   g09118(.A1(new_n10117_), .A2(new_n10120_), .ZN(new_n10121_));
  AOI21_X1   g09119(.A1(new_n10114_), .A2(new_n10121_), .B(new_n10081_), .ZN(new_n10122_));
  OAI21_X1   g09120(.A1(new_n9540_), .A2(new_n9624_), .B(new_n9607_), .ZN(new_n10123_));
  NOR2_X1    g09121(.A1(new_n10117_), .A2(new_n10120_), .ZN(new_n10124_));
  NOR2_X1    g09122(.A1(new_n10097_), .A2(new_n10113_), .ZN(new_n10125_));
  NOR3_X1    g09123(.A1(new_n10125_), .A2(new_n10124_), .A3(new_n10123_), .ZN(new_n10126_));
  NOR2_X1    g09124(.A1(new_n10126_), .A2(new_n10122_), .ZN(new_n10127_));
  NAND2_X1   g09125(.A1(new_n10080_), .A2(new_n10127_), .ZN(new_n10128_));
  AOI21_X1   g09126(.A1(new_n10077_), .A2(new_n10078_), .B(new_n10076_), .ZN(new_n10129_));
  NOR3_X1    g09127(.A1(new_n10068_), .A2(new_n10073_), .A3(new_n10039_), .ZN(new_n10130_));
  NOR2_X1    g09128(.A1(new_n10130_), .A2(new_n10129_), .ZN(new_n10131_));
  OAI21_X1   g09129(.A1(new_n10125_), .A2(new_n10124_), .B(new_n10123_), .ZN(new_n10132_));
  NAND3_X1   g09130(.A1(new_n10114_), .A2(new_n10121_), .A3(new_n10081_), .ZN(new_n10133_));
  NAND2_X1   g09131(.A1(new_n10132_), .A2(new_n10133_), .ZN(new_n10134_));
  NAND2_X1   g09132(.A1(new_n10131_), .A2(new_n10134_), .ZN(new_n10135_));
  AOI21_X1   g09133(.A1(new_n10128_), .A2(new_n10135_), .B(new_n10029_), .ZN(new_n10136_));
  OAI21_X1   g09134(.A1(new_n9635_), .A2(new_n9623_), .B(new_n9648_), .ZN(new_n10137_));
  NOR2_X1    g09135(.A1(new_n10131_), .A2(new_n10134_), .ZN(new_n10138_));
  NOR2_X1    g09136(.A1(new_n10080_), .A2(new_n10127_), .ZN(new_n10139_));
  NOR3_X1    g09137(.A1(new_n10139_), .A2(new_n10138_), .A3(new_n10137_), .ZN(new_n10140_));
  NOR2_X1    g09138(.A1(new_n10136_), .A2(new_n10140_), .ZN(new_n10141_));
  NAND2_X1   g09139(.A1(new_n10141_), .A2(new_n10028_), .ZN(new_n10142_));
  AOI21_X1   g09140(.A1(new_n10025_), .A2(new_n10026_), .B(new_n10024_), .ZN(new_n10143_));
  NOR3_X1    g09141(.A1(new_n10022_), .A2(new_n10015_), .A3(new_n9917_), .ZN(new_n10144_));
  NOR2_X1    g09142(.A1(new_n10143_), .A2(new_n10144_), .ZN(new_n10145_));
  OAI21_X1   g09143(.A1(new_n10139_), .A2(new_n10138_), .B(new_n10137_), .ZN(new_n10146_));
  NAND3_X1   g09144(.A1(new_n10128_), .A2(new_n10135_), .A3(new_n10029_), .ZN(new_n10147_));
  NAND2_X1   g09145(.A1(new_n10146_), .A2(new_n10147_), .ZN(new_n10148_));
  NAND2_X1   g09146(.A1(new_n10145_), .A2(new_n10148_), .ZN(new_n10149_));
  AOI21_X1   g09147(.A1(new_n10142_), .A2(new_n10149_), .B(new_n9915_), .ZN(new_n10150_));
  NOR3_X1    g09148(.A1(new_n9649_), .A2(new_n9650_), .A3(new_n9641_), .ZN(new_n10151_));
  OAI21_X1   g09149(.A1(new_n9379_), .A2(new_n10151_), .B(new_n9651_), .ZN(new_n10152_));
  NOR2_X1    g09150(.A1(new_n10145_), .A2(new_n10148_), .ZN(new_n10153_));
  NOR2_X1    g09151(.A1(new_n10141_), .A2(new_n10028_), .ZN(new_n10154_));
  NOR3_X1    g09152(.A1(new_n10154_), .A2(new_n10153_), .A3(new_n10152_), .ZN(new_n10155_));
  NOR2_X1    g09153(.A1(new_n10150_), .A2(new_n10155_), .ZN(new_n10156_));
  NAND2_X1   g09154(.A1(new_n10156_), .A2(new_n9914_), .ZN(new_n10157_));
  AOI21_X1   g09155(.A1(new_n9912_), .A2(new_n9911_), .B(new_n9910_), .ZN(new_n10158_));
  NOR3_X1    g09156(.A1(new_n9901_), .A2(new_n9908_), .A3(new_n9673_), .ZN(new_n10159_));
  NOR2_X1    g09157(.A1(new_n10158_), .A2(new_n10159_), .ZN(new_n10160_));
  OAI21_X1   g09158(.A1(new_n10154_), .A2(new_n10153_), .B(new_n10152_), .ZN(new_n10161_));
  NAND3_X1   g09159(.A1(new_n10142_), .A2(new_n10149_), .A3(new_n9915_), .ZN(new_n10162_));
  NAND2_X1   g09160(.A1(new_n10161_), .A2(new_n10162_), .ZN(new_n10163_));
  NAND2_X1   g09161(.A1(new_n10160_), .A2(new_n10163_), .ZN(new_n10164_));
  AOI21_X1   g09162(.A1(new_n10164_), .A2(new_n10157_), .B(new_n9671_), .ZN(new_n10165_));
  OAI21_X1   g09163(.A1(new_n9660_), .A2(new_n9662_), .B(new_n9661_), .ZN(new_n10166_));
  NOR2_X1    g09164(.A1(new_n10160_), .A2(new_n10163_), .ZN(new_n10167_));
  NOR2_X1    g09165(.A1(new_n10156_), .A2(new_n9914_), .ZN(new_n10168_));
  NOR3_X1    g09166(.A1(new_n10167_), .A2(new_n10168_), .A3(new_n10166_), .ZN(new_n10169_));
  NOR2_X1    g09167(.A1(new_n10165_), .A2(new_n10169_), .ZN(new_n10170_));
  NOR2_X1    g09168(.A1(new_n8525_), .A2(new_n8533_), .ZN(new_n10171_));
  OAI22_X1   g09169(.A1(new_n7970_), .A2(new_n8538_), .B1(new_n8534_), .B2(new_n10171_), .ZN(new_n10172_));
  AOI22_X1   g09170(.A1(new_n7675_), .A2(new_n7964_), .B1(new_n7961_), .B2(new_n7965_), .ZN(new_n10173_));
  NOR3_X1    g09171(.A1(new_n7652_), .A2(new_n7639_), .A3(new_n7653_), .ZN(new_n10174_));
  OAI21_X1   g09172(.A1(new_n7527_), .A2(new_n10174_), .B(new_n7672_), .ZN(new_n10175_));
  AOI21_X1   g09173(.A1(new_n7441_), .A2(new_n7524_), .B(new_n7668_), .ZN(new_n10176_));
  AOI21_X1   g09174(.A1(new_n7412_), .A2(new_n5689_), .B(new_n7418_), .ZN(new_n10177_));
  NOR2_X1    g09175(.A1(new_n7432_), .A2(new_n7431_), .ZN(new_n10178_));
  OAI21_X1   g09176(.A1(new_n10178_), .A2(new_n5728_), .B(new_n7395_), .ZN(new_n10179_));
  NOR2_X1    g09177(.A1(new_n10179_), .A2(new_n10177_), .ZN(new_n10180_));
  OAI21_X1   g09178(.A1(new_n7514_), .A2(new_n7415_), .B(new_n7425_), .ZN(new_n10181_));
  NAND2_X1   g09179(.A1(new_n7398_), .A2(new_n7399_), .ZN(new_n10182_));
  AOI21_X1   g09180(.A1(new_n10182_), .A2(new_n5742_), .B(new_n7430_), .ZN(new_n10183_));
  NOR2_X1    g09181(.A1(new_n10183_), .A2(new_n10181_), .ZN(new_n10184_));
  AOI21_X1   g09182(.A1(new_n7438_), .A2(new_n7436_), .B(new_n7433_), .ZN(new_n10185_));
  OAI22_X1   g09183(.A1(new_n10185_), .A2(new_n7420_), .B1(new_n10180_), .B2(new_n10184_), .ZN(new_n10186_));
  NAND2_X1   g09184(.A1(new_n10183_), .A2(new_n10181_), .ZN(new_n10187_));
  NAND2_X1   g09185(.A1(new_n10179_), .A2(new_n10177_), .ZN(new_n10188_));
  OAI21_X1   g09186(.A1(new_n7422_), .A2(new_n7426_), .B(new_n7400_), .ZN(new_n10189_));
  NAND4_X1   g09187(.A1(new_n10189_), .A2(new_n10187_), .A3(new_n10188_), .A4(new_n7517_), .ZN(new_n10190_));
  NAND2_X1   g09188(.A1(new_n10186_), .A2(new_n10190_), .ZN(new_n10191_));
  OAI21_X1   g09189(.A1(new_n7483_), .A2(new_n7472_), .B(new_n7502_), .ZN(new_n10192_));
  NAND2_X1   g09190(.A1(new_n7451_), .A2(new_n7450_), .ZN(new_n10193_));
  AOI21_X1   g09191(.A1(new_n10193_), .A2(new_n5650_), .B(new_n7491_), .ZN(new_n10194_));
  NAND2_X1   g09192(.A1(new_n10194_), .A2(new_n10192_), .ZN(new_n10195_));
  AOI21_X1   g09193(.A1(new_n7467_), .A2(new_n5596_), .B(new_n7475_), .ZN(new_n10196_));
  NOR2_X1    g09194(.A1(new_n7493_), .A2(new_n7492_), .ZN(new_n10197_));
  OAI21_X1   g09195(.A1(new_n10197_), .A2(new_n5636_), .B(new_n7447_), .ZN(new_n10198_));
  NAND2_X1   g09196(.A1(new_n10198_), .A2(new_n10196_), .ZN(new_n10199_));
  OAI21_X1   g09197(.A1(new_n7480_), .A2(new_n7487_), .B(new_n7452_), .ZN(new_n10200_));
  AOI22_X1   g09198(.A1(new_n10200_), .A2(new_n7504_), .B1(new_n10199_), .B2(new_n10195_), .ZN(new_n10201_));
  NOR2_X1    g09199(.A1(new_n10194_), .A2(new_n10192_), .ZN(new_n10202_));
  NAND2_X1   g09200(.A1(new_n7508_), .A2(new_n7467_), .ZN(new_n10203_));
  AOI21_X1   g09201(.A1(new_n7495_), .A2(new_n10203_), .B(new_n7494_), .ZN(new_n10204_));
  OAI22_X1   g09202(.A1(new_n10198_), .A2(new_n10196_), .B1(new_n7469_), .B2(new_n7476_), .ZN(new_n10205_));
  NOR3_X1    g09203(.A1(new_n10205_), .A2(new_n10204_), .A3(new_n10202_), .ZN(new_n10206_));
  NOR2_X1    g09204(.A1(new_n10201_), .A2(new_n10206_), .ZN(new_n10207_));
  NAND2_X1   g09205(.A1(new_n10191_), .A2(new_n10207_), .ZN(new_n10208_));
  AOI22_X1   g09206(.A1(new_n10189_), .A2(new_n7517_), .B1(new_n10188_), .B2(new_n10187_), .ZN(new_n10209_));
  OAI22_X1   g09207(.A1(new_n10179_), .A2(new_n10177_), .B1(new_n7414_), .B2(new_n7419_), .ZN(new_n10210_));
  NOR3_X1    g09208(.A1(new_n10210_), .A2(new_n10185_), .A3(new_n10184_), .ZN(new_n10211_));
  NOR2_X1    g09209(.A1(new_n10209_), .A2(new_n10211_), .ZN(new_n10212_));
  NOR2_X1    g09210(.A1(new_n10198_), .A2(new_n10196_), .ZN(new_n10213_));
  OAI22_X1   g09211(.A1(new_n10204_), .A2(new_n7477_), .B1(new_n10213_), .B2(new_n10202_), .ZN(new_n10214_));
  NAND4_X1   g09212(.A1(new_n10200_), .A2(new_n10195_), .A3(new_n10199_), .A4(new_n7504_), .ZN(new_n10215_));
  NAND2_X1   g09213(.A1(new_n10214_), .A2(new_n10215_), .ZN(new_n10216_));
  NAND2_X1   g09214(.A1(new_n10212_), .A2(new_n10216_), .ZN(new_n10217_));
  AOI21_X1   g09215(.A1(new_n10208_), .A2(new_n10217_), .B(new_n10176_), .ZN(new_n10218_));
  OAI21_X1   g09216(.A1(new_n7523_), .A2(new_n7667_), .B(new_n7525_), .ZN(new_n10219_));
  NOR2_X1    g09217(.A1(new_n10212_), .A2(new_n10216_), .ZN(new_n10220_));
  NOR2_X1    g09218(.A1(new_n10191_), .A2(new_n10207_), .ZN(new_n10221_));
  NOR3_X1    g09219(.A1(new_n10221_), .A2(new_n10220_), .A3(new_n10219_), .ZN(new_n10222_));
  NOR2_X1    g09220(.A1(new_n10218_), .A2(new_n10222_), .ZN(new_n10223_));
  OAI21_X1   g09221(.A1(new_n7581_), .A2(new_n7657_), .B(new_n7626_), .ZN(new_n10224_));
  OAI21_X1   g09222(.A1(new_n7552_), .A2(new_n5551_), .B(new_n7558_), .ZN(new_n10225_));
  AOI21_X1   g09223(.A1(new_n7544_), .A2(new_n5559_), .B(new_n7539_), .ZN(new_n10226_));
  NAND2_X1   g09224(.A1(new_n10226_), .A2(new_n10225_), .ZN(new_n10227_));
  AOI22_X1   g09225(.A1(new_n7564_), .A2(new_n5497_), .B1(new_n7555_), .B2(new_n7557_), .ZN(new_n10228_));
  OAI21_X1   g09226(.A1(new_n7575_), .A2(new_n5538_), .B(new_n7572_), .ZN(new_n10229_));
  NAND2_X1   g09227(.A1(new_n10228_), .A2(new_n10229_), .ZN(new_n10230_));
  OAI21_X1   g09228(.A1(new_n7643_), .A2(new_n7578_), .B(new_n7576_), .ZN(new_n10231_));
  AOI22_X1   g09229(.A1(new_n10231_), .A2(new_n7560_), .B1(new_n10227_), .B2(new_n10230_), .ZN(new_n10232_));
  NOR2_X1    g09230(.A1(new_n10228_), .A2(new_n10229_), .ZN(new_n10233_));
  NOR2_X1    g09231(.A1(new_n10226_), .A2(new_n10225_), .ZN(new_n10234_));
  AOI21_X1   g09232(.A1(new_n7561_), .A2(new_n7567_), .B(new_n7545_), .ZN(new_n10235_));
  NOR4_X1    g09233(.A1(new_n10235_), .A2(new_n10234_), .A3(new_n10233_), .A4(new_n7642_), .ZN(new_n10236_));
  NOR2_X1    g09234(.A1(new_n10232_), .A2(new_n10236_), .ZN(new_n10237_));
  AOI21_X1   g09235(.A1(new_n7610_), .A2(new_n5400_), .B(new_n7629_), .ZN(new_n10238_));
  NOR2_X1    g09236(.A1(new_n7590_), .A2(new_n7591_), .ZN(new_n10239_));
  OAI21_X1   g09237(.A1(new_n10239_), .A2(new_n5429_), .B(new_n7618_), .ZN(new_n10240_));
  NOR2_X1    g09238(.A1(new_n10238_), .A2(new_n10240_), .ZN(new_n10241_));
  OAI21_X1   g09239(.A1(new_n7599_), .A2(new_n5442_), .B(new_n7603_), .ZN(new_n10242_));
  NAND2_X1   g09240(.A1(new_n7620_), .A2(new_n7619_), .ZN(new_n10243_));
  AOI21_X1   g09241(.A1(new_n10243_), .A2(new_n5457_), .B(new_n7587_), .ZN(new_n10244_));
  NOR2_X1    g09242(.A1(new_n10244_), .A2(new_n10242_), .ZN(new_n10245_));
  AOI21_X1   g09243(.A1(new_n7607_), .A2(new_n7613_), .B(new_n7592_), .ZN(new_n10246_));
  OAI22_X1   g09244(.A1(new_n7631_), .A2(new_n10246_), .B1(new_n10241_), .B2(new_n10245_), .ZN(new_n10247_));
  NAND2_X1   g09245(.A1(new_n10244_), .A2(new_n10242_), .ZN(new_n10248_));
  NAND2_X1   g09246(.A1(new_n10238_), .A2(new_n10240_), .ZN(new_n10249_));
  NOR2_X1    g09247(.A1(new_n7635_), .A2(new_n7599_), .ZN(new_n10250_));
  OAI21_X1   g09248(.A1(new_n10250_), .A2(new_n7622_), .B(new_n7621_), .ZN(new_n10251_));
  NAND4_X1   g09249(.A1(new_n10251_), .A2(new_n10248_), .A3(new_n10249_), .A4(new_n7606_), .ZN(new_n10252_));
  NAND2_X1   g09250(.A1(new_n10247_), .A2(new_n10252_), .ZN(new_n10253_));
  NOR2_X1    g09251(.A1(new_n10237_), .A2(new_n10253_), .ZN(new_n10254_));
  OAI22_X1   g09252(.A1(new_n10235_), .A2(new_n7642_), .B1(new_n10234_), .B2(new_n10233_), .ZN(new_n10255_));
  NAND4_X1   g09253(.A1(new_n10231_), .A2(new_n10227_), .A3(new_n10230_), .A4(new_n7560_), .ZN(new_n10256_));
  NAND2_X1   g09254(.A1(new_n10256_), .A2(new_n10255_), .ZN(new_n10257_));
  AOI22_X1   g09255(.A1(new_n10251_), .A2(new_n7606_), .B1(new_n10248_), .B2(new_n10249_), .ZN(new_n10258_));
  NOR4_X1    g09256(.A1(new_n10246_), .A2(new_n10241_), .A3(new_n10245_), .A4(new_n7631_), .ZN(new_n10259_));
  NOR2_X1    g09257(.A1(new_n10258_), .A2(new_n10259_), .ZN(new_n10260_));
  NOR2_X1    g09258(.A1(new_n10257_), .A2(new_n10260_), .ZN(new_n10261_));
  OAI21_X1   g09259(.A1(new_n10254_), .A2(new_n10261_), .B(new_n10224_), .ZN(new_n10262_));
  AOI21_X1   g09260(.A1(new_n7649_), .A2(new_n7638_), .B(new_n7656_), .ZN(new_n10263_));
  NAND2_X1   g09261(.A1(new_n10257_), .A2(new_n10260_), .ZN(new_n10264_));
  NAND2_X1   g09262(.A1(new_n10237_), .A2(new_n10253_), .ZN(new_n10265_));
  NAND3_X1   g09263(.A1(new_n10265_), .A2(new_n10264_), .A3(new_n10263_), .ZN(new_n10266_));
  NAND2_X1   g09264(.A1(new_n10262_), .A2(new_n10266_), .ZN(new_n10267_));
  NOR2_X1    g09265(.A1(new_n10267_), .A2(new_n10223_), .ZN(new_n10268_));
  OAI21_X1   g09266(.A1(new_n10221_), .A2(new_n10220_), .B(new_n10219_), .ZN(new_n10269_));
  NAND3_X1   g09267(.A1(new_n10208_), .A2(new_n10217_), .A3(new_n10176_), .ZN(new_n10270_));
  NAND2_X1   g09268(.A1(new_n10270_), .A2(new_n10269_), .ZN(new_n10271_));
  AOI21_X1   g09269(.A1(new_n10265_), .A2(new_n10264_), .B(new_n10263_), .ZN(new_n10272_));
  NOR3_X1    g09270(.A1(new_n10254_), .A2(new_n10261_), .A3(new_n10224_), .ZN(new_n10273_));
  NOR2_X1    g09271(.A1(new_n10272_), .A2(new_n10273_), .ZN(new_n10274_));
  NOR2_X1    g09272(.A1(new_n10274_), .A2(new_n10271_), .ZN(new_n10275_));
  OAI21_X1   g09273(.A1(new_n10268_), .A2(new_n10275_), .B(new_n10175_), .ZN(new_n10276_));
  NAND2_X1   g09274(.A1(new_n7658_), .A2(new_n7661_), .ZN(new_n10277_));
  AOI22_X1   g09275(.A1(new_n7671_), .A2(new_n7670_), .B1(new_n10277_), .B2(new_n7653_), .ZN(new_n10278_));
  NAND2_X1   g09276(.A1(new_n10274_), .A2(new_n10271_), .ZN(new_n10279_));
  NAND2_X1   g09277(.A1(new_n10267_), .A2(new_n10223_), .ZN(new_n10280_));
  NAND3_X1   g09278(.A1(new_n10280_), .A2(new_n10279_), .A3(new_n10278_), .ZN(new_n10281_));
  NAND2_X1   g09279(.A1(new_n10276_), .A2(new_n10281_), .ZN(new_n10282_));
  NAND3_X1   g09280(.A1(new_n7936_), .A2(new_n7939_), .A3(new_n7943_), .ZN(new_n10283_));
  AOI21_X1   g09281(.A1(new_n7808_), .A2(new_n10283_), .B(new_n7944_), .ZN(new_n10284_));
  OAI21_X1   g09282(.A1(new_n7726_), .A2(new_n7805_), .B(new_n7951_), .ZN(new_n10285_));
  OAI22_X1   g09283(.A1(new_n7700_), .A2(new_n5351_), .B1(new_n7710_), .B2(new_n7703_), .ZN(new_n10286_));
  NAND2_X1   g09284(.A1(new_n7718_), .A2(new_n7719_), .ZN(new_n10287_));
  AOI21_X1   g09285(.A1(new_n10287_), .A2(new_n5357_), .B(new_n7681_), .ZN(new_n10288_));
  NAND2_X1   g09286(.A1(new_n10286_), .A2(new_n10288_), .ZN(new_n10289_));
  AOI21_X1   g09287(.A1(new_n7795_), .A2(new_n5305_), .B(new_n7711_), .ZN(new_n10290_));
  NOR2_X1    g09288(.A1(new_n7685_), .A2(new_n7684_), .ZN(new_n10291_));
  OAI21_X1   g09289(.A1(new_n10291_), .A2(new_n5334_), .B(new_n7717_), .ZN(new_n10292_));
  NAND2_X1   g09290(.A1(new_n10290_), .A2(new_n10292_), .ZN(new_n10293_));
  OAI21_X1   g09291(.A1(new_n7721_), .A2(new_n7723_), .B(new_n7720_), .ZN(new_n10294_));
  AOI22_X1   g09292(.A1(new_n10294_), .A2(new_n7707_), .B1(new_n10289_), .B2(new_n10293_), .ZN(new_n10295_));
  NOR2_X1    g09293(.A1(new_n10290_), .A2(new_n10292_), .ZN(new_n10296_));
  NOR2_X1    g09294(.A1(new_n10286_), .A2(new_n10288_), .ZN(new_n10297_));
  AOI21_X1   g09295(.A1(new_n7709_), .A2(new_n7712_), .B(new_n7686_), .ZN(new_n10298_));
  NOR4_X1    g09296(.A1(new_n10298_), .A2(new_n10297_), .A3(new_n10296_), .A4(new_n7798_), .ZN(new_n10299_));
  NOR2_X1    g09297(.A1(new_n10295_), .A2(new_n10299_), .ZN(new_n10300_));
  AOI21_X1   g09298(.A1(new_n7761_), .A2(new_n5261_), .B(new_n7780_), .ZN(new_n10301_));
  NOR2_X1    g09299(.A1(new_n7741_), .A2(new_n7740_), .ZN(new_n10302_));
  OAI21_X1   g09300(.A1(new_n10302_), .A2(new_n5273_), .B(new_n7769_), .ZN(new_n10303_));
  NOR2_X1    g09301(.A1(new_n10301_), .A2(new_n10303_), .ZN(new_n10304_));
  OAI21_X1   g09302(.A1(new_n7749_), .A2(new_n5206_), .B(new_n7753_), .ZN(new_n10305_));
  NAND2_X1   g09303(.A1(new_n7771_), .A2(new_n7770_), .ZN(new_n10306_));
  AOI21_X1   g09304(.A1(new_n10306_), .A2(new_n5247_), .B(new_n7737_), .ZN(new_n10307_));
  NOR2_X1    g09305(.A1(new_n10307_), .A2(new_n10305_), .ZN(new_n10308_));
  AOI21_X1   g09306(.A1(new_n7758_), .A2(new_n7764_), .B(new_n7742_), .ZN(new_n10309_));
  OAI22_X1   g09307(.A1(new_n7782_), .A2(new_n10309_), .B1(new_n10304_), .B2(new_n10308_), .ZN(new_n10310_));
  NAND2_X1   g09308(.A1(new_n10307_), .A2(new_n10305_), .ZN(new_n10311_));
  NAND2_X1   g09309(.A1(new_n10301_), .A2(new_n10303_), .ZN(new_n10312_));
  OAI21_X1   g09310(.A1(new_n7774_), .A2(new_n7784_), .B(new_n7772_), .ZN(new_n10313_));
  NAND4_X1   g09311(.A1(new_n10313_), .A2(new_n10311_), .A3(new_n10312_), .A4(new_n7756_), .ZN(new_n10314_));
  NAND2_X1   g09312(.A1(new_n10310_), .A2(new_n10314_), .ZN(new_n10315_));
  NOR2_X1    g09313(.A1(new_n10300_), .A2(new_n10315_), .ZN(new_n10316_));
  OAI22_X1   g09314(.A1(new_n10298_), .A2(new_n7798_), .B1(new_n10297_), .B2(new_n10296_), .ZN(new_n10317_));
  NAND4_X1   g09315(.A1(new_n7707_), .A2(new_n10294_), .A3(new_n10289_), .A4(new_n10293_), .ZN(new_n10318_));
  NAND2_X1   g09316(.A1(new_n10317_), .A2(new_n10318_), .ZN(new_n10319_));
  AOI22_X1   g09317(.A1(new_n10313_), .A2(new_n7756_), .B1(new_n10311_), .B2(new_n10312_), .ZN(new_n10320_));
  NOR4_X1    g09318(.A1(new_n10309_), .A2(new_n10304_), .A3(new_n10308_), .A4(new_n7782_), .ZN(new_n10321_));
  NOR2_X1    g09319(.A1(new_n10320_), .A2(new_n10321_), .ZN(new_n10322_));
  NOR2_X1    g09320(.A1(new_n10319_), .A2(new_n10322_), .ZN(new_n10323_));
  OAI21_X1   g09321(.A1(new_n10323_), .A2(new_n10316_), .B(new_n10285_), .ZN(new_n10324_));
  AOI21_X1   g09322(.A1(new_n7804_), .A2(new_n7950_), .B(new_n7806_), .ZN(new_n10325_));
  NAND2_X1   g09323(.A1(new_n10319_), .A2(new_n10322_), .ZN(new_n10326_));
  NAND2_X1   g09324(.A1(new_n10300_), .A2(new_n10315_), .ZN(new_n10327_));
  NAND3_X1   g09325(.A1(new_n10326_), .A2(new_n10327_), .A3(new_n10325_), .ZN(new_n10328_));
  NAND2_X1   g09326(.A1(new_n10328_), .A2(new_n10324_), .ZN(new_n10329_));
  AOI21_X1   g09327(.A1(new_n7928_), .A2(new_n7904_), .B(new_n7935_), .ZN(new_n10330_));
  AOI21_X1   g09328(.A1(new_n7832_), .A2(new_n5115_), .B(new_n7923_), .ZN(new_n10331_));
  NOR2_X1    g09329(.A1(new_n7852_), .A2(new_n7851_), .ZN(new_n10332_));
  OAI21_X1   g09330(.A1(new_n10332_), .A2(new_n5149_), .B(new_n7820_), .ZN(new_n10333_));
  NOR2_X1    g09331(.A1(new_n10331_), .A2(new_n10333_), .ZN(new_n10334_));
  OAI21_X1   g09332(.A1(new_n7841_), .A2(new_n5161_), .B(new_n7855_), .ZN(new_n10335_));
  NAND2_X1   g09333(.A1(new_n7824_), .A2(new_n7823_), .ZN(new_n10336_));
  AOI21_X1   g09334(.A1(new_n10336_), .A2(new_n5165_), .B(new_n7850_), .ZN(new_n10337_));
  NOR2_X1    g09335(.A1(new_n10337_), .A2(new_n10335_), .ZN(new_n10338_));
  NAND2_X1   g09336(.A1(new_n7837_), .A2(new_n7832_), .ZN(new_n10339_));
  AOI21_X1   g09337(.A1(new_n10339_), .A2(new_n7834_), .B(new_n7853_), .ZN(new_n10340_));
  OAI22_X1   g09338(.A1(new_n10340_), .A2(new_n7925_), .B1(new_n10338_), .B2(new_n10334_), .ZN(new_n10341_));
  NAND2_X1   g09339(.A1(new_n10337_), .A2(new_n10335_), .ZN(new_n10342_));
  NAND2_X1   g09340(.A1(new_n10331_), .A2(new_n10333_), .ZN(new_n10343_));
  OAI21_X1   g09341(.A1(new_n7919_), .A2(new_n7843_), .B(new_n7825_), .ZN(new_n10344_));
  NAND4_X1   g09342(.A1(new_n10344_), .A2(new_n10342_), .A3(new_n10343_), .A4(new_n7857_), .ZN(new_n10345_));
  NAND2_X1   g09343(.A1(new_n10341_), .A2(new_n10345_), .ZN(new_n10346_));
  OAI21_X1   g09344(.A1(new_n7895_), .A2(new_n5065_), .B(new_n7906_), .ZN(new_n10347_));
  NAND4_X1   g09345(.A1(new_n7868_), .A2(new_n7869_), .A3(new_n5042_), .A4(new_n5049_), .ZN(new_n10348_));
  OAI21_X1   g09346(.A1(new_n7862_), .A2(new_n7861_), .B(new_n5038_), .ZN(new_n10349_));
  NAND2_X1   g09347(.A1(new_n10348_), .A2(new_n10349_), .ZN(new_n10350_));
  AOI21_X1   g09348(.A1(new_n10350_), .A2(new_n5072_), .B(new_n7891_), .ZN(new_n10351_));
  NAND2_X1   g09349(.A1(new_n10351_), .A2(new_n10347_), .ZN(new_n10352_));
  AOI21_X1   g09350(.A1(new_n7879_), .A2(new_n5010_), .B(new_n7883_), .ZN(new_n10353_));
  OAI21_X1   g09351(.A1(new_n7871_), .A2(new_n5051_), .B(new_n7866_), .ZN(new_n10354_));
  NAND2_X1   g09352(.A1(new_n10353_), .A2(new_n10354_), .ZN(new_n10355_));
  NAND2_X1   g09353(.A1(new_n7909_), .A2(new_n7872_), .ZN(new_n10356_));
  AOI22_X1   g09354(.A1(new_n10356_), .A2(new_n7908_), .B1(new_n10355_), .B2(new_n10352_), .ZN(new_n10357_));
  NOR2_X1    g09355(.A1(new_n10353_), .A2(new_n10354_), .ZN(new_n10358_));
  NOR2_X1    g09356(.A1(new_n10351_), .A2(new_n10347_), .ZN(new_n10359_));
  AOI21_X1   g09357(.A1(new_n7900_), .A2(new_n7912_), .B(new_n7892_), .ZN(new_n10360_));
  NOR4_X1    g09358(.A1(new_n10360_), .A2(new_n10358_), .A3(new_n10359_), .A4(new_n7885_), .ZN(new_n10361_));
  NOR2_X1    g09359(.A1(new_n10357_), .A2(new_n10361_), .ZN(new_n10362_));
  NAND2_X1   g09360(.A1(new_n10346_), .A2(new_n10362_), .ZN(new_n10363_));
  AOI22_X1   g09361(.A1(new_n10344_), .A2(new_n7857_), .B1(new_n10342_), .B2(new_n10343_), .ZN(new_n10364_));
  OAI22_X1   g09362(.A1(new_n10331_), .A2(new_n10333_), .B1(new_n7922_), .B2(new_n7924_), .ZN(new_n10365_));
  NOR3_X1    g09363(.A1(new_n10365_), .A2(new_n10340_), .A3(new_n10338_), .ZN(new_n10366_));
  NOR2_X1    g09364(.A1(new_n10366_), .A2(new_n10364_), .ZN(new_n10367_));
  OAI22_X1   g09365(.A1(new_n10360_), .A2(new_n7885_), .B1(new_n10358_), .B2(new_n10359_), .ZN(new_n10368_));
  NAND4_X1   g09366(.A1(new_n10356_), .A2(new_n10352_), .A3(new_n10355_), .A4(new_n7908_), .ZN(new_n10369_));
  NAND2_X1   g09367(.A1(new_n10368_), .A2(new_n10369_), .ZN(new_n10370_));
  NAND2_X1   g09368(.A1(new_n10367_), .A2(new_n10370_), .ZN(new_n10371_));
  AOI21_X1   g09369(.A1(new_n10363_), .A2(new_n10371_), .B(new_n10330_), .ZN(new_n10372_));
  OAI21_X1   g09370(.A1(new_n7860_), .A2(new_n7934_), .B(new_n7916_), .ZN(new_n10373_));
  NOR2_X1    g09371(.A1(new_n10367_), .A2(new_n10370_), .ZN(new_n10374_));
  NOR2_X1    g09372(.A1(new_n10346_), .A2(new_n10362_), .ZN(new_n10375_));
  NOR3_X1    g09373(.A1(new_n10375_), .A2(new_n10374_), .A3(new_n10373_), .ZN(new_n10376_));
  NOR2_X1    g09374(.A1(new_n10372_), .A2(new_n10376_), .ZN(new_n10377_));
  NAND2_X1   g09375(.A1(new_n10329_), .A2(new_n10377_), .ZN(new_n10378_));
  AOI21_X1   g09376(.A1(new_n10326_), .A2(new_n10327_), .B(new_n10325_), .ZN(new_n10379_));
  NOR3_X1    g09377(.A1(new_n10323_), .A2(new_n10316_), .A3(new_n10285_), .ZN(new_n10380_));
  NOR2_X1    g09378(.A1(new_n10379_), .A2(new_n10380_), .ZN(new_n10381_));
  OAI21_X1   g09379(.A1(new_n10375_), .A2(new_n10374_), .B(new_n10373_), .ZN(new_n10382_));
  NAND3_X1   g09380(.A1(new_n10363_), .A2(new_n10371_), .A3(new_n10330_), .ZN(new_n10383_));
  NAND2_X1   g09381(.A1(new_n10382_), .A2(new_n10383_), .ZN(new_n10384_));
  NAND2_X1   g09382(.A1(new_n10381_), .A2(new_n10384_), .ZN(new_n10385_));
  AOI21_X1   g09383(.A1(new_n10378_), .A2(new_n10385_), .B(new_n10284_), .ZN(new_n10386_));
  OAI21_X1   g09384(.A1(new_n7931_), .A2(new_n7917_), .B(new_n7932_), .ZN(new_n10387_));
  OAI21_X1   g09385(.A1(new_n7953_), .A2(new_n7933_), .B(new_n10387_), .ZN(new_n10388_));
  NOR2_X1    g09386(.A1(new_n10381_), .A2(new_n10384_), .ZN(new_n10389_));
  NOR2_X1    g09387(.A1(new_n10329_), .A2(new_n10377_), .ZN(new_n10390_));
  NOR3_X1    g09388(.A1(new_n10390_), .A2(new_n10389_), .A3(new_n10388_), .ZN(new_n10391_));
  NOR2_X1    g09389(.A1(new_n10386_), .A2(new_n10391_), .ZN(new_n10392_));
  NAND2_X1   g09390(.A1(new_n10392_), .A2(new_n10282_), .ZN(new_n10393_));
  AOI21_X1   g09391(.A1(new_n10280_), .A2(new_n10279_), .B(new_n10278_), .ZN(new_n10394_));
  NOR3_X1    g09392(.A1(new_n10268_), .A2(new_n10275_), .A3(new_n10175_), .ZN(new_n10395_));
  NOR2_X1    g09393(.A1(new_n10394_), .A2(new_n10395_), .ZN(new_n10396_));
  OAI21_X1   g09394(.A1(new_n10390_), .A2(new_n10389_), .B(new_n10388_), .ZN(new_n10397_));
  NAND3_X1   g09395(.A1(new_n10378_), .A2(new_n10385_), .A3(new_n10284_), .ZN(new_n10398_));
  NAND2_X1   g09396(.A1(new_n10397_), .A2(new_n10398_), .ZN(new_n10399_));
  NAND2_X1   g09397(.A1(new_n10396_), .A2(new_n10399_), .ZN(new_n10400_));
  AOI21_X1   g09398(.A1(new_n10393_), .A2(new_n10400_), .B(new_n10173_), .ZN(new_n10401_));
  NAND2_X1   g09399(.A1(new_n7675_), .A2(new_n7964_), .ZN(new_n10402_));
  NAND2_X1   g09400(.A1(new_n10402_), .A2(new_n7966_), .ZN(new_n10403_));
  NOR2_X1    g09401(.A1(new_n10396_), .A2(new_n10399_), .ZN(new_n10404_));
  NOR2_X1    g09402(.A1(new_n10392_), .A2(new_n10282_), .ZN(new_n10405_));
  NOR3_X1    g09403(.A1(new_n10405_), .A2(new_n10404_), .A3(new_n10403_), .ZN(new_n10406_));
  NOR2_X1    g09404(.A1(new_n10401_), .A2(new_n10406_), .ZN(new_n10407_));
  NAND2_X1   g09405(.A1(new_n8521_), .A2(new_n8252_), .ZN(new_n10408_));
  NAND2_X1   g09406(.A1(new_n10408_), .A2(new_n8524_), .ZN(new_n10409_));
  NAND3_X1   g09407(.A1(new_n8217_), .A2(new_n8231_), .A3(new_n8233_), .ZN(new_n10410_));
  AOI21_X1   g09408(.A1(new_n8248_), .A2(new_n10410_), .B(new_n8249_), .ZN(new_n10411_));
  OAI21_X1   g09409(.A1(new_n8098_), .A2(new_n8245_), .B(new_n8100_), .ZN(new_n10412_));
  OAI21_X1   g09410(.A1(new_n8088_), .A2(new_n4494_), .B(new_n8085_), .ZN(new_n10413_));
  AOI21_X1   g09411(.A1(new_n8011_), .A2(new_n4532_), .B(new_n8010_), .ZN(new_n10414_));
  NAND2_X1   g09412(.A1(new_n10413_), .A2(new_n10414_), .ZN(new_n10415_));
  AOI22_X1   g09413(.A1(new_n7998_), .A2(new_n7984_), .B1(new_n8083_), .B2(new_n8084_), .ZN(new_n10416_));
  NOR3_X1    g09414(.A1(new_n7972_), .A2(new_n7971_), .A3(new_n4554_), .ZN(new_n10417_));
  AOI21_X1   g09415(.A1(new_n7977_), .A2(new_n7978_), .B(new_n4541_), .ZN(new_n10418_));
  NOR2_X1    g09416(.A1(new_n10418_), .A2(new_n10417_), .ZN(new_n10419_));
  OAI21_X1   g09417(.A1(new_n10419_), .A2(new_n4547_), .B(new_n7976_), .ZN(new_n10420_));
  NAND2_X1   g09418(.A1(new_n10416_), .A2(new_n10420_), .ZN(new_n10421_));
  NOR2_X1    g09419(.A1(new_n8090_), .A2(new_n8088_), .ZN(new_n10422_));
  OAI21_X1   g09420(.A1(new_n10422_), .A2(new_n8006_), .B(new_n7981_), .ZN(new_n10423_));
  AOI22_X1   g09421(.A1(new_n10423_), .A2(new_n8092_), .B1(new_n10415_), .B2(new_n10421_), .ZN(new_n10424_));
  NOR2_X1    g09422(.A1(new_n10416_), .A2(new_n10420_), .ZN(new_n10425_));
  NOR2_X1    g09423(.A1(new_n10413_), .A2(new_n10414_), .ZN(new_n10426_));
  NOR2_X1    g09424(.A1(new_n8007_), .A2(new_n8012_), .ZN(new_n10427_));
  NOR4_X1    g09425(.A1(new_n10427_), .A2(new_n10425_), .A3(new_n10426_), .A4(new_n8005_), .ZN(new_n10428_));
  NOR2_X1    g09426(.A1(new_n10424_), .A2(new_n10428_), .ZN(new_n10429_));
  AOI22_X1   g09427(.A1(new_n8043_), .A2(new_n4451_), .B1(new_n8063_), .B2(new_n8064_), .ZN(new_n10430_));
  NOR2_X1    g09428(.A1(new_n8055_), .A2(new_n8056_), .ZN(new_n10431_));
  OAI21_X1   g09429(.A1(new_n10431_), .A2(new_n4461_), .B(new_n8031_), .ZN(new_n10432_));
  NOR2_X1    g09430(.A1(new_n10430_), .A2(new_n10432_), .ZN(new_n10433_));
  OAI21_X1   g09431(.A1(new_n8062_), .A2(new_n4391_), .B(new_n8070_), .ZN(new_n10434_));
  NAND2_X1   g09432(.A1(new_n8035_), .A2(new_n8034_), .ZN(new_n10435_));
  AOI21_X1   g09433(.A1(new_n10435_), .A2(new_n4436_), .B(new_n8054_), .ZN(new_n10436_));
  NOR2_X1    g09434(.A1(new_n10436_), .A2(new_n10434_), .ZN(new_n10437_));
  AOI21_X1   g09435(.A1(new_n8058_), .A2(new_n8074_), .B(new_n8057_), .ZN(new_n10438_));
  OAI22_X1   g09436(.A1(new_n10438_), .A2(new_n8049_), .B1(new_n10433_), .B2(new_n10437_), .ZN(new_n10439_));
  NAND2_X1   g09437(.A1(new_n10436_), .A2(new_n10434_), .ZN(new_n10440_));
  NAND2_X1   g09438(.A1(new_n10430_), .A2(new_n10432_), .ZN(new_n10441_));
  NOR2_X1    g09439(.A1(new_n8065_), .A2(new_n8062_), .ZN(new_n10442_));
  OAI21_X1   g09440(.A1(new_n10442_), .A2(new_n8050_), .B(new_n8036_), .ZN(new_n10443_));
  NAND4_X1   g09441(.A1(new_n10443_), .A2(new_n10440_), .A3(new_n10441_), .A4(new_n8073_), .ZN(new_n10444_));
  NAND2_X1   g09442(.A1(new_n10439_), .A2(new_n10444_), .ZN(new_n10445_));
  NOR2_X1    g09443(.A1(new_n10429_), .A2(new_n10445_), .ZN(new_n10446_));
  OAI22_X1   g09444(.A1(new_n10427_), .A2(new_n8005_), .B1(new_n10426_), .B2(new_n10425_), .ZN(new_n10447_));
  NAND4_X1   g09445(.A1(new_n8092_), .A2(new_n10423_), .A3(new_n10415_), .A4(new_n10421_), .ZN(new_n10448_));
  NAND2_X1   g09446(.A1(new_n10447_), .A2(new_n10448_), .ZN(new_n10449_));
  AOI22_X1   g09447(.A1(new_n10443_), .A2(new_n8073_), .B1(new_n10441_), .B2(new_n10440_), .ZN(new_n10450_));
  NOR4_X1    g09448(.A1(new_n10438_), .A2(new_n10433_), .A3(new_n10437_), .A4(new_n8049_), .ZN(new_n10451_));
  NOR2_X1    g09449(.A1(new_n10450_), .A2(new_n10451_), .ZN(new_n10452_));
  NOR2_X1    g09450(.A1(new_n10449_), .A2(new_n10452_), .ZN(new_n10453_));
  OAI21_X1   g09451(.A1(new_n10453_), .A2(new_n10446_), .B(new_n10412_), .ZN(new_n10454_));
  AOI21_X1   g09452(.A1(new_n8018_), .A2(new_n8099_), .B(new_n8246_), .ZN(new_n10455_));
  NAND2_X1   g09453(.A1(new_n10449_), .A2(new_n10452_), .ZN(new_n10456_));
  NAND2_X1   g09454(.A1(new_n10429_), .A2(new_n10445_), .ZN(new_n10457_));
  NAND3_X1   g09455(.A1(new_n10456_), .A2(new_n10457_), .A3(new_n10455_), .ZN(new_n10458_));
  NAND2_X1   g09456(.A1(new_n10454_), .A2(new_n10458_), .ZN(new_n10459_));
  AOI21_X1   g09457(.A1(new_n8228_), .A2(new_n8237_), .B(new_n8230_), .ZN(new_n10460_));
  AOI21_X1   g09458(.A1(new_n8131_), .A2(new_n4314_), .B(new_n8223_), .ZN(new_n10461_));
  NOR2_X1    g09459(.A1(new_n8145_), .A2(new_n8146_), .ZN(new_n10462_));
  OAI21_X1   g09460(.A1(new_n10462_), .A2(new_n4341_), .B(new_n8119_), .ZN(new_n10463_));
  NOR2_X1    g09461(.A1(new_n10461_), .A2(new_n10463_), .ZN(new_n10464_));
  OAI21_X1   g09462(.A1(new_n8153_), .A2(new_n4369_), .B(new_n8150_), .ZN(new_n10465_));
  NAND2_X1   g09463(.A1(new_n8123_), .A2(new_n8122_), .ZN(new_n10466_));
  AOI21_X1   g09464(.A1(new_n10466_), .A2(new_n8106_), .B(new_n8144_), .ZN(new_n10467_));
  NOR2_X1    g09465(.A1(new_n10467_), .A2(new_n10465_), .ZN(new_n10468_));
  AOI21_X1   g09466(.A1(new_n8134_), .A2(new_n8140_), .B(new_n8147_), .ZN(new_n10469_));
  OAI22_X1   g09467(.A1(new_n10469_), .A2(new_n8225_), .B1(new_n10468_), .B2(new_n10464_), .ZN(new_n10470_));
  NAND2_X1   g09468(.A1(new_n10467_), .A2(new_n10465_), .ZN(new_n10471_));
  NAND2_X1   g09469(.A1(new_n10461_), .A2(new_n10463_), .ZN(new_n10472_));
  NOR2_X1    g09470(.A1(new_n8218_), .A2(new_n8153_), .ZN(new_n10473_));
  OAI21_X1   g09471(.A1(new_n8139_), .A2(new_n10473_), .B(new_n8124_), .ZN(new_n10474_));
  NAND4_X1   g09472(.A1(new_n10474_), .A2(new_n10471_), .A3(new_n10472_), .A4(new_n8156_), .ZN(new_n10475_));
  NAND2_X1   g09473(.A1(new_n10470_), .A2(new_n10475_), .ZN(new_n10476_));
  OAI21_X1   g09474(.A1(new_n8176_), .A2(new_n4260_), .B(new_n8182_), .ZN(new_n10477_));
  NAND4_X1   g09475(.A1(new_n8160_), .A2(new_n8161_), .A3(new_n4216_), .A4(new_n4234_), .ZN(new_n10478_));
  OAI21_X1   g09476(.A1(new_n8166_), .A2(new_n8165_), .B(new_n4246_), .ZN(new_n10479_));
  NAND2_X1   g09477(.A1(new_n10478_), .A2(new_n10479_), .ZN(new_n10480_));
  AOI21_X1   g09478(.A1(new_n10480_), .A2(new_n4264_), .B(new_n8164_), .ZN(new_n10481_));
  NAND2_X1   g09479(.A1(new_n10481_), .A2(new_n10477_), .ZN(new_n10482_));
  AOI21_X1   g09480(.A1(new_n8196_), .A2(new_n4209_), .B(new_n8207_), .ZN(new_n10483_));
  OAI21_X1   g09481(.A1(new_n8192_), .A2(new_n4236_), .B(new_n8191_), .ZN(new_n10484_));
  NAND2_X1   g09482(.A1(new_n10484_), .A2(new_n10483_), .ZN(new_n10485_));
  NAND2_X1   g09483(.A1(new_n8187_), .A2(new_n8193_), .ZN(new_n10486_));
  AOI22_X1   g09484(.A1(new_n10486_), .A2(new_n8184_), .B1(new_n10485_), .B2(new_n10482_), .ZN(new_n10487_));
  NOR2_X1    g09485(.A1(new_n10484_), .A2(new_n10483_), .ZN(new_n10488_));
  NOR2_X1    g09486(.A1(new_n10481_), .A2(new_n10477_), .ZN(new_n10489_));
  AOI21_X1   g09487(.A1(new_n8201_), .A2(new_n8186_), .B(new_n8169_), .ZN(new_n10490_));
  NOR4_X1    g09488(.A1(new_n10490_), .A2(new_n10488_), .A3(new_n10489_), .A4(new_n8209_), .ZN(new_n10491_));
  NOR2_X1    g09489(.A1(new_n10487_), .A2(new_n10491_), .ZN(new_n10492_));
  NAND2_X1   g09490(.A1(new_n10476_), .A2(new_n10492_), .ZN(new_n10493_));
  AOI22_X1   g09491(.A1(new_n10474_), .A2(new_n8156_), .B1(new_n10471_), .B2(new_n10472_), .ZN(new_n10494_));
  NOR4_X1    g09492(.A1(new_n10469_), .A2(new_n10468_), .A3(new_n10464_), .A4(new_n8225_), .ZN(new_n10495_));
  NOR2_X1    g09493(.A1(new_n10494_), .A2(new_n10495_), .ZN(new_n10496_));
  OAI22_X1   g09494(.A1(new_n10490_), .A2(new_n8209_), .B1(new_n10488_), .B2(new_n10489_), .ZN(new_n10497_));
  NAND4_X1   g09495(.A1(new_n10486_), .A2(new_n10482_), .A3(new_n10485_), .A4(new_n8184_), .ZN(new_n10498_));
  NAND2_X1   g09496(.A1(new_n10497_), .A2(new_n10498_), .ZN(new_n10499_));
  NAND2_X1   g09497(.A1(new_n10496_), .A2(new_n10499_), .ZN(new_n10500_));
  AOI21_X1   g09498(.A1(new_n10493_), .A2(new_n10500_), .B(new_n10460_), .ZN(new_n10501_));
  OAI21_X1   g09499(.A1(new_n8159_), .A2(new_n8229_), .B(new_n8238_), .ZN(new_n10502_));
  NOR2_X1    g09500(.A1(new_n10496_), .A2(new_n10499_), .ZN(new_n10503_));
  NOR2_X1    g09501(.A1(new_n10476_), .A2(new_n10492_), .ZN(new_n10504_));
  NOR3_X1    g09502(.A1(new_n10504_), .A2(new_n10503_), .A3(new_n10502_), .ZN(new_n10505_));
  NOR2_X1    g09503(.A1(new_n10501_), .A2(new_n10505_), .ZN(new_n10506_));
  NAND2_X1   g09504(.A1(new_n10459_), .A2(new_n10506_), .ZN(new_n10507_));
  AOI21_X1   g09505(.A1(new_n10456_), .A2(new_n10457_), .B(new_n10455_), .ZN(new_n10508_));
  NOR3_X1    g09506(.A1(new_n10453_), .A2(new_n10446_), .A3(new_n10412_), .ZN(new_n10509_));
  NOR2_X1    g09507(.A1(new_n10508_), .A2(new_n10509_), .ZN(new_n10510_));
  OAI21_X1   g09508(.A1(new_n10504_), .A2(new_n10503_), .B(new_n10502_), .ZN(new_n10511_));
  NAND3_X1   g09509(.A1(new_n10493_), .A2(new_n10500_), .A3(new_n10460_), .ZN(new_n10512_));
  NAND2_X1   g09510(.A1(new_n10511_), .A2(new_n10512_), .ZN(new_n10513_));
  NAND2_X1   g09511(.A1(new_n10510_), .A2(new_n10513_), .ZN(new_n10514_));
  AOI21_X1   g09512(.A1(new_n10507_), .A2(new_n10514_), .B(new_n10411_), .ZN(new_n10515_));
  NOR2_X1    g09513(.A1(new_n8239_), .A2(new_n8236_), .ZN(new_n10516_));
  OAI22_X1   g09514(.A1(new_n8102_), .A2(new_n8250_), .B1(new_n10516_), .B2(new_n8233_), .ZN(new_n10517_));
  NOR2_X1    g09515(.A1(new_n10510_), .A2(new_n10513_), .ZN(new_n10518_));
  NOR2_X1    g09516(.A1(new_n10459_), .A2(new_n10506_), .ZN(new_n10519_));
  NOR3_X1    g09517(.A1(new_n10519_), .A2(new_n10518_), .A3(new_n10517_), .ZN(new_n10520_));
  NOR2_X1    g09518(.A1(new_n10515_), .A2(new_n10520_), .ZN(new_n10521_));
  NOR2_X1    g09519(.A1(new_n8484_), .A2(new_n8498_), .ZN(new_n10522_));
  OAI22_X1   g09520(.A1(new_n8516_), .A2(new_n8500_), .B1(new_n10522_), .B2(new_n8507_), .ZN(new_n10523_));
  AOI21_X1   g09521(.A1(new_n8376_), .A2(new_n8513_), .B(new_n8378_), .ZN(new_n10524_));
  AOI21_X1   g09522(.A1(new_n8281_), .A2(new_n4946_), .B(new_n8367_), .ZN(new_n10525_));
  NOR2_X1    g09523(.A1(new_n8261_), .A2(new_n8262_), .ZN(new_n10526_));
  OAI21_X1   g09524(.A1(new_n10526_), .A2(new_n4956_), .B(new_n8289_), .ZN(new_n10527_));
  NOR2_X1    g09525(.A1(new_n10527_), .A2(new_n10525_), .ZN(new_n10528_));
  NAND2_X1   g09526(.A1(new_n8272_), .A2(new_n8274_), .ZN(new_n10529_));
  OAI21_X1   g09527(.A1(new_n8270_), .A2(new_n4893_), .B(new_n10529_), .ZN(new_n10530_));
  NAND2_X1   g09528(.A1(new_n8291_), .A2(new_n8290_), .ZN(new_n10531_));
  AOI21_X1   g09529(.A1(new_n10531_), .A2(new_n4931_), .B(new_n8258_), .ZN(new_n10532_));
  NOR2_X1    g09530(.A1(new_n10532_), .A2(new_n10530_), .ZN(new_n10533_));
  AOI21_X1   g09531(.A1(new_n8278_), .A2(new_n8284_), .B(new_n8263_), .ZN(new_n10534_));
  OAI22_X1   g09532(.A1(new_n10534_), .A2(new_n8370_), .B1(new_n10533_), .B2(new_n10528_), .ZN(new_n10535_));
  NAND2_X1   g09533(.A1(new_n10532_), .A2(new_n10530_), .ZN(new_n10536_));
  NAND2_X1   g09534(.A1(new_n10527_), .A2(new_n10525_), .ZN(new_n10537_));
  OAI21_X1   g09535(.A1(new_n8293_), .A2(new_n8295_), .B(new_n8292_), .ZN(new_n10538_));
  NAND4_X1   g09536(.A1(new_n10538_), .A2(new_n8277_), .A3(new_n10536_), .A4(new_n10537_), .ZN(new_n10539_));
  NAND2_X1   g09537(.A1(new_n10535_), .A2(new_n10539_), .ZN(new_n10540_));
  OAI21_X1   g09538(.A1(new_n8359_), .A2(new_n4800_), .B(new_n8332_), .ZN(new_n10541_));
  NAND2_X1   g09539(.A1(new_n8343_), .A2(new_n8342_), .ZN(new_n10542_));
  AOI21_X1   g09540(.A1(new_n10542_), .A2(new_n4838_), .B(new_n8313_), .ZN(new_n10543_));
  NAND2_X1   g09541(.A1(new_n10543_), .A2(new_n10541_), .ZN(new_n10544_));
  AOI21_X1   g09542(.A1(new_n8325_), .A2(new_n4849_), .B(new_n8328_), .ZN(new_n10545_));
  NOR2_X1    g09543(.A1(new_n8316_), .A2(new_n8317_), .ZN(new_n10546_));
  OAI21_X1   g09544(.A1(new_n10546_), .A2(new_n4860_), .B(new_n8341_), .ZN(new_n10547_));
  NAND2_X1   g09545(.A1(new_n10547_), .A2(new_n10545_), .ZN(new_n10548_));
  OAI21_X1   g09546(.A1(new_n8347_), .A2(new_n8345_), .B(new_n8344_), .ZN(new_n10549_));
  AOI22_X1   g09547(.A1(new_n10549_), .A2(new_n8334_), .B1(new_n10548_), .B2(new_n10544_), .ZN(new_n10550_));
  NOR2_X1    g09548(.A1(new_n10547_), .A2(new_n10545_), .ZN(new_n10551_));
  NOR2_X1    g09549(.A1(new_n10543_), .A2(new_n10541_), .ZN(new_n10552_));
  AOI21_X1   g09550(.A1(new_n8335_), .A2(new_n8336_), .B(new_n8318_), .ZN(new_n10553_));
  NOR4_X1    g09551(.A1(new_n10553_), .A2(new_n10551_), .A3(new_n10552_), .A4(new_n8354_), .ZN(new_n10554_));
  NOR2_X1    g09552(.A1(new_n10550_), .A2(new_n10554_), .ZN(new_n10555_));
  NAND2_X1   g09553(.A1(new_n10540_), .A2(new_n10555_), .ZN(new_n10556_));
  AOI22_X1   g09554(.A1(new_n10538_), .A2(new_n8277_), .B1(new_n10536_), .B2(new_n10537_), .ZN(new_n10557_));
  NOR4_X1    g09555(.A1(new_n10534_), .A2(new_n10528_), .A3(new_n10533_), .A4(new_n8370_), .ZN(new_n10558_));
  NOR2_X1    g09556(.A1(new_n10557_), .A2(new_n10558_), .ZN(new_n10559_));
  OAI22_X1   g09557(.A1(new_n10553_), .A2(new_n8354_), .B1(new_n10551_), .B2(new_n10552_), .ZN(new_n10560_));
  NAND4_X1   g09558(.A1(new_n10549_), .A2(new_n10544_), .A3(new_n10548_), .A4(new_n8334_), .ZN(new_n10561_));
  NAND2_X1   g09559(.A1(new_n10560_), .A2(new_n10561_), .ZN(new_n10562_));
  NAND2_X1   g09560(.A1(new_n10559_), .A2(new_n10562_), .ZN(new_n10563_));
  AOI21_X1   g09561(.A1(new_n10556_), .A2(new_n10563_), .B(new_n10524_), .ZN(new_n10564_));
  OAI21_X1   g09562(.A1(new_n8298_), .A2(new_n8377_), .B(new_n8514_), .ZN(new_n10565_));
  NOR2_X1    g09563(.A1(new_n10559_), .A2(new_n10562_), .ZN(new_n10566_));
  NOR2_X1    g09564(.A1(new_n10540_), .A2(new_n10555_), .ZN(new_n10567_));
  NOR3_X1    g09565(.A1(new_n10567_), .A2(new_n10566_), .A3(new_n10565_), .ZN(new_n10568_));
  NOR2_X1    g09566(.A1(new_n10564_), .A2(new_n10568_), .ZN(new_n10569_));
  OAI21_X1   g09567(.A1(new_n8426_), .A2(new_n8501_), .B(new_n8483_), .ZN(new_n10570_));
  OAI21_X1   g09568(.A1(new_n8417_), .A2(new_n4705_), .B(new_n8421_), .ZN(new_n10571_));
  NAND2_X1   g09569(.A1(new_n8390_), .A2(new_n8389_), .ZN(new_n10572_));
  AOI21_X1   g09570(.A1(new_n10572_), .A2(new_n4745_), .B(new_n8411_), .ZN(new_n10573_));
  NAND2_X1   g09571(.A1(new_n10573_), .A2(new_n10571_), .ZN(new_n10574_));
  AOI21_X1   g09572(.A1(new_n8398_), .A2(new_n4759_), .B(new_n8490_), .ZN(new_n10575_));
  NOR2_X1    g09573(.A1(new_n8412_), .A2(new_n8413_), .ZN(new_n10576_));
  OAI21_X1   g09574(.A1(new_n10576_), .A2(new_n4766_), .B(new_n8386_), .ZN(new_n10577_));
  NAND2_X1   g09575(.A1(new_n10575_), .A2(new_n10577_), .ZN(new_n10578_));
  NOR2_X1    g09576(.A1(new_n8485_), .A2(new_n8417_), .ZN(new_n10579_));
  OAI21_X1   g09577(.A1(new_n8406_), .A2(new_n10579_), .B(new_n8391_), .ZN(new_n10580_));
  AOI22_X1   g09578(.A1(new_n10580_), .A2(new_n8423_), .B1(new_n10574_), .B2(new_n10578_), .ZN(new_n10581_));
  NOR2_X1    g09579(.A1(new_n10575_), .A2(new_n10577_), .ZN(new_n10582_));
  NOR2_X1    g09580(.A1(new_n10573_), .A2(new_n10571_), .ZN(new_n10583_));
  AOI21_X1   g09581(.A1(new_n8400_), .A2(new_n8407_), .B(new_n8414_), .ZN(new_n10584_));
  NOR4_X1    g09582(.A1(new_n10584_), .A2(new_n10582_), .A3(new_n10583_), .A4(new_n8492_), .ZN(new_n10585_));
  NOR2_X1    g09583(.A1(new_n10581_), .A2(new_n10585_), .ZN(new_n10586_));
  AOI21_X1   g09584(.A1(new_n8444_), .A2(new_n4598_), .B(new_n8448_), .ZN(new_n10587_));
  NOR3_X1    g09585(.A1(new_n8427_), .A2(new_n8428_), .A3(new_n4625_), .ZN(new_n10588_));
  AOI21_X1   g09586(.A1(new_n8433_), .A2(new_n8434_), .B(new_n4661_), .ZN(new_n10589_));
  NOR2_X1    g09587(.A1(new_n10589_), .A2(new_n10588_), .ZN(new_n10590_));
  OAI21_X1   g09588(.A1(new_n10590_), .A2(new_n4640_), .B(new_n8432_), .ZN(new_n10591_));
  NOR2_X1    g09589(.A1(new_n10587_), .A2(new_n10591_), .ZN(new_n10592_));
  OAI21_X1   g09590(.A1(new_n8462_), .A2(new_n4655_), .B(new_n8473_), .ZN(new_n10593_));
  AOI22_X1   g09591(.A1(new_n8456_), .A2(new_n4665_), .B1(new_n8429_), .B2(new_n8431_), .ZN(new_n10594_));
  NOR2_X1    g09592(.A1(new_n10594_), .A2(new_n10593_), .ZN(new_n10595_));
  AOI21_X1   g09593(.A1(new_n8467_), .A2(new_n8476_), .B(new_n8459_), .ZN(new_n10596_));
  OAI22_X1   g09594(.A1(new_n8450_), .A2(new_n10596_), .B1(new_n10592_), .B2(new_n10595_), .ZN(new_n10597_));
  NAND2_X1   g09595(.A1(new_n10594_), .A2(new_n10593_), .ZN(new_n10598_));
  NAND2_X1   g09596(.A1(new_n10587_), .A2(new_n10591_), .ZN(new_n10599_));
  NOR2_X1    g09597(.A1(new_n8465_), .A2(new_n8462_), .ZN(new_n10600_));
  OAI21_X1   g09598(.A1(new_n8453_), .A2(new_n10600_), .B(new_n8437_), .ZN(new_n10601_));
  NAND4_X1   g09599(.A1(new_n10601_), .A2(new_n10598_), .A3(new_n10599_), .A4(new_n8475_), .ZN(new_n10602_));
  NAND2_X1   g09600(.A1(new_n10597_), .A2(new_n10602_), .ZN(new_n10603_));
  NOR2_X1    g09601(.A1(new_n10586_), .A2(new_n10603_), .ZN(new_n10604_));
  OAI22_X1   g09602(.A1(new_n8492_), .A2(new_n10584_), .B1(new_n10582_), .B2(new_n10583_), .ZN(new_n10605_));
  NAND4_X1   g09603(.A1(new_n10580_), .A2(new_n10574_), .A3(new_n10578_), .A4(new_n8423_), .ZN(new_n10606_));
  NAND2_X1   g09604(.A1(new_n10605_), .A2(new_n10606_), .ZN(new_n10607_));
  AOI22_X1   g09605(.A1(new_n10601_), .A2(new_n8475_), .B1(new_n10598_), .B2(new_n10599_), .ZN(new_n10608_));
  NOR4_X1    g09606(.A1(new_n10596_), .A2(new_n10592_), .A3(new_n10595_), .A4(new_n8450_), .ZN(new_n10609_));
  NOR2_X1    g09607(.A1(new_n10608_), .A2(new_n10609_), .ZN(new_n10610_));
  NOR2_X1    g09608(.A1(new_n10607_), .A2(new_n10610_), .ZN(new_n10611_));
  OAI21_X1   g09609(.A1(new_n10611_), .A2(new_n10604_), .B(new_n10570_), .ZN(new_n10612_));
  AOI21_X1   g09610(.A1(new_n8495_), .A2(new_n8471_), .B(new_n8502_), .ZN(new_n10613_));
  NAND2_X1   g09611(.A1(new_n10607_), .A2(new_n10610_), .ZN(new_n10614_));
  NAND3_X1   g09612(.A1(new_n10603_), .A2(new_n10605_), .A3(new_n10606_), .ZN(new_n10615_));
  NAND3_X1   g09613(.A1(new_n10614_), .A2(new_n10615_), .A3(new_n10613_), .ZN(new_n10616_));
  NAND2_X1   g09614(.A1(new_n10612_), .A2(new_n10616_), .ZN(new_n10617_));
  NOR2_X1    g09615(.A1(new_n10569_), .A2(new_n10617_), .ZN(new_n10618_));
  OAI21_X1   g09616(.A1(new_n10567_), .A2(new_n10566_), .B(new_n10565_), .ZN(new_n10619_));
  NAND3_X1   g09617(.A1(new_n10556_), .A2(new_n10563_), .A3(new_n10524_), .ZN(new_n10620_));
  NAND2_X1   g09618(.A1(new_n10619_), .A2(new_n10620_), .ZN(new_n10621_));
  AOI21_X1   g09619(.A1(new_n10614_), .A2(new_n10615_), .B(new_n10613_), .ZN(new_n10622_));
  NOR3_X1    g09620(.A1(new_n10611_), .A2(new_n10604_), .A3(new_n10570_), .ZN(new_n10623_));
  NOR2_X1    g09621(.A1(new_n10623_), .A2(new_n10622_), .ZN(new_n10624_));
  NOR2_X1    g09622(.A1(new_n10621_), .A2(new_n10624_), .ZN(new_n10625_));
  OAI21_X1   g09623(.A1(new_n10625_), .A2(new_n10618_), .B(new_n10523_), .ZN(new_n10626_));
  NAND3_X1   g09624(.A1(new_n8506_), .A2(new_n8503_), .A3(new_n8507_), .ZN(new_n10627_));
  AOI21_X1   g09625(.A1(new_n8380_), .A2(new_n10627_), .B(new_n8508_), .ZN(new_n10628_));
  NAND2_X1   g09626(.A1(new_n10621_), .A2(new_n10624_), .ZN(new_n10629_));
  NAND3_X1   g09627(.A1(new_n10617_), .A2(new_n10619_), .A3(new_n10620_), .ZN(new_n10630_));
  NAND3_X1   g09628(.A1(new_n10629_), .A2(new_n10630_), .A3(new_n10628_), .ZN(new_n10631_));
  NAND2_X1   g09629(.A1(new_n10626_), .A2(new_n10631_), .ZN(new_n10632_));
  NOR2_X1    g09630(.A1(new_n10521_), .A2(new_n10632_), .ZN(new_n10633_));
  OAI21_X1   g09631(.A1(new_n10519_), .A2(new_n10518_), .B(new_n10517_), .ZN(new_n10634_));
  NAND3_X1   g09632(.A1(new_n10507_), .A2(new_n10514_), .A3(new_n10411_), .ZN(new_n10635_));
  NAND2_X1   g09633(.A1(new_n10634_), .A2(new_n10635_), .ZN(new_n10636_));
  AOI21_X1   g09634(.A1(new_n10629_), .A2(new_n10630_), .B(new_n10628_), .ZN(new_n10637_));
  NOR3_X1    g09635(.A1(new_n10625_), .A2(new_n10618_), .A3(new_n10523_), .ZN(new_n10638_));
  NOR2_X1    g09636(.A1(new_n10638_), .A2(new_n10637_), .ZN(new_n10639_));
  NOR2_X1    g09637(.A1(new_n10636_), .A2(new_n10639_), .ZN(new_n10640_));
  OAI21_X1   g09638(.A1(new_n10640_), .A2(new_n10633_), .B(new_n10409_), .ZN(new_n10641_));
  AOI22_X1   g09639(.A1(new_n8521_), .A2(new_n8252_), .B1(new_n8523_), .B2(new_n8522_), .ZN(new_n10642_));
  NAND2_X1   g09640(.A1(new_n10636_), .A2(new_n10639_), .ZN(new_n10643_));
  NAND3_X1   g09641(.A1(new_n10632_), .A2(new_n10634_), .A3(new_n10635_), .ZN(new_n10644_));
  NAND3_X1   g09642(.A1(new_n10643_), .A2(new_n10644_), .A3(new_n10642_), .ZN(new_n10645_));
  NAND2_X1   g09643(.A1(new_n10641_), .A2(new_n10645_), .ZN(new_n10646_));
  NOR2_X1    g09644(.A1(new_n10407_), .A2(new_n10646_), .ZN(new_n10647_));
  OAI21_X1   g09645(.A1(new_n10405_), .A2(new_n10404_), .B(new_n10403_), .ZN(new_n10648_));
  NAND3_X1   g09646(.A1(new_n10393_), .A2(new_n10400_), .A3(new_n10173_), .ZN(new_n10649_));
  NAND2_X1   g09647(.A1(new_n10648_), .A2(new_n10649_), .ZN(new_n10650_));
  AOI21_X1   g09648(.A1(new_n10643_), .A2(new_n10644_), .B(new_n10642_), .ZN(new_n10651_));
  NOR3_X1    g09649(.A1(new_n10640_), .A2(new_n10633_), .A3(new_n10409_), .ZN(new_n10652_));
  NOR2_X1    g09650(.A1(new_n10652_), .A2(new_n10651_), .ZN(new_n10653_));
  NOR2_X1    g09651(.A1(new_n10650_), .A2(new_n10653_), .ZN(new_n10654_));
  OAI21_X1   g09652(.A1(new_n10654_), .A2(new_n10647_), .B(new_n10172_), .ZN(new_n10655_));
  INV_X1     g09653(.I(new_n8538_), .ZN(new_n10656_));
  AOI21_X1   g09654(.A1(new_n7969_), .A2(new_n10656_), .B(new_n8539_), .ZN(new_n10657_));
  NAND2_X1   g09655(.A1(new_n10650_), .A2(new_n10653_), .ZN(new_n10658_));
  NAND3_X1   g09656(.A1(new_n10646_), .A2(new_n10648_), .A3(new_n10649_), .ZN(new_n10659_));
  NAND3_X1   g09657(.A1(new_n10658_), .A2(new_n10659_), .A3(new_n10657_), .ZN(new_n10660_));
  NAND2_X1   g09658(.A1(new_n10655_), .A2(new_n10660_), .ZN(new_n10661_));
  NOR2_X1    g09659(.A1(new_n10170_), .A2(new_n10661_), .ZN(new_n10662_));
  OAI21_X1   g09660(.A1(new_n10167_), .A2(new_n10168_), .B(new_n10166_), .ZN(new_n10663_));
  NAND3_X1   g09661(.A1(new_n10164_), .A2(new_n10157_), .A3(new_n9671_), .ZN(new_n10664_));
  NAND2_X1   g09662(.A1(new_n10663_), .A2(new_n10664_), .ZN(new_n10665_));
  AOI21_X1   g09663(.A1(new_n10658_), .A2(new_n10659_), .B(new_n10657_), .ZN(new_n10666_));
  NOR3_X1    g09664(.A1(new_n10654_), .A2(new_n10647_), .A3(new_n10172_), .ZN(new_n10667_));
  NOR2_X1    g09665(.A1(new_n10667_), .A2(new_n10666_), .ZN(new_n10668_));
  NOR2_X1    g09666(.A1(new_n10668_), .A2(new_n10665_), .ZN(new_n10669_));
  OAI21_X1   g09667(.A1(new_n10669_), .A2(new_n10662_), .B(new_n9669_), .ZN(new_n10670_));
  AOI21_X1   g09668(.A1(new_n8537_), .A2(new_n8540_), .B(new_n9666_), .ZN(new_n10671_));
  INV_X1     g09669(.I(new_n9665_), .ZN(new_n10672_));
  AOI21_X1   g09670(.A1(new_n10672_), .A2(new_n9667_), .B(new_n10671_), .ZN(new_n10673_));
  NAND2_X1   g09671(.A1(new_n10668_), .A2(new_n10665_), .ZN(new_n10674_));
  NAND3_X1   g09672(.A1(new_n10661_), .A2(new_n10663_), .A3(new_n10664_), .ZN(new_n10675_));
  NAND3_X1   g09673(.A1(new_n10674_), .A2(new_n10675_), .A3(new_n10673_), .ZN(new_n10676_));
  NAND3_X1   g09674(.A1(new_n10670_), .A2(new_n10676_), .A3(new_n4171_), .ZN(new_n10677_));
  XNOR2_X1   g09675(.A1(new_n7383_), .A2(new_n5752_), .ZN(new_n10678_));
  INV_X1     g09676(.I(new_n2344_), .ZN(new_n10679_));
  NOR3_X1    g09677(.A1(new_n2342_), .A2(new_n1523_), .A3(new_n2343_), .ZN(new_n10680_));
  AOI21_X1   g09678(.A1(new_n10679_), .A2(new_n1523_), .B(new_n10680_), .ZN(new_n10681_));
  NOR2_X1    g09679(.A1(new_n10678_), .A2(new_n10681_), .ZN(new_n10682_));
  NAND3_X1   g09680(.A1(new_n8537_), .A2(new_n7384_), .A3(new_n8540_), .ZN(new_n10683_));
  NAND2_X1   g09681(.A1(new_n8541_), .A2(new_n9666_), .ZN(new_n10684_));
  AOI21_X1   g09682(.A1(new_n10684_), .A2(new_n10683_), .B(new_n10672_), .ZN(new_n10685_));
  AOI21_X1   g09683(.A1(new_n8542_), .A2(new_n9667_), .B(new_n9665_), .ZN(new_n10686_));
  OAI21_X1   g09684(.A1(new_n10685_), .A2(new_n10686_), .B(new_n10682_), .ZN(new_n10687_));
  NOR3_X1    g09685(.A1(new_n4158_), .A2(new_n4163_), .A3(new_n2346_), .ZN(new_n10688_));
  NOR2_X1    g09686(.A1(new_n4164_), .A2(new_n2345_), .ZN(new_n10689_));
  OAI21_X1   g09687(.A1(new_n10689_), .A2(new_n10688_), .B(new_n4165_), .ZN(new_n10690_));
  OAI21_X1   g09688(.A1(new_n3032_), .A2(new_n4166_), .B(new_n3560_), .ZN(new_n10691_));
  NAND2_X1   g09689(.A1(new_n10690_), .A2(new_n10691_), .ZN(new_n10692_));
  INV_X1     g09690(.I(new_n10692_), .ZN(new_n10693_));
  NOR3_X1    g09691(.A1(new_n10685_), .A2(new_n10686_), .A3(new_n10682_), .ZN(new_n10694_));
  OAI21_X1   g09692(.A1(new_n10693_), .A2(new_n10694_), .B(new_n10687_), .ZN(new_n10695_));
  OR2_X2     g09693(.A1(new_n4156_), .A2(new_n4170_), .Z(new_n10696_));
  AOI21_X1   g09694(.A1(new_n10674_), .A2(new_n10675_), .B(new_n10673_), .ZN(new_n10697_));
  NOR3_X1    g09695(.A1(new_n10669_), .A2(new_n10662_), .A3(new_n9669_), .ZN(new_n10698_));
  OAI21_X1   g09696(.A1(new_n10698_), .A2(new_n10697_), .B(new_n10696_), .ZN(new_n10699_));
  NAND2_X1   g09697(.A1(new_n10699_), .A2(new_n10695_), .ZN(new_n10700_));
  NOR4_X1    g09698(.A1(new_n10165_), .A2(new_n10169_), .A3(new_n10667_), .A4(new_n10666_), .ZN(new_n10701_));
  OAI22_X1   g09699(.A1(new_n10165_), .A2(new_n10169_), .B1(new_n10667_), .B2(new_n10666_), .ZN(new_n10702_));
  AOI21_X1   g09700(.A1(new_n9669_), .A2(new_n10702_), .B(new_n10701_), .ZN(new_n10703_));
  NAND4_X1   g09701(.A1(new_n10648_), .A2(new_n10649_), .A3(new_n10641_), .A4(new_n10645_), .ZN(new_n10704_));
  AOI22_X1   g09702(.A1(new_n10648_), .A2(new_n10649_), .B1(new_n10641_), .B2(new_n10645_), .ZN(new_n10705_));
  OAI21_X1   g09703(.A1(new_n10657_), .A2(new_n10705_), .B(new_n10704_), .ZN(new_n10706_));
  NAND4_X1   g09704(.A1(new_n10634_), .A2(new_n10626_), .A3(new_n10635_), .A4(new_n10631_), .ZN(new_n10707_));
  OAI21_X1   g09705(.A1(new_n10521_), .A2(new_n10639_), .B(new_n10409_), .ZN(new_n10708_));
  NAND4_X1   g09706(.A1(new_n10619_), .A2(new_n10612_), .A3(new_n10620_), .A4(new_n10616_), .ZN(new_n10709_));
  INV_X1     g09707(.I(new_n10709_), .ZN(new_n10710_));
  AOI21_X1   g09708(.A1(new_n10621_), .A2(new_n10617_), .B(new_n10628_), .ZN(new_n10711_));
  OAI21_X1   g09709(.A1(new_n10553_), .A2(new_n8354_), .B(new_n10545_), .ZN(new_n10712_));
  OAI21_X1   g09710(.A1(new_n8352_), .A2(new_n8353_), .B(new_n10541_), .ZN(new_n10713_));
  OAI21_X1   g09711(.A1(new_n10553_), .A2(new_n10713_), .B(new_n10543_), .ZN(new_n10714_));
  NAND2_X1   g09712(.A1(new_n10714_), .A2(new_n10712_), .ZN(new_n10715_));
  NAND2_X1   g09713(.A1(new_n10538_), .A2(new_n8277_), .ZN(new_n10716_));
  AOI21_X1   g09714(.A1(new_n8276_), .A2(new_n8271_), .B(new_n10525_), .ZN(new_n10717_));
  NAND2_X1   g09715(.A1(new_n10717_), .A2(new_n10538_), .ZN(new_n10718_));
  AOI22_X1   g09716(.A1(new_n10718_), .A2(new_n10532_), .B1(new_n10716_), .B2(new_n10525_), .ZN(new_n10719_));
  NAND2_X1   g09717(.A1(new_n10719_), .A2(new_n10715_), .ZN(new_n10720_));
  AND2_X2    g09718(.A1(new_n10714_), .A2(new_n10712_), .Z(new_n10721_));
  NOR2_X1    g09719(.A1(new_n10534_), .A2(new_n8370_), .ZN(new_n10722_));
  OAI21_X1   g09720(.A1(new_n8368_), .A2(new_n8369_), .B(new_n10530_), .ZN(new_n10723_));
  NOR2_X1    g09721(.A1(new_n10534_), .A2(new_n10723_), .ZN(new_n10724_));
  OAI22_X1   g09722(.A1(new_n10724_), .A2(new_n10527_), .B1(new_n10722_), .B2(new_n10530_), .ZN(new_n10725_));
  NAND2_X1   g09723(.A1(new_n10721_), .A2(new_n10725_), .ZN(new_n10726_));
  NAND2_X1   g09724(.A1(new_n10726_), .A2(new_n10720_), .ZN(new_n10727_));
  AOI22_X1   g09725(.A1(new_n10535_), .A2(new_n10539_), .B1(new_n10560_), .B2(new_n10561_), .ZN(new_n10728_));
  INV_X1     g09726(.I(new_n10728_), .ZN(new_n10729_));
  NAND2_X1   g09727(.A1(new_n10729_), .A2(new_n10565_), .ZN(new_n10730_));
  NAND4_X1   g09728(.A1(new_n10535_), .A2(new_n10539_), .A3(new_n10560_), .A4(new_n10561_), .ZN(new_n10731_));
  OAI21_X1   g09729(.A1(new_n10524_), .A2(new_n10728_), .B(new_n10731_), .ZN(new_n10732_));
  NOR2_X1    g09730(.A1(new_n10721_), .A2(new_n10725_), .ZN(new_n10733_));
  NOR2_X1    g09731(.A1(new_n10719_), .A2(new_n10715_), .ZN(new_n10734_));
  NOR4_X1    g09732(.A1(new_n10557_), .A2(new_n10558_), .A3(new_n10550_), .A4(new_n10554_), .ZN(new_n10735_));
  NOR3_X1    g09733(.A1(new_n10733_), .A2(new_n10734_), .A3(new_n10735_), .ZN(new_n10736_));
  AOI22_X1   g09734(.A1(new_n10736_), .A2(new_n10730_), .B1(new_n10727_), .B2(new_n10732_), .ZN(new_n10737_));
  NAND2_X1   g09735(.A1(new_n10601_), .A2(new_n8475_), .ZN(new_n10738_));
  AOI21_X1   g09736(.A1(new_n8472_), .A2(new_n8474_), .B(new_n10587_), .ZN(new_n10739_));
  NAND2_X1   g09737(.A1(new_n10739_), .A2(new_n10601_), .ZN(new_n10740_));
  AOI22_X1   g09738(.A1(new_n10740_), .A2(new_n10594_), .B1(new_n10738_), .B2(new_n10587_), .ZN(new_n10741_));
  OAI21_X1   g09739(.A1(new_n10584_), .A2(new_n8492_), .B(new_n10575_), .ZN(new_n10742_));
  NAND2_X1   g09740(.A1(new_n8423_), .A2(new_n10571_), .ZN(new_n10743_));
  OAI21_X1   g09741(.A1(new_n10743_), .A2(new_n10584_), .B(new_n10573_), .ZN(new_n10744_));
  NAND2_X1   g09742(.A1(new_n10744_), .A2(new_n10742_), .ZN(new_n10745_));
  NOR2_X1    g09743(.A1(new_n10745_), .A2(new_n10741_), .ZN(new_n10746_));
  OAI21_X1   g09744(.A1(new_n10596_), .A2(new_n8450_), .B(new_n10587_), .ZN(new_n10747_));
  OAI21_X1   g09745(.A1(new_n8445_), .A2(new_n8449_), .B(new_n10593_), .ZN(new_n10748_));
  OAI21_X1   g09746(.A1(new_n10748_), .A2(new_n10596_), .B(new_n10594_), .ZN(new_n10749_));
  NAND2_X1   g09747(.A1(new_n10749_), .A2(new_n10747_), .ZN(new_n10750_));
  AOI21_X1   g09748(.A1(new_n10580_), .A2(new_n8423_), .B(new_n10571_), .ZN(new_n10751_));
  AOI21_X1   g09749(.A1(new_n8418_), .A2(new_n8422_), .B(new_n10575_), .ZN(new_n10752_));
  AOI21_X1   g09750(.A1(new_n10752_), .A2(new_n10580_), .B(new_n10577_), .ZN(new_n10753_));
  NOR2_X1    g09751(.A1(new_n10753_), .A2(new_n10751_), .ZN(new_n10754_));
  NOR2_X1    g09752(.A1(new_n10754_), .A2(new_n10750_), .ZN(new_n10755_));
  NOR2_X1    g09753(.A1(new_n10746_), .A2(new_n10755_), .ZN(new_n10756_));
  AOI22_X1   g09754(.A1(new_n10605_), .A2(new_n10606_), .B1(new_n10597_), .B2(new_n10602_), .ZN(new_n10757_));
  NOR2_X1    g09755(.A1(new_n10613_), .A2(new_n10757_), .ZN(new_n10758_));
  NAND2_X1   g09756(.A1(new_n10607_), .A2(new_n10603_), .ZN(new_n10759_));
  NOR4_X1    g09757(.A1(new_n10581_), .A2(new_n10585_), .A3(new_n10608_), .A4(new_n10609_), .ZN(new_n10760_));
  AOI21_X1   g09758(.A1(new_n10759_), .A2(new_n10570_), .B(new_n10760_), .ZN(new_n10761_));
  NAND2_X1   g09759(.A1(new_n10754_), .A2(new_n10750_), .ZN(new_n10762_));
  NAND2_X1   g09760(.A1(new_n10745_), .A2(new_n10741_), .ZN(new_n10763_));
  NAND4_X1   g09761(.A1(new_n10605_), .A2(new_n10597_), .A3(new_n10606_), .A4(new_n10602_), .ZN(new_n10764_));
  NAND3_X1   g09762(.A1(new_n10763_), .A2(new_n10762_), .A3(new_n10764_), .ZN(new_n10765_));
  OAI22_X1   g09763(.A1(new_n10756_), .A2(new_n10761_), .B1(new_n10765_), .B2(new_n10758_), .ZN(new_n10766_));
  NOR2_X1    g09764(.A1(new_n10737_), .A2(new_n10766_), .ZN(new_n10767_));
  NOR2_X1    g09765(.A1(new_n10733_), .A2(new_n10734_), .ZN(new_n10768_));
  NOR2_X1    g09766(.A1(new_n10524_), .A2(new_n10728_), .ZN(new_n10769_));
  AOI21_X1   g09767(.A1(new_n10729_), .A2(new_n10565_), .B(new_n10735_), .ZN(new_n10770_));
  NAND3_X1   g09768(.A1(new_n10726_), .A2(new_n10720_), .A3(new_n10731_), .ZN(new_n10771_));
  OAI22_X1   g09769(.A1(new_n10768_), .A2(new_n10770_), .B1(new_n10771_), .B2(new_n10769_), .ZN(new_n10772_));
  NAND2_X1   g09770(.A1(new_n10763_), .A2(new_n10762_), .ZN(new_n10773_));
  NAND2_X1   g09771(.A1(new_n10759_), .A2(new_n10570_), .ZN(new_n10774_));
  OAI21_X1   g09772(.A1(new_n10613_), .A2(new_n10757_), .B(new_n10764_), .ZN(new_n10775_));
  NOR3_X1    g09773(.A1(new_n10746_), .A2(new_n10755_), .A3(new_n10760_), .ZN(new_n10776_));
  AOI22_X1   g09774(.A1(new_n10776_), .A2(new_n10774_), .B1(new_n10773_), .B2(new_n10775_), .ZN(new_n10777_));
  NOR2_X1    g09775(.A1(new_n10772_), .A2(new_n10777_), .ZN(new_n10778_));
  OAI22_X1   g09776(.A1(new_n10778_), .A2(new_n10767_), .B1(new_n10711_), .B2(new_n10710_), .ZN(new_n10779_));
  OAI21_X1   g09777(.A1(new_n10569_), .A2(new_n10624_), .B(new_n10523_), .ZN(new_n10780_));
  NAND2_X1   g09778(.A1(new_n10772_), .A2(new_n10777_), .ZN(new_n10781_));
  NAND2_X1   g09779(.A1(new_n10737_), .A2(new_n10766_), .ZN(new_n10782_));
  NAND4_X1   g09780(.A1(new_n10780_), .A2(new_n10781_), .A3(new_n10782_), .A4(new_n10709_), .ZN(new_n10783_));
  NAND2_X1   g09781(.A1(new_n10779_), .A2(new_n10783_), .ZN(new_n10784_));
  NAND4_X1   g09782(.A1(new_n10454_), .A2(new_n10458_), .A3(new_n10511_), .A4(new_n10512_), .ZN(new_n10785_));
  OAI21_X1   g09783(.A1(new_n10510_), .A2(new_n10506_), .B(new_n10517_), .ZN(new_n10786_));
  NAND2_X1   g09784(.A1(new_n10486_), .A2(new_n8184_), .ZN(new_n10787_));
  NAND3_X1   g09785(.A1(new_n10486_), .A2(new_n8184_), .A3(new_n10477_), .ZN(new_n10788_));
  AOI22_X1   g09786(.A1(new_n10788_), .A2(new_n10481_), .B1(new_n10787_), .B2(new_n10483_), .ZN(new_n10789_));
  OAI21_X1   g09787(.A1(new_n10469_), .A2(new_n8225_), .B(new_n10461_), .ZN(new_n10790_));
  OAI21_X1   g09788(.A1(new_n8222_), .A2(new_n8224_), .B(new_n10465_), .ZN(new_n10791_));
  OAI21_X1   g09789(.A1(new_n10791_), .A2(new_n10469_), .B(new_n10467_), .ZN(new_n10792_));
  NAND2_X1   g09790(.A1(new_n10792_), .A2(new_n10790_), .ZN(new_n10793_));
  NOR2_X1    g09791(.A1(new_n10789_), .A2(new_n10793_), .ZN(new_n10794_));
  OAI21_X1   g09792(.A1(new_n10490_), .A2(new_n8209_), .B(new_n10483_), .ZN(new_n10795_));
  OAI21_X1   g09793(.A1(new_n8206_), .A2(new_n8208_), .B(new_n10477_), .ZN(new_n10796_));
  OAI21_X1   g09794(.A1(new_n10490_), .A2(new_n10796_), .B(new_n10481_), .ZN(new_n10797_));
  NAND2_X1   g09795(.A1(new_n10797_), .A2(new_n10795_), .ZN(new_n10798_));
  AOI21_X1   g09796(.A1(new_n10474_), .A2(new_n8156_), .B(new_n10465_), .ZN(new_n10799_));
  AOI21_X1   g09797(.A1(new_n8154_), .A2(new_n8155_), .B(new_n10461_), .ZN(new_n10800_));
  AOI21_X1   g09798(.A1(new_n10800_), .A2(new_n10474_), .B(new_n10463_), .ZN(new_n10801_));
  NOR2_X1    g09799(.A1(new_n10801_), .A2(new_n10799_), .ZN(new_n10802_));
  NOR2_X1    g09800(.A1(new_n10802_), .A2(new_n10798_), .ZN(new_n10803_));
  NOR2_X1    g09801(.A1(new_n10794_), .A2(new_n10803_), .ZN(new_n10804_));
  AOI22_X1   g09802(.A1(new_n10470_), .A2(new_n10475_), .B1(new_n10497_), .B2(new_n10498_), .ZN(new_n10805_));
  NOR2_X1    g09803(.A1(new_n10460_), .A2(new_n10805_), .ZN(new_n10806_));
  OAI22_X1   g09804(.A1(new_n10494_), .A2(new_n10495_), .B1(new_n10487_), .B2(new_n10491_), .ZN(new_n10807_));
  NOR4_X1    g09805(.A1(new_n10494_), .A2(new_n10495_), .A3(new_n10487_), .A4(new_n10491_), .ZN(new_n10808_));
  AOI21_X1   g09806(.A1(new_n10502_), .A2(new_n10807_), .B(new_n10808_), .ZN(new_n10809_));
  NAND2_X1   g09807(.A1(new_n10802_), .A2(new_n10798_), .ZN(new_n10810_));
  NAND2_X1   g09808(.A1(new_n10789_), .A2(new_n10793_), .ZN(new_n10811_));
  NAND4_X1   g09809(.A1(new_n10470_), .A2(new_n10475_), .A3(new_n10497_), .A4(new_n10498_), .ZN(new_n10812_));
  NAND3_X1   g09810(.A1(new_n10811_), .A2(new_n10810_), .A3(new_n10812_), .ZN(new_n10813_));
  OAI22_X1   g09811(.A1(new_n10806_), .A2(new_n10813_), .B1(new_n10804_), .B2(new_n10809_), .ZN(new_n10814_));
  OAI21_X1   g09812(.A1(new_n10438_), .A2(new_n8049_), .B(new_n10430_), .ZN(new_n10815_));
  OAI21_X1   g09813(.A1(new_n8044_), .A2(new_n8048_), .B(new_n10434_), .ZN(new_n10816_));
  OAI21_X1   g09814(.A1(new_n10438_), .A2(new_n10816_), .B(new_n10436_), .ZN(new_n10817_));
  NAND2_X1   g09815(.A1(new_n10817_), .A2(new_n10815_), .ZN(new_n10818_));
  AOI21_X1   g09816(.A1(new_n10423_), .A2(new_n8092_), .B(new_n10413_), .ZN(new_n10819_));
  AOI21_X1   g09817(.A1(new_n8089_), .A2(new_n8091_), .B(new_n10416_), .ZN(new_n10820_));
  AOI21_X1   g09818(.A1(new_n10820_), .A2(new_n10423_), .B(new_n10420_), .ZN(new_n10821_));
  NOR2_X1    g09819(.A1(new_n10821_), .A2(new_n10819_), .ZN(new_n10822_));
  NAND2_X1   g09820(.A1(new_n10822_), .A2(new_n10818_), .ZN(new_n10823_));
  NAND2_X1   g09821(.A1(new_n10443_), .A2(new_n8073_), .ZN(new_n10824_));
  NAND3_X1   g09822(.A1(new_n10443_), .A2(new_n8073_), .A3(new_n10434_), .ZN(new_n10825_));
  AOI22_X1   g09823(.A1(new_n10825_), .A2(new_n10436_), .B1(new_n10824_), .B2(new_n10430_), .ZN(new_n10826_));
  OAI21_X1   g09824(.A1(new_n10427_), .A2(new_n8005_), .B(new_n10416_), .ZN(new_n10827_));
  OAI21_X1   g09825(.A1(new_n8000_), .A2(new_n8004_), .B(new_n10413_), .ZN(new_n10828_));
  OAI21_X1   g09826(.A1(new_n10828_), .A2(new_n10427_), .B(new_n10414_), .ZN(new_n10829_));
  NAND2_X1   g09827(.A1(new_n10829_), .A2(new_n10827_), .ZN(new_n10830_));
  NAND2_X1   g09828(.A1(new_n10826_), .A2(new_n10830_), .ZN(new_n10831_));
  NAND2_X1   g09829(.A1(new_n10831_), .A2(new_n10823_), .ZN(new_n10832_));
  OAI22_X1   g09830(.A1(new_n10424_), .A2(new_n10428_), .B1(new_n10450_), .B2(new_n10451_), .ZN(new_n10833_));
  NAND2_X1   g09831(.A1(new_n10412_), .A2(new_n10833_), .ZN(new_n10834_));
  AOI22_X1   g09832(.A1(new_n10447_), .A2(new_n10448_), .B1(new_n10439_), .B2(new_n10444_), .ZN(new_n10835_));
  NAND4_X1   g09833(.A1(new_n10447_), .A2(new_n10439_), .A3(new_n10448_), .A4(new_n10444_), .ZN(new_n10836_));
  OAI21_X1   g09834(.A1(new_n10455_), .A2(new_n10835_), .B(new_n10836_), .ZN(new_n10837_));
  NOR2_X1    g09835(.A1(new_n10826_), .A2(new_n10830_), .ZN(new_n10838_));
  NOR2_X1    g09836(.A1(new_n10822_), .A2(new_n10818_), .ZN(new_n10839_));
  NOR4_X1    g09837(.A1(new_n10424_), .A2(new_n10428_), .A3(new_n10450_), .A4(new_n10451_), .ZN(new_n10840_));
  NOR3_X1    g09838(.A1(new_n10838_), .A2(new_n10839_), .A3(new_n10840_), .ZN(new_n10841_));
  AOI22_X1   g09839(.A1(new_n10841_), .A2(new_n10834_), .B1(new_n10837_), .B2(new_n10832_), .ZN(new_n10842_));
  NAND2_X1   g09840(.A1(new_n10842_), .A2(new_n10814_), .ZN(new_n10843_));
  NAND2_X1   g09841(.A1(new_n10811_), .A2(new_n10810_), .ZN(new_n10844_));
  NAND2_X1   g09842(.A1(new_n10502_), .A2(new_n10807_), .ZN(new_n10845_));
  OAI21_X1   g09843(.A1(new_n10460_), .A2(new_n10805_), .B(new_n10812_), .ZN(new_n10846_));
  NOR3_X1    g09844(.A1(new_n10794_), .A2(new_n10803_), .A3(new_n10808_), .ZN(new_n10847_));
  AOI22_X1   g09845(.A1(new_n10847_), .A2(new_n10845_), .B1(new_n10844_), .B2(new_n10846_), .ZN(new_n10848_));
  NOR2_X1    g09846(.A1(new_n10838_), .A2(new_n10839_), .ZN(new_n10849_));
  NOR2_X1    g09847(.A1(new_n10455_), .A2(new_n10835_), .ZN(new_n10850_));
  AOI21_X1   g09848(.A1(new_n10412_), .A2(new_n10833_), .B(new_n10840_), .ZN(new_n10851_));
  NAND3_X1   g09849(.A1(new_n10831_), .A2(new_n10823_), .A3(new_n10836_), .ZN(new_n10852_));
  OAI22_X1   g09850(.A1(new_n10850_), .A2(new_n10852_), .B1(new_n10849_), .B2(new_n10851_), .ZN(new_n10853_));
  NAND2_X1   g09851(.A1(new_n10853_), .A2(new_n10848_), .ZN(new_n10854_));
  AOI22_X1   g09852(.A1(new_n10843_), .A2(new_n10854_), .B1(new_n10786_), .B2(new_n10785_), .ZN(new_n10855_));
  NOR2_X1    g09853(.A1(new_n10459_), .A2(new_n10513_), .ZN(new_n10856_));
  AOI21_X1   g09854(.A1(new_n10459_), .A2(new_n10513_), .B(new_n10411_), .ZN(new_n10857_));
  NOR2_X1    g09855(.A1(new_n10853_), .A2(new_n10848_), .ZN(new_n10858_));
  NOR2_X1    g09856(.A1(new_n10842_), .A2(new_n10814_), .ZN(new_n10859_));
  NOR4_X1    g09857(.A1(new_n10858_), .A2(new_n10859_), .A3(new_n10857_), .A4(new_n10856_), .ZN(new_n10860_));
  NOR2_X1    g09858(.A1(new_n10855_), .A2(new_n10860_), .ZN(new_n10861_));
  NAND2_X1   g09859(.A1(new_n10784_), .A2(new_n10861_), .ZN(new_n10862_));
  AOI22_X1   g09860(.A1(new_n10781_), .A2(new_n10782_), .B1(new_n10780_), .B2(new_n10709_), .ZN(new_n10863_));
  AOI22_X1   g09861(.A1(new_n10619_), .A2(new_n10620_), .B1(new_n10612_), .B2(new_n10616_), .ZN(new_n10864_));
  OAI21_X1   g09862(.A1(new_n10864_), .A2(new_n10628_), .B(new_n10709_), .ZN(new_n10865_));
  NOR3_X1    g09863(.A1(new_n10865_), .A2(new_n10778_), .A3(new_n10767_), .ZN(new_n10866_));
  NOR2_X1    g09864(.A1(new_n10863_), .A2(new_n10866_), .ZN(new_n10867_));
  OAI22_X1   g09865(.A1(new_n10858_), .A2(new_n10859_), .B1(new_n10857_), .B2(new_n10856_), .ZN(new_n10868_));
  NAND4_X1   g09866(.A1(new_n10786_), .A2(new_n10843_), .A3(new_n10854_), .A4(new_n10785_), .ZN(new_n10869_));
  NAND2_X1   g09867(.A1(new_n10868_), .A2(new_n10869_), .ZN(new_n10870_));
  NAND2_X1   g09868(.A1(new_n10867_), .A2(new_n10870_), .ZN(new_n10871_));
  AOI22_X1   g09869(.A1(new_n10862_), .A2(new_n10871_), .B1(new_n10708_), .B2(new_n10707_), .ZN(new_n10872_));
  AOI22_X1   g09870(.A1(new_n10634_), .A2(new_n10635_), .B1(new_n10626_), .B2(new_n10631_), .ZN(new_n10873_));
  OAI21_X1   g09871(.A1(new_n10873_), .A2(new_n10642_), .B(new_n10707_), .ZN(new_n10874_));
  NOR2_X1    g09872(.A1(new_n10867_), .A2(new_n10870_), .ZN(new_n10875_));
  NOR2_X1    g09873(.A1(new_n10784_), .A2(new_n10861_), .ZN(new_n10876_));
  NOR3_X1    g09874(.A1(new_n10874_), .A2(new_n10876_), .A3(new_n10875_), .ZN(new_n10877_));
  NOR2_X1    g09875(.A1(new_n10872_), .A2(new_n10877_), .ZN(new_n10878_));
  NOR2_X1    g09876(.A1(new_n10282_), .A2(new_n10399_), .ZN(new_n10879_));
  AOI21_X1   g09877(.A1(new_n10282_), .A2(new_n10399_), .B(new_n10173_), .ZN(new_n10880_));
  NAND4_X1   g09878(.A1(new_n10324_), .A2(new_n10328_), .A3(new_n10382_), .A4(new_n10383_), .ZN(new_n10881_));
  OAI21_X1   g09879(.A1(new_n10381_), .A2(new_n10377_), .B(new_n10388_), .ZN(new_n10882_));
  NAND2_X1   g09880(.A1(new_n10313_), .A2(new_n7756_), .ZN(new_n10883_));
  NAND3_X1   g09881(.A1(new_n10313_), .A2(new_n7756_), .A3(new_n10305_), .ZN(new_n10884_));
  AOI22_X1   g09882(.A1(new_n10884_), .A2(new_n10307_), .B1(new_n10883_), .B2(new_n10301_), .ZN(new_n10885_));
  NOR2_X1    g09883(.A1(new_n10298_), .A2(new_n7798_), .ZN(new_n10886_));
  NOR3_X1    g09884(.A1(new_n10298_), .A2(new_n7798_), .A3(new_n10290_), .ZN(new_n10887_));
  OAI22_X1   g09885(.A1(new_n10887_), .A2(new_n10292_), .B1(new_n10886_), .B2(new_n10286_), .ZN(new_n10888_));
  NOR2_X1    g09886(.A1(new_n10888_), .A2(new_n10885_), .ZN(new_n10889_));
  OAI21_X1   g09887(.A1(new_n10309_), .A2(new_n7782_), .B(new_n10301_), .ZN(new_n10890_));
  OAI21_X1   g09888(.A1(new_n7779_), .A2(new_n7781_), .B(new_n10305_), .ZN(new_n10891_));
  OAI21_X1   g09889(.A1(new_n10891_), .A2(new_n10309_), .B(new_n10307_), .ZN(new_n10892_));
  NAND2_X1   g09890(.A1(new_n10892_), .A2(new_n10890_), .ZN(new_n10893_));
  AOI21_X1   g09891(.A1(new_n10294_), .A2(new_n7707_), .B(new_n10286_), .ZN(new_n10894_));
  AOI21_X1   g09892(.A1(new_n7701_), .A2(new_n7706_), .B(new_n10290_), .ZN(new_n10895_));
  AOI21_X1   g09893(.A1(new_n10895_), .A2(new_n10294_), .B(new_n10292_), .ZN(new_n10896_));
  NOR2_X1    g09894(.A1(new_n10896_), .A2(new_n10894_), .ZN(new_n10897_));
  NOR2_X1    g09895(.A1(new_n10897_), .A2(new_n10893_), .ZN(new_n10898_));
  NOR2_X1    g09896(.A1(new_n10889_), .A2(new_n10898_), .ZN(new_n10899_));
  AOI22_X1   g09897(.A1(new_n10317_), .A2(new_n10318_), .B1(new_n10310_), .B2(new_n10314_), .ZN(new_n10900_));
  NOR2_X1    g09898(.A1(new_n10325_), .A2(new_n10900_), .ZN(new_n10901_));
  OAI22_X1   g09899(.A1(new_n10295_), .A2(new_n10299_), .B1(new_n10320_), .B2(new_n10321_), .ZN(new_n10902_));
  NOR4_X1    g09900(.A1(new_n10295_), .A2(new_n10320_), .A3(new_n10299_), .A4(new_n10321_), .ZN(new_n10903_));
  AOI21_X1   g09901(.A1(new_n10285_), .A2(new_n10902_), .B(new_n10903_), .ZN(new_n10904_));
  NAND2_X1   g09902(.A1(new_n10897_), .A2(new_n10893_), .ZN(new_n10905_));
  NAND2_X1   g09903(.A1(new_n10888_), .A2(new_n10885_), .ZN(new_n10906_));
  NAND4_X1   g09904(.A1(new_n10317_), .A2(new_n10310_), .A3(new_n10318_), .A4(new_n10314_), .ZN(new_n10907_));
  NAND3_X1   g09905(.A1(new_n10906_), .A2(new_n10905_), .A3(new_n10907_), .ZN(new_n10908_));
  OAI22_X1   g09906(.A1(new_n10901_), .A2(new_n10908_), .B1(new_n10899_), .B2(new_n10904_), .ZN(new_n10909_));
  OAI21_X1   g09907(.A1(new_n10360_), .A2(new_n7885_), .B(new_n10353_), .ZN(new_n10910_));
  OAI21_X1   g09908(.A1(new_n7880_), .A2(new_n7884_), .B(new_n10347_), .ZN(new_n10911_));
  OAI21_X1   g09909(.A1(new_n10911_), .A2(new_n10360_), .B(new_n10351_), .ZN(new_n10912_));
  NAND2_X1   g09910(.A1(new_n10912_), .A2(new_n10910_), .ZN(new_n10913_));
  AOI21_X1   g09911(.A1(new_n10344_), .A2(new_n7857_), .B(new_n10335_), .ZN(new_n10914_));
  AOI21_X1   g09912(.A1(new_n7854_), .A2(new_n7856_), .B(new_n10331_), .ZN(new_n10915_));
  AOI21_X1   g09913(.A1(new_n10915_), .A2(new_n10344_), .B(new_n10333_), .ZN(new_n10916_));
  NOR2_X1    g09914(.A1(new_n10916_), .A2(new_n10914_), .ZN(new_n10917_));
  NAND2_X1   g09915(.A1(new_n10917_), .A2(new_n10913_), .ZN(new_n10918_));
  NAND2_X1   g09916(.A1(new_n10356_), .A2(new_n7908_), .ZN(new_n10919_));
  NAND3_X1   g09917(.A1(new_n10356_), .A2(new_n7908_), .A3(new_n10347_), .ZN(new_n10920_));
  AOI22_X1   g09918(.A1(new_n10920_), .A2(new_n10351_), .B1(new_n10919_), .B2(new_n10353_), .ZN(new_n10921_));
  OAI21_X1   g09919(.A1(new_n10340_), .A2(new_n7925_), .B(new_n10331_), .ZN(new_n10922_));
  OAI21_X1   g09920(.A1(new_n7922_), .A2(new_n7924_), .B(new_n10335_), .ZN(new_n10923_));
  OAI21_X1   g09921(.A1(new_n10340_), .A2(new_n10923_), .B(new_n10337_), .ZN(new_n10924_));
  NAND2_X1   g09922(.A1(new_n10924_), .A2(new_n10922_), .ZN(new_n10925_));
  NAND2_X1   g09923(.A1(new_n10921_), .A2(new_n10925_), .ZN(new_n10926_));
  NAND2_X1   g09924(.A1(new_n10926_), .A2(new_n10918_), .ZN(new_n10927_));
  OAI22_X1   g09925(.A1(new_n10364_), .A2(new_n10366_), .B1(new_n10357_), .B2(new_n10361_), .ZN(new_n10928_));
  NAND2_X1   g09926(.A1(new_n10373_), .A2(new_n10928_), .ZN(new_n10929_));
  AOI22_X1   g09927(.A1(new_n10341_), .A2(new_n10345_), .B1(new_n10368_), .B2(new_n10369_), .ZN(new_n10930_));
  NAND4_X1   g09928(.A1(new_n10341_), .A2(new_n10368_), .A3(new_n10345_), .A4(new_n10369_), .ZN(new_n10931_));
  OAI21_X1   g09929(.A1(new_n10330_), .A2(new_n10930_), .B(new_n10931_), .ZN(new_n10932_));
  NOR2_X1    g09930(.A1(new_n10921_), .A2(new_n10925_), .ZN(new_n10933_));
  NOR2_X1    g09931(.A1(new_n10917_), .A2(new_n10913_), .ZN(new_n10934_));
  NOR4_X1    g09932(.A1(new_n10364_), .A2(new_n10366_), .A3(new_n10357_), .A4(new_n10361_), .ZN(new_n10935_));
  NOR3_X1    g09933(.A1(new_n10933_), .A2(new_n10934_), .A3(new_n10935_), .ZN(new_n10936_));
  AOI22_X1   g09934(.A1(new_n10936_), .A2(new_n10929_), .B1(new_n10927_), .B2(new_n10932_), .ZN(new_n10937_));
  NAND2_X1   g09935(.A1(new_n10909_), .A2(new_n10937_), .ZN(new_n10938_));
  NAND2_X1   g09936(.A1(new_n10906_), .A2(new_n10905_), .ZN(new_n10939_));
  NAND2_X1   g09937(.A1(new_n10285_), .A2(new_n10902_), .ZN(new_n10940_));
  OAI21_X1   g09938(.A1(new_n10325_), .A2(new_n10900_), .B(new_n10907_), .ZN(new_n10941_));
  NOR3_X1    g09939(.A1(new_n10889_), .A2(new_n10898_), .A3(new_n10903_), .ZN(new_n10942_));
  AOI22_X1   g09940(.A1(new_n10942_), .A2(new_n10940_), .B1(new_n10941_), .B2(new_n10939_), .ZN(new_n10943_));
  NOR2_X1    g09941(.A1(new_n10933_), .A2(new_n10934_), .ZN(new_n10944_));
  NOR2_X1    g09942(.A1(new_n10330_), .A2(new_n10930_), .ZN(new_n10945_));
  AOI21_X1   g09943(.A1(new_n10373_), .A2(new_n10928_), .B(new_n10935_), .ZN(new_n10946_));
  NAND3_X1   g09944(.A1(new_n10926_), .A2(new_n10918_), .A3(new_n10931_), .ZN(new_n10947_));
  OAI22_X1   g09945(.A1(new_n10945_), .A2(new_n10947_), .B1(new_n10944_), .B2(new_n10946_), .ZN(new_n10948_));
  NAND2_X1   g09946(.A1(new_n10943_), .A2(new_n10948_), .ZN(new_n10949_));
  AOI22_X1   g09947(.A1(new_n10938_), .A2(new_n10949_), .B1(new_n10882_), .B2(new_n10881_), .ZN(new_n10950_));
  AOI22_X1   g09948(.A1(new_n10328_), .A2(new_n10324_), .B1(new_n10382_), .B2(new_n10383_), .ZN(new_n10951_));
  OAI21_X1   g09949(.A1(new_n10284_), .A2(new_n10951_), .B(new_n10881_), .ZN(new_n10952_));
  NOR2_X1    g09950(.A1(new_n10943_), .A2(new_n10948_), .ZN(new_n10953_));
  NOR2_X1    g09951(.A1(new_n10909_), .A2(new_n10937_), .ZN(new_n10954_));
  NOR3_X1    g09952(.A1(new_n10952_), .A2(new_n10953_), .A3(new_n10954_), .ZN(new_n10955_));
  NOR2_X1    g09953(.A1(new_n10955_), .A2(new_n10950_), .ZN(new_n10956_));
  NOR2_X1    g09954(.A1(new_n10267_), .A2(new_n10271_), .ZN(new_n10957_));
  AOI22_X1   g09955(.A1(new_n10262_), .A2(new_n10266_), .B1(new_n10270_), .B2(new_n10269_), .ZN(new_n10958_));
  NOR2_X1    g09956(.A1(new_n10958_), .A2(new_n10278_), .ZN(new_n10959_));
  OAI21_X1   g09957(.A1(new_n10246_), .A2(new_n7631_), .B(new_n10238_), .ZN(new_n10960_));
  OAI21_X1   g09958(.A1(new_n7628_), .A2(new_n7630_), .B(new_n10242_), .ZN(new_n10961_));
  OAI21_X1   g09959(.A1(new_n10961_), .A2(new_n10246_), .B(new_n10244_), .ZN(new_n10962_));
  NAND2_X1   g09960(.A1(new_n10962_), .A2(new_n10960_), .ZN(new_n10963_));
  AOI21_X1   g09961(.A1(new_n10231_), .A2(new_n7560_), .B(new_n10225_), .ZN(new_n10964_));
  AOI21_X1   g09962(.A1(new_n7554_), .A2(new_n7559_), .B(new_n10228_), .ZN(new_n10965_));
  AOI21_X1   g09963(.A1(new_n10231_), .A2(new_n10965_), .B(new_n10229_), .ZN(new_n10966_));
  NOR2_X1    g09964(.A1(new_n10966_), .A2(new_n10964_), .ZN(new_n10967_));
  NAND2_X1   g09965(.A1(new_n10967_), .A2(new_n10963_), .ZN(new_n10968_));
  NAND2_X1   g09966(.A1(new_n10251_), .A2(new_n7606_), .ZN(new_n10969_));
  NAND3_X1   g09967(.A1(new_n10251_), .A2(new_n7606_), .A3(new_n10242_), .ZN(new_n10970_));
  AOI22_X1   g09968(.A1(new_n10970_), .A2(new_n10244_), .B1(new_n10969_), .B2(new_n10238_), .ZN(new_n10971_));
  OAI21_X1   g09969(.A1(new_n10235_), .A2(new_n7642_), .B(new_n10228_), .ZN(new_n10972_));
  NAND2_X1   g09970(.A1(new_n7560_), .A2(new_n10225_), .ZN(new_n10973_));
  OAI21_X1   g09971(.A1(new_n10973_), .A2(new_n10235_), .B(new_n10226_), .ZN(new_n10974_));
  NAND2_X1   g09972(.A1(new_n10974_), .A2(new_n10972_), .ZN(new_n10975_));
  NAND2_X1   g09973(.A1(new_n10975_), .A2(new_n10971_), .ZN(new_n10976_));
  NAND2_X1   g09974(.A1(new_n10976_), .A2(new_n10968_), .ZN(new_n10977_));
  OAI22_X1   g09975(.A1(new_n10232_), .A2(new_n10236_), .B1(new_n10258_), .B2(new_n10259_), .ZN(new_n10978_));
  NAND2_X1   g09976(.A1(new_n10224_), .A2(new_n10978_), .ZN(new_n10979_));
  AOI22_X1   g09977(.A1(new_n10256_), .A2(new_n10255_), .B1(new_n10247_), .B2(new_n10252_), .ZN(new_n10980_));
  NAND4_X1   g09978(.A1(new_n10255_), .A2(new_n10256_), .A3(new_n10247_), .A4(new_n10252_), .ZN(new_n10981_));
  OAI21_X1   g09979(.A1(new_n10263_), .A2(new_n10980_), .B(new_n10981_), .ZN(new_n10982_));
  NOR2_X1    g09980(.A1(new_n10975_), .A2(new_n10971_), .ZN(new_n10983_));
  NOR2_X1    g09981(.A1(new_n10967_), .A2(new_n10963_), .ZN(new_n10984_));
  NOR4_X1    g09982(.A1(new_n10232_), .A2(new_n10236_), .A3(new_n10258_), .A4(new_n10259_), .ZN(new_n10985_));
  NOR3_X1    g09983(.A1(new_n10983_), .A2(new_n10984_), .A3(new_n10985_), .ZN(new_n10986_));
  AOI22_X1   g09984(.A1(new_n10986_), .A2(new_n10979_), .B1(new_n10977_), .B2(new_n10982_), .ZN(new_n10987_));
  AOI21_X1   g09985(.A1(new_n10200_), .A2(new_n7504_), .B(new_n10192_), .ZN(new_n10988_));
  AOI21_X1   g09986(.A1(new_n7501_), .A2(new_n7503_), .B(new_n10196_), .ZN(new_n10989_));
  AOI21_X1   g09987(.A1(new_n10989_), .A2(new_n10200_), .B(new_n10198_), .ZN(new_n10990_));
  NOR2_X1    g09988(.A1(new_n10990_), .A2(new_n10988_), .ZN(new_n10991_));
  OAI21_X1   g09989(.A1(new_n10185_), .A2(new_n7420_), .B(new_n10177_), .ZN(new_n10992_));
  OAI21_X1   g09990(.A1(new_n7414_), .A2(new_n7419_), .B(new_n10181_), .ZN(new_n10993_));
  OAI21_X1   g09991(.A1(new_n10185_), .A2(new_n10993_), .B(new_n10183_), .ZN(new_n10994_));
  NAND2_X1   g09992(.A1(new_n10994_), .A2(new_n10992_), .ZN(new_n10995_));
  NOR2_X1    g09993(.A1(new_n10995_), .A2(new_n10991_), .ZN(new_n10996_));
  OAI21_X1   g09994(.A1(new_n10204_), .A2(new_n7477_), .B(new_n10196_), .ZN(new_n10997_));
  OAI21_X1   g09995(.A1(new_n7469_), .A2(new_n7476_), .B(new_n10192_), .ZN(new_n10998_));
  OAI21_X1   g09996(.A1(new_n10204_), .A2(new_n10998_), .B(new_n10194_), .ZN(new_n10999_));
  NAND2_X1   g09997(.A1(new_n10999_), .A2(new_n10997_), .ZN(new_n11000_));
  AOI21_X1   g09998(.A1(new_n10189_), .A2(new_n7517_), .B(new_n10181_), .ZN(new_n11001_));
  AOI21_X1   g09999(.A1(new_n7515_), .A2(new_n7516_), .B(new_n10177_), .ZN(new_n11002_));
  AOI21_X1   g10000(.A1(new_n11002_), .A2(new_n10189_), .B(new_n10179_), .ZN(new_n11003_));
  NOR2_X1    g10001(.A1(new_n11003_), .A2(new_n11001_), .ZN(new_n11004_));
  NOR2_X1    g10002(.A1(new_n11004_), .A2(new_n11000_), .ZN(new_n11005_));
  NOR2_X1    g10003(.A1(new_n10996_), .A2(new_n11005_), .ZN(new_n11006_));
  AOI22_X1   g10004(.A1(new_n10186_), .A2(new_n10190_), .B1(new_n10214_), .B2(new_n10215_), .ZN(new_n11007_));
  NOR2_X1    g10005(.A1(new_n10176_), .A2(new_n11007_), .ZN(new_n11008_));
  OAI22_X1   g10006(.A1(new_n10209_), .A2(new_n10211_), .B1(new_n10201_), .B2(new_n10206_), .ZN(new_n11009_));
  NOR4_X1    g10007(.A1(new_n10209_), .A2(new_n10201_), .A3(new_n10211_), .A4(new_n10206_), .ZN(new_n11010_));
  AOI21_X1   g10008(.A1(new_n10219_), .A2(new_n11009_), .B(new_n11010_), .ZN(new_n11011_));
  NAND2_X1   g10009(.A1(new_n11004_), .A2(new_n11000_), .ZN(new_n11012_));
  NAND2_X1   g10010(.A1(new_n10995_), .A2(new_n10991_), .ZN(new_n11013_));
  NAND4_X1   g10011(.A1(new_n10186_), .A2(new_n10214_), .A3(new_n10190_), .A4(new_n10215_), .ZN(new_n11014_));
  NAND3_X1   g10012(.A1(new_n11013_), .A2(new_n11012_), .A3(new_n11014_), .ZN(new_n11015_));
  OAI22_X1   g10013(.A1(new_n11008_), .A2(new_n11015_), .B1(new_n11006_), .B2(new_n11011_), .ZN(new_n11016_));
  NOR2_X1    g10014(.A1(new_n10987_), .A2(new_n11016_), .ZN(new_n11017_));
  NOR2_X1    g10015(.A1(new_n10983_), .A2(new_n10984_), .ZN(new_n11018_));
  NOR2_X1    g10016(.A1(new_n10263_), .A2(new_n10980_), .ZN(new_n11019_));
  AOI21_X1   g10017(.A1(new_n10224_), .A2(new_n10978_), .B(new_n10985_), .ZN(new_n11020_));
  NAND3_X1   g10018(.A1(new_n10976_), .A2(new_n10968_), .A3(new_n10981_), .ZN(new_n11021_));
  OAI22_X1   g10019(.A1(new_n11019_), .A2(new_n11021_), .B1(new_n11018_), .B2(new_n11020_), .ZN(new_n11022_));
  NAND2_X1   g10020(.A1(new_n11013_), .A2(new_n11012_), .ZN(new_n11023_));
  NAND2_X1   g10021(.A1(new_n10219_), .A2(new_n11009_), .ZN(new_n11024_));
  OAI21_X1   g10022(.A1(new_n10176_), .A2(new_n11007_), .B(new_n11014_), .ZN(new_n11025_));
  NOR3_X1    g10023(.A1(new_n10996_), .A2(new_n11005_), .A3(new_n11010_), .ZN(new_n11026_));
  AOI22_X1   g10024(.A1(new_n11024_), .A2(new_n11026_), .B1(new_n11025_), .B2(new_n11023_), .ZN(new_n11027_));
  NOR2_X1    g10025(.A1(new_n11022_), .A2(new_n11027_), .ZN(new_n11028_));
  OAI22_X1   g10026(.A1(new_n10959_), .A2(new_n10957_), .B1(new_n11028_), .B2(new_n11017_), .ZN(new_n11029_));
  NAND4_X1   g10027(.A1(new_n10270_), .A2(new_n10262_), .A3(new_n10266_), .A4(new_n10269_), .ZN(new_n11030_));
  OAI21_X1   g10028(.A1(new_n10274_), .A2(new_n10223_), .B(new_n10175_), .ZN(new_n11031_));
  NAND2_X1   g10029(.A1(new_n11022_), .A2(new_n11027_), .ZN(new_n11032_));
  NAND2_X1   g10030(.A1(new_n10987_), .A2(new_n11016_), .ZN(new_n11033_));
  NAND4_X1   g10031(.A1(new_n11031_), .A2(new_n11032_), .A3(new_n11033_), .A4(new_n11030_), .ZN(new_n11034_));
  NAND2_X1   g10032(.A1(new_n11029_), .A2(new_n11034_), .ZN(new_n11035_));
  NOR2_X1    g10033(.A1(new_n10956_), .A2(new_n11035_), .ZN(new_n11036_));
  INV_X1     g10034(.I(new_n10881_), .ZN(new_n11037_));
  AOI21_X1   g10035(.A1(new_n10329_), .A2(new_n10384_), .B(new_n10284_), .ZN(new_n11038_));
  OAI22_X1   g10036(.A1(new_n10953_), .A2(new_n10954_), .B1(new_n11038_), .B2(new_n11037_), .ZN(new_n11039_));
  NAND4_X1   g10037(.A1(new_n10949_), .A2(new_n10882_), .A3(new_n10938_), .A4(new_n10881_), .ZN(new_n11040_));
  NAND2_X1   g10038(.A1(new_n11039_), .A2(new_n11040_), .ZN(new_n11041_));
  AOI22_X1   g10039(.A1(new_n11032_), .A2(new_n11033_), .B1(new_n11031_), .B2(new_n11030_), .ZN(new_n11042_));
  NOR4_X1    g10040(.A1(new_n10959_), .A2(new_n11028_), .A3(new_n11017_), .A4(new_n10957_), .ZN(new_n11043_));
  NOR2_X1    g10041(.A1(new_n11042_), .A2(new_n11043_), .ZN(new_n11044_));
  NOR2_X1    g10042(.A1(new_n11044_), .A2(new_n11041_), .ZN(new_n11045_));
  OAI22_X1   g10043(.A1(new_n11036_), .A2(new_n11045_), .B1(new_n10879_), .B2(new_n10880_), .ZN(new_n11046_));
  NAND4_X1   g10044(.A1(new_n10276_), .A2(new_n10281_), .A3(new_n10397_), .A4(new_n10398_), .ZN(new_n11047_));
  OAI21_X1   g10045(.A1(new_n10396_), .A2(new_n10392_), .B(new_n10403_), .ZN(new_n11048_));
  NAND2_X1   g10046(.A1(new_n11044_), .A2(new_n11041_), .ZN(new_n11049_));
  NAND2_X1   g10047(.A1(new_n10956_), .A2(new_n11035_), .ZN(new_n11050_));
  NAND4_X1   g10048(.A1(new_n11050_), .A2(new_n11049_), .A3(new_n11048_), .A4(new_n11047_), .ZN(new_n11051_));
  NAND2_X1   g10049(.A1(new_n11046_), .A2(new_n11051_), .ZN(new_n11052_));
  NOR2_X1    g10050(.A1(new_n10878_), .A2(new_n11052_), .ZN(new_n11053_));
  OAI21_X1   g10051(.A1(new_n10875_), .A2(new_n10876_), .B(new_n10874_), .ZN(new_n11054_));
  NAND4_X1   g10052(.A1(new_n10862_), .A2(new_n10871_), .A3(new_n10708_), .A4(new_n10707_), .ZN(new_n11055_));
  NAND2_X1   g10053(.A1(new_n11054_), .A2(new_n11055_), .ZN(new_n11056_));
  AOI22_X1   g10054(.A1(new_n11050_), .A2(new_n11049_), .B1(new_n11048_), .B2(new_n11047_), .ZN(new_n11057_));
  AOI22_X1   g10055(.A1(new_n10276_), .A2(new_n10281_), .B1(new_n10397_), .B2(new_n10398_), .ZN(new_n11058_));
  OAI21_X1   g10056(.A1(new_n10173_), .A2(new_n11058_), .B(new_n11047_), .ZN(new_n11059_));
  NOR3_X1    g10057(.A1(new_n11059_), .A2(new_n11036_), .A3(new_n11045_), .ZN(new_n11060_));
  NOR2_X1    g10058(.A1(new_n11057_), .A2(new_n11060_), .ZN(new_n11061_));
  NOR2_X1    g10059(.A1(new_n11061_), .A2(new_n11056_), .ZN(new_n11062_));
  OAI21_X1   g10060(.A1(new_n11053_), .A2(new_n11062_), .B(new_n10706_), .ZN(new_n11063_));
  NOR4_X1    g10061(.A1(new_n10401_), .A2(new_n10406_), .A3(new_n10652_), .A4(new_n10651_), .ZN(new_n11064_));
  OAI22_X1   g10062(.A1(new_n10401_), .A2(new_n10406_), .B1(new_n10652_), .B2(new_n10651_), .ZN(new_n11065_));
  AOI21_X1   g10063(.A1(new_n10172_), .A2(new_n11065_), .B(new_n11064_), .ZN(new_n11066_));
  NAND2_X1   g10064(.A1(new_n11061_), .A2(new_n11056_), .ZN(new_n11067_));
  NAND2_X1   g10065(.A1(new_n10878_), .A2(new_n11052_), .ZN(new_n11068_));
  NAND3_X1   g10066(.A1(new_n11066_), .A2(new_n11067_), .A3(new_n11068_), .ZN(new_n11069_));
  NAND2_X1   g10067(.A1(new_n11063_), .A2(new_n11069_), .ZN(new_n11070_));
  NOR4_X1    g10068(.A1(new_n10158_), .A2(new_n10150_), .A3(new_n10155_), .A4(new_n10159_), .ZN(new_n11071_));
  OAI22_X1   g10069(.A1(new_n10150_), .A2(new_n10155_), .B1(new_n10158_), .B2(new_n10159_), .ZN(new_n11072_));
  AOI21_X1   g10070(.A1(new_n10166_), .A2(new_n11072_), .B(new_n11071_), .ZN(new_n11073_));
  NAND4_X1   g10071(.A1(new_n10023_), .A2(new_n10027_), .A3(new_n10146_), .A4(new_n10147_), .ZN(new_n11074_));
  AOI22_X1   g10072(.A1(new_n10023_), .A2(new_n10027_), .B1(new_n10146_), .B2(new_n10147_), .ZN(new_n11075_));
  OAI21_X1   g10073(.A1(new_n9915_), .A2(new_n11075_), .B(new_n11074_), .ZN(new_n11076_));
  NAND4_X1   g10074(.A1(new_n10074_), .A2(new_n10079_), .A3(new_n10132_), .A4(new_n10133_), .ZN(new_n11077_));
  OAI22_X1   g10075(.A1(new_n10130_), .A2(new_n10129_), .B1(new_n10122_), .B2(new_n10126_), .ZN(new_n11078_));
  NAND2_X1   g10076(.A1(new_n10137_), .A2(new_n11078_), .ZN(new_n11079_));
  NAND2_X1   g10077(.A1(new_n10065_), .A2(new_n9479_), .ZN(new_n11080_));
  NAND3_X1   g10078(.A1(new_n10065_), .A2(new_n9479_), .A3(new_n10057_), .ZN(new_n11081_));
  AOI22_X1   g10079(.A1(new_n11081_), .A2(new_n10059_), .B1(new_n11080_), .B2(new_n10052_), .ZN(new_n11082_));
  OAI21_X1   g10080(.A1(new_n10046_), .A2(new_n9405_), .B(new_n10040_), .ZN(new_n11083_));
  OAI21_X1   g10081(.A1(new_n9404_), .A2(new_n9400_), .B(new_n10043_), .ZN(new_n11084_));
  OAI21_X1   g10082(.A1(new_n10046_), .A2(new_n11084_), .B(new_n10044_), .ZN(new_n11085_));
  NAND2_X1   g10083(.A1(new_n11085_), .A2(new_n11083_), .ZN(new_n11086_));
  NOR2_X1    g10084(.A1(new_n11082_), .A2(new_n11086_), .ZN(new_n11087_));
  OAI21_X1   g10085(.A1(new_n10061_), .A2(new_n9449_), .B(new_n10052_), .ZN(new_n11088_));
  OAI21_X1   g10086(.A1(new_n9444_), .A2(new_n9448_), .B(new_n10057_), .ZN(new_n11089_));
  OAI21_X1   g10087(.A1(new_n11089_), .A2(new_n10061_), .B(new_n10059_), .ZN(new_n11090_));
  NAND2_X1   g10088(.A1(new_n11090_), .A2(new_n11088_), .ZN(new_n11091_));
  AOI21_X1   g10089(.A1(new_n10050_), .A2(new_n10033_), .B(new_n10043_), .ZN(new_n11092_));
  AOI21_X1   g10090(.A1(new_n10031_), .A2(new_n10032_), .B(new_n10040_), .ZN(new_n11093_));
  AOI21_X1   g10091(.A1(new_n11093_), .A2(new_n10050_), .B(new_n10041_), .ZN(new_n11094_));
  NOR2_X1    g10092(.A1(new_n11094_), .A2(new_n11092_), .ZN(new_n11095_));
  NOR2_X1    g10093(.A1(new_n11095_), .A2(new_n11091_), .ZN(new_n11096_));
  NOR2_X1    g10094(.A1(new_n11087_), .A2(new_n11096_), .ZN(new_n11097_));
  AOI22_X1   g10095(.A1(new_n10047_), .A2(new_n10051_), .B1(new_n10062_), .B2(new_n10066_), .ZN(new_n11098_));
  NOR2_X1    g10096(.A1(new_n10076_), .A2(new_n11098_), .ZN(new_n11099_));
  AOI22_X1   g10097(.A1(new_n10050_), .A2(new_n10033_), .B1(new_n10048_), .B2(new_n10049_), .ZN(new_n11100_));
  NOR4_X1    g10098(.A1(new_n10046_), .A2(new_n10042_), .A3(new_n10045_), .A4(new_n9405_), .ZN(new_n11101_));
  OAI22_X1   g10099(.A1(new_n11100_), .A2(new_n11101_), .B1(new_n10070_), .B2(new_n10071_), .ZN(new_n11102_));
  NOR4_X1    g10100(.A1(new_n11100_), .A2(new_n11101_), .A3(new_n10070_), .A4(new_n10071_), .ZN(new_n11103_));
  AOI21_X1   g10101(.A1(new_n10039_), .A2(new_n11102_), .B(new_n11103_), .ZN(new_n11104_));
  NAND2_X1   g10102(.A1(new_n11095_), .A2(new_n11091_), .ZN(new_n11105_));
  NAND2_X1   g10103(.A1(new_n11082_), .A2(new_n11086_), .ZN(new_n11106_));
  NAND4_X1   g10104(.A1(new_n10047_), .A2(new_n10062_), .A3(new_n10051_), .A4(new_n10066_), .ZN(new_n11107_));
  NAND3_X1   g10105(.A1(new_n11106_), .A2(new_n11105_), .A3(new_n11107_), .ZN(new_n11108_));
  OAI22_X1   g10106(.A1(new_n11099_), .A2(new_n11108_), .B1(new_n11104_), .B2(new_n11097_), .ZN(new_n11109_));
  OAI21_X1   g10107(.A1(new_n10111_), .A2(new_n9574_), .B(new_n10102_), .ZN(new_n11110_));
  OAI21_X1   g10108(.A1(new_n9569_), .A2(new_n9573_), .B(new_n10098_), .ZN(new_n11111_));
  OAI21_X1   g10109(.A1(new_n11111_), .A2(new_n10111_), .B(new_n10100_), .ZN(new_n11112_));
  NAND2_X1   g10110(.A1(new_n11112_), .A2(new_n11110_), .ZN(new_n11113_));
  AOI21_X1   g10111(.A1(new_n10095_), .A2(new_n9537_), .B(new_n10086_), .ZN(new_n11114_));
  AOI21_X1   g10112(.A1(new_n9535_), .A2(new_n9536_), .B(new_n10082_), .ZN(new_n11115_));
  AOI21_X1   g10113(.A1(new_n11115_), .A2(new_n10095_), .B(new_n10084_), .ZN(new_n11116_));
  NOR2_X1    g10114(.A1(new_n11116_), .A2(new_n11114_), .ZN(new_n11117_));
  NAND2_X1   g10115(.A1(new_n11117_), .A2(new_n11113_), .ZN(new_n11118_));
  NAND2_X1   g10116(.A1(new_n10107_), .A2(new_n9599_), .ZN(new_n11119_));
  NAND3_X1   g10117(.A1(new_n10107_), .A2(new_n9599_), .A3(new_n10098_), .ZN(new_n11120_));
  AOI22_X1   g10118(.A1(new_n11120_), .A2(new_n10100_), .B1(new_n11119_), .B2(new_n10102_), .ZN(new_n11121_));
  OAI21_X1   g10119(.A1(new_n10090_), .A2(new_n9615_), .B(new_n10082_), .ZN(new_n11122_));
  OAI21_X1   g10120(.A1(new_n9612_), .A2(new_n9614_), .B(new_n10086_), .ZN(new_n11123_));
  OAI21_X1   g10121(.A1(new_n11123_), .A2(new_n10090_), .B(new_n10088_), .ZN(new_n11124_));
  NAND2_X1   g10122(.A1(new_n11124_), .A2(new_n11122_), .ZN(new_n11125_));
  NAND2_X1   g10123(.A1(new_n11121_), .A2(new_n11125_), .ZN(new_n11126_));
  NAND2_X1   g10124(.A1(new_n11126_), .A2(new_n11118_), .ZN(new_n11127_));
  OAI22_X1   g10125(.A1(new_n10115_), .A2(new_n10116_), .B1(new_n10108_), .B2(new_n10112_), .ZN(new_n11128_));
  NAND2_X1   g10126(.A1(new_n10123_), .A2(new_n11128_), .ZN(new_n11129_));
  AOI22_X1   g10127(.A1(new_n10091_), .A2(new_n10096_), .B1(new_n10118_), .B2(new_n10119_), .ZN(new_n11130_));
  NAND4_X1   g10128(.A1(new_n10091_), .A2(new_n10096_), .A3(new_n10118_), .A4(new_n10119_), .ZN(new_n11131_));
  OAI21_X1   g10129(.A1(new_n10081_), .A2(new_n11130_), .B(new_n11131_), .ZN(new_n11132_));
  NOR2_X1    g10130(.A1(new_n11121_), .A2(new_n11125_), .ZN(new_n11133_));
  NOR2_X1    g10131(.A1(new_n11117_), .A2(new_n11113_), .ZN(new_n11134_));
  NOR4_X1    g10132(.A1(new_n10115_), .A2(new_n10116_), .A3(new_n10108_), .A4(new_n10112_), .ZN(new_n11135_));
  NOR3_X1    g10133(.A1(new_n11133_), .A2(new_n11134_), .A3(new_n11135_), .ZN(new_n11136_));
  AOI22_X1   g10134(.A1(new_n11136_), .A2(new_n11129_), .B1(new_n11132_), .B2(new_n11127_), .ZN(new_n11137_));
  NAND2_X1   g10135(.A1(new_n11109_), .A2(new_n11137_), .ZN(new_n11138_));
  NAND2_X1   g10136(.A1(new_n11106_), .A2(new_n11105_), .ZN(new_n11139_));
  NAND2_X1   g10137(.A1(new_n10039_), .A2(new_n11102_), .ZN(new_n11140_));
  OAI21_X1   g10138(.A1(new_n10076_), .A2(new_n11098_), .B(new_n11107_), .ZN(new_n11141_));
  NOR3_X1    g10139(.A1(new_n11087_), .A2(new_n11096_), .A3(new_n11103_), .ZN(new_n11142_));
  AOI22_X1   g10140(.A1(new_n11142_), .A2(new_n11140_), .B1(new_n11141_), .B2(new_n11139_), .ZN(new_n11143_));
  NOR2_X1    g10141(.A1(new_n11133_), .A2(new_n11134_), .ZN(new_n11144_));
  NOR2_X1    g10142(.A1(new_n10081_), .A2(new_n11130_), .ZN(new_n11145_));
  AOI21_X1   g10143(.A1(new_n10123_), .A2(new_n11128_), .B(new_n11135_), .ZN(new_n11146_));
  NAND3_X1   g10144(.A1(new_n11126_), .A2(new_n11118_), .A3(new_n11131_), .ZN(new_n11147_));
  OAI22_X1   g10145(.A1(new_n11144_), .A2(new_n11146_), .B1(new_n11147_), .B2(new_n11145_), .ZN(new_n11148_));
  NAND2_X1   g10146(.A1(new_n11143_), .A2(new_n11148_), .ZN(new_n11149_));
  AOI22_X1   g10147(.A1(new_n11079_), .A2(new_n11077_), .B1(new_n11138_), .B2(new_n11149_), .ZN(new_n11150_));
  AOI22_X1   g10148(.A1(new_n10074_), .A2(new_n10079_), .B1(new_n10132_), .B2(new_n10133_), .ZN(new_n11151_));
  OAI21_X1   g10149(.A1(new_n10029_), .A2(new_n11151_), .B(new_n11077_), .ZN(new_n11152_));
  NOR2_X1    g10150(.A1(new_n11143_), .A2(new_n11148_), .ZN(new_n11153_));
  NOR2_X1    g10151(.A1(new_n11109_), .A2(new_n11137_), .ZN(new_n11154_));
  NOR3_X1    g10152(.A1(new_n11152_), .A2(new_n11153_), .A3(new_n11154_), .ZN(new_n11155_));
  NOR2_X1    g10153(.A1(new_n11150_), .A2(new_n11155_), .ZN(new_n11156_));
  NOR2_X1    g10154(.A1(new_n10018_), .A2(new_n10014_), .ZN(new_n11157_));
  AOI21_X1   g10155(.A1(new_n10018_), .A2(new_n10014_), .B(new_n10024_), .ZN(new_n11158_));
  OAI21_X1   g10156(.A1(new_n9994_), .A2(new_n9335_), .B(new_n9983_), .ZN(new_n11159_));
  OAI21_X1   g10157(.A1(new_n9332_), .A2(new_n9334_), .B(new_n9987_), .ZN(new_n11160_));
  OAI21_X1   g10158(.A1(new_n11160_), .A2(new_n9994_), .B(new_n9991_), .ZN(new_n11161_));
  NAND2_X1   g10159(.A1(new_n11161_), .A2(new_n11159_), .ZN(new_n11162_));
  AOI21_X1   g10160(.A1(new_n9976_), .A2(new_n9281_), .B(new_n9967_), .ZN(new_n11163_));
  AOI21_X1   g10161(.A1(new_n9279_), .A2(new_n9280_), .B(new_n9971_), .ZN(new_n11164_));
  AOI21_X1   g10162(.A1(new_n11164_), .A2(new_n9976_), .B(new_n9973_), .ZN(new_n11165_));
  NOR2_X1    g10163(.A1(new_n11165_), .A2(new_n11163_), .ZN(new_n11166_));
  NAND2_X1   g10164(.A1(new_n11166_), .A2(new_n11162_), .ZN(new_n11167_));
  AOI21_X1   g10165(.A1(new_n9998_), .A2(new_n9307_), .B(new_n9987_), .ZN(new_n11168_));
  NOR2_X1    g10166(.A1(new_n9335_), .A2(new_n9983_), .ZN(new_n11169_));
  AOI21_X1   g10167(.A1(new_n11169_), .A2(new_n9998_), .B(new_n9984_), .ZN(new_n11170_));
  NOR2_X1    g10168(.A1(new_n11170_), .A2(new_n11168_), .ZN(new_n11171_));
  OAI21_X1   g10169(.A1(new_n9980_), .A2(new_n9351_), .B(new_n9971_), .ZN(new_n11172_));
  OAI21_X1   g10170(.A1(new_n9348_), .A2(new_n9350_), .B(new_n9967_), .ZN(new_n11173_));
  OAI21_X1   g10171(.A1(new_n11173_), .A2(new_n9980_), .B(new_n9969_), .ZN(new_n11174_));
  NAND2_X1   g10172(.A1(new_n11174_), .A2(new_n11172_), .ZN(new_n11175_));
  NAND2_X1   g10173(.A1(new_n11171_), .A2(new_n11175_), .ZN(new_n11176_));
  NAND2_X1   g10174(.A1(new_n11176_), .A2(new_n11167_), .ZN(new_n11177_));
  OAI22_X1   g10175(.A1(new_n9977_), .A2(new_n9981_), .B1(new_n10005_), .B2(new_n10006_), .ZN(new_n11178_));
  NAND2_X1   g10176(.A1(new_n9966_), .A2(new_n11178_), .ZN(new_n11179_));
  AOI22_X1   g10177(.A1(new_n10002_), .A2(new_n10003_), .B1(new_n9995_), .B2(new_n9999_), .ZN(new_n11180_));
  NAND4_X1   g10178(.A1(new_n10002_), .A2(new_n10003_), .A3(new_n9995_), .A4(new_n9999_), .ZN(new_n11181_));
  OAI21_X1   g10179(.A1(new_n10010_), .A2(new_n11180_), .B(new_n11181_), .ZN(new_n11182_));
  NOR2_X1    g10180(.A1(new_n11171_), .A2(new_n11175_), .ZN(new_n11183_));
  NOR2_X1    g10181(.A1(new_n11166_), .A2(new_n11162_), .ZN(new_n11184_));
  NOR4_X1    g10182(.A1(new_n9977_), .A2(new_n9981_), .A3(new_n10005_), .A4(new_n10006_), .ZN(new_n11185_));
  NOR3_X1    g10183(.A1(new_n11183_), .A2(new_n11184_), .A3(new_n11185_), .ZN(new_n11186_));
  AOI22_X1   g10184(.A1(new_n11186_), .A2(new_n11179_), .B1(new_n11177_), .B2(new_n11182_), .ZN(new_n11187_));
  NAND2_X1   g10185(.A1(new_n9945_), .A2(new_n9187_), .ZN(new_n11188_));
  NOR2_X1    g10186(.A1(new_n9211_), .A2(new_n9940_), .ZN(new_n11189_));
  NAND2_X1   g10187(.A1(new_n11189_), .A2(new_n9945_), .ZN(new_n11190_));
  AOI22_X1   g10188(.A1(new_n11190_), .A2(new_n9938_), .B1(new_n11188_), .B2(new_n9940_), .ZN(new_n11191_));
  OAI21_X1   g10189(.A1(new_n9928_), .A2(new_n9227_), .B(new_n9919_), .ZN(new_n11192_));
  OAI21_X1   g10190(.A1(new_n9224_), .A2(new_n9226_), .B(new_n9925_), .ZN(new_n11193_));
  OAI21_X1   g10191(.A1(new_n9928_), .A2(new_n11193_), .B(new_n9926_), .ZN(new_n11194_));
  NAND2_X1   g10192(.A1(new_n11194_), .A2(new_n11192_), .ZN(new_n11195_));
  NOR2_X1    g10193(.A1(new_n11191_), .A2(new_n11195_), .ZN(new_n11196_));
  OAI21_X1   g10194(.A1(new_n9949_), .A2(new_n9211_), .B(new_n9940_), .ZN(new_n11197_));
  OAI21_X1   g10195(.A1(new_n9209_), .A2(new_n9210_), .B(new_n9936_), .ZN(new_n11198_));
  OAI21_X1   g10196(.A1(new_n9949_), .A2(new_n11198_), .B(new_n9938_), .ZN(new_n11199_));
  NAND2_X1   g10197(.A1(new_n11199_), .A2(new_n11197_), .ZN(new_n11200_));
  AOI21_X1   g10198(.A1(new_n9933_), .A2(new_n9138_), .B(new_n9925_), .ZN(new_n11201_));
  AOI21_X1   g10199(.A1(new_n9136_), .A2(new_n9137_), .B(new_n9919_), .ZN(new_n11202_));
  AOI21_X1   g10200(.A1(new_n11202_), .A2(new_n9933_), .B(new_n9923_), .ZN(new_n11203_));
  NOR2_X1    g10201(.A1(new_n11203_), .A2(new_n11201_), .ZN(new_n11204_));
  NOR2_X1    g10202(.A1(new_n11204_), .A2(new_n11200_), .ZN(new_n11205_));
  NOR2_X1    g10203(.A1(new_n11196_), .A2(new_n11205_), .ZN(new_n11206_));
  AOI22_X1   g10204(.A1(new_n9929_), .A2(new_n9934_), .B1(new_n9956_), .B2(new_n9957_), .ZN(new_n11207_));
  NOR2_X1    g10205(.A1(new_n9918_), .A2(new_n11207_), .ZN(new_n11208_));
  OAI22_X1   g10206(.A1(new_n9953_), .A2(new_n9954_), .B1(new_n9946_), .B2(new_n9950_), .ZN(new_n11209_));
  NOR4_X1    g10207(.A1(new_n9953_), .A2(new_n9946_), .A3(new_n9954_), .A4(new_n9950_), .ZN(new_n11210_));
  AOI21_X1   g10208(.A1(new_n9961_), .A2(new_n11209_), .B(new_n11210_), .ZN(new_n11211_));
  NAND2_X1   g10209(.A1(new_n11204_), .A2(new_n11200_), .ZN(new_n11212_));
  NAND2_X1   g10210(.A1(new_n11191_), .A2(new_n11195_), .ZN(new_n11213_));
  NAND4_X1   g10211(.A1(new_n9929_), .A2(new_n9956_), .A3(new_n9934_), .A4(new_n9957_), .ZN(new_n11214_));
  NAND3_X1   g10212(.A1(new_n11213_), .A2(new_n11212_), .A3(new_n11214_), .ZN(new_n11215_));
  OAI22_X1   g10213(.A1(new_n11208_), .A2(new_n11215_), .B1(new_n11206_), .B2(new_n11211_), .ZN(new_n11216_));
  NOR2_X1    g10214(.A1(new_n11216_), .A2(new_n11187_), .ZN(new_n11217_));
  NOR2_X1    g10215(.A1(new_n11183_), .A2(new_n11184_), .ZN(new_n11218_));
  NOR2_X1    g10216(.A1(new_n10010_), .A2(new_n11180_), .ZN(new_n11219_));
  AOI21_X1   g10217(.A1(new_n9966_), .A2(new_n11178_), .B(new_n11185_), .ZN(new_n11220_));
  NAND3_X1   g10218(.A1(new_n11176_), .A2(new_n11167_), .A3(new_n11181_), .ZN(new_n11221_));
  OAI22_X1   g10219(.A1(new_n11219_), .A2(new_n11221_), .B1(new_n11218_), .B2(new_n11220_), .ZN(new_n11222_));
  NAND2_X1   g10220(.A1(new_n11213_), .A2(new_n11212_), .ZN(new_n11223_));
  NAND2_X1   g10221(.A1(new_n9961_), .A2(new_n11209_), .ZN(new_n11224_));
  OAI21_X1   g10222(.A1(new_n9918_), .A2(new_n11207_), .B(new_n11214_), .ZN(new_n11225_));
  NOR3_X1    g10223(.A1(new_n11196_), .A2(new_n11205_), .A3(new_n11210_), .ZN(new_n11226_));
  AOI22_X1   g10224(.A1(new_n11226_), .A2(new_n11224_), .B1(new_n11223_), .B2(new_n11225_), .ZN(new_n11227_));
  NOR2_X1    g10225(.A1(new_n11227_), .A2(new_n11222_), .ZN(new_n11228_));
  OAI22_X1   g10226(.A1(new_n11217_), .A2(new_n11228_), .B1(new_n11158_), .B2(new_n11157_), .ZN(new_n11229_));
  NAND4_X1   g10227(.A1(new_n10016_), .A2(new_n10017_), .A3(new_n10009_), .A4(new_n10013_), .ZN(new_n11230_));
  OAI21_X1   g10228(.A1(new_n9965_), .A2(new_n10021_), .B(new_n9917_), .ZN(new_n11231_));
  NAND2_X1   g10229(.A1(new_n11227_), .A2(new_n11222_), .ZN(new_n11232_));
  NAND2_X1   g10230(.A1(new_n11216_), .A2(new_n11187_), .ZN(new_n11233_));
  NAND4_X1   g10231(.A1(new_n11231_), .A2(new_n11233_), .A3(new_n11232_), .A4(new_n11230_), .ZN(new_n11234_));
  NAND2_X1   g10232(.A1(new_n11229_), .A2(new_n11234_), .ZN(new_n11235_));
  NOR2_X1    g10233(.A1(new_n11156_), .A2(new_n11235_), .ZN(new_n11236_));
  NOR4_X1    g10234(.A1(new_n10130_), .A2(new_n10129_), .A3(new_n10122_), .A4(new_n10126_), .ZN(new_n11237_));
  NOR2_X1    g10235(.A1(new_n11151_), .A2(new_n10029_), .ZN(new_n11238_));
  OAI22_X1   g10236(.A1(new_n11153_), .A2(new_n11154_), .B1(new_n11238_), .B2(new_n11237_), .ZN(new_n11239_));
  NAND4_X1   g10237(.A1(new_n11079_), .A2(new_n11138_), .A3(new_n11149_), .A4(new_n11077_), .ZN(new_n11240_));
  NAND2_X1   g10238(.A1(new_n11239_), .A2(new_n11240_), .ZN(new_n11241_));
  AOI22_X1   g10239(.A1(new_n11232_), .A2(new_n11233_), .B1(new_n11231_), .B2(new_n11230_), .ZN(new_n11242_));
  NOR4_X1    g10240(.A1(new_n11217_), .A2(new_n11228_), .A3(new_n11158_), .A4(new_n11157_), .ZN(new_n11243_));
  NOR2_X1    g10241(.A1(new_n11242_), .A2(new_n11243_), .ZN(new_n11244_));
  NOR2_X1    g10242(.A1(new_n11241_), .A2(new_n11244_), .ZN(new_n11245_));
  OAI21_X1   g10243(.A1(new_n11236_), .A2(new_n11245_), .B(new_n11076_), .ZN(new_n11246_));
  OAI21_X1   g10244(.A1(new_n10145_), .A2(new_n10141_), .B(new_n10152_), .ZN(new_n11247_));
  NAND2_X1   g10245(.A1(new_n11241_), .A2(new_n11244_), .ZN(new_n11248_));
  NAND2_X1   g10246(.A1(new_n11156_), .A2(new_n11235_), .ZN(new_n11249_));
  NAND4_X1   g10247(.A1(new_n11248_), .A2(new_n11249_), .A3(new_n11247_), .A4(new_n11074_), .ZN(new_n11250_));
  NAND2_X1   g10248(.A1(new_n11246_), .A2(new_n11250_), .ZN(new_n11251_));
  NAND4_X1   g10249(.A1(new_n9902_), .A2(new_n9894_), .A3(new_n9899_), .A4(new_n9903_), .ZN(new_n11252_));
  OAI21_X1   g10250(.A1(new_n9907_), .A2(new_n9788_), .B(new_n9673_), .ZN(new_n11253_));
  NAND4_X1   g10251(.A1(new_n9887_), .A2(new_n9880_), .A3(new_n9884_), .A4(new_n9888_), .ZN(new_n11254_));
  INV_X1     g10252(.I(new_n11254_), .ZN(new_n11255_));
  AOI21_X1   g10253(.A1(new_n9889_), .A2(new_n9885_), .B(new_n9896_), .ZN(new_n11256_));
  OAI21_X1   g10254(.A1(new_n9864_), .A2(new_n9050_), .B(new_n9855_), .ZN(new_n11257_));
  OAI21_X1   g10255(.A1(new_n9048_), .A2(new_n9049_), .B(new_n9861_), .ZN(new_n11258_));
  OAI21_X1   g10256(.A1(new_n9864_), .A2(new_n11258_), .B(new_n9862_), .ZN(new_n11259_));
  NAND2_X1   g10257(.A1(new_n11259_), .A2(new_n11257_), .ZN(new_n11260_));
  NAND2_X1   g10258(.A1(new_n9848_), .A2(new_n8980_), .ZN(new_n11261_));
  NAND3_X1   g10259(.A1(new_n9848_), .A2(new_n8980_), .A3(new_n9839_), .ZN(new_n11262_));
  AOI22_X1   g10260(.A1(new_n11262_), .A2(new_n9843_), .B1(new_n11261_), .B2(new_n9845_), .ZN(new_n11263_));
  NAND2_X1   g10261(.A1(new_n11263_), .A2(new_n11260_), .ZN(new_n11264_));
  NAND2_X1   g10262(.A1(new_n9869_), .A2(new_n9028_), .ZN(new_n11265_));
  NAND3_X1   g10263(.A1(new_n9869_), .A2(new_n9028_), .A3(new_n9861_), .ZN(new_n11266_));
  AOI22_X1   g10264(.A1(new_n11266_), .A2(new_n9862_), .B1(new_n11265_), .B2(new_n9855_), .ZN(new_n11267_));
  NOR2_X1    g10265(.A1(new_n9852_), .A2(new_n9063_), .ZN(new_n11268_));
  NOR3_X1    g10266(.A1(new_n9852_), .A2(new_n9063_), .A3(new_n9845_), .ZN(new_n11269_));
  OAI22_X1   g10267(.A1(new_n11269_), .A2(new_n9846_), .B1(new_n11268_), .B2(new_n9839_), .ZN(new_n11270_));
  NAND2_X1   g10268(.A1(new_n11270_), .A2(new_n11267_), .ZN(new_n11271_));
  NAND2_X1   g10269(.A1(new_n11271_), .A2(new_n11264_), .ZN(new_n11272_));
  OAI22_X1   g10270(.A1(new_n9849_), .A2(new_n9853_), .B1(new_n9877_), .B2(new_n9876_), .ZN(new_n11273_));
  NAND2_X1   g10271(.A1(new_n9838_), .A2(new_n11273_), .ZN(new_n11274_));
  AOI22_X1   g10272(.A1(new_n9873_), .A2(new_n9874_), .B1(new_n9865_), .B2(new_n9870_), .ZN(new_n11275_));
  NAND4_X1   g10273(.A1(new_n9873_), .A2(new_n9865_), .A3(new_n9870_), .A4(new_n9874_), .ZN(new_n11276_));
  OAI21_X1   g10274(.A1(new_n9881_), .A2(new_n11275_), .B(new_n11276_), .ZN(new_n11277_));
  NOR2_X1    g10275(.A1(new_n11270_), .A2(new_n11267_), .ZN(new_n11278_));
  NOR2_X1    g10276(.A1(new_n11263_), .A2(new_n11260_), .ZN(new_n11279_));
  NOR4_X1    g10277(.A1(new_n9849_), .A2(new_n9853_), .A3(new_n9877_), .A4(new_n9876_), .ZN(new_n11280_));
  NOR3_X1    g10278(.A1(new_n11278_), .A2(new_n11279_), .A3(new_n11280_), .ZN(new_n11281_));
  AOI22_X1   g10279(.A1(new_n11281_), .A2(new_n11274_), .B1(new_n11272_), .B2(new_n11277_), .ZN(new_n11282_));
  AOI21_X1   g10280(.A1(new_n9817_), .A2(new_n8898_), .B(new_n9808_), .ZN(new_n11283_));
  NOR2_X1    g10281(.A1(new_n8922_), .A2(new_n9812_), .ZN(new_n11284_));
  AOI21_X1   g10282(.A1(new_n11284_), .A2(new_n9817_), .B(new_n9814_), .ZN(new_n11285_));
  NOR2_X1    g10283(.A1(new_n11285_), .A2(new_n11283_), .ZN(new_n11286_));
  OAI21_X1   g10284(.A1(new_n9800_), .A2(new_n8937_), .B(new_n9792_), .ZN(new_n11287_));
  OAI21_X1   g10285(.A1(new_n8935_), .A2(new_n8936_), .B(new_n9796_), .ZN(new_n11288_));
  OAI21_X1   g10286(.A1(new_n11288_), .A2(new_n9800_), .B(new_n9798_), .ZN(new_n11289_));
  NAND2_X1   g10287(.A1(new_n11289_), .A2(new_n11287_), .ZN(new_n11290_));
  NOR2_X1    g10288(.A1(new_n11286_), .A2(new_n11290_), .ZN(new_n11291_));
  OAI21_X1   g10289(.A1(new_n9821_), .A2(new_n8922_), .B(new_n9812_), .ZN(new_n11292_));
  OAI21_X1   g10290(.A1(new_n8919_), .A2(new_n8921_), .B(new_n9808_), .ZN(new_n11293_));
  OAI21_X1   g10291(.A1(new_n9821_), .A2(new_n11293_), .B(new_n9810_), .ZN(new_n11294_));
  NAND2_X1   g10292(.A1(new_n11294_), .A2(new_n11292_), .ZN(new_n11295_));
  AOI21_X1   g10293(.A1(new_n9804_), .A2(new_n8854_), .B(new_n9796_), .ZN(new_n11296_));
  AOI21_X1   g10294(.A1(new_n8852_), .A2(new_n8853_), .B(new_n9792_), .ZN(new_n11297_));
  AOI21_X1   g10295(.A1(new_n11297_), .A2(new_n9804_), .B(new_n9794_), .ZN(new_n11298_));
  NOR2_X1    g10296(.A1(new_n11298_), .A2(new_n11296_), .ZN(new_n11299_));
  NOR2_X1    g10297(.A1(new_n11299_), .A2(new_n11295_), .ZN(new_n11300_));
  NOR2_X1    g10298(.A1(new_n11291_), .A2(new_n11300_), .ZN(new_n11301_));
  AOI22_X1   g10299(.A1(new_n9801_), .A2(new_n9805_), .B1(new_n9828_), .B2(new_n9829_), .ZN(new_n11302_));
  NOR2_X1    g10300(.A1(new_n9791_), .A2(new_n11302_), .ZN(new_n11303_));
  OAI22_X1   g10301(.A1(new_n9825_), .A2(new_n9826_), .B1(new_n9818_), .B2(new_n9822_), .ZN(new_n11304_));
  NOR4_X1    g10302(.A1(new_n9825_), .A2(new_n9818_), .A3(new_n9826_), .A4(new_n9822_), .ZN(new_n11305_));
  AOI21_X1   g10303(.A1(new_n9833_), .A2(new_n11304_), .B(new_n11305_), .ZN(new_n11306_));
  NAND2_X1   g10304(.A1(new_n11299_), .A2(new_n11295_), .ZN(new_n11307_));
  NAND2_X1   g10305(.A1(new_n11286_), .A2(new_n11290_), .ZN(new_n11308_));
  NAND4_X1   g10306(.A1(new_n9801_), .A2(new_n9805_), .A3(new_n9828_), .A4(new_n9829_), .ZN(new_n11309_));
  NAND3_X1   g10307(.A1(new_n11308_), .A2(new_n11307_), .A3(new_n11309_), .ZN(new_n11310_));
  OAI22_X1   g10308(.A1(new_n11301_), .A2(new_n11306_), .B1(new_n11310_), .B2(new_n11303_), .ZN(new_n11311_));
  NOR2_X1    g10309(.A1(new_n11282_), .A2(new_n11311_), .ZN(new_n11312_));
  NOR2_X1    g10310(.A1(new_n11278_), .A2(new_n11279_), .ZN(new_n11313_));
  INV_X1     g10311(.I(new_n11274_), .ZN(new_n11314_));
  AOI21_X1   g10312(.A1(new_n9838_), .A2(new_n11273_), .B(new_n11280_), .ZN(new_n11315_));
  NAND3_X1   g10313(.A1(new_n11271_), .A2(new_n11264_), .A3(new_n11276_), .ZN(new_n11316_));
  OAI22_X1   g10314(.A1(new_n11314_), .A2(new_n11316_), .B1(new_n11313_), .B2(new_n11315_), .ZN(new_n11317_));
  NAND2_X1   g10315(.A1(new_n11308_), .A2(new_n11307_), .ZN(new_n11318_));
  NAND2_X1   g10316(.A1(new_n9833_), .A2(new_n11304_), .ZN(new_n11319_));
  OAI21_X1   g10317(.A1(new_n9791_), .A2(new_n11302_), .B(new_n11309_), .ZN(new_n11320_));
  NOR3_X1    g10318(.A1(new_n11291_), .A2(new_n11300_), .A3(new_n11305_), .ZN(new_n11321_));
  AOI22_X1   g10319(.A1(new_n11319_), .A2(new_n11321_), .B1(new_n11320_), .B2(new_n11318_), .ZN(new_n11322_));
  NOR2_X1    g10320(.A1(new_n11317_), .A2(new_n11322_), .ZN(new_n11323_));
  OAI22_X1   g10321(.A1(new_n11312_), .A2(new_n11323_), .B1(new_n11256_), .B2(new_n11255_), .ZN(new_n11324_));
  OAI21_X1   g10322(.A1(new_n9892_), .A2(new_n9837_), .B(new_n9790_), .ZN(new_n11325_));
  NAND2_X1   g10323(.A1(new_n11317_), .A2(new_n11322_), .ZN(new_n11326_));
  NAND2_X1   g10324(.A1(new_n11282_), .A2(new_n11311_), .ZN(new_n11327_));
  NAND4_X1   g10325(.A1(new_n11326_), .A2(new_n11327_), .A3(new_n11325_), .A4(new_n11254_), .ZN(new_n11328_));
  NAND2_X1   g10326(.A1(new_n11324_), .A2(new_n11328_), .ZN(new_n11329_));
  NAND4_X1   g10327(.A1(new_n9720_), .A2(new_n9778_), .A3(new_n9779_), .A4(new_n9724_), .ZN(new_n11330_));
  OAI21_X1   g10328(.A1(new_n9773_), .A2(new_n9777_), .B(new_n9784_), .ZN(new_n11331_));
  AOI21_X1   g10329(.A1(new_n9753_), .A2(new_n8760_), .B(new_n9743_), .ZN(new_n11332_));
  AOI21_X1   g10330(.A1(new_n8758_), .A2(new_n8759_), .B(new_n9746_), .ZN(new_n11333_));
  AOI21_X1   g10331(.A1(new_n11333_), .A2(new_n9753_), .B(new_n9750_), .ZN(new_n11334_));
  NOR2_X1    g10332(.A1(new_n11334_), .A2(new_n11332_), .ZN(new_n11335_));
  NOR2_X1    g10333(.A1(new_n9736_), .A2(new_n8795_), .ZN(new_n11336_));
  OAI21_X1   g10334(.A1(new_n8793_), .A2(new_n8794_), .B(new_n9730_), .ZN(new_n11337_));
  NOR2_X1    g10335(.A1(new_n11337_), .A2(new_n9736_), .ZN(new_n11338_));
  OAI22_X1   g10336(.A1(new_n11338_), .A2(new_n9728_), .B1(new_n11336_), .B2(new_n9730_), .ZN(new_n11339_));
  NOR2_X1    g10337(.A1(new_n11339_), .A2(new_n11335_), .ZN(new_n11340_));
  NOR2_X1    g10338(.A1(new_n9757_), .A2(new_n8785_), .ZN(new_n11341_));
  OAI21_X1   g10339(.A1(new_n8782_), .A2(new_n8784_), .B(new_n9743_), .ZN(new_n11342_));
  NOR2_X1    g10340(.A1(new_n9757_), .A2(new_n11342_), .ZN(new_n11343_));
  OAI22_X1   g10341(.A1(new_n9750_), .A2(new_n11343_), .B1(new_n11341_), .B2(new_n9743_), .ZN(new_n11344_));
  NAND2_X1   g10342(.A1(new_n9740_), .A2(new_n8699_), .ZN(new_n11345_));
  NAND3_X1   g10343(.A1(new_n9740_), .A2(new_n8699_), .A3(new_n9730_), .ZN(new_n11346_));
  AOI22_X1   g10344(.A1(new_n11346_), .A2(new_n9734_), .B1(new_n11345_), .B2(new_n9727_), .ZN(new_n11347_));
  NOR2_X1    g10345(.A1(new_n11344_), .A2(new_n11347_), .ZN(new_n11348_));
  NOR2_X1    g10346(.A1(new_n11348_), .A2(new_n11340_), .ZN(new_n11349_));
  AOI22_X1   g10347(.A1(new_n9764_), .A2(new_n9765_), .B1(new_n9737_), .B2(new_n9741_), .ZN(new_n11350_));
  NOR2_X1    g10348(.A1(new_n9726_), .A2(new_n11350_), .ZN(new_n11351_));
  OAI22_X1   g10349(.A1(new_n9754_), .A2(new_n9758_), .B1(new_n9761_), .B2(new_n9762_), .ZN(new_n11352_));
  NOR4_X1    g10350(.A1(new_n9761_), .A2(new_n9754_), .A3(new_n9758_), .A4(new_n9762_), .ZN(new_n11353_));
  AOI21_X1   g10351(.A1(new_n9769_), .A2(new_n11352_), .B(new_n11353_), .ZN(new_n11354_));
  NAND2_X1   g10352(.A1(new_n11344_), .A2(new_n11347_), .ZN(new_n11355_));
  NAND2_X1   g10353(.A1(new_n11339_), .A2(new_n11335_), .ZN(new_n11356_));
  NAND4_X1   g10354(.A1(new_n9764_), .A2(new_n9737_), .A3(new_n9765_), .A4(new_n9741_), .ZN(new_n11357_));
  NAND3_X1   g10355(.A1(new_n11355_), .A2(new_n11356_), .A3(new_n11357_), .ZN(new_n11358_));
  OAI22_X1   g10356(.A1(new_n11351_), .A2(new_n11358_), .B1(new_n11349_), .B2(new_n11354_), .ZN(new_n11359_));
  OAI21_X1   g10357(.A1(new_n9702_), .A2(new_n8642_), .B(new_n9693_), .ZN(new_n11360_));
  OAI21_X1   g10358(.A1(new_n8640_), .A2(new_n8641_), .B(new_n9697_), .ZN(new_n11361_));
  OAI21_X1   g10359(.A1(new_n11361_), .A2(new_n9702_), .B(new_n9699_), .ZN(new_n11362_));
  NAND2_X1   g10360(.A1(new_n11362_), .A2(new_n11360_), .ZN(new_n11363_));
  AOI21_X1   g10361(.A1(new_n9686_), .A2(new_n8654_), .B(new_n9677_), .ZN(new_n11364_));
  AOI21_X1   g10362(.A1(new_n8652_), .A2(new_n8653_), .B(new_n9680_), .ZN(new_n11365_));
  AOI21_X1   g10363(.A1(new_n11365_), .A2(new_n9686_), .B(new_n9684_), .ZN(new_n11366_));
  NOR2_X1    g10364(.A1(new_n11366_), .A2(new_n11364_), .ZN(new_n11367_));
  NAND2_X1   g10365(.A1(new_n11367_), .A2(new_n11363_), .ZN(new_n11368_));
  NAND2_X1   g10366(.A1(new_n9707_), .A2(new_n8619_), .ZN(new_n11369_));
  NAND3_X1   g10367(.A1(new_n9707_), .A2(new_n8619_), .A3(new_n9697_), .ZN(new_n11370_));
  AOI22_X1   g10368(.A1(new_n11370_), .A2(new_n9699_), .B1(new_n11369_), .B2(new_n9693_), .ZN(new_n11371_));
  OAI21_X1   g10369(.A1(new_n9689_), .A2(new_n8572_), .B(new_n9680_), .ZN(new_n11372_));
  OAI21_X1   g10370(.A1(new_n8567_), .A2(new_n8571_), .B(new_n9677_), .ZN(new_n11373_));
  OAI21_X1   g10371(.A1(new_n11373_), .A2(new_n9689_), .B(new_n9678_), .ZN(new_n11374_));
  NAND2_X1   g10372(.A1(new_n11374_), .A2(new_n11372_), .ZN(new_n11375_));
  NAND2_X1   g10373(.A1(new_n11371_), .A2(new_n11375_), .ZN(new_n11376_));
  NAND2_X1   g10374(.A1(new_n11376_), .A2(new_n11368_), .ZN(new_n11377_));
  OAI22_X1   g10375(.A1(new_n9687_), .A2(new_n9691_), .B1(new_n9715_), .B2(new_n9717_), .ZN(new_n11378_));
  NAND2_X1   g10376(.A1(new_n9676_), .A2(new_n11378_), .ZN(new_n11379_));
  AOI22_X1   g10377(.A1(new_n9712_), .A2(new_n9713_), .B1(new_n9703_), .B2(new_n9708_), .ZN(new_n11380_));
  NAND4_X1   g10378(.A1(new_n9712_), .A2(new_n9703_), .A3(new_n9713_), .A4(new_n9708_), .ZN(new_n11381_));
  OAI21_X1   g10379(.A1(new_n9721_), .A2(new_n11380_), .B(new_n11381_), .ZN(new_n11382_));
  NOR2_X1    g10380(.A1(new_n11371_), .A2(new_n11375_), .ZN(new_n11383_));
  NOR2_X1    g10381(.A1(new_n11367_), .A2(new_n11363_), .ZN(new_n11384_));
  NOR4_X1    g10382(.A1(new_n9687_), .A2(new_n9715_), .A3(new_n9691_), .A4(new_n9717_), .ZN(new_n11385_));
  NOR3_X1    g10383(.A1(new_n11383_), .A2(new_n11384_), .A3(new_n11385_), .ZN(new_n11386_));
  AOI22_X1   g10384(.A1(new_n11386_), .A2(new_n11379_), .B1(new_n11382_), .B2(new_n11377_), .ZN(new_n11387_));
  NAND2_X1   g10385(.A1(new_n11359_), .A2(new_n11387_), .ZN(new_n11388_));
  NAND2_X1   g10386(.A1(new_n11355_), .A2(new_n11356_), .ZN(new_n11389_));
  NAND2_X1   g10387(.A1(new_n9769_), .A2(new_n11352_), .ZN(new_n11390_));
  OAI21_X1   g10388(.A1(new_n9726_), .A2(new_n11350_), .B(new_n11357_), .ZN(new_n11391_));
  NOR3_X1    g10389(.A1(new_n11348_), .A2(new_n11340_), .A3(new_n11353_), .ZN(new_n11392_));
  AOI22_X1   g10390(.A1(new_n11392_), .A2(new_n11390_), .B1(new_n11389_), .B2(new_n11391_), .ZN(new_n11393_));
  NOR2_X1    g10391(.A1(new_n11383_), .A2(new_n11384_), .ZN(new_n11394_));
  NOR2_X1    g10392(.A1(new_n9721_), .A2(new_n11380_), .ZN(new_n11395_));
  AOI21_X1   g10393(.A1(new_n9676_), .A2(new_n11378_), .B(new_n11385_), .ZN(new_n11396_));
  NAND3_X1   g10394(.A1(new_n11376_), .A2(new_n11368_), .A3(new_n11381_), .ZN(new_n11397_));
  OAI22_X1   g10395(.A1(new_n11395_), .A2(new_n11397_), .B1(new_n11394_), .B2(new_n11396_), .ZN(new_n11398_));
  NAND2_X1   g10396(.A1(new_n11393_), .A2(new_n11398_), .ZN(new_n11399_));
  AOI22_X1   g10397(.A1(new_n11331_), .A2(new_n11330_), .B1(new_n11388_), .B2(new_n11399_), .ZN(new_n11400_));
  AOI22_X1   g10398(.A1(new_n9778_), .A2(new_n9779_), .B1(new_n9720_), .B2(new_n9724_), .ZN(new_n11401_));
  OAI21_X1   g10399(.A1(new_n9675_), .A2(new_n11401_), .B(new_n11330_), .ZN(new_n11402_));
  NOR2_X1    g10400(.A1(new_n11393_), .A2(new_n11398_), .ZN(new_n11403_));
  NOR2_X1    g10401(.A1(new_n11359_), .A2(new_n11387_), .ZN(new_n11404_));
  NOR3_X1    g10402(.A1(new_n11402_), .A2(new_n11403_), .A3(new_n11404_), .ZN(new_n11405_));
  NOR2_X1    g10403(.A1(new_n11400_), .A2(new_n11405_), .ZN(new_n11406_));
  NAND2_X1   g10404(.A1(new_n11406_), .A2(new_n11329_), .ZN(new_n11407_));
  AOI22_X1   g10405(.A1(new_n11326_), .A2(new_n11327_), .B1(new_n11325_), .B2(new_n11254_), .ZN(new_n11408_));
  AOI22_X1   g10406(.A1(new_n9880_), .A2(new_n9884_), .B1(new_n9887_), .B2(new_n9888_), .ZN(new_n11409_));
  OAI21_X1   g10407(.A1(new_n9896_), .A2(new_n11409_), .B(new_n11254_), .ZN(new_n11410_));
  NOR3_X1    g10408(.A1(new_n11410_), .A2(new_n11312_), .A3(new_n11323_), .ZN(new_n11411_));
  NOR2_X1    g10409(.A1(new_n11411_), .A2(new_n11408_), .ZN(new_n11412_));
  INV_X1     g10410(.I(new_n11330_), .ZN(new_n11413_));
  AOI21_X1   g10411(.A1(new_n9725_), .A2(new_n9780_), .B(new_n9675_), .ZN(new_n11414_));
  OAI22_X1   g10412(.A1(new_n11403_), .A2(new_n11404_), .B1(new_n11414_), .B2(new_n11413_), .ZN(new_n11415_));
  NAND4_X1   g10413(.A1(new_n11331_), .A2(new_n11388_), .A3(new_n11399_), .A4(new_n11330_), .ZN(new_n11416_));
  NAND2_X1   g10414(.A1(new_n11415_), .A2(new_n11416_), .ZN(new_n11417_));
  NAND2_X1   g10415(.A1(new_n11412_), .A2(new_n11417_), .ZN(new_n11418_));
  AOI22_X1   g10416(.A1(new_n11407_), .A2(new_n11418_), .B1(new_n11253_), .B2(new_n11252_), .ZN(new_n11419_));
  AOI22_X1   g10417(.A1(new_n9894_), .A2(new_n9899_), .B1(new_n9902_), .B2(new_n9903_), .ZN(new_n11420_));
  OAI21_X1   g10418(.A1(new_n9910_), .A2(new_n11420_), .B(new_n11252_), .ZN(new_n11421_));
  NOR2_X1    g10419(.A1(new_n11412_), .A2(new_n11417_), .ZN(new_n11422_));
  NOR2_X1    g10420(.A1(new_n11406_), .A2(new_n11329_), .ZN(new_n11423_));
  NOR3_X1    g10421(.A1(new_n11421_), .A2(new_n11423_), .A3(new_n11422_), .ZN(new_n11424_));
  NOR2_X1    g10422(.A1(new_n11419_), .A2(new_n11424_), .ZN(new_n11425_));
  NAND2_X1   g10423(.A1(new_n11251_), .A2(new_n11425_), .ZN(new_n11426_));
  AOI22_X1   g10424(.A1(new_n11248_), .A2(new_n11249_), .B1(new_n11074_), .B2(new_n11247_), .ZN(new_n11427_));
  NOR3_X1    g10425(.A1(new_n11076_), .A2(new_n11245_), .A3(new_n11236_), .ZN(new_n11428_));
  NOR2_X1    g10426(.A1(new_n11427_), .A2(new_n11428_), .ZN(new_n11429_));
  INV_X1     g10427(.I(new_n11252_), .ZN(new_n11430_));
  AOI21_X1   g10428(.A1(new_n9900_), .A2(new_n9904_), .B(new_n9910_), .ZN(new_n11431_));
  OAI22_X1   g10429(.A1(new_n11423_), .A2(new_n11422_), .B1(new_n11430_), .B2(new_n11431_), .ZN(new_n11432_));
  NAND4_X1   g10430(.A1(new_n11407_), .A2(new_n11418_), .A3(new_n11253_), .A4(new_n11252_), .ZN(new_n11433_));
  NAND2_X1   g10431(.A1(new_n11432_), .A2(new_n11433_), .ZN(new_n11434_));
  NAND2_X1   g10432(.A1(new_n11429_), .A2(new_n11434_), .ZN(new_n11435_));
  AOI21_X1   g10433(.A1(new_n11426_), .A2(new_n11435_), .B(new_n11073_), .ZN(new_n11436_));
  NAND4_X1   g10434(.A1(new_n9909_), .A2(new_n10161_), .A3(new_n10162_), .A4(new_n9913_), .ZN(new_n11437_));
  AOI22_X1   g10435(.A1(new_n10161_), .A2(new_n10162_), .B1(new_n9909_), .B2(new_n9913_), .ZN(new_n11438_));
  OAI21_X1   g10436(.A1(new_n9671_), .A2(new_n11438_), .B(new_n11437_), .ZN(new_n11439_));
  NOR2_X1    g10437(.A1(new_n11429_), .A2(new_n11434_), .ZN(new_n11440_));
  NOR2_X1    g10438(.A1(new_n11251_), .A2(new_n11425_), .ZN(new_n11441_));
  NOR3_X1    g10439(.A1(new_n11439_), .A2(new_n11441_), .A3(new_n11440_), .ZN(new_n11442_));
  NOR2_X1    g10440(.A1(new_n11436_), .A2(new_n11442_), .ZN(new_n11443_));
  NAND2_X1   g10441(.A1(new_n11443_), .A2(new_n11070_), .ZN(new_n11444_));
  AOI21_X1   g10442(.A1(new_n11067_), .A2(new_n11068_), .B(new_n11066_), .ZN(new_n11445_));
  NOR3_X1    g10443(.A1(new_n10706_), .A2(new_n11062_), .A3(new_n11053_), .ZN(new_n11446_));
  NOR2_X1    g10444(.A1(new_n11445_), .A2(new_n11446_), .ZN(new_n11447_));
  OAI21_X1   g10445(.A1(new_n11440_), .A2(new_n11441_), .B(new_n11439_), .ZN(new_n11448_));
  NAND3_X1   g10446(.A1(new_n11073_), .A2(new_n11426_), .A3(new_n11435_), .ZN(new_n11449_));
  NAND2_X1   g10447(.A1(new_n11448_), .A2(new_n11449_), .ZN(new_n11450_));
  NAND2_X1   g10448(.A1(new_n11447_), .A2(new_n11450_), .ZN(new_n11451_));
  AOI21_X1   g10449(.A1(new_n11444_), .A2(new_n11451_), .B(new_n10703_), .ZN(new_n11452_));
  NAND4_X1   g10450(.A1(new_n10663_), .A2(new_n10664_), .A3(new_n10655_), .A4(new_n10660_), .ZN(new_n11453_));
  AOI22_X1   g10451(.A1(new_n10663_), .A2(new_n10664_), .B1(new_n10655_), .B2(new_n10660_), .ZN(new_n11454_));
  OAI21_X1   g10452(.A1(new_n10673_), .A2(new_n11454_), .B(new_n11453_), .ZN(new_n11455_));
  NOR2_X1    g10453(.A1(new_n11447_), .A2(new_n11450_), .ZN(new_n11456_));
  NOR2_X1    g10454(.A1(new_n11443_), .A2(new_n11070_), .ZN(new_n11457_));
  NOR3_X1    g10455(.A1(new_n11456_), .A2(new_n11457_), .A3(new_n11455_), .ZN(new_n11458_));
  OAI21_X1   g10456(.A1(new_n4151_), .A2(new_n4150_), .B(new_n4148_), .ZN(new_n11459_));
  NOR2_X1    g10457(.A1(new_n4151_), .A2(new_n4148_), .ZN(new_n11460_));
  AOI22_X1   g10458(.A1(new_n11459_), .A2(new_n4167_), .B1(new_n11460_), .B2(new_n3894_), .ZN(new_n11461_));
  NOR2_X1    g10459(.A1(new_n4137_), .A2(new_n4133_), .ZN(new_n11462_));
  NAND2_X1   g10460(.A1(new_n4137_), .A2(new_n4133_), .ZN(new_n11463_));
  AOI21_X1   g10461(.A1(new_n3899_), .A2(new_n11463_), .B(new_n11462_), .ZN(new_n11464_));
  NOR2_X1    g10462(.A1(new_n4122_), .A2(new_n4120_), .ZN(new_n11465_));
  AOI21_X1   g10463(.A1(new_n4122_), .A2(new_n4120_), .B(new_n4129_), .ZN(new_n11466_));
  OAI21_X1   g10464(.A1(new_n4098_), .A2(new_n3526_), .B(new_n4089_), .ZN(new_n11467_));
  NAND2_X1   g10465(.A1(new_n3508_), .A2(new_n4096_), .ZN(new_n11468_));
  OAI21_X1   g10466(.A1(new_n11468_), .A2(new_n4098_), .B(new_n4090_), .ZN(new_n11469_));
  NAND2_X1   g10467(.A1(new_n11469_), .A2(new_n11467_), .ZN(new_n11470_));
  AOI21_X1   g10468(.A1(new_n4081_), .A2(new_n4071_), .B(new_n4072_), .ZN(new_n11471_));
  NOR2_X1    g10469(.A1(new_n3449_), .A2(new_n4076_), .ZN(new_n11472_));
  AOI21_X1   g10470(.A1(new_n11472_), .A2(new_n4081_), .B(new_n4078_), .ZN(new_n11473_));
  NOR2_X1    g10471(.A1(new_n11473_), .A2(new_n11471_), .ZN(new_n11474_));
  NAND2_X1   g10472(.A1(new_n11474_), .A2(new_n11470_), .ZN(new_n11475_));
  NOR2_X1    g10473(.A1(new_n11474_), .A2(new_n11470_), .ZN(new_n11476_));
  INV_X1     g10474(.I(new_n11476_), .ZN(new_n11477_));
  NAND2_X1   g10475(.A1(new_n11477_), .A2(new_n11475_), .ZN(new_n11478_));
  NAND2_X1   g10476(.A1(new_n4109_), .A2(new_n4105_), .ZN(new_n11479_));
  NAND2_X1   g10477(.A1(new_n11479_), .A2(new_n4069_), .ZN(new_n11480_));
  NOR4_X1    g10478(.A1(new_n4087_), .A2(new_n4082_), .A3(new_n4110_), .A4(new_n4111_), .ZN(new_n11481_));
  INV_X1     g10479(.I(new_n11481_), .ZN(new_n11482_));
  NAND2_X1   g10480(.A1(new_n11480_), .A2(new_n11482_), .ZN(new_n11483_));
  INV_X1     g10481(.I(new_n11475_), .ZN(new_n11484_));
  NOR3_X1    g10482(.A1(new_n11484_), .A2(new_n11476_), .A3(new_n11481_), .ZN(new_n11485_));
  AOI22_X1   g10483(.A1(new_n11483_), .A2(new_n11478_), .B1(new_n11485_), .B2(new_n11480_), .ZN(new_n11486_));
  OAI21_X1   g10484(.A1(new_n4045_), .A2(new_n3398_), .B(new_n4039_), .ZN(new_n11487_));
  NOR2_X1    g10485(.A1(new_n3398_), .A2(new_n4039_), .ZN(new_n11488_));
  INV_X1     g10486(.I(new_n11488_), .ZN(new_n11489_));
  OAI21_X1   g10487(.A1(new_n11489_), .A2(new_n4045_), .B(new_n4043_), .ZN(new_n11490_));
  NAND2_X1   g10488(.A1(new_n11490_), .A2(new_n11487_), .ZN(new_n11491_));
  NAND3_X1   g10489(.A1(new_n4031_), .A2(new_n4033_), .A3(new_n4023_), .ZN(new_n11492_));
  AOI22_X1   g10490(.A1(new_n11492_), .A2(new_n4025_), .B1(new_n4034_), .B2(new_n4027_), .ZN(new_n11493_));
  NAND2_X1   g10491(.A1(new_n11491_), .A2(new_n11493_), .ZN(new_n11494_));
  NAND2_X1   g10492(.A1(new_n4049_), .A2(new_n11488_), .ZN(new_n11495_));
  AOI22_X1   g10493(.A1(new_n11495_), .A2(new_n4043_), .B1(new_n4058_), .B2(new_n4039_), .ZN(new_n11496_));
  NAND2_X1   g10494(.A1(new_n4034_), .A2(new_n4027_), .ZN(new_n11497_));
  NAND2_X1   g10495(.A1(new_n11492_), .A2(new_n4025_), .ZN(new_n11498_));
  NAND2_X1   g10496(.A1(new_n11498_), .A2(new_n11497_), .ZN(new_n11499_));
  NAND2_X1   g10497(.A1(new_n11499_), .A2(new_n11496_), .ZN(new_n11500_));
  NAND2_X1   g10498(.A1(new_n11494_), .A2(new_n11500_), .ZN(new_n11501_));
  NOR2_X1    g10499(.A1(new_n4038_), .A2(new_n4060_), .ZN(new_n11502_));
  NAND4_X1   g10500(.A1(new_n4054_), .A2(new_n4046_), .A3(new_n4050_), .A4(new_n4055_), .ZN(new_n11503_));
  OAI21_X1   g10501(.A1(new_n11502_), .A2(new_n4064_), .B(new_n11503_), .ZN(new_n11504_));
  NAND2_X1   g10502(.A1(new_n11501_), .A2(new_n11504_), .ZN(new_n11505_));
  NAND2_X1   g10503(.A1(new_n4056_), .A2(new_n4051_), .ZN(new_n11506_));
  NAND2_X1   g10504(.A1(new_n11506_), .A2(new_n4021_), .ZN(new_n11507_));
  NOR2_X1    g10505(.A1(new_n11499_), .A2(new_n11496_), .ZN(new_n11508_));
  NOR2_X1    g10506(.A1(new_n11491_), .A2(new_n11493_), .ZN(new_n11509_));
  INV_X1     g10507(.I(new_n11503_), .ZN(new_n11510_));
  NOR3_X1    g10508(.A1(new_n11509_), .A2(new_n11508_), .A3(new_n11510_), .ZN(new_n11511_));
  NAND2_X1   g10509(.A1(new_n11511_), .A2(new_n11507_), .ZN(new_n11512_));
  NAND2_X1   g10510(.A1(new_n11512_), .A2(new_n11505_), .ZN(new_n11513_));
  NOR2_X1    g10511(.A1(new_n11513_), .A2(new_n11486_), .ZN(new_n11514_));
  NOR2_X1    g10512(.A1(new_n11484_), .A2(new_n11476_), .ZN(new_n11515_));
  AOI21_X1   g10513(.A1(new_n4109_), .A2(new_n4105_), .B(new_n4116_), .ZN(new_n11516_));
  NOR2_X1    g10514(.A1(new_n11516_), .A2(new_n11481_), .ZN(new_n11517_));
  NAND3_X1   g10515(.A1(new_n11477_), .A2(new_n11475_), .A3(new_n11482_), .ZN(new_n11518_));
  OAI22_X1   g10516(.A1(new_n11517_), .A2(new_n11515_), .B1(new_n11516_), .B2(new_n11518_), .ZN(new_n11519_));
  AOI22_X1   g10517(.A1(new_n11511_), .A2(new_n11507_), .B1(new_n11501_), .B2(new_n11504_), .ZN(new_n11520_));
  NOR2_X1    g10518(.A1(new_n11519_), .A2(new_n11520_), .ZN(new_n11521_));
  OAI22_X1   g10519(.A1(new_n11514_), .A2(new_n11521_), .B1(new_n11466_), .B2(new_n11465_), .ZN(new_n11522_));
  INV_X1     g10520(.I(new_n11465_), .ZN(new_n11523_));
  NAND2_X1   g10521(.A1(new_n4122_), .A2(new_n4120_), .ZN(new_n11524_));
  NAND2_X1   g10522(.A1(new_n11524_), .A2(new_n4019_), .ZN(new_n11525_));
  NAND2_X1   g10523(.A1(new_n11519_), .A2(new_n11520_), .ZN(new_n11526_));
  NAND2_X1   g10524(.A1(new_n11513_), .A2(new_n11486_), .ZN(new_n11527_));
  NAND4_X1   g10525(.A1(new_n11527_), .A2(new_n11525_), .A3(new_n11526_), .A4(new_n11523_), .ZN(new_n11528_));
  NAND2_X1   g10526(.A1(new_n11522_), .A2(new_n11528_), .ZN(new_n11529_));
  NAND2_X1   g10527(.A1(new_n4006_), .A2(new_n4002_), .ZN(new_n11530_));
  NAND2_X1   g10528(.A1(new_n3949_), .A2(new_n4009_), .ZN(new_n11531_));
  NAND2_X1   g10529(.A1(new_n11531_), .A2(new_n4013_), .ZN(new_n11532_));
  OAI21_X1   g10530(.A1(new_n3985_), .A2(new_n3952_), .B(new_n3978_), .ZN(new_n11533_));
  NAND2_X1   g10531(.A1(new_n3247_), .A2(new_n3975_), .ZN(new_n11534_));
  OAI21_X1   g10532(.A1(new_n11534_), .A2(new_n3985_), .B(new_n3976_), .ZN(new_n11535_));
  NAND2_X1   g10533(.A1(new_n11535_), .A2(new_n11533_), .ZN(new_n11536_));
  NAND3_X1   g10534(.A1(new_n3971_), .A2(new_n3271_), .A3(new_n3965_), .ZN(new_n11537_));
  AOI22_X1   g10535(.A1(new_n11537_), .A2(new_n3962_), .B1(new_n3990_), .B2(new_n3961_), .ZN(new_n11538_));
  NAND2_X1   g10536(.A1(new_n11538_), .A2(new_n11536_), .ZN(new_n11539_));
  INV_X1     g10537(.I(new_n11539_), .ZN(new_n11540_));
  NOR2_X1    g10538(.A1(new_n11538_), .A2(new_n11536_), .ZN(new_n11541_));
  NOR2_X1    g10539(.A1(new_n11540_), .A2(new_n11541_), .ZN(new_n11542_));
  AOI21_X1   g10540(.A1(new_n3973_), .A2(new_n3995_), .B(new_n3960_), .ZN(new_n11543_));
  NAND2_X1   g10541(.A1(new_n3973_), .A2(new_n3995_), .ZN(new_n11544_));
  NAND4_X1   g10542(.A1(new_n3968_), .A2(new_n3994_), .A3(new_n3972_), .A4(new_n3993_), .ZN(new_n11545_));
  INV_X1     g10543(.I(new_n11545_), .ZN(new_n11546_));
  AOI21_X1   g10544(.A1(new_n3998_), .A2(new_n11544_), .B(new_n11546_), .ZN(new_n11547_));
  INV_X1     g10545(.I(new_n11536_), .ZN(new_n11548_));
  NAND2_X1   g10546(.A1(new_n3990_), .A2(new_n3961_), .ZN(new_n11549_));
  NAND2_X1   g10547(.A1(new_n11537_), .A2(new_n3962_), .ZN(new_n11550_));
  NAND2_X1   g10548(.A1(new_n11550_), .A2(new_n11549_), .ZN(new_n11551_));
  NAND2_X1   g10549(.A1(new_n11551_), .A2(new_n11548_), .ZN(new_n11552_));
  NAND3_X1   g10550(.A1(new_n11552_), .A2(new_n11539_), .A3(new_n11545_), .ZN(new_n11553_));
  OAI22_X1   g10551(.A1(new_n11542_), .A2(new_n11547_), .B1(new_n11553_), .B2(new_n11543_), .ZN(new_n11554_));
  NOR2_X1    g10552(.A1(new_n3928_), .A2(new_n3142_), .ZN(new_n11555_));
  NAND2_X1   g10553(.A1(new_n3108_), .A2(new_n3924_), .ZN(new_n11556_));
  NOR2_X1    g10554(.A1(new_n11556_), .A2(new_n3928_), .ZN(new_n11557_));
  OAI22_X1   g10555(.A1(new_n11557_), .A2(new_n3921_), .B1(new_n11555_), .B2(new_n3924_), .ZN(new_n11558_));
  NAND2_X1   g10556(.A1(new_n3911_), .A2(new_n3061_), .ZN(new_n11559_));
  NAND3_X1   g10557(.A1(new_n3911_), .A2(new_n3061_), .A3(new_n3902_), .ZN(new_n11560_));
  AOI22_X1   g10558(.A1(new_n11560_), .A2(new_n3905_), .B1(new_n11559_), .B2(new_n3907_), .ZN(new_n11561_));
  NAND2_X1   g10559(.A1(new_n11558_), .A2(new_n11561_), .ZN(new_n11562_));
  NAND2_X1   g10560(.A1(new_n3932_), .A2(new_n3108_), .ZN(new_n11563_));
  NAND3_X1   g10561(.A1(new_n3932_), .A2(new_n3108_), .A3(new_n3924_), .ZN(new_n11564_));
  AOI22_X1   g10562(.A1(new_n11564_), .A2(new_n3926_), .B1(new_n11563_), .B2(new_n3918_), .ZN(new_n11565_));
  OAI21_X1   g10563(.A1(new_n3915_), .A2(new_n3133_), .B(new_n3907_), .ZN(new_n11566_));
  NAND2_X1   g10564(.A1(new_n3061_), .A2(new_n3902_), .ZN(new_n11567_));
  OAI21_X1   g10565(.A1(new_n11567_), .A2(new_n3915_), .B(new_n3905_), .ZN(new_n11568_));
  NAND2_X1   g10566(.A1(new_n11568_), .A2(new_n11566_), .ZN(new_n11569_));
  NAND2_X1   g10567(.A1(new_n11569_), .A2(new_n11565_), .ZN(new_n11570_));
  NAND2_X1   g10568(.A1(new_n11562_), .A2(new_n11570_), .ZN(new_n11571_));
  NAND2_X1   g10569(.A1(new_n3938_), .A2(new_n3934_), .ZN(new_n11572_));
  NAND2_X1   g10570(.A1(new_n3901_), .A2(new_n11572_), .ZN(new_n11573_));
  NOR2_X1    g10571(.A1(new_n3917_), .A2(new_n3941_), .ZN(new_n11574_));
  NAND4_X1   g10572(.A1(new_n3936_), .A2(new_n3937_), .A3(new_n3929_), .A4(new_n3933_), .ZN(new_n11575_));
  OAI21_X1   g10573(.A1(new_n11574_), .A2(new_n3945_), .B(new_n11575_), .ZN(new_n11576_));
  NOR2_X1    g10574(.A1(new_n11569_), .A2(new_n11565_), .ZN(new_n11577_));
  NOR2_X1    g10575(.A1(new_n11558_), .A2(new_n11561_), .ZN(new_n11578_));
  NOR4_X1    g10576(.A1(new_n3916_), .A2(new_n3912_), .A3(new_n3939_), .A4(new_n3940_), .ZN(new_n11579_));
  NOR3_X1    g10577(.A1(new_n11578_), .A2(new_n11577_), .A3(new_n11579_), .ZN(new_n11580_));
  AOI22_X1   g10578(.A1(new_n11580_), .A2(new_n11573_), .B1(new_n11571_), .B2(new_n11576_), .ZN(new_n11581_));
  NAND2_X1   g10579(.A1(new_n11554_), .A2(new_n11581_), .ZN(new_n11582_));
  NAND2_X1   g10580(.A1(new_n11552_), .A2(new_n11539_), .ZN(new_n11583_));
  NAND2_X1   g10581(.A1(new_n11544_), .A2(new_n3998_), .ZN(new_n11584_));
  NAND2_X1   g10582(.A1(new_n11584_), .A2(new_n11545_), .ZN(new_n11585_));
  NOR3_X1    g10583(.A1(new_n11540_), .A2(new_n11541_), .A3(new_n11546_), .ZN(new_n11586_));
  AOI22_X1   g10584(.A1(new_n11585_), .A2(new_n11583_), .B1(new_n11586_), .B2(new_n11584_), .ZN(new_n11587_));
  NOR2_X1    g10585(.A1(new_n11578_), .A2(new_n11577_), .ZN(new_n11588_));
  NOR2_X1    g10586(.A1(new_n11574_), .A2(new_n3945_), .ZN(new_n11589_));
  AOI21_X1   g10587(.A1(new_n3901_), .A2(new_n11572_), .B(new_n11579_), .ZN(new_n11590_));
  NAND3_X1   g10588(.A1(new_n11562_), .A2(new_n11570_), .A3(new_n11575_), .ZN(new_n11591_));
  OAI22_X1   g10589(.A1(new_n11588_), .A2(new_n11590_), .B1(new_n11591_), .B2(new_n11589_), .ZN(new_n11592_));
  NAND2_X1   g10590(.A1(new_n11587_), .A2(new_n11592_), .ZN(new_n11593_));
  AOI22_X1   g10591(.A1(new_n11532_), .A2(new_n11530_), .B1(new_n11593_), .B2(new_n11582_), .ZN(new_n11594_));
  NOR2_X1    g10592(.A1(new_n3949_), .A2(new_n4009_), .ZN(new_n11595_));
  AOI21_X1   g10593(.A1(new_n3949_), .A2(new_n4009_), .B(new_n3900_), .ZN(new_n11596_));
  NOR2_X1    g10594(.A1(new_n11587_), .A2(new_n11592_), .ZN(new_n11597_));
  NOR2_X1    g10595(.A1(new_n11554_), .A2(new_n11581_), .ZN(new_n11598_));
  NOR4_X1    g10596(.A1(new_n11597_), .A2(new_n11596_), .A3(new_n11598_), .A4(new_n11595_), .ZN(new_n11599_));
  NOR2_X1    g10597(.A1(new_n11594_), .A2(new_n11599_), .ZN(new_n11600_));
  NAND2_X1   g10598(.A1(new_n11529_), .A2(new_n11600_), .ZN(new_n11601_));
  AOI22_X1   g10599(.A1(new_n11527_), .A2(new_n11526_), .B1(new_n11525_), .B2(new_n11523_), .ZN(new_n11602_));
  NOR4_X1    g10600(.A1(new_n11514_), .A2(new_n11466_), .A3(new_n11521_), .A4(new_n11465_), .ZN(new_n11603_));
  NOR2_X1    g10601(.A1(new_n11602_), .A2(new_n11603_), .ZN(new_n11604_));
  OAI22_X1   g10602(.A1(new_n11597_), .A2(new_n11598_), .B1(new_n11596_), .B2(new_n11595_), .ZN(new_n11605_));
  NAND4_X1   g10603(.A1(new_n11532_), .A2(new_n11593_), .A3(new_n11582_), .A4(new_n11530_), .ZN(new_n11606_));
  NAND2_X1   g10604(.A1(new_n11605_), .A2(new_n11606_), .ZN(new_n11607_));
  NAND2_X1   g10605(.A1(new_n11604_), .A2(new_n11607_), .ZN(new_n11608_));
  AOI21_X1   g10606(.A1(new_n11601_), .A2(new_n11608_), .B(new_n11464_), .ZN(new_n11609_));
  NAND2_X1   g10607(.A1(new_n4017_), .A2(new_n4140_), .ZN(new_n11610_));
  NOR2_X1    g10608(.A1(new_n4017_), .A2(new_n4140_), .ZN(new_n11611_));
  OAI21_X1   g10609(.A1(new_n4144_), .A2(new_n11611_), .B(new_n11610_), .ZN(new_n11612_));
  NOR2_X1    g10610(.A1(new_n11604_), .A2(new_n11607_), .ZN(new_n11613_));
  NOR2_X1    g10611(.A1(new_n11529_), .A2(new_n11600_), .ZN(new_n11614_));
  NOR3_X1    g10612(.A1(new_n11612_), .A2(new_n11614_), .A3(new_n11613_), .ZN(new_n11615_));
  NOR2_X1    g10613(.A1(new_n11609_), .A2(new_n11615_), .ZN(new_n11616_));
  NAND2_X1   g10614(.A1(new_n3665_), .A2(new_n3661_), .ZN(new_n11617_));
  NOR2_X1    g10615(.A1(new_n3665_), .A2(new_n3661_), .ZN(new_n11618_));
  OAI21_X1   g10616(.A1(new_n3564_), .A2(new_n11618_), .B(new_n11617_), .ZN(new_n11619_));
  OAI21_X1   g10617(.A1(new_n3643_), .A2(new_n2490_), .B(new_n3636_), .ZN(new_n11620_));
  NAND2_X1   g10618(.A1(new_n2516_), .A2(new_n3633_), .ZN(new_n11621_));
  OAI21_X1   g10619(.A1(new_n11621_), .A2(new_n3643_), .B(new_n3634_), .ZN(new_n11622_));
  NAND2_X1   g10620(.A1(new_n11622_), .A2(new_n11620_), .ZN(new_n11623_));
  NAND2_X1   g10621(.A1(new_n3648_), .A2(new_n3616_), .ZN(new_n11624_));
  NAND2_X1   g10622(.A1(new_n2528_), .A2(new_n3623_), .ZN(new_n11625_));
  OAI21_X1   g10623(.A1(new_n11625_), .A2(new_n3626_), .B(new_n3624_), .ZN(new_n11626_));
  NAND2_X1   g10624(.A1(new_n11624_), .A2(new_n11626_), .ZN(new_n11627_));
  INV_X1     g10625(.I(new_n11627_), .ZN(new_n11628_));
  NAND2_X1   g10626(.A1(new_n11628_), .A2(new_n11623_), .ZN(new_n11629_));
  INV_X1     g10627(.I(new_n11623_), .ZN(new_n11630_));
  NAND2_X1   g10628(.A1(new_n11630_), .A2(new_n11627_), .ZN(new_n11631_));
  NAND2_X1   g10629(.A1(new_n11629_), .A2(new_n11631_), .ZN(new_n11632_));
  NAND2_X1   g10630(.A1(new_n3632_), .A2(new_n3653_), .ZN(new_n11633_));
  NAND2_X1   g10631(.A1(new_n11633_), .A2(new_n3657_), .ZN(new_n11634_));
  NAND4_X1   g10632(.A1(new_n3627_), .A2(new_n3651_), .A3(new_n3631_), .A4(new_n3652_), .ZN(new_n11635_));
  NAND2_X1   g10633(.A1(new_n11634_), .A2(new_n11635_), .ZN(new_n11636_));
  NOR2_X1    g10634(.A1(new_n11630_), .A2(new_n11627_), .ZN(new_n11637_));
  NOR2_X1    g10635(.A1(new_n11628_), .A2(new_n11623_), .ZN(new_n11638_));
  INV_X1     g10636(.I(new_n11635_), .ZN(new_n11639_));
  NOR3_X1    g10637(.A1(new_n11638_), .A2(new_n11637_), .A3(new_n11639_), .ZN(new_n11640_));
  AOI22_X1   g10638(.A1(new_n11640_), .A2(new_n11634_), .B1(new_n11636_), .B2(new_n11632_), .ZN(new_n11641_));
  NAND2_X1   g10639(.A1(new_n3604_), .A2(new_n3582_), .ZN(new_n11642_));
  NAND2_X1   g10640(.A1(new_n2426_), .A2(new_n3588_), .ZN(new_n11643_));
  OAI21_X1   g10641(.A1(new_n11643_), .A2(new_n3591_), .B(new_n3589_), .ZN(new_n11644_));
  NAND2_X1   g10642(.A1(new_n11642_), .A2(new_n11644_), .ZN(new_n11645_));
  INV_X1     g10643(.I(new_n11645_), .ZN(new_n11646_));
  NAND2_X1   g10644(.A1(new_n3577_), .A2(new_n3571_), .ZN(new_n11647_));
  NAND2_X1   g10645(.A1(new_n2366_), .A2(new_n3568_), .ZN(new_n11648_));
  OAI21_X1   g10646(.A1(new_n11648_), .A2(new_n3599_), .B(new_n3569_), .ZN(new_n11649_));
  NAND2_X1   g10647(.A1(new_n11647_), .A2(new_n11649_), .ZN(new_n11650_));
  NOR2_X1    g10648(.A1(new_n11646_), .A2(new_n11650_), .ZN(new_n11651_));
  AND2_X2    g10649(.A1(new_n11647_), .A2(new_n11649_), .Z(new_n11652_));
  NOR2_X1    g10650(.A1(new_n11652_), .A2(new_n11645_), .ZN(new_n11653_));
  NOR2_X1    g10651(.A1(new_n11651_), .A2(new_n11653_), .ZN(new_n11654_));
  NAND2_X1   g10652(.A1(new_n3597_), .A2(new_n3602_), .ZN(new_n11655_));
  NAND2_X1   g10653(.A1(new_n3566_), .A2(new_n11655_), .ZN(new_n11656_));
  INV_X1     g10654(.I(new_n11656_), .ZN(new_n11657_));
  NAND4_X1   g10655(.A1(new_n3592_), .A2(new_n3600_), .A3(new_n3601_), .A4(new_n3596_), .ZN(new_n11658_));
  INV_X1     g10656(.I(new_n11658_), .ZN(new_n11659_));
  AOI21_X1   g10657(.A1(new_n3566_), .A2(new_n11655_), .B(new_n11659_), .ZN(new_n11660_));
  NAND2_X1   g10658(.A1(new_n11652_), .A2(new_n11645_), .ZN(new_n11661_));
  NAND2_X1   g10659(.A1(new_n11646_), .A2(new_n11650_), .ZN(new_n11662_));
  NAND3_X1   g10660(.A1(new_n11662_), .A2(new_n11661_), .A3(new_n11658_), .ZN(new_n11663_));
  OAI22_X1   g10661(.A1(new_n11663_), .A2(new_n11657_), .B1(new_n11654_), .B2(new_n11660_), .ZN(new_n11664_));
  NOR2_X1    g10662(.A1(new_n11664_), .A2(new_n11641_), .ZN(new_n11665_));
  NAND2_X1   g10663(.A1(new_n11636_), .A2(new_n11632_), .ZN(new_n11666_));
  NAND4_X1   g10664(.A1(new_n11634_), .A2(new_n11629_), .A3(new_n11631_), .A4(new_n11635_), .ZN(new_n11667_));
  NAND2_X1   g10665(.A1(new_n11666_), .A2(new_n11667_), .ZN(new_n11668_));
  NAND2_X1   g10666(.A1(new_n11662_), .A2(new_n11661_), .ZN(new_n11669_));
  NAND2_X1   g10667(.A1(new_n11656_), .A2(new_n11658_), .ZN(new_n11670_));
  NOR3_X1    g10668(.A1(new_n11651_), .A2(new_n11653_), .A3(new_n11659_), .ZN(new_n11671_));
  AOI22_X1   g10669(.A1(new_n11669_), .A2(new_n11670_), .B1(new_n11671_), .B2(new_n11656_), .ZN(new_n11672_));
  NOR2_X1    g10670(.A1(new_n11668_), .A2(new_n11672_), .ZN(new_n11673_));
  OAI21_X1   g10671(.A1(new_n11665_), .A2(new_n11673_), .B(new_n11619_), .ZN(new_n11674_));
  NOR2_X1    g10672(.A1(new_n3613_), .A2(new_n3668_), .ZN(new_n11675_));
  NAND2_X1   g10673(.A1(new_n3613_), .A2(new_n3668_), .ZN(new_n11676_));
  AOI21_X1   g10674(.A1(new_n3563_), .A2(new_n11676_), .B(new_n11675_), .ZN(new_n11677_));
  NAND2_X1   g10675(.A1(new_n11668_), .A2(new_n11672_), .ZN(new_n11678_));
  NAND2_X1   g10676(.A1(new_n11664_), .A2(new_n11641_), .ZN(new_n11679_));
  NAND3_X1   g10677(.A1(new_n11677_), .A2(new_n11678_), .A3(new_n11679_), .ZN(new_n11680_));
  NAND2_X1   g10678(.A1(new_n11674_), .A2(new_n11680_), .ZN(new_n11681_));
  NAND4_X1   g10679(.A1(new_n3715_), .A2(new_n3719_), .A3(new_n3772_), .A4(new_n3773_), .ZN(new_n11682_));
  INV_X1     g10680(.I(new_n11682_), .ZN(new_n11683_));
  AOI22_X1   g10681(.A1(new_n3719_), .A2(new_n3715_), .B1(new_n3772_), .B2(new_n3773_), .ZN(new_n11684_));
  NOR2_X1    g10682(.A1(new_n11684_), .A2(new_n3677_), .ZN(new_n11685_));
  OAI21_X1   g10683(.A1(new_n3754_), .A2(new_n2946_), .B(new_n3746_), .ZN(new_n11686_));
  NAND2_X1   g10684(.A1(new_n2969_), .A2(new_n3742_), .ZN(new_n11687_));
  OAI21_X1   g10685(.A1(new_n11687_), .A2(new_n3754_), .B(new_n3744_), .ZN(new_n11688_));
  NAND2_X1   g10686(.A1(new_n11688_), .A2(new_n11686_), .ZN(new_n11689_));
  AOI21_X1   g10687(.A1(new_n3736_), .A2(new_n2918_), .B(new_n3725_), .ZN(new_n11690_));
  NOR2_X1    g10688(.A1(new_n2984_), .A2(new_n3722_), .ZN(new_n11691_));
  AOI21_X1   g10689(.A1(new_n11691_), .A2(new_n3736_), .B(new_n3723_), .ZN(new_n11692_));
  NOR2_X1    g10690(.A1(new_n11692_), .A2(new_n11690_), .ZN(new_n11693_));
  NAND2_X1   g10691(.A1(new_n11693_), .A2(new_n11689_), .ZN(new_n11694_));
  OAI21_X1   g10692(.A1(new_n3732_), .A2(new_n2984_), .B(new_n3722_), .ZN(new_n11695_));
  OAI21_X1   g10693(.A1(new_n2982_), .A2(new_n2983_), .B(new_n3725_), .ZN(new_n11696_));
  OAI21_X1   g10694(.A1(new_n11696_), .A2(new_n3732_), .B(new_n3729_), .ZN(new_n11697_));
  NAND2_X1   g10695(.A1(new_n11697_), .A2(new_n11695_), .ZN(new_n11698_));
  NAND3_X1   g10696(.A1(new_n11698_), .A2(new_n11686_), .A3(new_n11688_), .ZN(new_n11699_));
  NAND2_X1   g10697(.A1(new_n11694_), .A2(new_n11699_), .ZN(new_n11700_));
  AOI22_X1   g10698(.A1(new_n3733_), .A2(new_n3737_), .B1(new_n3761_), .B2(new_n3762_), .ZN(new_n11701_));
  INV_X1     g10699(.I(new_n11701_), .ZN(new_n11702_));
  NAND2_X1   g10700(.A1(new_n11702_), .A2(new_n3766_), .ZN(new_n11703_));
  NAND4_X1   g10701(.A1(new_n3733_), .A2(new_n3737_), .A3(new_n3761_), .A4(new_n3762_), .ZN(new_n11704_));
  OAI21_X1   g10702(.A1(new_n3721_), .A2(new_n11701_), .B(new_n11704_), .ZN(new_n11705_));
  AOI21_X1   g10703(.A1(new_n11686_), .A2(new_n11688_), .B(new_n11698_), .ZN(new_n11706_));
  NOR2_X1    g10704(.A1(new_n11693_), .A2(new_n11689_), .ZN(new_n11707_));
  NOR4_X1    g10705(.A1(new_n3758_), .A2(new_n3759_), .A3(new_n3751_), .A4(new_n3755_), .ZN(new_n11708_));
  NOR3_X1    g10706(.A1(new_n11707_), .A2(new_n11706_), .A3(new_n11708_), .ZN(new_n11709_));
  AOI22_X1   g10707(.A1(new_n11709_), .A2(new_n11703_), .B1(new_n11700_), .B2(new_n11705_), .ZN(new_n11710_));
  NAND2_X1   g10708(.A1(new_n3698_), .A2(new_n2836_), .ZN(new_n11711_));
  OAI21_X1   g10709(.A1(new_n2853_), .A2(new_n2854_), .B(new_n3692_), .ZN(new_n11712_));
  INV_X1     g10710(.I(new_n11712_), .ZN(new_n11713_));
  NAND2_X1   g10711(.A1(new_n11713_), .A2(new_n3698_), .ZN(new_n11714_));
  AOI22_X1   g10712(.A1(new_n11714_), .A2(new_n3693_), .B1(new_n3695_), .B2(new_n11711_), .ZN(new_n11715_));
  OAI21_X1   g10713(.A1(new_n3684_), .A2(new_n2871_), .B(new_n3678_), .ZN(new_n11716_));
  NAND2_X1   g10714(.A1(new_n2795_), .A2(new_n3681_), .ZN(new_n11717_));
  OAI21_X1   g10715(.A1(new_n11717_), .A2(new_n3684_), .B(new_n3682_), .ZN(new_n11718_));
  NAND2_X1   g10716(.A1(new_n11718_), .A2(new_n11716_), .ZN(new_n11719_));
  NOR2_X1    g10717(.A1(new_n11715_), .A2(new_n11719_), .ZN(new_n11720_));
  OAI21_X1   g10718(.A1(new_n3703_), .A2(new_n2855_), .B(new_n3695_), .ZN(new_n11721_));
  OAI21_X1   g10719(.A1(new_n3703_), .A2(new_n11712_), .B(new_n3693_), .ZN(new_n11722_));
  NAND2_X1   g10720(.A1(new_n11722_), .A2(new_n11721_), .ZN(new_n11723_));
  NAND2_X1   g10721(.A1(new_n3689_), .A2(new_n2795_), .ZN(new_n11724_));
  AOI21_X1   g10722(.A1(new_n2790_), .A2(new_n2794_), .B(new_n3678_), .ZN(new_n11725_));
  NAND2_X1   g10723(.A1(new_n11725_), .A2(new_n3689_), .ZN(new_n11726_));
  AOI22_X1   g10724(.A1(new_n11726_), .A2(new_n3682_), .B1(new_n11724_), .B2(new_n3678_), .ZN(new_n11727_));
  NOR2_X1    g10725(.A1(new_n11727_), .A2(new_n11723_), .ZN(new_n11728_));
  NOR2_X1    g10726(.A1(new_n11720_), .A2(new_n11728_), .ZN(new_n11729_));
  AOI22_X1   g10727(.A1(new_n3685_), .A2(new_n3690_), .B1(new_n3710_), .B2(new_n3711_), .ZN(new_n11730_));
  NOR2_X1    g10728(.A1(new_n3714_), .A2(new_n11730_), .ZN(new_n11731_));
  OAI22_X1   g10729(.A1(new_n3707_), .A2(new_n3708_), .B1(new_n3704_), .B2(new_n3699_), .ZN(new_n11732_));
  NOR4_X1    g10730(.A1(new_n3707_), .A2(new_n3708_), .A3(new_n3704_), .A4(new_n3699_), .ZN(new_n11733_));
  AOI21_X1   g10731(.A1(new_n3718_), .A2(new_n11732_), .B(new_n11733_), .ZN(new_n11734_));
  NAND2_X1   g10732(.A1(new_n11727_), .A2(new_n11723_), .ZN(new_n11735_));
  NAND2_X1   g10733(.A1(new_n11715_), .A2(new_n11719_), .ZN(new_n11736_));
  NAND4_X1   g10734(.A1(new_n3685_), .A2(new_n3690_), .A3(new_n3710_), .A4(new_n3711_), .ZN(new_n11737_));
  NAND3_X1   g10735(.A1(new_n11736_), .A2(new_n11735_), .A3(new_n11737_), .ZN(new_n11738_));
  OAI22_X1   g10736(.A1(new_n11731_), .A2(new_n11738_), .B1(new_n11729_), .B2(new_n11734_), .ZN(new_n11739_));
  NOR2_X1    g10737(.A1(new_n11739_), .A2(new_n11710_), .ZN(new_n11740_));
  NOR2_X1    g10738(.A1(new_n11707_), .A2(new_n11706_), .ZN(new_n11741_));
  NOR2_X1    g10739(.A1(new_n3721_), .A2(new_n11701_), .ZN(new_n11742_));
  AOI21_X1   g10740(.A1(new_n11702_), .A2(new_n3766_), .B(new_n11708_), .ZN(new_n11743_));
  NAND3_X1   g10741(.A1(new_n11694_), .A2(new_n11699_), .A3(new_n11704_), .ZN(new_n11744_));
  OAI22_X1   g10742(.A1(new_n11741_), .A2(new_n11743_), .B1(new_n11744_), .B2(new_n11742_), .ZN(new_n11745_));
  NAND2_X1   g10743(.A1(new_n11736_), .A2(new_n11735_), .ZN(new_n11746_));
  NAND2_X1   g10744(.A1(new_n3718_), .A2(new_n11732_), .ZN(new_n11747_));
  OAI21_X1   g10745(.A1(new_n3714_), .A2(new_n11730_), .B(new_n11737_), .ZN(new_n11748_));
  NOR3_X1    g10746(.A1(new_n11720_), .A2(new_n11728_), .A3(new_n11733_), .ZN(new_n11749_));
  AOI22_X1   g10747(.A1(new_n11749_), .A2(new_n11747_), .B1(new_n11746_), .B2(new_n11748_), .ZN(new_n11750_));
  NOR2_X1    g10748(.A1(new_n11750_), .A2(new_n11745_), .ZN(new_n11751_));
  OAI22_X1   g10749(.A1(new_n11740_), .A2(new_n11751_), .B1(new_n11685_), .B2(new_n11683_), .ZN(new_n11752_));
  OAI21_X1   g10750(.A1(new_n3781_), .A2(new_n3770_), .B(new_n3778_), .ZN(new_n11753_));
  NAND2_X1   g10751(.A1(new_n11750_), .A2(new_n11745_), .ZN(new_n11754_));
  NAND2_X1   g10752(.A1(new_n11739_), .A2(new_n11710_), .ZN(new_n11755_));
  NAND4_X1   g10753(.A1(new_n11754_), .A2(new_n11755_), .A3(new_n11753_), .A4(new_n11682_), .ZN(new_n11756_));
  AOI21_X1   g10754(.A1(new_n3851_), .A2(new_n3855_), .B(new_n3859_), .ZN(new_n11757_));
  NAND2_X1   g10755(.A1(new_n3851_), .A2(new_n3859_), .ZN(new_n11758_));
  OAI22_X1   g10756(.A1(new_n11757_), .A2(new_n3786_), .B1(new_n11758_), .B2(new_n3861_), .ZN(new_n11759_));
  AOI21_X1   g10757(.A1(new_n3791_), .A2(new_n2577_), .B(new_n3793_), .ZN(new_n11760_));
  INV_X1     g10758(.I(new_n11760_), .ZN(new_n11761_));
  NAND3_X1   g10759(.A1(new_n2595_), .A2(new_n3798_), .A3(new_n3799_), .ZN(new_n11762_));
  OAI21_X1   g10760(.A1(new_n11762_), .A2(new_n3788_), .B(new_n3797_), .ZN(new_n11763_));
  OAI21_X1   g10761(.A1(new_n3788_), .A2(new_n3802_), .B(new_n3804_), .ZN(new_n11764_));
  AOI21_X1   g10762(.A1(new_n11763_), .A2(new_n11764_), .B(new_n11761_), .ZN(new_n11765_));
  NAND2_X1   g10763(.A1(new_n2596_), .A2(new_n2553_), .ZN(new_n11766_));
  NOR3_X1    g10764(.A1(new_n3802_), .A2(new_n3792_), .A3(new_n3795_), .ZN(new_n11767_));
  AOI21_X1   g10765(.A1(new_n11767_), .A2(new_n11766_), .B(new_n3789_), .ZN(new_n11768_));
  AOI22_X1   g10766(.A1(new_n11766_), .A2(new_n2595_), .B1(new_n3798_), .B2(new_n3799_), .ZN(new_n11769_));
  NOR3_X1    g10767(.A1(new_n11768_), .A2(new_n11769_), .A3(new_n11760_), .ZN(new_n11770_));
  NOR2_X1    g10768(.A1(new_n11765_), .A2(new_n11770_), .ZN(new_n11771_));
  NAND2_X1   g10769(.A1(new_n3835_), .A2(new_n2697_), .ZN(new_n11772_));
  NAND3_X1   g10770(.A1(new_n3835_), .A2(new_n2697_), .A3(new_n3824_), .ZN(new_n11773_));
  AOI22_X1   g10771(.A1(new_n11773_), .A2(new_n3826_), .B1(new_n11772_), .B2(new_n3830_), .ZN(new_n11774_));
  OAI21_X1   g10772(.A1(new_n3817_), .A2(new_n2645_), .B(new_n3808_), .ZN(new_n11775_));
  NAND2_X1   g10773(.A1(new_n2714_), .A2(new_n3814_), .ZN(new_n11776_));
  OAI21_X1   g10774(.A1(new_n11776_), .A2(new_n3817_), .B(new_n3815_), .ZN(new_n11777_));
  NAND2_X1   g10775(.A1(new_n11777_), .A2(new_n11775_), .ZN(new_n11778_));
  NOR2_X1    g10776(.A1(new_n11778_), .A2(new_n11774_), .ZN(new_n11779_));
  OAI21_X1   g10777(.A1(new_n3839_), .A2(new_n2672_), .B(new_n3830_), .ZN(new_n11780_));
  NAND2_X1   g10778(.A1(new_n2697_), .A2(new_n3824_), .ZN(new_n11781_));
  OAI21_X1   g10779(.A1(new_n11781_), .A2(new_n3839_), .B(new_n3826_), .ZN(new_n11782_));
  NAND2_X1   g10780(.A1(new_n11782_), .A2(new_n11780_), .ZN(new_n11783_));
  NAND2_X1   g10781(.A1(new_n3821_), .A2(new_n2714_), .ZN(new_n11784_));
  NAND3_X1   g10782(.A1(new_n3821_), .A2(new_n2714_), .A3(new_n3814_), .ZN(new_n11785_));
  AOI22_X1   g10783(.A1(new_n11785_), .A2(new_n3815_), .B1(new_n11784_), .B2(new_n3808_), .ZN(new_n11786_));
  NOR2_X1    g10784(.A1(new_n11783_), .A2(new_n11786_), .ZN(new_n11787_));
  NAND2_X1   g10785(.A1(new_n2691_), .A2(new_n2706_), .ZN(new_n11788_));
  OAI22_X1   g10786(.A1(new_n11788_), .A2(new_n2700_), .B1(new_n2712_), .B2(new_n2716_), .ZN(new_n11789_));
  AOI22_X1   g10787(.A1(new_n11789_), .A2(new_n2719_), .B1(new_n3823_), .B2(new_n3848_), .ZN(new_n11790_));
  NOR4_X1    g10788(.A1(new_n3844_), .A2(new_n3843_), .A3(new_n3836_), .A4(new_n3840_), .ZN(new_n11791_));
  OAI22_X1   g10789(.A1(new_n11790_), .A2(new_n11791_), .B1(new_n11779_), .B2(new_n11787_), .ZN(new_n11792_));
  NAND2_X1   g10790(.A1(new_n11783_), .A2(new_n11786_), .ZN(new_n11793_));
  NAND2_X1   g10791(.A1(new_n11778_), .A2(new_n11774_), .ZN(new_n11794_));
  NOR2_X1    g10792(.A1(new_n2703_), .A2(new_n2692_), .ZN(new_n11795_));
  AOI22_X1   g10793(.A1(new_n11795_), .A2(new_n2676_), .B1(new_n2637_), .B2(new_n2647_), .ZN(new_n11796_));
  OAI22_X1   g10794(.A1(new_n11796_), .A2(new_n2727_), .B1(new_n3845_), .B2(new_n3841_), .ZN(new_n11797_));
  INV_X1     g10795(.I(new_n11791_), .ZN(new_n11798_));
  NAND4_X1   g10796(.A1(new_n11797_), .A2(new_n11793_), .A3(new_n11794_), .A4(new_n11798_), .ZN(new_n11799_));
  NAND3_X1   g10797(.A1(new_n11799_), .A2(new_n11792_), .A3(new_n11771_), .ZN(new_n11800_));
  OAI21_X1   g10798(.A1(new_n11768_), .A2(new_n11769_), .B(new_n11760_), .ZN(new_n11801_));
  NAND3_X1   g10799(.A1(new_n11763_), .A2(new_n11764_), .A3(new_n11761_), .ZN(new_n11802_));
  NAND2_X1   g10800(.A1(new_n11801_), .A2(new_n11802_), .ZN(new_n11803_));
  AOI22_X1   g10801(.A1(new_n11797_), .A2(new_n11798_), .B1(new_n11793_), .B2(new_n11794_), .ZN(new_n11804_));
  NOR4_X1    g10802(.A1(new_n11790_), .A2(new_n11779_), .A3(new_n11787_), .A4(new_n11791_), .ZN(new_n11805_));
  OAI21_X1   g10803(.A1(new_n11804_), .A2(new_n11805_), .B(new_n11803_), .ZN(new_n11806_));
  NAND3_X1   g10804(.A1(new_n11759_), .A2(new_n11800_), .A3(new_n11806_), .ZN(new_n11807_));
  OAI21_X1   g10805(.A1(new_n3860_), .A2(new_n3861_), .B(new_n3807_), .ZN(new_n11808_));
  NOR2_X1    g10806(.A1(new_n3860_), .A2(new_n3807_), .ZN(new_n11809_));
  AOI22_X1   g10807(.A1(new_n11808_), .A2(new_n3865_), .B1(new_n11809_), .B2(new_n3855_), .ZN(new_n11810_));
  NAND2_X1   g10808(.A1(new_n11806_), .A2(new_n11800_), .ZN(new_n11811_));
  NAND2_X1   g10809(.A1(new_n11811_), .A2(new_n11810_), .ZN(new_n11812_));
  NAND2_X1   g10810(.A1(new_n11812_), .A2(new_n11807_), .ZN(new_n11813_));
  NAND3_X1   g10811(.A1(new_n11813_), .A2(new_n11752_), .A3(new_n11756_), .ZN(new_n11814_));
  NAND2_X1   g10812(.A1(new_n11752_), .A2(new_n11756_), .ZN(new_n11815_));
  NOR2_X1    g10813(.A1(new_n11811_), .A2(new_n11810_), .ZN(new_n11816_));
  AOI21_X1   g10814(.A1(new_n11800_), .A2(new_n11806_), .B(new_n11759_), .ZN(new_n11817_));
  NOR2_X1    g10815(.A1(new_n11817_), .A2(new_n11816_), .ZN(new_n11818_));
  NAND2_X1   g10816(.A1(new_n11815_), .A2(new_n11818_), .ZN(new_n11819_));
  NOR3_X1    g10817(.A1(new_n3875_), .A2(new_n3784_), .A3(new_n3776_), .ZN(new_n11820_));
  OAI21_X1   g10818(.A1(new_n3776_), .A2(new_n3784_), .B(new_n3875_), .ZN(new_n11821_));
  AOI21_X1   g10819(.A1(new_n11821_), .A2(new_n3881_), .B(new_n11820_), .ZN(new_n11822_));
  NAND3_X1   g10820(.A1(new_n11822_), .A2(new_n11819_), .A3(new_n11814_), .ZN(new_n11823_));
  NOR2_X1    g10821(.A1(new_n11815_), .A2(new_n11818_), .ZN(new_n11824_));
  AOI22_X1   g10822(.A1(new_n11754_), .A2(new_n11755_), .B1(new_n11753_), .B2(new_n11682_), .ZN(new_n11825_));
  OAI21_X1   g10823(.A1(new_n3677_), .A2(new_n11684_), .B(new_n11682_), .ZN(new_n11826_));
  NOR3_X1    g10824(.A1(new_n11826_), .A2(new_n11751_), .A3(new_n11740_), .ZN(new_n11827_));
  NOR2_X1    g10825(.A1(new_n11825_), .A2(new_n11827_), .ZN(new_n11828_));
  NOR2_X1    g10826(.A1(new_n11828_), .A2(new_n11813_), .ZN(new_n11829_));
  NAND3_X1   g10827(.A1(new_n3869_), .A2(new_n3871_), .A3(new_n3872_), .ZN(new_n11830_));
  AOI21_X1   g10828(.A1(new_n3871_), .A2(new_n3872_), .B(new_n3869_), .ZN(new_n11831_));
  OAI21_X1   g10829(.A1(new_n11831_), .A2(new_n3675_), .B(new_n11830_), .ZN(new_n11832_));
  OAI21_X1   g10830(.A1(new_n11824_), .A2(new_n11829_), .B(new_n11832_), .ZN(new_n11833_));
  AOI21_X1   g10831(.A1(new_n11833_), .A2(new_n11823_), .B(new_n11681_), .ZN(new_n11834_));
  AOI21_X1   g10832(.A1(new_n11678_), .A2(new_n11679_), .B(new_n11677_), .ZN(new_n11835_));
  NOR3_X1    g10833(.A1(new_n11619_), .A2(new_n11673_), .A3(new_n11665_), .ZN(new_n11836_));
  NOR2_X1    g10834(.A1(new_n11835_), .A2(new_n11836_), .ZN(new_n11837_));
  NOR3_X1    g10835(.A1(new_n11824_), .A2(new_n11829_), .A3(new_n11832_), .ZN(new_n11838_));
  AOI21_X1   g10836(.A1(new_n11814_), .A2(new_n11819_), .B(new_n11822_), .ZN(new_n11839_));
  NOR3_X1    g10837(.A1(new_n11839_), .A2(new_n11838_), .A3(new_n11837_), .ZN(new_n11840_));
  NAND3_X1   g10838(.A1(new_n3889_), .A2(new_n3890_), .A3(new_n3674_), .ZN(new_n11841_));
  AOI21_X1   g10839(.A1(new_n3889_), .A2(new_n3890_), .B(new_n3674_), .ZN(new_n11842_));
  OAI21_X1   g10840(.A1(new_n3893_), .A2(new_n11842_), .B(new_n11841_), .ZN(new_n11843_));
  NOR3_X1    g10841(.A1(new_n11840_), .A2(new_n11843_), .A3(new_n11834_), .ZN(new_n11844_));
  OAI21_X1   g10842(.A1(new_n11839_), .A2(new_n11838_), .B(new_n11837_), .ZN(new_n11845_));
  NAND3_X1   g10843(.A1(new_n11833_), .A2(new_n11823_), .A3(new_n11681_), .ZN(new_n11846_));
  NOR2_X1    g10844(.A1(new_n3877_), .A2(new_n3888_), .ZN(new_n11847_));
  OAI21_X1   g10845(.A1(new_n3877_), .A2(new_n3884_), .B(new_n3888_), .ZN(new_n11848_));
  AOI22_X1   g10846(.A1(new_n11848_), .A2(new_n3892_), .B1(new_n11847_), .B2(new_n3890_), .ZN(new_n11849_));
  AOI21_X1   g10847(.A1(new_n11845_), .A2(new_n11846_), .B(new_n11849_), .ZN(new_n11850_));
  OAI21_X1   g10848(.A1(new_n11850_), .A2(new_n11844_), .B(new_n11616_), .ZN(new_n11851_));
  OAI21_X1   g10849(.A1(new_n11613_), .A2(new_n11614_), .B(new_n11612_), .ZN(new_n11852_));
  NAND3_X1   g10850(.A1(new_n11464_), .A2(new_n11601_), .A3(new_n11608_), .ZN(new_n11853_));
  NAND2_X1   g10851(.A1(new_n11852_), .A2(new_n11853_), .ZN(new_n11854_));
  NAND3_X1   g10852(.A1(new_n11845_), .A2(new_n11849_), .A3(new_n11846_), .ZN(new_n11855_));
  OAI21_X1   g10853(.A1(new_n11840_), .A2(new_n11834_), .B(new_n11843_), .ZN(new_n11856_));
  NAND3_X1   g10854(.A1(new_n11856_), .A2(new_n11855_), .A3(new_n11854_), .ZN(new_n11857_));
  AOI21_X1   g10855(.A1(new_n11851_), .A2(new_n11857_), .B(new_n11461_), .ZN(new_n11858_));
  AOI21_X1   g10856(.A1(new_n3894_), .A2(new_n3897_), .B(new_n4154_), .ZN(new_n11859_));
  NAND3_X1   g10857(.A1(new_n3894_), .A2(new_n3897_), .A3(new_n4154_), .ZN(new_n11860_));
  OAI21_X1   g10858(.A1(new_n3562_), .A2(new_n11859_), .B(new_n11860_), .ZN(new_n11861_));
  AOI21_X1   g10859(.A1(new_n11856_), .A2(new_n11855_), .B(new_n11854_), .ZN(new_n11862_));
  NOR3_X1    g10860(.A1(new_n11850_), .A2(new_n11844_), .A3(new_n11616_), .ZN(new_n11863_));
  NOR3_X1    g10861(.A1(new_n11863_), .A2(new_n11861_), .A3(new_n11862_), .ZN(new_n11864_));
  NOR2_X1    g10862(.A1(new_n11858_), .A2(new_n11864_), .ZN(new_n11865_));
  OAI21_X1   g10863(.A1(new_n11452_), .A2(new_n11458_), .B(new_n11865_), .ZN(new_n11866_));
  OAI21_X1   g10864(.A1(new_n11456_), .A2(new_n11457_), .B(new_n11455_), .ZN(new_n11867_));
  NAND3_X1   g10865(.A1(new_n10703_), .A2(new_n11451_), .A3(new_n11444_), .ZN(new_n11868_));
  OAI21_X1   g10866(.A1(new_n11863_), .A2(new_n11862_), .B(new_n11861_), .ZN(new_n11869_));
  NAND3_X1   g10867(.A1(new_n11461_), .A2(new_n11851_), .A3(new_n11857_), .ZN(new_n11870_));
  NAND2_X1   g10868(.A1(new_n11869_), .A2(new_n11870_), .ZN(new_n11871_));
  NAND3_X1   g10869(.A1(new_n11868_), .A2(new_n11867_), .A3(new_n11871_), .ZN(new_n11872_));
  AOI22_X1   g10870(.A1(new_n11866_), .A2(new_n11872_), .B1(new_n10700_), .B2(new_n10677_), .ZN(new_n11873_));
  INV_X1     g10871(.I(new_n10695_), .ZN(new_n11874_));
  AOI21_X1   g10872(.A1(new_n10670_), .A2(new_n10676_), .B(new_n4171_), .ZN(new_n11875_));
  OAI21_X1   g10873(.A1(new_n11874_), .A2(new_n11875_), .B(new_n10677_), .ZN(new_n11876_));
  AOI21_X1   g10874(.A1(new_n11868_), .A2(new_n11867_), .B(new_n11871_), .ZN(new_n11877_));
  NOR3_X1    g10875(.A1(new_n11452_), .A2(new_n11458_), .A3(new_n11865_), .ZN(new_n11878_));
  NOR3_X1    g10876(.A1(new_n11876_), .A2(new_n11877_), .A3(new_n11878_), .ZN(new_n11879_));
  INV_X1     g10877(.I(\A[471] ), .ZN(new_n11880_));
  INV_X1     g10878(.I(\A[469] ), .ZN(new_n11881_));
  NAND2_X1   g10879(.A1(new_n11881_), .A2(\A[470] ), .ZN(new_n11882_));
  NOR2_X1    g10880(.A1(new_n11881_), .A2(\A[470] ), .ZN(new_n11883_));
  NOR2_X1    g10881(.A1(new_n11883_), .A2(new_n11880_), .ZN(new_n11884_));
  INV_X1     g10882(.I(\A[470] ), .ZN(new_n11885_));
  NAND2_X1   g10883(.A1(new_n11885_), .A2(\A[469] ), .ZN(new_n11886_));
  NAND2_X1   g10884(.A1(new_n11882_), .A2(new_n11886_), .ZN(new_n11887_));
  AOI22_X1   g10885(.A1(new_n11887_), .A2(new_n11880_), .B1(new_n11884_), .B2(new_n11882_), .ZN(new_n11888_));
  INV_X1     g10886(.I(\A[474] ), .ZN(new_n11889_));
  INV_X1     g10887(.I(\A[472] ), .ZN(new_n11890_));
  NAND2_X1   g10888(.A1(new_n11890_), .A2(\A[473] ), .ZN(new_n11891_));
  NOR2_X1    g10889(.A1(new_n11890_), .A2(\A[473] ), .ZN(new_n11892_));
  NOR2_X1    g10890(.A1(new_n11892_), .A2(new_n11889_), .ZN(new_n11893_));
  INV_X1     g10891(.I(\A[473] ), .ZN(new_n11894_));
  NAND2_X1   g10892(.A1(new_n11894_), .A2(\A[472] ), .ZN(new_n11895_));
  NAND2_X1   g10893(.A1(new_n11891_), .A2(new_n11895_), .ZN(new_n11896_));
  AOI22_X1   g10894(.A1(new_n11896_), .A2(new_n11889_), .B1(new_n11893_), .B2(new_n11891_), .ZN(new_n11897_));
  XOR2_X1    g10895(.A1(new_n11888_), .A2(new_n11897_), .Z(new_n11898_));
  NOR2_X1    g10896(.A1(new_n11894_), .A2(\A[472] ), .ZN(new_n11899_));
  NOR2_X1    g10897(.A1(new_n11899_), .A2(new_n11892_), .ZN(new_n11900_));
  NOR2_X1    g10898(.A1(new_n11890_), .A2(new_n11894_), .ZN(new_n11901_));
  INV_X1     g10899(.I(new_n11901_), .ZN(new_n11902_));
  OAI21_X1   g10900(.A1(new_n11900_), .A2(new_n11889_), .B(new_n11902_), .ZN(new_n11903_));
  NOR2_X1    g10901(.A1(new_n11881_), .A2(new_n11885_), .ZN(new_n11904_));
  AOI21_X1   g10902(.A1(new_n11887_), .A2(\A[471] ), .B(new_n11904_), .ZN(new_n11905_));
  INV_X1     g10903(.I(new_n11905_), .ZN(new_n11906_));
  NOR2_X1    g10904(.A1(new_n11888_), .A2(new_n11897_), .ZN(new_n11907_));
  NAND3_X1   g10905(.A1(new_n11907_), .A2(new_n11903_), .A3(new_n11906_), .ZN(new_n11908_));
  NAND2_X1   g10906(.A1(new_n11898_), .A2(new_n11908_), .ZN(new_n11909_));
  INV_X1     g10907(.I(\A[467] ), .ZN(new_n11910_));
  NOR2_X1    g10908(.A1(new_n11910_), .A2(\A[466] ), .ZN(new_n11911_));
  NAND2_X1   g10909(.A1(new_n11910_), .A2(\A[466] ), .ZN(new_n11912_));
  NAND2_X1   g10910(.A1(new_n11912_), .A2(\A[468] ), .ZN(new_n11913_));
  INV_X1     g10911(.I(\A[466] ), .ZN(new_n11914_));
  NOR2_X1    g10912(.A1(new_n11914_), .A2(\A[467] ), .ZN(new_n11915_));
  NOR2_X1    g10913(.A1(new_n11911_), .A2(new_n11915_), .ZN(new_n11916_));
  OAI22_X1   g10914(.A1(new_n11916_), .A2(\A[468] ), .B1(new_n11913_), .B2(new_n11911_), .ZN(new_n11917_));
  INV_X1     g10915(.I(\A[465] ), .ZN(new_n11918_));
  INV_X1     g10916(.I(\A[463] ), .ZN(new_n11919_));
  NAND2_X1   g10917(.A1(new_n11919_), .A2(\A[464] ), .ZN(new_n11920_));
  NOR2_X1    g10918(.A1(new_n11919_), .A2(\A[464] ), .ZN(new_n11921_));
  NOR2_X1    g10919(.A1(new_n11921_), .A2(new_n11918_), .ZN(new_n11922_));
  INV_X1     g10920(.I(\A[464] ), .ZN(new_n11923_));
  NAND2_X1   g10921(.A1(new_n11923_), .A2(\A[463] ), .ZN(new_n11924_));
  NAND2_X1   g10922(.A1(new_n11920_), .A2(new_n11924_), .ZN(new_n11925_));
  AOI22_X1   g10923(.A1(new_n11925_), .A2(new_n11918_), .B1(new_n11922_), .B2(new_n11920_), .ZN(new_n11926_));
  XNOR2_X1   g10924(.A1(new_n11926_), .A2(new_n11917_), .ZN(new_n11927_));
  INV_X1     g10925(.I(\A[468] ), .ZN(new_n11928_));
  NOR2_X1    g10926(.A1(new_n11914_), .A2(new_n11910_), .ZN(new_n11929_));
  INV_X1     g10927(.I(new_n11929_), .ZN(new_n11930_));
  OAI21_X1   g10928(.A1(new_n11916_), .A2(new_n11928_), .B(new_n11930_), .ZN(new_n11931_));
  NOR2_X1    g10929(.A1(new_n11919_), .A2(new_n11923_), .ZN(new_n11932_));
  AOI21_X1   g10930(.A1(new_n11925_), .A2(\A[465] ), .B(new_n11932_), .ZN(new_n11933_));
  INV_X1     g10931(.I(new_n11933_), .ZN(new_n11934_));
  INV_X1     g10932(.I(new_n11917_), .ZN(new_n11935_));
  NOR2_X1    g10933(.A1(new_n11935_), .A2(new_n11926_), .ZN(new_n11936_));
  NAND3_X1   g10934(.A1(new_n11936_), .A2(new_n11931_), .A3(new_n11934_), .ZN(new_n11937_));
  NAND2_X1   g10935(.A1(new_n11937_), .A2(new_n11927_), .ZN(new_n11938_));
  XOR2_X1    g10936(.A1(new_n11938_), .A2(new_n11909_), .Z(new_n11939_));
  INV_X1     g10937(.I(\A[482] ), .ZN(new_n11940_));
  NOR2_X1    g10938(.A1(new_n11940_), .A2(\A[481] ), .ZN(new_n11941_));
  NAND2_X1   g10939(.A1(new_n11940_), .A2(\A[481] ), .ZN(new_n11942_));
  NAND2_X1   g10940(.A1(new_n11942_), .A2(\A[483] ), .ZN(new_n11943_));
  INV_X1     g10941(.I(\A[481] ), .ZN(new_n11944_));
  NOR2_X1    g10942(.A1(new_n11944_), .A2(\A[482] ), .ZN(new_n11945_));
  NOR2_X1    g10943(.A1(new_n11941_), .A2(new_n11945_), .ZN(new_n11946_));
  OAI22_X1   g10944(.A1(new_n11946_), .A2(\A[483] ), .B1(new_n11943_), .B2(new_n11941_), .ZN(new_n11947_));
  INV_X1     g10945(.I(\A[486] ), .ZN(new_n11948_));
  INV_X1     g10946(.I(\A[484] ), .ZN(new_n11949_));
  NAND2_X1   g10947(.A1(new_n11949_), .A2(\A[485] ), .ZN(new_n11950_));
  NOR2_X1    g10948(.A1(new_n11949_), .A2(\A[485] ), .ZN(new_n11951_));
  NOR2_X1    g10949(.A1(new_n11951_), .A2(new_n11948_), .ZN(new_n11952_));
  INV_X1     g10950(.I(\A[485] ), .ZN(new_n11953_));
  NAND2_X1   g10951(.A1(new_n11953_), .A2(\A[484] ), .ZN(new_n11954_));
  NAND2_X1   g10952(.A1(new_n11950_), .A2(new_n11954_), .ZN(new_n11955_));
  AOI22_X1   g10953(.A1(new_n11955_), .A2(new_n11948_), .B1(new_n11952_), .B2(new_n11950_), .ZN(new_n11956_));
  XNOR2_X1   g10954(.A1(new_n11956_), .A2(new_n11947_), .ZN(new_n11957_));
  NOR2_X1    g10955(.A1(new_n11953_), .A2(\A[484] ), .ZN(new_n11958_));
  NOR2_X1    g10956(.A1(new_n11958_), .A2(new_n11951_), .ZN(new_n11959_));
  NOR2_X1    g10957(.A1(new_n11949_), .A2(new_n11953_), .ZN(new_n11960_));
  INV_X1     g10958(.I(new_n11960_), .ZN(new_n11961_));
  OAI21_X1   g10959(.A1(new_n11959_), .A2(new_n11948_), .B(new_n11961_), .ZN(new_n11962_));
  NAND2_X1   g10960(.A1(new_n11944_), .A2(\A[482] ), .ZN(new_n11963_));
  NAND2_X1   g10961(.A1(new_n11963_), .A2(new_n11942_), .ZN(new_n11964_));
  NOR2_X1    g10962(.A1(new_n11944_), .A2(new_n11940_), .ZN(new_n11965_));
  AOI21_X1   g10963(.A1(new_n11964_), .A2(\A[483] ), .B(new_n11965_), .ZN(new_n11966_));
  INV_X1     g10964(.I(new_n11966_), .ZN(new_n11967_));
  INV_X1     g10965(.I(new_n11947_), .ZN(new_n11968_));
  NOR2_X1    g10966(.A1(new_n11968_), .A2(new_n11956_), .ZN(new_n11969_));
  NAND3_X1   g10967(.A1(new_n11969_), .A2(new_n11962_), .A3(new_n11967_), .ZN(new_n11970_));
  NAND2_X1   g10968(.A1(new_n11970_), .A2(new_n11957_), .ZN(new_n11971_));
  INV_X1     g10969(.I(\A[476] ), .ZN(new_n11972_));
  NOR2_X1    g10970(.A1(new_n11972_), .A2(\A[475] ), .ZN(new_n11973_));
  NAND2_X1   g10971(.A1(new_n11972_), .A2(\A[475] ), .ZN(new_n11974_));
  NAND2_X1   g10972(.A1(new_n11974_), .A2(\A[477] ), .ZN(new_n11975_));
  INV_X1     g10973(.I(\A[475] ), .ZN(new_n11976_));
  NOR2_X1    g10974(.A1(new_n11976_), .A2(\A[476] ), .ZN(new_n11977_));
  NOR2_X1    g10975(.A1(new_n11973_), .A2(new_n11977_), .ZN(new_n11978_));
  OAI22_X1   g10976(.A1(new_n11978_), .A2(\A[477] ), .B1(new_n11975_), .B2(new_n11973_), .ZN(new_n11979_));
  INV_X1     g10977(.I(\A[480] ), .ZN(new_n11980_));
  INV_X1     g10978(.I(\A[478] ), .ZN(new_n11981_));
  NAND2_X1   g10979(.A1(new_n11981_), .A2(\A[479] ), .ZN(new_n11982_));
  NOR2_X1    g10980(.A1(new_n11981_), .A2(\A[479] ), .ZN(new_n11983_));
  NOR2_X1    g10981(.A1(new_n11983_), .A2(new_n11980_), .ZN(new_n11984_));
  INV_X1     g10982(.I(\A[479] ), .ZN(new_n11985_));
  NAND2_X1   g10983(.A1(new_n11985_), .A2(\A[478] ), .ZN(new_n11986_));
  NAND2_X1   g10984(.A1(new_n11982_), .A2(new_n11986_), .ZN(new_n11987_));
  AOI22_X1   g10985(.A1(new_n11987_), .A2(new_n11980_), .B1(new_n11984_), .B2(new_n11982_), .ZN(new_n11988_));
  XNOR2_X1   g10986(.A1(new_n11988_), .A2(new_n11979_), .ZN(new_n11989_));
  INV_X1     g10987(.I(new_n11982_), .ZN(new_n11990_));
  NOR2_X1    g10988(.A1(new_n11990_), .A2(new_n11983_), .ZN(new_n11991_));
  NOR2_X1    g10989(.A1(new_n11981_), .A2(new_n11985_), .ZN(new_n11992_));
  INV_X1     g10990(.I(new_n11992_), .ZN(new_n11993_));
  OAI21_X1   g10991(.A1(new_n11991_), .A2(new_n11980_), .B(new_n11993_), .ZN(new_n11994_));
  NAND2_X1   g10992(.A1(new_n11976_), .A2(\A[476] ), .ZN(new_n11995_));
  NAND2_X1   g10993(.A1(new_n11995_), .A2(new_n11974_), .ZN(new_n11996_));
  NOR2_X1    g10994(.A1(new_n11976_), .A2(new_n11972_), .ZN(new_n11997_));
  AOI21_X1   g10995(.A1(new_n11996_), .A2(\A[477] ), .B(new_n11997_), .ZN(new_n11998_));
  INV_X1     g10996(.I(new_n11998_), .ZN(new_n11999_));
  INV_X1     g10997(.I(new_n11979_), .ZN(new_n12000_));
  NOR2_X1    g10998(.A1(new_n12000_), .A2(new_n11988_), .ZN(new_n12001_));
  NAND3_X1   g10999(.A1(new_n12001_), .A2(new_n11994_), .A3(new_n11999_), .ZN(new_n12002_));
  NAND2_X1   g11000(.A1(new_n12002_), .A2(new_n11989_), .ZN(new_n12003_));
  XOR2_X1    g11001(.A1(new_n11971_), .A2(new_n12003_), .Z(new_n12004_));
  XOR2_X1    g11002(.A1(new_n12004_), .A2(new_n11939_), .Z(new_n12005_));
  INV_X1     g11003(.I(\A[506] ), .ZN(new_n12006_));
  NOR2_X1    g11004(.A1(new_n12006_), .A2(\A[505] ), .ZN(new_n12007_));
  NAND2_X1   g11005(.A1(new_n12006_), .A2(\A[505] ), .ZN(new_n12008_));
  NAND2_X1   g11006(.A1(new_n12008_), .A2(\A[507] ), .ZN(new_n12009_));
  INV_X1     g11007(.I(\A[505] ), .ZN(new_n12010_));
  NOR2_X1    g11008(.A1(new_n12010_), .A2(\A[506] ), .ZN(new_n12011_));
  NOR2_X1    g11009(.A1(new_n12007_), .A2(new_n12011_), .ZN(new_n12012_));
  OAI22_X1   g11010(.A1(new_n12012_), .A2(\A[507] ), .B1(new_n12009_), .B2(new_n12007_), .ZN(new_n12013_));
  INV_X1     g11011(.I(\A[510] ), .ZN(new_n12014_));
  INV_X1     g11012(.I(\A[508] ), .ZN(new_n12015_));
  NAND2_X1   g11013(.A1(new_n12015_), .A2(\A[509] ), .ZN(new_n12016_));
  NOR2_X1    g11014(.A1(new_n12015_), .A2(\A[509] ), .ZN(new_n12017_));
  NOR2_X1    g11015(.A1(new_n12017_), .A2(new_n12014_), .ZN(new_n12018_));
  INV_X1     g11016(.I(\A[509] ), .ZN(new_n12019_));
  NAND2_X1   g11017(.A1(new_n12019_), .A2(\A[508] ), .ZN(new_n12020_));
  NAND2_X1   g11018(.A1(new_n12016_), .A2(new_n12020_), .ZN(new_n12021_));
  AOI22_X1   g11019(.A1(new_n12021_), .A2(new_n12014_), .B1(new_n12018_), .B2(new_n12016_), .ZN(new_n12022_));
  XNOR2_X1   g11020(.A1(new_n12022_), .A2(new_n12013_), .ZN(new_n12023_));
  NOR2_X1    g11021(.A1(new_n12019_), .A2(\A[508] ), .ZN(new_n12024_));
  NOR2_X1    g11022(.A1(new_n12024_), .A2(new_n12017_), .ZN(new_n12025_));
  NOR2_X1    g11023(.A1(new_n12015_), .A2(new_n12019_), .ZN(new_n12026_));
  INV_X1     g11024(.I(new_n12026_), .ZN(new_n12027_));
  OAI21_X1   g11025(.A1(new_n12025_), .A2(new_n12014_), .B(new_n12027_), .ZN(new_n12028_));
  NAND2_X1   g11026(.A1(new_n12010_), .A2(\A[506] ), .ZN(new_n12029_));
  NAND2_X1   g11027(.A1(new_n12029_), .A2(new_n12008_), .ZN(new_n12030_));
  NOR2_X1    g11028(.A1(new_n12010_), .A2(new_n12006_), .ZN(new_n12031_));
  AOI21_X1   g11029(.A1(new_n12030_), .A2(\A[507] ), .B(new_n12031_), .ZN(new_n12032_));
  INV_X1     g11030(.I(new_n12032_), .ZN(new_n12033_));
  INV_X1     g11031(.I(new_n12013_), .ZN(new_n12034_));
  NOR2_X1    g11032(.A1(new_n12034_), .A2(new_n12022_), .ZN(new_n12035_));
  NAND3_X1   g11033(.A1(new_n12035_), .A2(new_n12028_), .A3(new_n12033_), .ZN(new_n12036_));
  NAND2_X1   g11034(.A1(new_n12036_), .A2(new_n12023_), .ZN(new_n12037_));
  INV_X1     g11035(.I(\A[500] ), .ZN(new_n12038_));
  NOR2_X1    g11036(.A1(new_n12038_), .A2(\A[499] ), .ZN(new_n12039_));
  NAND2_X1   g11037(.A1(new_n12038_), .A2(\A[499] ), .ZN(new_n12040_));
  NAND2_X1   g11038(.A1(new_n12040_), .A2(\A[501] ), .ZN(new_n12041_));
  INV_X1     g11039(.I(\A[499] ), .ZN(new_n12042_));
  NOR2_X1    g11040(.A1(new_n12042_), .A2(\A[500] ), .ZN(new_n12043_));
  NOR2_X1    g11041(.A1(new_n12039_), .A2(new_n12043_), .ZN(new_n12044_));
  OAI22_X1   g11042(.A1(new_n12044_), .A2(\A[501] ), .B1(new_n12041_), .B2(new_n12039_), .ZN(new_n12045_));
  INV_X1     g11043(.I(\A[504] ), .ZN(new_n12046_));
  INV_X1     g11044(.I(\A[502] ), .ZN(new_n12047_));
  NAND2_X1   g11045(.A1(new_n12047_), .A2(\A[503] ), .ZN(new_n12048_));
  NOR2_X1    g11046(.A1(new_n12047_), .A2(\A[503] ), .ZN(new_n12049_));
  NOR2_X1    g11047(.A1(new_n12049_), .A2(new_n12046_), .ZN(new_n12050_));
  INV_X1     g11048(.I(\A[503] ), .ZN(new_n12051_));
  NAND2_X1   g11049(.A1(new_n12051_), .A2(\A[502] ), .ZN(new_n12052_));
  NAND2_X1   g11050(.A1(new_n12048_), .A2(new_n12052_), .ZN(new_n12053_));
  AOI22_X1   g11051(.A1(new_n12053_), .A2(new_n12046_), .B1(new_n12050_), .B2(new_n12048_), .ZN(new_n12054_));
  XNOR2_X1   g11052(.A1(new_n12054_), .A2(new_n12045_), .ZN(new_n12055_));
  NOR2_X1    g11053(.A1(new_n12051_), .A2(\A[502] ), .ZN(new_n12056_));
  NOR2_X1    g11054(.A1(new_n12056_), .A2(new_n12049_), .ZN(new_n12057_));
  NOR2_X1    g11055(.A1(new_n12047_), .A2(new_n12051_), .ZN(new_n12058_));
  INV_X1     g11056(.I(new_n12058_), .ZN(new_n12059_));
  OAI21_X1   g11057(.A1(new_n12057_), .A2(new_n12046_), .B(new_n12059_), .ZN(new_n12060_));
  NAND2_X1   g11058(.A1(new_n12042_), .A2(\A[500] ), .ZN(new_n12061_));
  NAND2_X1   g11059(.A1(new_n12061_), .A2(new_n12040_), .ZN(new_n12062_));
  NOR2_X1    g11060(.A1(new_n12042_), .A2(new_n12038_), .ZN(new_n12063_));
  AOI21_X1   g11061(.A1(new_n12062_), .A2(\A[501] ), .B(new_n12063_), .ZN(new_n12064_));
  INV_X1     g11062(.I(new_n12064_), .ZN(new_n12065_));
  INV_X1     g11063(.I(new_n12045_), .ZN(new_n12066_));
  NOR2_X1    g11064(.A1(new_n12066_), .A2(new_n12054_), .ZN(new_n12067_));
  NAND3_X1   g11065(.A1(new_n12067_), .A2(new_n12060_), .A3(new_n12065_), .ZN(new_n12068_));
  NAND2_X1   g11066(.A1(new_n12068_), .A2(new_n12055_), .ZN(new_n12069_));
  XOR2_X1    g11067(.A1(new_n12037_), .A2(new_n12069_), .Z(new_n12070_));
  INV_X1     g11068(.I(\A[495] ), .ZN(new_n12071_));
  INV_X1     g11069(.I(\A[493] ), .ZN(new_n12072_));
  NAND2_X1   g11070(.A1(new_n12072_), .A2(\A[494] ), .ZN(new_n12073_));
  NOR2_X1    g11071(.A1(new_n12072_), .A2(\A[494] ), .ZN(new_n12074_));
  NOR2_X1    g11072(.A1(new_n12074_), .A2(new_n12071_), .ZN(new_n12075_));
  INV_X1     g11073(.I(\A[494] ), .ZN(new_n12076_));
  NAND2_X1   g11074(.A1(new_n12076_), .A2(\A[493] ), .ZN(new_n12077_));
  NAND2_X1   g11075(.A1(new_n12073_), .A2(new_n12077_), .ZN(new_n12078_));
  AOI22_X1   g11076(.A1(new_n12078_), .A2(new_n12071_), .B1(new_n12075_), .B2(new_n12073_), .ZN(new_n12079_));
  INV_X1     g11077(.I(\A[498] ), .ZN(new_n12080_));
  INV_X1     g11078(.I(\A[496] ), .ZN(new_n12081_));
  NAND2_X1   g11079(.A1(new_n12081_), .A2(\A[497] ), .ZN(new_n12082_));
  NOR2_X1    g11080(.A1(new_n12081_), .A2(\A[497] ), .ZN(new_n12083_));
  NOR2_X1    g11081(.A1(new_n12083_), .A2(new_n12080_), .ZN(new_n12084_));
  INV_X1     g11082(.I(\A[497] ), .ZN(new_n12085_));
  NAND2_X1   g11083(.A1(new_n12085_), .A2(\A[496] ), .ZN(new_n12086_));
  NAND2_X1   g11084(.A1(new_n12082_), .A2(new_n12086_), .ZN(new_n12087_));
  AOI22_X1   g11085(.A1(new_n12087_), .A2(new_n12080_), .B1(new_n12084_), .B2(new_n12082_), .ZN(new_n12088_));
  XOR2_X1    g11086(.A1(new_n12079_), .A2(new_n12088_), .Z(new_n12089_));
  NOR2_X1    g11087(.A1(new_n12085_), .A2(\A[496] ), .ZN(new_n12090_));
  NOR2_X1    g11088(.A1(new_n12090_), .A2(new_n12083_), .ZN(new_n12091_));
  NOR2_X1    g11089(.A1(new_n12081_), .A2(new_n12085_), .ZN(new_n12092_));
  INV_X1     g11090(.I(new_n12092_), .ZN(new_n12093_));
  OAI21_X1   g11091(.A1(new_n12091_), .A2(new_n12080_), .B(new_n12093_), .ZN(new_n12094_));
  NOR2_X1    g11092(.A1(new_n12072_), .A2(new_n12076_), .ZN(new_n12095_));
  AOI21_X1   g11093(.A1(new_n12078_), .A2(\A[495] ), .B(new_n12095_), .ZN(new_n12096_));
  INV_X1     g11094(.I(new_n12096_), .ZN(new_n12097_));
  NOR2_X1    g11095(.A1(new_n12079_), .A2(new_n12088_), .ZN(new_n12098_));
  NAND3_X1   g11096(.A1(new_n12098_), .A2(new_n12094_), .A3(new_n12097_), .ZN(new_n12099_));
  NAND2_X1   g11097(.A1(new_n12089_), .A2(new_n12099_), .ZN(new_n12100_));
  INV_X1     g11098(.I(\A[489] ), .ZN(new_n12101_));
  INV_X1     g11099(.I(\A[487] ), .ZN(new_n12102_));
  NAND2_X1   g11100(.A1(new_n12102_), .A2(\A[488] ), .ZN(new_n12103_));
  NOR2_X1    g11101(.A1(new_n12102_), .A2(\A[488] ), .ZN(new_n12104_));
  NOR2_X1    g11102(.A1(new_n12104_), .A2(new_n12101_), .ZN(new_n12105_));
  INV_X1     g11103(.I(\A[488] ), .ZN(new_n12106_));
  NAND2_X1   g11104(.A1(new_n12106_), .A2(\A[487] ), .ZN(new_n12107_));
  NAND2_X1   g11105(.A1(new_n12103_), .A2(new_n12107_), .ZN(new_n12108_));
  AOI22_X1   g11106(.A1(new_n12108_), .A2(new_n12101_), .B1(new_n12105_), .B2(new_n12103_), .ZN(new_n12109_));
  INV_X1     g11107(.I(\A[492] ), .ZN(new_n12110_));
  INV_X1     g11108(.I(\A[490] ), .ZN(new_n12111_));
  NAND2_X1   g11109(.A1(new_n12111_), .A2(\A[491] ), .ZN(new_n12112_));
  NOR2_X1    g11110(.A1(new_n12111_), .A2(\A[491] ), .ZN(new_n12113_));
  NOR2_X1    g11111(.A1(new_n12113_), .A2(new_n12110_), .ZN(new_n12114_));
  INV_X1     g11112(.I(\A[491] ), .ZN(new_n12115_));
  NAND2_X1   g11113(.A1(new_n12115_), .A2(\A[490] ), .ZN(new_n12116_));
  NAND2_X1   g11114(.A1(new_n12112_), .A2(new_n12116_), .ZN(new_n12117_));
  AOI22_X1   g11115(.A1(new_n12117_), .A2(new_n12110_), .B1(new_n12114_), .B2(new_n12112_), .ZN(new_n12118_));
  XOR2_X1    g11116(.A1(new_n12109_), .A2(new_n12118_), .Z(new_n12119_));
  NOR2_X1    g11117(.A1(new_n12115_), .A2(\A[490] ), .ZN(new_n12120_));
  NOR2_X1    g11118(.A1(new_n12120_), .A2(new_n12113_), .ZN(new_n12121_));
  NOR2_X1    g11119(.A1(new_n12111_), .A2(new_n12115_), .ZN(new_n12122_));
  INV_X1     g11120(.I(new_n12122_), .ZN(new_n12123_));
  OAI21_X1   g11121(.A1(new_n12121_), .A2(new_n12110_), .B(new_n12123_), .ZN(new_n12124_));
  NOR2_X1    g11122(.A1(new_n12102_), .A2(new_n12106_), .ZN(new_n12125_));
  AOI21_X1   g11123(.A1(new_n12108_), .A2(\A[489] ), .B(new_n12125_), .ZN(new_n12126_));
  INV_X1     g11124(.I(new_n12126_), .ZN(new_n12127_));
  NOR2_X1    g11125(.A1(new_n12109_), .A2(new_n12118_), .ZN(new_n12128_));
  NAND3_X1   g11126(.A1(new_n12128_), .A2(new_n12124_), .A3(new_n12127_), .ZN(new_n12129_));
  NAND2_X1   g11127(.A1(new_n12119_), .A2(new_n12129_), .ZN(new_n12130_));
  XOR2_X1    g11128(.A1(new_n12100_), .A2(new_n12130_), .Z(new_n12131_));
  XOR2_X1    g11129(.A1(new_n12070_), .A2(new_n12131_), .Z(new_n12132_));
  XOR2_X1    g11130(.A1(new_n12005_), .A2(new_n12132_), .Z(new_n12133_));
  INV_X1     g11131(.I(\A[554] ), .ZN(new_n12134_));
  NOR2_X1    g11132(.A1(new_n12134_), .A2(\A[553] ), .ZN(new_n12135_));
  NAND2_X1   g11133(.A1(new_n12134_), .A2(\A[553] ), .ZN(new_n12136_));
  NAND2_X1   g11134(.A1(new_n12136_), .A2(\A[555] ), .ZN(new_n12137_));
  INV_X1     g11135(.I(\A[553] ), .ZN(new_n12138_));
  NOR2_X1    g11136(.A1(new_n12138_), .A2(\A[554] ), .ZN(new_n12139_));
  NOR2_X1    g11137(.A1(new_n12135_), .A2(new_n12139_), .ZN(new_n12140_));
  OAI22_X1   g11138(.A1(new_n12140_), .A2(\A[555] ), .B1(new_n12137_), .B2(new_n12135_), .ZN(new_n12141_));
  INV_X1     g11139(.I(\A[558] ), .ZN(new_n12142_));
  INV_X1     g11140(.I(\A[556] ), .ZN(new_n12143_));
  NAND2_X1   g11141(.A1(new_n12143_), .A2(\A[557] ), .ZN(new_n12144_));
  NOR2_X1    g11142(.A1(new_n12143_), .A2(\A[557] ), .ZN(new_n12145_));
  NOR2_X1    g11143(.A1(new_n12145_), .A2(new_n12142_), .ZN(new_n12146_));
  INV_X1     g11144(.I(\A[557] ), .ZN(new_n12147_));
  NAND2_X1   g11145(.A1(new_n12147_), .A2(\A[556] ), .ZN(new_n12148_));
  NAND2_X1   g11146(.A1(new_n12144_), .A2(new_n12148_), .ZN(new_n12149_));
  AOI22_X1   g11147(.A1(new_n12149_), .A2(new_n12142_), .B1(new_n12146_), .B2(new_n12144_), .ZN(new_n12150_));
  XNOR2_X1   g11148(.A1(new_n12150_), .A2(new_n12141_), .ZN(new_n12151_));
  NOR2_X1    g11149(.A1(new_n12147_), .A2(\A[556] ), .ZN(new_n12152_));
  NOR2_X1    g11150(.A1(new_n12152_), .A2(new_n12145_), .ZN(new_n12153_));
  NOR2_X1    g11151(.A1(new_n12143_), .A2(new_n12147_), .ZN(new_n12154_));
  INV_X1     g11152(.I(new_n12154_), .ZN(new_n12155_));
  OAI21_X1   g11153(.A1(new_n12153_), .A2(new_n12142_), .B(new_n12155_), .ZN(new_n12156_));
  NAND2_X1   g11154(.A1(new_n12138_), .A2(\A[554] ), .ZN(new_n12157_));
  NAND2_X1   g11155(.A1(new_n12157_), .A2(new_n12136_), .ZN(new_n12158_));
  NOR2_X1    g11156(.A1(new_n12138_), .A2(new_n12134_), .ZN(new_n12159_));
  AOI21_X1   g11157(.A1(new_n12158_), .A2(\A[555] ), .B(new_n12159_), .ZN(new_n12160_));
  INV_X1     g11158(.I(new_n12160_), .ZN(new_n12161_));
  INV_X1     g11159(.I(new_n12141_), .ZN(new_n12162_));
  NOR2_X1    g11160(.A1(new_n12162_), .A2(new_n12150_), .ZN(new_n12163_));
  NAND3_X1   g11161(.A1(new_n12163_), .A2(new_n12156_), .A3(new_n12161_), .ZN(new_n12164_));
  NAND2_X1   g11162(.A1(new_n12164_), .A2(new_n12151_), .ZN(new_n12165_));
  INV_X1     g11163(.I(\A[548] ), .ZN(new_n12166_));
  NOR2_X1    g11164(.A1(new_n12166_), .A2(\A[547] ), .ZN(new_n12167_));
  NAND2_X1   g11165(.A1(new_n12166_), .A2(\A[547] ), .ZN(new_n12168_));
  NAND2_X1   g11166(.A1(new_n12168_), .A2(\A[549] ), .ZN(new_n12169_));
  INV_X1     g11167(.I(\A[547] ), .ZN(new_n12170_));
  NOR2_X1    g11168(.A1(new_n12170_), .A2(\A[548] ), .ZN(new_n12171_));
  NOR2_X1    g11169(.A1(new_n12167_), .A2(new_n12171_), .ZN(new_n12172_));
  OAI22_X1   g11170(.A1(new_n12172_), .A2(\A[549] ), .B1(new_n12169_), .B2(new_n12167_), .ZN(new_n12173_));
  INV_X1     g11171(.I(\A[552] ), .ZN(new_n12174_));
  INV_X1     g11172(.I(\A[550] ), .ZN(new_n12175_));
  NAND2_X1   g11173(.A1(new_n12175_), .A2(\A[551] ), .ZN(new_n12176_));
  NOR2_X1    g11174(.A1(new_n12175_), .A2(\A[551] ), .ZN(new_n12177_));
  NOR2_X1    g11175(.A1(new_n12177_), .A2(new_n12174_), .ZN(new_n12178_));
  INV_X1     g11176(.I(\A[551] ), .ZN(new_n12179_));
  NAND2_X1   g11177(.A1(new_n12179_), .A2(\A[550] ), .ZN(new_n12180_));
  NAND2_X1   g11178(.A1(new_n12176_), .A2(new_n12180_), .ZN(new_n12181_));
  AOI22_X1   g11179(.A1(new_n12181_), .A2(new_n12174_), .B1(new_n12178_), .B2(new_n12176_), .ZN(new_n12182_));
  XNOR2_X1   g11180(.A1(new_n12182_), .A2(new_n12173_), .ZN(new_n12183_));
  NOR2_X1    g11181(.A1(new_n12179_), .A2(\A[550] ), .ZN(new_n12184_));
  NOR2_X1    g11182(.A1(new_n12184_), .A2(new_n12177_), .ZN(new_n12185_));
  NOR2_X1    g11183(.A1(new_n12175_), .A2(new_n12179_), .ZN(new_n12186_));
  INV_X1     g11184(.I(new_n12186_), .ZN(new_n12187_));
  OAI21_X1   g11185(.A1(new_n12185_), .A2(new_n12174_), .B(new_n12187_), .ZN(new_n12188_));
  NAND2_X1   g11186(.A1(new_n12170_), .A2(\A[548] ), .ZN(new_n12189_));
  NAND2_X1   g11187(.A1(new_n12189_), .A2(new_n12168_), .ZN(new_n12190_));
  NOR2_X1    g11188(.A1(new_n12170_), .A2(new_n12166_), .ZN(new_n12191_));
  AOI21_X1   g11189(.A1(new_n12190_), .A2(\A[549] ), .B(new_n12191_), .ZN(new_n12192_));
  INV_X1     g11190(.I(new_n12192_), .ZN(new_n12193_));
  INV_X1     g11191(.I(new_n12173_), .ZN(new_n12194_));
  NOR2_X1    g11192(.A1(new_n12194_), .A2(new_n12182_), .ZN(new_n12195_));
  NAND3_X1   g11193(.A1(new_n12195_), .A2(new_n12188_), .A3(new_n12193_), .ZN(new_n12196_));
  NAND2_X1   g11194(.A1(new_n12196_), .A2(new_n12183_), .ZN(new_n12197_));
  XOR2_X1    g11195(.A1(new_n12165_), .A2(new_n12197_), .Z(new_n12198_));
  INV_X1     g11196(.I(\A[542] ), .ZN(new_n12199_));
  NOR2_X1    g11197(.A1(new_n12199_), .A2(\A[541] ), .ZN(new_n12200_));
  NAND2_X1   g11198(.A1(new_n12199_), .A2(\A[541] ), .ZN(new_n12201_));
  NAND2_X1   g11199(.A1(new_n12201_), .A2(\A[543] ), .ZN(new_n12202_));
  INV_X1     g11200(.I(\A[541] ), .ZN(new_n12203_));
  NOR2_X1    g11201(.A1(new_n12203_), .A2(\A[542] ), .ZN(new_n12204_));
  NOR2_X1    g11202(.A1(new_n12200_), .A2(new_n12204_), .ZN(new_n12205_));
  OAI22_X1   g11203(.A1(new_n12205_), .A2(\A[543] ), .B1(new_n12202_), .B2(new_n12200_), .ZN(new_n12206_));
  INV_X1     g11204(.I(\A[546] ), .ZN(new_n12207_));
  INV_X1     g11205(.I(\A[544] ), .ZN(new_n12208_));
  NAND2_X1   g11206(.A1(new_n12208_), .A2(\A[545] ), .ZN(new_n12209_));
  NOR2_X1    g11207(.A1(new_n12208_), .A2(\A[545] ), .ZN(new_n12210_));
  NOR2_X1    g11208(.A1(new_n12210_), .A2(new_n12207_), .ZN(new_n12211_));
  INV_X1     g11209(.I(\A[545] ), .ZN(new_n12212_));
  NAND2_X1   g11210(.A1(new_n12212_), .A2(\A[544] ), .ZN(new_n12213_));
  NAND2_X1   g11211(.A1(new_n12209_), .A2(new_n12213_), .ZN(new_n12214_));
  AOI22_X1   g11212(.A1(new_n12214_), .A2(new_n12207_), .B1(new_n12211_), .B2(new_n12209_), .ZN(new_n12215_));
  XNOR2_X1   g11213(.A1(new_n12215_), .A2(new_n12206_), .ZN(new_n12216_));
  NOR2_X1    g11214(.A1(new_n12212_), .A2(\A[544] ), .ZN(new_n12217_));
  NOR2_X1    g11215(.A1(new_n12217_), .A2(new_n12210_), .ZN(new_n12218_));
  NOR2_X1    g11216(.A1(new_n12208_), .A2(new_n12212_), .ZN(new_n12219_));
  INV_X1     g11217(.I(new_n12219_), .ZN(new_n12220_));
  OAI21_X1   g11218(.A1(new_n12218_), .A2(new_n12207_), .B(new_n12220_), .ZN(new_n12221_));
  NAND2_X1   g11219(.A1(new_n12203_), .A2(\A[542] ), .ZN(new_n12222_));
  NAND2_X1   g11220(.A1(new_n12222_), .A2(new_n12201_), .ZN(new_n12223_));
  NOR2_X1    g11221(.A1(new_n12203_), .A2(new_n12199_), .ZN(new_n12224_));
  AOI21_X1   g11222(.A1(new_n12223_), .A2(\A[543] ), .B(new_n12224_), .ZN(new_n12225_));
  INV_X1     g11223(.I(new_n12225_), .ZN(new_n12226_));
  INV_X1     g11224(.I(new_n12206_), .ZN(new_n12227_));
  NOR2_X1    g11225(.A1(new_n12227_), .A2(new_n12215_), .ZN(new_n12228_));
  NAND3_X1   g11226(.A1(new_n12228_), .A2(new_n12221_), .A3(new_n12226_), .ZN(new_n12229_));
  NAND2_X1   g11227(.A1(new_n12229_), .A2(new_n12216_), .ZN(new_n12230_));
  INV_X1     g11228(.I(\A[537] ), .ZN(new_n12231_));
  INV_X1     g11229(.I(\A[535] ), .ZN(new_n12232_));
  NAND2_X1   g11230(.A1(new_n12232_), .A2(\A[536] ), .ZN(new_n12233_));
  NOR2_X1    g11231(.A1(new_n12232_), .A2(\A[536] ), .ZN(new_n12234_));
  NOR2_X1    g11232(.A1(new_n12234_), .A2(new_n12231_), .ZN(new_n12235_));
  INV_X1     g11233(.I(\A[536] ), .ZN(new_n12236_));
  NAND2_X1   g11234(.A1(new_n12236_), .A2(\A[535] ), .ZN(new_n12237_));
  NAND2_X1   g11235(.A1(new_n12233_), .A2(new_n12237_), .ZN(new_n12238_));
  AOI22_X1   g11236(.A1(new_n12238_), .A2(new_n12231_), .B1(new_n12235_), .B2(new_n12233_), .ZN(new_n12239_));
  INV_X1     g11237(.I(\A[540] ), .ZN(new_n12240_));
  INV_X1     g11238(.I(\A[538] ), .ZN(new_n12241_));
  NAND2_X1   g11239(.A1(new_n12241_), .A2(\A[539] ), .ZN(new_n12242_));
  NOR2_X1    g11240(.A1(new_n12241_), .A2(\A[539] ), .ZN(new_n12243_));
  NOR2_X1    g11241(.A1(new_n12243_), .A2(new_n12240_), .ZN(new_n12244_));
  INV_X1     g11242(.I(\A[539] ), .ZN(new_n12245_));
  NAND2_X1   g11243(.A1(new_n12245_), .A2(\A[538] ), .ZN(new_n12246_));
  NAND2_X1   g11244(.A1(new_n12242_), .A2(new_n12246_), .ZN(new_n12247_));
  AOI22_X1   g11245(.A1(new_n12247_), .A2(new_n12240_), .B1(new_n12244_), .B2(new_n12242_), .ZN(new_n12248_));
  XOR2_X1    g11246(.A1(new_n12239_), .A2(new_n12248_), .Z(new_n12249_));
  NOR2_X1    g11247(.A1(new_n12245_), .A2(\A[538] ), .ZN(new_n12250_));
  NOR2_X1    g11248(.A1(new_n12250_), .A2(new_n12243_), .ZN(new_n12251_));
  NOR2_X1    g11249(.A1(new_n12241_), .A2(new_n12245_), .ZN(new_n12252_));
  INV_X1     g11250(.I(new_n12252_), .ZN(new_n12253_));
  OAI21_X1   g11251(.A1(new_n12251_), .A2(new_n12240_), .B(new_n12253_), .ZN(new_n12254_));
  NOR2_X1    g11252(.A1(new_n12232_), .A2(new_n12236_), .ZN(new_n12255_));
  AOI21_X1   g11253(.A1(new_n12238_), .A2(\A[537] ), .B(new_n12255_), .ZN(new_n12256_));
  INV_X1     g11254(.I(new_n12256_), .ZN(new_n12257_));
  NOR2_X1    g11255(.A1(new_n12239_), .A2(new_n12248_), .ZN(new_n12258_));
  NAND3_X1   g11256(.A1(new_n12258_), .A2(new_n12254_), .A3(new_n12257_), .ZN(new_n12259_));
  NAND2_X1   g11257(.A1(new_n12249_), .A2(new_n12259_), .ZN(new_n12260_));
  XOR2_X1    g11258(.A1(new_n12230_), .A2(new_n12260_), .Z(new_n12261_));
  XOR2_X1    g11259(.A1(new_n12198_), .A2(new_n12261_), .Z(new_n12262_));
  INV_X1     g11260(.I(\A[530] ), .ZN(new_n12263_));
  NOR2_X1    g11261(.A1(new_n12263_), .A2(\A[529] ), .ZN(new_n12264_));
  NAND2_X1   g11262(.A1(new_n12263_), .A2(\A[529] ), .ZN(new_n12265_));
  NAND2_X1   g11263(.A1(new_n12265_), .A2(\A[531] ), .ZN(new_n12266_));
  INV_X1     g11264(.I(\A[529] ), .ZN(new_n12267_));
  NOR2_X1    g11265(.A1(new_n12267_), .A2(\A[530] ), .ZN(new_n12268_));
  NOR2_X1    g11266(.A1(new_n12264_), .A2(new_n12268_), .ZN(new_n12269_));
  OAI22_X1   g11267(.A1(new_n12269_), .A2(\A[531] ), .B1(new_n12266_), .B2(new_n12264_), .ZN(new_n12270_));
  INV_X1     g11268(.I(\A[534] ), .ZN(new_n12271_));
  INV_X1     g11269(.I(\A[532] ), .ZN(new_n12272_));
  NAND2_X1   g11270(.A1(new_n12272_), .A2(\A[533] ), .ZN(new_n12273_));
  NOR2_X1    g11271(.A1(new_n12272_), .A2(\A[533] ), .ZN(new_n12274_));
  NOR2_X1    g11272(.A1(new_n12274_), .A2(new_n12271_), .ZN(new_n12275_));
  INV_X1     g11273(.I(\A[533] ), .ZN(new_n12276_));
  NAND2_X1   g11274(.A1(new_n12276_), .A2(\A[532] ), .ZN(new_n12277_));
  NAND2_X1   g11275(.A1(new_n12273_), .A2(new_n12277_), .ZN(new_n12278_));
  AOI22_X1   g11276(.A1(new_n12278_), .A2(new_n12271_), .B1(new_n12275_), .B2(new_n12273_), .ZN(new_n12279_));
  XNOR2_X1   g11277(.A1(new_n12279_), .A2(new_n12270_), .ZN(new_n12280_));
  NOR2_X1    g11278(.A1(new_n12276_), .A2(\A[532] ), .ZN(new_n12281_));
  NOR2_X1    g11279(.A1(new_n12281_), .A2(new_n12274_), .ZN(new_n12282_));
  NOR2_X1    g11280(.A1(new_n12272_), .A2(new_n12276_), .ZN(new_n12283_));
  INV_X1     g11281(.I(new_n12283_), .ZN(new_n12284_));
  OAI21_X1   g11282(.A1(new_n12282_), .A2(new_n12271_), .B(new_n12284_), .ZN(new_n12285_));
  NAND2_X1   g11283(.A1(new_n12267_), .A2(\A[530] ), .ZN(new_n12286_));
  NAND2_X1   g11284(.A1(new_n12286_), .A2(new_n12265_), .ZN(new_n12287_));
  NOR2_X1    g11285(.A1(new_n12267_), .A2(new_n12263_), .ZN(new_n12288_));
  AOI21_X1   g11286(.A1(new_n12287_), .A2(\A[531] ), .B(new_n12288_), .ZN(new_n12289_));
  INV_X1     g11287(.I(new_n12289_), .ZN(new_n12290_));
  INV_X1     g11288(.I(new_n12270_), .ZN(new_n12291_));
  NOR2_X1    g11289(.A1(new_n12291_), .A2(new_n12279_), .ZN(new_n12292_));
  NAND3_X1   g11290(.A1(new_n12292_), .A2(new_n12285_), .A3(new_n12290_), .ZN(new_n12293_));
  NAND2_X1   g11291(.A1(new_n12293_), .A2(new_n12280_), .ZN(new_n12294_));
  INV_X1     g11292(.I(\A[524] ), .ZN(new_n12295_));
  NOR2_X1    g11293(.A1(new_n12295_), .A2(\A[523] ), .ZN(new_n12296_));
  NAND2_X1   g11294(.A1(new_n12295_), .A2(\A[523] ), .ZN(new_n12297_));
  NAND2_X1   g11295(.A1(new_n12297_), .A2(\A[525] ), .ZN(new_n12298_));
  INV_X1     g11296(.I(\A[523] ), .ZN(new_n12299_));
  NOR2_X1    g11297(.A1(new_n12299_), .A2(\A[524] ), .ZN(new_n12300_));
  NOR2_X1    g11298(.A1(new_n12296_), .A2(new_n12300_), .ZN(new_n12301_));
  OAI22_X1   g11299(.A1(new_n12301_), .A2(\A[525] ), .B1(new_n12298_), .B2(new_n12296_), .ZN(new_n12302_));
  INV_X1     g11300(.I(\A[528] ), .ZN(new_n12303_));
  INV_X1     g11301(.I(\A[526] ), .ZN(new_n12304_));
  NAND2_X1   g11302(.A1(new_n12304_), .A2(\A[527] ), .ZN(new_n12305_));
  NOR2_X1    g11303(.A1(new_n12304_), .A2(\A[527] ), .ZN(new_n12306_));
  NOR2_X1    g11304(.A1(new_n12306_), .A2(new_n12303_), .ZN(new_n12307_));
  INV_X1     g11305(.I(\A[527] ), .ZN(new_n12308_));
  NAND2_X1   g11306(.A1(new_n12308_), .A2(\A[526] ), .ZN(new_n12309_));
  NAND2_X1   g11307(.A1(new_n12305_), .A2(new_n12309_), .ZN(new_n12310_));
  AOI22_X1   g11308(.A1(new_n12310_), .A2(new_n12303_), .B1(new_n12307_), .B2(new_n12305_), .ZN(new_n12311_));
  XNOR2_X1   g11309(.A1(new_n12311_), .A2(new_n12302_), .ZN(new_n12312_));
  NOR2_X1    g11310(.A1(new_n12308_), .A2(\A[526] ), .ZN(new_n12313_));
  NOR2_X1    g11311(.A1(new_n12313_), .A2(new_n12306_), .ZN(new_n12314_));
  NOR2_X1    g11312(.A1(new_n12304_), .A2(new_n12308_), .ZN(new_n12315_));
  INV_X1     g11313(.I(new_n12315_), .ZN(new_n12316_));
  OAI21_X1   g11314(.A1(new_n12314_), .A2(new_n12303_), .B(new_n12316_), .ZN(new_n12317_));
  NAND2_X1   g11315(.A1(new_n12299_), .A2(\A[524] ), .ZN(new_n12318_));
  NAND2_X1   g11316(.A1(new_n12318_), .A2(new_n12297_), .ZN(new_n12319_));
  NOR2_X1    g11317(.A1(new_n12299_), .A2(new_n12295_), .ZN(new_n12320_));
  AOI21_X1   g11318(.A1(new_n12319_), .A2(\A[525] ), .B(new_n12320_), .ZN(new_n12321_));
  INV_X1     g11319(.I(new_n12321_), .ZN(new_n12322_));
  INV_X1     g11320(.I(new_n12302_), .ZN(new_n12323_));
  NOR2_X1    g11321(.A1(new_n12323_), .A2(new_n12311_), .ZN(new_n12324_));
  NAND3_X1   g11322(.A1(new_n12324_), .A2(new_n12317_), .A3(new_n12322_), .ZN(new_n12325_));
  NAND2_X1   g11323(.A1(new_n12325_), .A2(new_n12312_), .ZN(new_n12326_));
  XOR2_X1    g11324(.A1(new_n12294_), .A2(new_n12326_), .Z(new_n12327_));
  INV_X1     g11325(.I(\A[518] ), .ZN(new_n12328_));
  NOR2_X1    g11326(.A1(new_n12328_), .A2(\A[517] ), .ZN(new_n12329_));
  NAND2_X1   g11327(.A1(new_n12328_), .A2(\A[517] ), .ZN(new_n12330_));
  NAND2_X1   g11328(.A1(new_n12330_), .A2(\A[519] ), .ZN(new_n12331_));
  INV_X1     g11329(.I(\A[517] ), .ZN(new_n12332_));
  NOR2_X1    g11330(.A1(new_n12332_), .A2(\A[518] ), .ZN(new_n12333_));
  NOR2_X1    g11331(.A1(new_n12329_), .A2(new_n12333_), .ZN(new_n12334_));
  OAI22_X1   g11332(.A1(new_n12334_), .A2(\A[519] ), .B1(new_n12331_), .B2(new_n12329_), .ZN(new_n12335_));
  INV_X1     g11333(.I(\A[522] ), .ZN(new_n12336_));
  INV_X1     g11334(.I(\A[520] ), .ZN(new_n12337_));
  NAND2_X1   g11335(.A1(new_n12337_), .A2(\A[521] ), .ZN(new_n12338_));
  NOR2_X1    g11336(.A1(new_n12337_), .A2(\A[521] ), .ZN(new_n12339_));
  NOR2_X1    g11337(.A1(new_n12339_), .A2(new_n12336_), .ZN(new_n12340_));
  INV_X1     g11338(.I(\A[521] ), .ZN(new_n12341_));
  NAND2_X1   g11339(.A1(new_n12341_), .A2(\A[520] ), .ZN(new_n12342_));
  NAND2_X1   g11340(.A1(new_n12338_), .A2(new_n12342_), .ZN(new_n12343_));
  AOI22_X1   g11341(.A1(new_n12343_), .A2(new_n12336_), .B1(new_n12340_), .B2(new_n12338_), .ZN(new_n12344_));
  XNOR2_X1   g11342(.A1(new_n12344_), .A2(new_n12335_), .ZN(new_n12345_));
  NOR2_X1    g11343(.A1(new_n12341_), .A2(\A[520] ), .ZN(new_n12346_));
  NOR2_X1    g11344(.A1(new_n12346_), .A2(new_n12339_), .ZN(new_n12347_));
  NOR2_X1    g11345(.A1(new_n12337_), .A2(new_n12341_), .ZN(new_n12348_));
  INV_X1     g11346(.I(new_n12348_), .ZN(new_n12349_));
  OAI21_X1   g11347(.A1(new_n12347_), .A2(new_n12336_), .B(new_n12349_), .ZN(new_n12350_));
  NAND2_X1   g11348(.A1(new_n12332_), .A2(\A[518] ), .ZN(new_n12351_));
  NAND2_X1   g11349(.A1(new_n12351_), .A2(new_n12330_), .ZN(new_n12352_));
  NOR2_X1    g11350(.A1(new_n12332_), .A2(new_n12328_), .ZN(new_n12353_));
  AOI21_X1   g11351(.A1(new_n12352_), .A2(\A[519] ), .B(new_n12353_), .ZN(new_n12354_));
  INV_X1     g11352(.I(new_n12354_), .ZN(new_n12355_));
  INV_X1     g11353(.I(new_n12335_), .ZN(new_n12356_));
  NOR2_X1    g11354(.A1(new_n12356_), .A2(new_n12344_), .ZN(new_n12357_));
  NAND3_X1   g11355(.A1(new_n12357_), .A2(new_n12350_), .A3(new_n12355_), .ZN(new_n12358_));
  NAND2_X1   g11356(.A1(new_n12358_), .A2(new_n12345_), .ZN(new_n12359_));
  INV_X1     g11357(.I(\A[512] ), .ZN(new_n12360_));
  NOR2_X1    g11358(.A1(new_n12360_), .A2(\A[511] ), .ZN(new_n12361_));
  NAND2_X1   g11359(.A1(new_n12360_), .A2(\A[511] ), .ZN(new_n12362_));
  NAND2_X1   g11360(.A1(new_n12362_), .A2(\A[513] ), .ZN(new_n12363_));
  INV_X1     g11361(.I(\A[511] ), .ZN(new_n12364_));
  NOR2_X1    g11362(.A1(new_n12364_), .A2(\A[512] ), .ZN(new_n12365_));
  NOR2_X1    g11363(.A1(new_n12361_), .A2(new_n12365_), .ZN(new_n12366_));
  OAI22_X1   g11364(.A1(new_n12366_), .A2(\A[513] ), .B1(new_n12363_), .B2(new_n12361_), .ZN(new_n12367_));
  INV_X1     g11365(.I(\A[516] ), .ZN(new_n12368_));
  INV_X1     g11366(.I(\A[514] ), .ZN(new_n12369_));
  NAND2_X1   g11367(.A1(new_n12369_), .A2(\A[515] ), .ZN(new_n12370_));
  NOR2_X1    g11368(.A1(new_n12369_), .A2(\A[515] ), .ZN(new_n12371_));
  NOR2_X1    g11369(.A1(new_n12371_), .A2(new_n12368_), .ZN(new_n12372_));
  INV_X1     g11370(.I(\A[515] ), .ZN(new_n12373_));
  NAND2_X1   g11371(.A1(new_n12373_), .A2(\A[514] ), .ZN(new_n12374_));
  NAND2_X1   g11372(.A1(new_n12370_), .A2(new_n12374_), .ZN(new_n12375_));
  AOI22_X1   g11373(.A1(new_n12375_), .A2(new_n12368_), .B1(new_n12372_), .B2(new_n12370_), .ZN(new_n12376_));
  XNOR2_X1   g11374(.A1(new_n12376_), .A2(new_n12367_), .ZN(new_n12377_));
  NOR2_X1    g11375(.A1(new_n12373_), .A2(\A[514] ), .ZN(new_n12378_));
  NOR2_X1    g11376(.A1(new_n12378_), .A2(new_n12371_), .ZN(new_n12379_));
  NOR2_X1    g11377(.A1(new_n12369_), .A2(new_n12373_), .ZN(new_n12380_));
  INV_X1     g11378(.I(new_n12380_), .ZN(new_n12381_));
  OAI21_X1   g11379(.A1(new_n12379_), .A2(new_n12368_), .B(new_n12381_), .ZN(new_n12382_));
  NAND2_X1   g11380(.A1(new_n12364_), .A2(\A[512] ), .ZN(new_n12383_));
  NAND2_X1   g11381(.A1(new_n12383_), .A2(new_n12362_), .ZN(new_n12384_));
  NOR2_X1    g11382(.A1(new_n12364_), .A2(new_n12360_), .ZN(new_n12385_));
  AOI21_X1   g11383(.A1(new_n12384_), .A2(\A[513] ), .B(new_n12385_), .ZN(new_n12386_));
  INV_X1     g11384(.I(new_n12386_), .ZN(new_n12387_));
  INV_X1     g11385(.I(new_n12367_), .ZN(new_n12388_));
  NOR2_X1    g11386(.A1(new_n12388_), .A2(new_n12376_), .ZN(new_n12389_));
  NAND3_X1   g11387(.A1(new_n12389_), .A2(new_n12382_), .A3(new_n12387_), .ZN(new_n12390_));
  NAND2_X1   g11388(.A1(new_n12390_), .A2(new_n12377_), .ZN(new_n12391_));
  XOR2_X1    g11389(.A1(new_n12359_), .A2(new_n12391_), .Z(new_n12392_));
  XOR2_X1    g11390(.A1(new_n12327_), .A2(new_n12392_), .Z(new_n12393_));
  XOR2_X1    g11391(.A1(new_n12393_), .A2(new_n12262_), .Z(new_n12394_));
  XOR2_X1    g11392(.A1(new_n12133_), .A2(new_n12394_), .Z(new_n12395_));
  INV_X1     g11393(.I(\A[650] ), .ZN(new_n12396_));
  NOR2_X1    g11394(.A1(new_n12396_), .A2(\A[649] ), .ZN(new_n12397_));
  NAND2_X1   g11395(.A1(new_n12396_), .A2(\A[649] ), .ZN(new_n12398_));
  NAND2_X1   g11396(.A1(new_n12398_), .A2(\A[651] ), .ZN(new_n12399_));
  INV_X1     g11397(.I(\A[649] ), .ZN(new_n12400_));
  NOR2_X1    g11398(.A1(new_n12400_), .A2(\A[650] ), .ZN(new_n12401_));
  NOR2_X1    g11399(.A1(new_n12397_), .A2(new_n12401_), .ZN(new_n12402_));
  OAI22_X1   g11400(.A1(new_n12402_), .A2(\A[651] ), .B1(new_n12399_), .B2(new_n12397_), .ZN(new_n12403_));
  INV_X1     g11401(.I(\A[654] ), .ZN(new_n12404_));
  INV_X1     g11402(.I(\A[652] ), .ZN(new_n12405_));
  NAND2_X1   g11403(.A1(new_n12405_), .A2(\A[653] ), .ZN(new_n12406_));
  NOR2_X1    g11404(.A1(new_n12405_), .A2(\A[653] ), .ZN(new_n12407_));
  NOR2_X1    g11405(.A1(new_n12407_), .A2(new_n12404_), .ZN(new_n12408_));
  INV_X1     g11406(.I(\A[653] ), .ZN(new_n12409_));
  NAND2_X1   g11407(.A1(new_n12409_), .A2(\A[652] ), .ZN(new_n12410_));
  NAND2_X1   g11408(.A1(new_n12406_), .A2(new_n12410_), .ZN(new_n12411_));
  AOI22_X1   g11409(.A1(new_n12411_), .A2(new_n12404_), .B1(new_n12408_), .B2(new_n12406_), .ZN(new_n12412_));
  XNOR2_X1   g11410(.A1(new_n12412_), .A2(new_n12403_), .ZN(new_n12413_));
  NOR2_X1    g11411(.A1(new_n12409_), .A2(\A[652] ), .ZN(new_n12414_));
  NOR2_X1    g11412(.A1(new_n12414_), .A2(new_n12407_), .ZN(new_n12415_));
  NOR2_X1    g11413(.A1(new_n12405_), .A2(new_n12409_), .ZN(new_n12416_));
  INV_X1     g11414(.I(new_n12416_), .ZN(new_n12417_));
  OAI21_X1   g11415(.A1(new_n12415_), .A2(new_n12404_), .B(new_n12417_), .ZN(new_n12418_));
  INV_X1     g11416(.I(\A[651] ), .ZN(new_n12419_));
  NOR2_X1    g11417(.A1(new_n12400_), .A2(new_n12396_), .ZN(new_n12420_));
  INV_X1     g11418(.I(new_n12420_), .ZN(new_n12421_));
  OAI21_X1   g11419(.A1(new_n12402_), .A2(new_n12419_), .B(new_n12421_), .ZN(new_n12422_));
  INV_X1     g11420(.I(new_n12403_), .ZN(new_n12423_));
  NOR2_X1    g11421(.A1(new_n12423_), .A2(new_n12412_), .ZN(new_n12424_));
  NAND3_X1   g11422(.A1(new_n12424_), .A2(new_n12418_), .A3(new_n12422_), .ZN(new_n12425_));
  NAND2_X1   g11423(.A1(new_n12425_), .A2(new_n12413_), .ZN(new_n12426_));
  INV_X1     g11424(.I(\A[644] ), .ZN(new_n12427_));
  NOR2_X1    g11425(.A1(new_n12427_), .A2(\A[643] ), .ZN(new_n12428_));
  NAND2_X1   g11426(.A1(new_n12427_), .A2(\A[643] ), .ZN(new_n12429_));
  NAND2_X1   g11427(.A1(new_n12429_), .A2(\A[645] ), .ZN(new_n12430_));
  INV_X1     g11428(.I(\A[643] ), .ZN(new_n12431_));
  NOR2_X1    g11429(.A1(new_n12431_), .A2(\A[644] ), .ZN(new_n12432_));
  NOR2_X1    g11430(.A1(new_n12428_), .A2(new_n12432_), .ZN(new_n12433_));
  OAI22_X1   g11431(.A1(new_n12433_), .A2(\A[645] ), .B1(new_n12430_), .B2(new_n12428_), .ZN(new_n12434_));
  INV_X1     g11432(.I(\A[648] ), .ZN(new_n12435_));
  INV_X1     g11433(.I(\A[646] ), .ZN(new_n12436_));
  NAND2_X1   g11434(.A1(new_n12436_), .A2(\A[647] ), .ZN(new_n12437_));
  INV_X1     g11435(.I(\A[647] ), .ZN(new_n12438_));
  AOI21_X1   g11436(.A1(\A[646] ), .A2(new_n12438_), .B(new_n12435_), .ZN(new_n12439_));
  NAND2_X1   g11437(.A1(new_n12438_), .A2(\A[646] ), .ZN(new_n12440_));
  NAND2_X1   g11438(.A1(new_n12437_), .A2(new_n12440_), .ZN(new_n12441_));
  AOI22_X1   g11439(.A1(new_n12441_), .A2(new_n12435_), .B1(new_n12437_), .B2(new_n12439_), .ZN(new_n12442_));
  XNOR2_X1   g11440(.A1(new_n12434_), .A2(new_n12442_), .ZN(new_n12443_));
  NOR2_X1    g11441(.A1(new_n12436_), .A2(new_n12438_), .ZN(new_n12444_));
  INV_X1     g11442(.I(new_n12444_), .ZN(new_n12445_));
  NAND2_X1   g11443(.A1(new_n12441_), .A2(\A[648] ), .ZN(new_n12446_));
  NAND2_X1   g11444(.A1(new_n12446_), .A2(new_n12445_), .ZN(new_n12447_));
  INV_X1     g11445(.I(\A[645] ), .ZN(new_n12448_));
  NOR2_X1    g11446(.A1(new_n12431_), .A2(new_n12427_), .ZN(new_n12449_));
  INV_X1     g11447(.I(new_n12449_), .ZN(new_n12450_));
  OAI21_X1   g11448(.A1(new_n12433_), .A2(new_n12448_), .B(new_n12450_), .ZN(new_n12451_));
  INV_X1     g11449(.I(new_n12434_), .ZN(new_n12452_));
  NOR2_X1    g11450(.A1(new_n12452_), .A2(new_n12442_), .ZN(new_n12453_));
  NAND3_X1   g11451(.A1(new_n12453_), .A2(new_n12447_), .A3(new_n12451_), .ZN(new_n12454_));
  NAND2_X1   g11452(.A1(new_n12454_), .A2(new_n12443_), .ZN(new_n12455_));
  XOR2_X1    g11453(.A1(new_n12426_), .A2(new_n12455_), .Z(new_n12456_));
  INV_X1     g11454(.I(\A[638] ), .ZN(new_n12457_));
  NOR2_X1    g11455(.A1(new_n12457_), .A2(\A[637] ), .ZN(new_n12458_));
  NAND2_X1   g11456(.A1(new_n12457_), .A2(\A[637] ), .ZN(new_n12459_));
  NAND2_X1   g11457(.A1(new_n12459_), .A2(\A[639] ), .ZN(new_n12460_));
  INV_X1     g11458(.I(\A[637] ), .ZN(new_n12461_));
  NOR2_X1    g11459(.A1(new_n12461_), .A2(\A[638] ), .ZN(new_n12462_));
  NOR2_X1    g11460(.A1(new_n12458_), .A2(new_n12462_), .ZN(new_n12463_));
  OAI22_X1   g11461(.A1(new_n12463_), .A2(\A[639] ), .B1(new_n12460_), .B2(new_n12458_), .ZN(new_n12464_));
  INV_X1     g11462(.I(\A[642] ), .ZN(new_n12465_));
  INV_X1     g11463(.I(\A[640] ), .ZN(new_n12466_));
  NAND2_X1   g11464(.A1(new_n12466_), .A2(\A[641] ), .ZN(new_n12467_));
  NOR2_X1    g11465(.A1(new_n12466_), .A2(\A[641] ), .ZN(new_n12468_));
  NOR2_X1    g11466(.A1(new_n12468_), .A2(new_n12465_), .ZN(new_n12469_));
  INV_X1     g11467(.I(\A[641] ), .ZN(new_n12470_));
  NAND2_X1   g11468(.A1(new_n12470_), .A2(\A[640] ), .ZN(new_n12471_));
  NAND2_X1   g11469(.A1(new_n12467_), .A2(new_n12471_), .ZN(new_n12472_));
  AOI22_X1   g11470(.A1(new_n12472_), .A2(new_n12465_), .B1(new_n12469_), .B2(new_n12467_), .ZN(new_n12473_));
  XNOR2_X1   g11471(.A1(new_n12473_), .A2(new_n12464_), .ZN(new_n12474_));
  NOR2_X1    g11472(.A1(new_n12470_), .A2(\A[640] ), .ZN(new_n12475_));
  NOR2_X1    g11473(.A1(new_n12475_), .A2(new_n12468_), .ZN(new_n12476_));
  NOR2_X1    g11474(.A1(new_n12466_), .A2(new_n12470_), .ZN(new_n12477_));
  INV_X1     g11475(.I(new_n12477_), .ZN(new_n12478_));
  OAI21_X1   g11476(.A1(new_n12476_), .A2(new_n12465_), .B(new_n12478_), .ZN(new_n12479_));
  NAND2_X1   g11477(.A1(new_n12461_), .A2(\A[638] ), .ZN(new_n12480_));
  NAND2_X1   g11478(.A1(new_n12480_), .A2(new_n12459_), .ZN(new_n12481_));
  NOR2_X1    g11479(.A1(new_n12461_), .A2(new_n12457_), .ZN(new_n12482_));
  AOI21_X1   g11480(.A1(new_n12481_), .A2(\A[639] ), .B(new_n12482_), .ZN(new_n12483_));
  INV_X1     g11481(.I(new_n12483_), .ZN(new_n12484_));
  INV_X1     g11482(.I(new_n12464_), .ZN(new_n12485_));
  NOR2_X1    g11483(.A1(new_n12485_), .A2(new_n12473_), .ZN(new_n12486_));
  NAND3_X1   g11484(.A1(new_n12486_), .A2(new_n12479_), .A3(new_n12484_), .ZN(new_n12487_));
  NAND2_X1   g11485(.A1(new_n12487_), .A2(new_n12474_), .ZN(new_n12488_));
  INV_X1     g11486(.I(\A[633] ), .ZN(new_n12489_));
  INV_X1     g11487(.I(\A[631] ), .ZN(new_n12490_));
  NAND2_X1   g11488(.A1(new_n12490_), .A2(\A[632] ), .ZN(new_n12491_));
  NOR2_X1    g11489(.A1(new_n12490_), .A2(\A[632] ), .ZN(new_n12492_));
  NOR2_X1    g11490(.A1(new_n12492_), .A2(new_n12489_), .ZN(new_n12493_));
  INV_X1     g11491(.I(\A[632] ), .ZN(new_n12494_));
  NAND2_X1   g11492(.A1(new_n12494_), .A2(\A[631] ), .ZN(new_n12495_));
  NAND2_X1   g11493(.A1(new_n12491_), .A2(new_n12495_), .ZN(new_n12496_));
  AOI22_X1   g11494(.A1(new_n12496_), .A2(new_n12489_), .B1(new_n12493_), .B2(new_n12491_), .ZN(new_n12497_));
  INV_X1     g11495(.I(\A[636] ), .ZN(new_n12498_));
  INV_X1     g11496(.I(\A[634] ), .ZN(new_n12499_));
  NAND2_X1   g11497(.A1(new_n12499_), .A2(\A[635] ), .ZN(new_n12500_));
  NOR2_X1    g11498(.A1(new_n12499_), .A2(\A[635] ), .ZN(new_n12501_));
  NOR2_X1    g11499(.A1(new_n12501_), .A2(new_n12498_), .ZN(new_n12502_));
  INV_X1     g11500(.I(\A[635] ), .ZN(new_n12503_));
  NAND2_X1   g11501(.A1(new_n12503_), .A2(\A[634] ), .ZN(new_n12504_));
  NAND2_X1   g11502(.A1(new_n12500_), .A2(new_n12504_), .ZN(new_n12505_));
  AOI22_X1   g11503(.A1(new_n12505_), .A2(new_n12498_), .B1(new_n12502_), .B2(new_n12500_), .ZN(new_n12506_));
  XOR2_X1    g11504(.A1(new_n12497_), .A2(new_n12506_), .Z(new_n12507_));
  NOR2_X1    g11505(.A1(new_n12503_), .A2(\A[634] ), .ZN(new_n12508_));
  NOR2_X1    g11506(.A1(new_n12508_), .A2(new_n12501_), .ZN(new_n12509_));
  NOR2_X1    g11507(.A1(new_n12499_), .A2(new_n12503_), .ZN(new_n12510_));
  INV_X1     g11508(.I(new_n12510_), .ZN(new_n12511_));
  OAI21_X1   g11509(.A1(new_n12509_), .A2(new_n12498_), .B(new_n12511_), .ZN(new_n12512_));
  NOR2_X1    g11510(.A1(new_n12490_), .A2(new_n12494_), .ZN(new_n12513_));
  AOI21_X1   g11511(.A1(new_n12496_), .A2(\A[633] ), .B(new_n12513_), .ZN(new_n12514_));
  INV_X1     g11512(.I(new_n12514_), .ZN(new_n12515_));
  NOR2_X1    g11513(.A1(new_n12497_), .A2(new_n12506_), .ZN(new_n12516_));
  NAND3_X1   g11514(.A1(new_n12516_), .A2(new_n12512_), .A3(new_n12515_), .ZN(new_n12517_));
  NAND2_X1   g11515(.A1(new_n12507_), .A2(new_n12517_), .ZN(new_n12518_));
  XOR2_X1    g11516(.A1(new_n12488_), .A2(new_n12518_), .Z(new_n12519_));
  XOR2_X1    g11517(.A1(new_n12456_), .A2(new_n12519_), .Z(new_n12520_));
  INV_X1     g11518(.I(\A[626] ), .ZN(new_n12521_));
  NOR2_X1    g11519(.A1(new_n12521_), .A2(\A[625] ), .ZN(new_n12522_));
  NAND2_X1   g11520(.A1(new_n12521_), .A2(\A[625] ), .ZN(new_n12523_));
  NAND2_X1   g11521(.A1(new_n12523_), .A2(\A[627] ), .ZN(new_n12524_));
  INV_X1     g11522(.I(\A[625] ), .ZN(new_n12525_));
  NOR2_X1    g11523(.A1(new_n12525_), .A2(\A[626] ), .ZN(new_n12526_));
  NOR2_X1    g11524(.A1(new_n12522_), .A2(new_n12526_), .ZN(new_n12527_));
  OAI22_X1   g11525(.A1(new_n12527_), .A2(\A[627] ), .B1(new_n12524_), .B2(new_n12522_), .ZN(new_n12528_));
  INV_X1     g11526(.I(\A[630] ), .ZN(new_n12529_));
  INV_X1     g11527(.I(\A[628] ), .ZN(new_n12530_));
  NAND2_X1   g11528(.A1(new_n12530_), .A2(\A[629] ), .ZN(new_n12531_));
  NOR2_X1    g11529(.A1(new_n12530_), .A2(\A[629] ), .ZN(new_n12532_));
  NOR2_X1    g11530(.A1(new_n12532_), .A2(new_n12529_), .ZN(new_n12533_));
  INV_X1     g11531(.I(\A[629] ), .ZN(new_n12534_));
  NAND2_X1   g11532(.A1(new_n12534_), .A2(\A[628] ), .ZN(new_n12535_));
  NAND2_X1   g11533(.A1(new_n12531_), .A2(new_n12535_), .ZN(new_n12536_));
  AOI22_X1   g11534(.A1(new_n12536_), .A2(new_n12529_), .B1(new_n12533_), .B2(new_n12531_), .ZN(new_n12537_));
  XNOR2_X1   g11535(.A1(new_n12537_), .A2(new_n12528_), .ZN(new_n12538_));
  NOR2_X1    g11536(.A1(new_n12534_), .A2(\A[628] ), .ZN(new_n12539_));
  NOR2_X1    g11537(.A1(new_n12539_), .A2(new_n12532_), .ZN(new_n12540_));
  NOR2_X1    g11538(.A1(new_n12530_), .A2(new_n12534_), .ZN(new_n12541_));
  INV_X1     g11539(.I(new_n12541_), .ZN(new_n12542_));
  OAI21_X1   g11540(.A1(new_n12540_), .A2(new_n12529_), .B(new_n12542_), .ZN(new_n12543_));
  NAND2_X1   g11541(.A1(new_n12525_), .A2(\A[626] ), .ZN(new_n12544_));
  NAND2_X1   g11542(.A1(new_n12544_), .A2(new_n12523_), .ZN(new_n12545_));
  NOR2_X1    g11543(.A1(new_n12525_), .A2(new_n12521_), .ZN(new_n12546_));
  AOI21_X1   g11544(.A1(new_n12545_), .A2(\A[627] ), .B(new_n12546_), .ZN(new_n12547_));
  INV_X1     g11545(.I(new_n12547_), .ZN(new_n12548_));
  INV_X1     g11546(.I(new_n12528_), .ZN(new_n12549_));
  NOR2_X1    g11547(.A1(new_n12549_), .A2(new_n12537_), .ZN(new_n12550_));
  NAND3_X1   g11548(.A1(new_n12550_), .A2(new_n12543_), .A3(new_n12548_), .ZN(new_n12551_));
  NAND2_X1   g11549(.A1(new_n12551_), .A2(new_n12538_), .ZN(new_n12552_));
  INV_X1     g11550(.I(\A[620] ), .ZN(new_n12553_));
  NOR2_X1    g11551(.A1(new_n12553_), .A2(\A[619] ), .ZN(new_n12554_));
  NAND2_X1   g11552(.A1(new_n12553_), .A2(\A[619] ), .ZN(new_n12555_));
  NAND2_X1   g11553(.A1(new_n12555_), .A2(\A[621] ), .ZN(new_n12556_));
  INV_X1     g11554(.I(\A[619] ), .ZN(new_n12557_));
  NOR2_X1    g11555(.A1(new_n12557_), .A2(\A[620] ), .ZN(new_n12558_));
  NOR2_X1    g11556(.A1(new_n12554_), .A2(new_n12558_), .ZN(new_n12559_));
  OAI22_X1   g11557(.A1(new_n12559_), .A2(\A[621] ), .B1(new_n12556_), .B2(new_n12554_), .ZN(new_n12560_));
  INV_X1     g11558(.I(\A[624] ), .ZN(new_n12561_));
  INV_X1     g11559(.I(\A[622] ), .ZN(new_n12562_));
  NAND2_X1   g11560(.A1(new_n12562_), .A2(\A[623] ), .ZN(new_n12563_));
  NOR2_X1    g11561(.A1(new_n12562_), .A2(\A[623] ), .ZN(new_n12564_));
  NOR2_X1    g11562(.A1(new_n12564_), .A2(new_n12561_), .ZN(new_n12565_));
  INV_X1     g11563(.I(\A[623] ), .ZN(new_n12566_));
  NAND2_X1   g11564(.A1(new_n12566_), .A2(\A[622] ), .ZN(new_n12567_));
  NAND2_X1   g11565(.A1(new_n12563_), .A2(new_n12567_), .ZN(new_n12568_));
  AOI22_X1   g11566(.A1(new_n12568_), .A2(new_n12561_), .B1(new_n12565_), .B2(new_n12563_), .ZN(new_n12569_));
  XNOR2_X1   g11567(.A1(new_n12569_), .A2(new_n12560_), .ZN(new_n12570_));
  NOR2_X1    g11568(.A1(new_n12566_), .A2(\A[622] ), .ZN(new_n12571_));
  NOR2_X1    g11569(.A1(new_n12571_), .A2(new_n12564_), .ZN(new_n12572_));
  NOR2_X1    g11570(.A1(new_n12562_), .A2(new_n12566_), .ZN(new_n12573_));
  INV_X1     g11571(.I(new_n12573_), .ZN(new_n12574_));
  OAI21_X1   g11572(.A1(new_n12572_), .A2(new_n12561_), .B(new_n12574_), .ZN(new_n12575_));
  NAND2_X1   g11573(.A1(new_n12557_), .A2(\A[620] ), .ZN(new_n12576_));
  NAND2_X1   g11574(.A1(new_n12576_), .A2(new_n12555_), .ZN(new_n12577_));
  NOR2_X1    g11575(.A1(new_n12557_), .A2(new_n12553_), .ZN(new_n12578_));
  AOI21_X1   g11576(.A1(new_n12577_), .A2(\A[621] ), .B(new_n12578_), .ZN(new_n12579_));
  INV_X1     g11577(.I(new_n12579_), .ZN(new_n12580_));
  INV_X1     g11578(.I(new_n12560_), .ZN(new_n12581_));
  NOR2_X1    g11579(.A1(new_n12581_), .A2(new_n12569_), .ZN(new_n12582_));
  NAND3_X1   g11580(.A1(new_n12582_), .A2(new_n12575_), .A3(new_n12580_), .ZN(new_n12583_));
  NAND2_X1   g11581(.A1(new_n12583_), .A2(new_n12570_), .ZN(new_n12584_));
  XOR2_X1    g11582(.A1(new_n12552_), .A2(new_n12584_), .Z(new_n12585_));
  INV_X1     g11583(.I(\A[614] ), .ZN(new_n12586_));
  NOR2_X1    g11584(.A1(new_n12586_), .A2(\A[613] ), .ZN(new_n12587_));
  NAND2_X1   g11585(.A1(new_n12586_), .A2(\A[613] ), .ZN(new_n12588_));
  NAND2_X1   g11586(.A1(new_n12588_), .A2(\A[615] ), .ZN(new_n12589_));
  INV_X1     g11587(.I(\A[613] ), .ZN(new_n12590_));
  NOR2_X1    g11588(.A1(new_n12590_), .A2(\A[614] ), .ZN(new_n12591_));
  NOR2_X1    g11589(.A1(new_n12587_), .A2(new_n12591_), .ZN(new_n12592_));
  OAI22_X1   g11590(.A1(new_n12592_), .A2(\A[615] ), .B1(new_n12589_), .B2(new_n12587_), .ZN(new_n12593_));
  INV_X1     g11591(.I(\A[618] ), .ZN(new_n12594_));
  INV_X1     g11592(.I(\A[616] ), .ZN(new_n12595_));
  NAND2_X1   g11593(.A1(new_n12595_), .A2(\A[617] ), .ZN(new_n12596_));
  NOR2_X1    g11594(.A1(new_n12595_), .A2(\A[617] ), .ZN(new_n12597_));
  NOR2_X1    g11595(.A1(new_n12597_), .A2(new_n12594_), .ZN(new_n12598_));
  INV_X1     g11596(.I(\A[617] ), .ZN(new_n12599_));
  NAND2_X1   g11597(.A1(new_n12599_), .A2(\A[616] ), .ZN(new_n12600_));
  NAND2_X1   g11598(.A1(new_n12596_), .A2(new_n12600_), .ZN(new_n12601_));
  AOI22_X1   g11599(.A1(new_n12601_), .A2(new_n12594_), .B1(new_n12598_), .B2(new_n12596_), .ZN(new_n12602_));
  XNOR2_X1   g11600(.A1(new_n12602_), .A2(new_n12593_), .ZN(new_n12603_));
  NOR2_X1    g11601(.A1(new_n12599_), .A2(\A[616] ), .ZN(new_n12604_));
  NOR2_X1    g11602(.A1(new_n12604_), .A2(new_n12597_), .ZN(new_n12605_));
  NOR2_X1    g11603(.A1(new_n12595_), .A2(new_n12599_), .ZN(new_n12606_));
  INV_X1     g11604(.I(new_n12606_), .ZN(new_n12607_));
  OAI21_X1   g11605(.A1(new_n12605_), .A2(new_n12594_), .B(new_n12607_), .ZN(new_n12608_));
  NAND2_X1   g11606(.A1(new_n12590_), .A2(\A[614] ), .ZN(new_n12609_));
  NAND2_X1   g11607(.A1(new_n12609_), .A2(new_n12588_), .ZN(new_n12610_));
  NOR2_X1    g11608(.A1(new_n12590_), .A2(new_n12586_), .ZN(new_n12611_));
  AOI21_X1   g11609(.A1(new_n12610_), .A2(\A[615] ), .B(new_n12611_), .ZN(new_n12612_));
  INV_X1     g11610(.I(new_n12612_), .ZN(new_n12613_));
  INV_X1     g11611(.I(new_n12593_), .ZN(new_n12614_));
  NOR2_X1    g11612(.A1(new_n12614_), .A2(new_n12602_), .ZN(new_n12615_));
  NAND3_X1   g11613(.A1(new_n12615_), .A2(new_n12608_), .A3(new_n12613_), .ZN(new_n12616_));
  NAND2_X1   g11614(.A1(new_n12616_), .A2(new_n12603_), .ZN(new_n12617_));
  INV_X1     g11615(.I(\A[608] ), .ZN(new_n12618_));
  NOR2_X1    g11616(.A1(new_n12618_), .A2(\A[607] ), .ZN(new_n12619_));
  NAND2_X1   g11617(.A1(new_n12618_), .A2(\A[607] ), .ZN(new_n12620_));
  NAND2_X1   g11618(.A1(new_n12620_), .A2(\A[609] ), .ZN(new_n12621_));
  INV_X1     g11619(.I(\A[607] ), .ZN(new_n12622_));
  NOR2_X1    g11620(.A1(new_n12622_), .A2(\A[608] ), .ZN(new_n12623_));
  NOR2_X1    g11621(.A1(new_n12619_), .A2(new_n12623_), .ZN(new_n12624_));
  OAI22_X1   g11622(.A1(new_n12624_), .A2(\A[609] ), .B1(new_n12621_), .B2(new_n12619_), .ZN(new_n12625_));
  INV_X1     g11623(.I(\A[612] ), .ZN(new_n12626_));
  INV_X1     g11624(.I(\A[610] ), .ZN(new_n12627_));
  NAND2_X1   g11625(.A1(new_n12627_), .A2(\A[611] ), .ZN(new_n12628_));
  NOR2_X1    g11626(.A1(new_n12627_), .A2(\A[611] ), .ZN(new_n12629_));
  NOR2_X1    g11627(.A1(new_n12629_), .A2(new_n12626_), .ZN(new_n12630_));
  INV_X1     g11628(.I(\A[611] ), .ZN(new_n12631_));
  NAND2_X1   g11629(.A1(new_n12631_), .A2(\A[610] ), .ZN(new_n12632_));
  NAND2_X1   g11630(.A1(new_n12628_), .A2(new_n12632_), .ZN(new_n12633_));
  AOI22_X1   g11631(.A1(new_n12633_), .A2(new_n12626_), .B1(new_n12630_), .B2(new_n12628_), .ZN(new_n12634_));
  XNOR2_X1   g11632(.A1(new_n12634_), .A2(new_n12625_), .ZN(new_n12635_));
  NOR2_X1    g11633(.A1(new_n12631_), .A2(\A[610] ), .ZN(new_n12636_));
  NOR2_X1    g11634(.A1(new_n12636_), .A2(new_n12629_), .ZN(new_n12637_));
  NOR2_X1    g11635(.A1(new_n12627_), .A2(new_n12631_), .ZN(new_n12638_));
  INV_X1     g11636(.I(new_n12638_), .ZN(new_n12639_));
  OAI21_X1   g11637(.A1(new_n12637_), .A2(new_n12626_), .B(new_n12639_), .ZN(new_n12640_));
  NAND2_X1   g11638(.A1(new_n12622_), .A2(\A[608] ), .ZN(new_n12641_));
  NAND2_X1   g11639(.A1(new_n12641_), .A2(new_n12620_), .ZN(new_n12642_));
  NOR2_X1    g11640(.A1(new_n12622_), .A2(new_n12618_), .ZN(new_n12643_));
  AOI21_X1   g11641(.A1(new_n12642_), .A2(\A[609] ), .B(new_n12643_), .ZN(new_n12644_));
  INV_X1     g11642(.I(new_n12644_), .ZN(new_n12645_));
  INV_X1     g11643(.I(new_n12625_), .ZN(new_n12646_));
  NOR2_X1    g11644(.A1(new_n12646_), .A2(new_n12634_), .ZN(new_n12647_));
  NAND3_X1   g11645(.A1(new_n12647_), .A2(new_n12640_), .A3(new_n12645_), .ZN(new_n12648_));
  NAND2_X1   g11646(.A1(new_n12648_), .A2(new_n12635_), .ZN(new_n12649_));
  XOR2_X1    g11647(.A1(new_n12617_), .A2(new_n12649_), .Z(new_n12650_));
  XOR2_X1    g11648(.A1(new_n12585_), .A2(new_n12650_), .Z(new_n12651_));
  XOR2_X1    g11649(.A1(new_n12651_), .A2(new_n12520_), .Z(new_n12652_));
  INV_X1     g11650(.I(\A[602] ), .ZN(new_n12653_));
  NOR2_X1    g11651(.A1(new_n12653_), .A2(\A[601] ), .ZN(new_n12654_));
  NAND2_X1   g11652(.A1(new_n12653_), .A2(\A[601] ), .ZN(new_n12655_));
  NAND2_X1   g11653(.A1(new_n12655_), .A2(\A[603] ), .ZN(new_n12656_));
  INV_X1     g11654(.I(\A[601] ), .ZN(new_n12657_));
  NOR2_X1    g11655(.A1(new_n12657_), .A2(\A[602] ), .ZN(new_n12658_));
  NOR2_X1    g11656(.A1(new_n12654_), .A2(new_n12658_), .ZN(new_n12659_));
  OAI22_X1   g11657(.A1(new_n12659_), .A2(\A[603] ), .B1(new_n12656_), .B2(new_n12654_), .ZN(new_n12660_));
  INV_X1     g11658(.I(\A[606] ), .ZN(new_n12661_));
  INV_X1     g11659(.I(\A[604] ), .ZN(new_n12662_));
  NAND2_X1   g11660(.A1(new_n12662_), .A2(\A[605] ), .ZN(new_n12663_));
  NOR2_X1    g11661(.A1(new_n12662_), .A2(\A[605] ), .ZN(new_n12664_));
  NOR2_X1    g11662(.A1(new_n12664_), .A2(new_n12661_), .ZN(new_n12665_));
  INV_X1     g11663(.I(\A[605] ), .ZN(new_n12666_));
  NAND2_X1   g11664(.A1(new_n12666_), .A2(\A[604] ), .ZN(new_n12667_));
  NAND2_X1   g11665(.A1(new_n12663_), .A2(new_n12667_), .ZN(new_n12668_));
  AOI22_X1   g11666(.A1(new_n12668_), .A2(new_n12661_), .B1(new_n12665_), .B2(new_n12663_), .ZN(new_n12669_));
  XNOR2_X1   g11667(.A1(new_n12669_), .A2(new_n12660_), .ZN(new_n12670_));
  NOR2_X1    g11668(.A1(new_n12666_), .A2(\A[604] ), .ZN(new_n12671_));
  NOR2_X1    g11669(.A1(new_n12671_), .A2(new_n12664_), .ZN(new_n12672_));
  NOR2_X1    g11670(.A1(new_n12662_), .A2(new_n12666_), .ZN(new_n12673_));
  INV_X1     g11671(.I(new_n12673_), .ZN(new_n12674_));
  OAI21_X1   g11672(.A1(new_n12672_), .A2(new_n12661_), .B(new_n12674_), .ZN(new_n12675_));
  NAND2_X1   g11673(.A1(new_n12657_), .A2(\A[602] ), .ZN(new_n12676_));
  NAND2_X1   g11674(.A1(new_n12676_), .A2(new_n12655_), .ZN(new_n12677_));
  NOR2_X1    g11675(.A1(new_n12657_), .A2(new_n12653_), .ZN(new_n12678_));
  AOI21_X1   g11676(.A1(new_n12677_), .A2(\A[603] ), .B(new_n12678_), .ZN(new_n12679_));
  INV_X1     g11677(.I(new_n12679_), .ZN(new_n12680_));
  INV_X1     g11678(.I(new_n12660_), .ZN(new_n12681_));
  NOR2_X1    g11679(.A1(new_n12681_), .A2(new_n12669_), .ZN(new_n12682_));
  NAND3_X1   g11680(.A1(new_n12682_), .A2(new_n12675_), .A3(new_n12680_), .ZN(new_n12683_));
  NAND2_X1   g11681(.A1(new_n12683_), .A2(new_n12670_), .ZN(new_n12684_));
  INV_X1     g11682(.I(\A[596] ), .ZN(new_n12685_));
  NOR2_X1    g11683(.A1(new_n12685_), .A2(\A[595] ), .ZN(new_n12686_));
  NAND2_X1   g11684(.A1(new_n12685_), .A2(\A[595] ), .ZN(new_n12687_));
  NAND2_X1   g11685(.A1(new_n12687_), .A2(\A[597] ), .ZN(new_n12688_));
  INV_X1     g11686(.I(\A[595] ), .ZN(new_n12689_));
  NOR2_X1    g11687(.A1(new_n12689_), .A2(\A[596] ), .ZN(new_n12690_));
  NOR2_X1    g11688(.A1(new_n12686_), .A2(new_n12690_), .ZN(new_n12691_));
  OAI22_X1   g11689(.A1(new_n12691_), .A2(\A[597] ), .B1(new_n12688_), .B2(new_n12686_), .ZN(new_n12692_));
  INV_X1     g11690(.I(\A[600] ), .ZN(new_n12693_));
  INV_X1     g11691(.I(\A[598] ), .ZN(new_n12694_));
  NAND2_X1   g11692(.A1(new_n12694_), .A2(\A[599] ), .ZN(new_n12695_));
  NOR2_X1    g11693(.A1(new_n12694_), .A2(\A[599] ), .ZN(new_n12696_));
  NOR2_X1    g11694(.A1(new_n12696_), .A2(new_n12693_), .ZN(new_n12697_));
  INV_X1     g11695(.I(\A[599] ), .ZN(new_n12698_));
  NAND2_X1   g11696(.A1(new_n12698_), .A2(\A[598] ), .ZN(new_n12699_));
  NAND2_X1   g11697(.A1(new_n12695_), .A2(new_n12699_), .ZN(new_n12700_));
  AOI22_X1   g11698(.A1(new_n12700_), .A2(new_n12693_), .B1(new_n12697_), .B2(new_n12695_), .ZN(new_n12701_));
  XNOR2_X1   g11699(.A1(new_n12701_), .A2(new_n12692_), .ZN(new_n12702_));
  NOR2_X1    g11700(.A1(new_n12698_), .A2(\A[598] ), .ZN(new_n12703_));
  NOR2_X1    g11701(.A1(new_n12703_), .A2(new_n12696_), .ZN(new_n12704_));
  NOR2_X1    g11702(.A1(new_n12694_), .A2(new_n12698_), .ZN(new_n12705_));
  INV_X1     g11703(.I(new_n12705_), .ZN(new_n12706_));
  OAI21_X1   g11704(.A1(new_n12704_), .A2(new_n12693_), .B(new_n12706_), .ZN(new_n12707_));
  NAND2_X1   g11705(.A1(new_n12689_), .A2(\A[596] ), .ZN(new_n12708_));
  NAND2_X1   g11706(.A1(new_n12708_), .A2(new_n12687_), .ZN(new_n12709_));
  NOR2_X1    g11707(.A1(new_n12689_), .A2(new_n12685_), .ZN(new_n12710_));
  AOI21_X1   g11708(.A1(new_n12709_), .A2(\A[597] ), .B(new_n12710_), .ZN(new_n12711_));
  INV_X1     g11709(.I(new_n12711_), .ZN(new_n12712_));
  INV_X1     g11710(.I(new_n12692_), .ZN(new_n12713_));
  NOR2_X1    g11711(.A1(new_n12713_), .A2(new_n12701_), .ZN(new_n12714_));
  NAND3_X1   g11712(.A1(new_n12714_), .A2(new_n12707_), .A3(new_n12712_), .ZN(new_n12715_));
  NAND2_X1   g11713(.A1(new_n12715_), .A2(new_n12702_), .ZN(new_n12716_));
  XOR2_X1    g11714(.A1(new_n12684_), .A2(new_n12716_), .Z(new_n12717_));
  INV_X1     g11715(.I(\A[590] ), .ZN(new_n12718_));
  NOR2_X1    g11716(.A1(new_n12718_), .A2(\A[589] ), .ZN(new_n12719_));
  NAND2_X1   g11717(.A1(new_n12718_), .A2(\A[589] ), .ZN(new_n12720_));
  NAND2_X1   g11718(.A1(new_n12720_), .A2(\A[591] ), .ZN(new_n12721_));
  INV_X1     g11719(.I(\A[589] ), .ZN(new_n12722_));
  NOR2_X1    g11720(.A1(new_n12722_), .A2(\A[590] ), .ZN(new_n12723_));
  NOR2_X1    g11721(.A1(new_n12719_), .A2(new_n12723_), .ZN(new_n12724_));
  OAI22_X1   g11722(.A1(new_n12724_), .A2(\A[591] ), .B1(new_n12721_), .B2(new_n12719_), .ZN(new_n12725_));
  INV_X1     g11723(.I(\A[594] ), .ZN(new_n12726_));
  INV_X1     g11724(.I(\A[592] ), .ZN(new_n12727_));
  NAND2_X1   g11725(.A1(new_n12727_), .A2(\A[593] ), .ZN(new_n12728_));
  NOR2_X1    g11726(.A1(new_n12727_), .A2(\A[593] ), .ZN(new_n12729_));
  NOR2_X1    g11727(.A1(new_n12729_), .A2(new_n12726_), .ZN(new_n12730_));
  INV_X1     g11728(.I(\A[593] ), .ZN(new_n12731_));
  NAND2_X1   g11729(.A1(new_n12731_), .A2(\A[592] ), .ZN(new_n12732_));
  NAND2_X1   g11730(.A1(new_n12728_), .A2(new_n12732_), .ZN(new_n12733_));
  AOI22_X1   g11731(.A1(new_n12733_), .A2(new_n12726_), .B1(new_n12730_), .B2(new_n12728_), .ZN(new_n12734_));
  XNOR2_X1   g11732(.A1(new_n12734_), .A2(new_n12725_), .ZN(new_n12735_));
  NOR2_X1    g11733(.A1(new_n12731_), .A2(\A[592] ), .ZN(new_n12736_));
  NOR2_X1    g11734(.A1(new_n12736_), .A2(new_n12729_), .ZN(new_n12737_));
  NOR2_X1    g11735(.A1(new_n12727_), .A2(new_n12731_), .ZN(new_n12738_));
  INV_X1     g11736(.I(new_n12738_), .ZN(new_n12739_));
  OAI21_X1   g11737(.A1(new_n12737_), .A2(new_n12726_), .B(new_n12739_), .ZN(new_n12740_));
  NAND2_X1   g11738(.A1(new_n12722_), .A2(\A[590] ), .ZN(new_n12741_));
  NAND2_X1   g11739(.A1(new_n12741_), .A2(new_n12720_), .ZN(new_n12742_));
  NOR2_X1    g11740(.A1(new_n12722_), .A2(new_n12718_), .ZN(new_n12743_));
  AOI21_X1   g11741(.A1(new_n12742_), .A2(\A[591] ), .B(new_n12743_), .ZN(new_n12744_));
  INV_X1     g11742(.I(new_n12744_), .ZN(new_n12745_));
  INV_X1     g11743(.I(new_n12725_), .ZN(new_n12746_));
  NOR2_X1    g11744(.A1(new_n12746_), .A2(new_n12734_), .ZN(new_n12747_));
  NAND3_X1   g11745(.A1(new_n12747_), .A2(new_n12740_), .A3(new_n12745_), .ZN(new_n12748_));
  NAND2_X1   g11746(.A1(new_n12748_), .A2(new_n12735_), .ZN(new_n12749_));
  INV_X1     g11747(.I(\A[585] ), .ZN(new_n12750_));
  INV_X1     g11748(.I(\A[583] ), .ZN(new_n12751_));
  NAND2_X1   g11749(.A1(new_n12751_), .A2(\A[584] ), .ZN(new_n12752_));
  NOR2_X1    g11750(.A1(new_n12751_), .A2(\A[584] ), .ZN(new_n12753_));
  NOR2_X1    g11751(.A1(new_n12753_), .A2(new_n12750_), .ZN(new_n12754_));
  INV_X1     g11752(.I(\A[584] ), .ZN(new_n12755_));
  NAND2_X1   g11753(.A1(new_n12755_), .A2(\A[583] ), .ZN(new_n12756_));
  NAND2_X1   g11754(.A1(new_n12752_), .A2(new_n12756_), .ZN(new_n12757_));
  AOI22_X1   g11755(.A1(new_n12757_), .A2(new_n12750_), .B1(new_n12754_), .B2(new_n12752_), .ZN(new_n12758_));
  INV_X1     g11756(.I(\A[588] ), .ZN(new_n12759_));
  INV_X1     g11757(.I(\A[586] ), .ZN(new_n12760_));
  NAND2_X1   g11758(.A1(new_n12760_), .A2(\A[587] ), .ZN(new_n12761_));
  NOR2_X1    g11759(.A1(new_n12760_), .A2(\A[587] ), .ZN(new_n12762_));
  NOR2_X1    g11760(.A1(new_n12762_), .A2(new_n12759_), .ZN(new_n12763_));
  INV_X1     g11761(.I(\A[587] ), .ZN(new_n12764_));
  NAND2_X1   g11762(.A1(new_n12764_), .A2(\A[586] ), .ZN(new_n12765_));
  NAND2_X1   g11763(.A1(new_n12761_), .A2(new_n12765_), .ZN(new_n12766_));
  AOI22_X1   g11764(.A1(new_n12766_), .A2(new_n12759_), .B1(new_n12763_), .B2(new_n12761_), .ZN(new_n12767_));
  XOR2_X1    g11765(.A1(new_n12758_), .A2(new_n12767_), .Z(new_n12768_));
  NOR2_X1    g11766(.A1(new_n12764_), .A2(\A[586] ), .ZN(new_n12769_));
  NOR2_X1    g11767(.A1(new_n12769_), .A2(new_n12762_), .ZN(new_n12770_));
  NOR2_X1    g11768(.A1(new_n12760_), .A2(new_n12764_), .ZN(new_n12771_));
  INV_X1     g11769(.I(new_n12771_), .ZN(new_n12772_));
  OAI21_X1   g11770(.A1(new_n12770_), .A2(new_n12759_), .B(new_n12772_), .ZN(new_n12773_));
  NOR2_X1    g11771(.A1(new_n12751_), .A2(new_n12755_), .ZN(new_n12774_));
  AOI21_X1   g11772(.A1(new_n12757_), .A2(\A[585] ), .B(new_n12774_), .ZN(new_n12775_));
  INV_X1     g11773(.I(new_n12775_), .ZN(new_n12776_));
  NOR2_X1    g11774(.A1(new_n12758_), .A2(new_n12767_), .ZN(new_n12777_));
  NAND3_X1   g11775(.A1(new_n12777_), .A2(new_n12773_), .A3(new_n12776_), .ZN(new_n12778_));
  NAND2_X1   g11776(.A1(new_n12768_), .A2(new_n12778_), .ZN(new_n12779_));
  XOR2_X1    g11777(.A1(new_n12749_), .A2(new_n12779_), .Z(new_n12780_));
  XOR2_X1    g11778(.A1(new_n12717_), .A2(new_n12780_), .Z(new_n12781_));
  INV_X1     g11779(.I(\A[578] ), .ZN(new_n12782_));
  NOR2_X1    g11780(.A1(new_n12782_), .A2(\A[577] ), .ZN(new_n12783_));
  NAND2_X1   g11781(.A1(new_n12782_), .A2(\A[577] ), .ZN(new_n12784_));
  NAND2_X1   g11782(.A1(new_n12784_), .A2(\A[579] ), .ZN(new_n12785_));
  INV_X1     g11783(.I(\A[577] ), .ZN(new_n12786_));
  NOR2_X1    g11784(.A1(new_n12786_), .A2(\A[578] ), .ZN(new_n12787_));
  NOR2_X1    g11785(.A1(new_n12783_), .A2(new_n12787_), .ZN(new_n12788_));
  OAI22_X1   g11786(.A1(new_n12788_), .A2(\A[579] ), .B1(new_n12785_), .B2(new_n12783_), .ZN(new_n12789_));
  INV_X1     g11787(.I(\A[582] ), .ZN(new_n12790_));
  INV_X1     g11788(.I(\A[580] ), .ZN(new_n12791_));
  NAND2_X1   g11789(.A1(new_n12791_), .A2(\A[581] ), .ZN(new_n12792_));
  NOR2_X1    g11790(.A1(new_n12791_), .A2(\A[581] ), .ZN(new_n12793_));
  NOR2_X1    g11791(.A1(new_n12793_), .A2(new_n12790_), .ZN(new_n12794_));
  INV_X1     g11792(.I(\A[581] ), .ZN(new_n12795_));
  NAND2_X1   g11793(.A1(new_n12795_), .A2(\A[580] ), .ZN(new_n12796_));
  NAND2_X1   g11794(.A1(new_n12792_), .A2(new_n12796_), .ZN(new_n12797_));
  AOI22_X1   g11795(.A1(new_n12797_), .A2(new_n12790_), .B1(new_n12794_), .B2(new_n12792_), .ZN(new_n12798_));
  XNOR2_X1   g11796(.A1(new_n12798_), .A2(new_n12789_), .ZN(new_n12799_));
  NOR2_X1    g11797(.A1(new_n12795_), .A2(\A[580] ), .ZN(new_n12800_));
  NOR2_X1    g11798(.A1(new_n12800_), .A2(new_n12793_), .ZN(new_n12801_));
  NOR2_X1    g11799(.A1(new_n12791_), .A2(new_n12795_), .ZN(new_n12802_));
  INV_X1     g11800(.I(new_n12802_), .ZN(new_n12803_));
  OAI21_X1   g11801(.A1(new_n12801_), .A2(new_n12790_), .B(new_n12803_), .ZN(new_n12804_));
  NAND2_X1   g11802(.A1(new_n12786_), .A2(\A[578] ), .ZN(new_n12805_));
  NAND2_X1   g11803(.A1(new_n12805_), .A2(new_n12784_), .ZN(new_n12806_));
  NOR2_X1    g11804(.A1(new_n12786_), .A2(new_n12782_), .ZN(new_n12807_));
  AOI21_X1   g11805(.A1(new_n12806_), .A2(\A[579] ), .B(new_n12807_), .ZN(new_n12808_));
  INV_X1     g11806(.I(new_n12808_), .ZN(new_n12809_));
  INV_X1     g11807(.I(new_n12789_), .ZN(new_n12810_));
  NOR2_X1    g11808(.A1(new_n12810_), .A2(new_n12798_), .ZN(new_n12811_));
  NAND3_X1   g11809(.A1(new_n12811_), .A2(new_n12804_), .A3(new_n12809_), .ZN(new_n12812_));
  NAND2_X1   g11810(.A1(new_n12812_), .A2(new_n12799_), .ZN(new_n12813_));
  INV_X1     g11811(.I(\A[572] ), .ZN(new_n12814_));
  NOR2_X1    g11812(.A1(new_n12814_), .A2(\A[571] ), .ZN(new_n12815_));
  NAND2_X1   g11813(.A1(new_n12814_), .A2(\A[571] ), .ZN(new_n12816_));
  NAND2_X1   g11814(.A1(new_n12816_), .A2(\A[573] ), .ZN(new_n12817_));
  INV_X1     g11815(.I(\A[571] ), .ZN(new_n12818_));
  NOR2_X1    g11816(.A1(new_n12818_), .A2(\A[572] ), .ZN(new_n12819_));
  NOR2_X1    g11817(.A1(new_n12815_), .A2(new_n12819_), .ZN(new_n12820_));
  OAI22_X1   g11818(.A1(new_n12820_), .A2(\A[573] ), .B1(new_n12817_), .B2(new_n12815_), .ZN(new_n12821_));
  INV_X1     g11819(.I(\A[576] ), .ZN(new_n12822_));
  INV_X1     g11820(.I(\A[574] ), .ZN(new_n12823_));
  NAND2_X1   g11821(.A1(new_n12823_), .A2(\A[575] ), .ZN(new_n12824_));
  NOR2_X1    g11822(.A1(new_n12823_), .A2(\A[575] ), .ZN(new_n12825_));
  NOR2_X1    g11823(.A1(new_n12825_), .A2(new_n12822_), .ZN(new_n12826_));
  INV_X1     g11824(.I(\A[575] ), .ZN(new_n12827_));
  NAND2_X1   g11825(.A1(new_n12827_), .A2(\A[574] ), .ZN(new_n12828_));
  NAND2_X1   g11826(.A1(new_n12824_), .A2(new_n12828_), .ZN(new_n12829_));
  AOI22_X1   g11827(.A1(new_n12829_), .A2(new_n12822_), .B1(new_n12826_), .B2(new_n12824_), .ZN(new_n12830_));
  XNOR2_X1   g11828(.A1(new_n12830_), .A2(new_n12821_), .ZN(new_n12831_));
  NOR2_X1    g11829(.A1(new_n12827_), .A2(\A[574] ), .ZN(new_n12832_));
  NOR2_X1    g11830(.A1(new_n12832_), .A2(new_n12825_), .ZN(new_n12833_));
  NOR2_X1    g11831(.A1(new_n12823_), .A2(new_n12827_), .ZN(new_n12834_));
  INV_X1     g11832(.I(new_n12834_), .ZN(new_n12835_));
  OAI21_X1   g11833(.A1(new_n12833_), .A2(new_n12822_), .B(new_n12835_), .ZN(new_n12836_));
  NAND2_X1   g11834(.A1(new_n12818_), .A2(\A[572] ), .ZN(new_n12837_));
  NAND2_X1   g11835(.A1(new_n12837_), .A2(new_n12816_), .ZN(new_n12838_));
  NOR2_X1    g11836(.A1(new_n12818_), .A2(new_n12814_), .ZN(new_n12839_));
  AOI21_X1   g11837(.A1(new_n12838_), .A2(\A[573] ), .B(new_n12839_), .ZN(new_n12840_));
  INV_X1     g11838(.I(new_n12840_), .ZN(new_n12841_));
  INV_X1     g11839(.I(new_n12821_), .ZN(new_n12842_));
  NOR2_X1    g11840(.A1(new_n12842_), .A2(new_n12830_), .ZN(new_n12843_));
  NAND3_X1   g11841(.A1(new_n12843_), .A2(new_n12836_), .A3(new_n12841_), .ZN(new_n12844_));
  NAND2_X1   g11842(.A1(new_n12844_), .A2(new_n12831_), .ZN(new_n12845_));
  XOR2_X1    g11843(.A1(new_n12813_), .A2(new_n12845_), .Z(new_n12846_));
  INV_X1     g11844(.I(\A[566] ), .ZN(new_n12847_));
  NOR2_X1    g11845(.A1(new_n12847_), .A2(\A[565] ), .ZN(new_n12848_));
  NAND2_X1   g11846(.A1(new_n12847_), .A2(\A[565] ), .ZN(new_n12849_));
  NAND2_X1   g11847(.A1(new_n12849_), .A2(\A[567] ), .ZN(new_n12850_));
  INV_X1     g11848(.I(\A[565] ), .ZN(new_n12851_));
  NOR2_X1    g11849(.A1(new_n12851_), .A2(\A[566] ), .ZN(new_n12852_));
  NOR2_X1    g11850(.A1(new_n12848_), .A2(new_n12852_), .ZN(new_n12853_));
  OAI22_X1   g11851(.A1(new_n12853_), .A2(\A[567] ), .B1(new_n12850_), .B2(new_n12848_), .ZN(new_n12854_));
  INV_X1     g11852(.I(\A[570] ), .ZN(new_n12855_));
  INV_X1     g11853(.I(\A[568] ), .ZN(new_n12856_));
  NAND2_X1   g11854(.A1(new_n12856_), .A2(\A[569] ), .ZN(new_n12857_));
  NOR2_X1    g11855(.A1(new_n12856_), .A2(\A[569] ), .ZN(new_n12858_));
  NOR2_X1    g11856(.A1(new_n12858_), .A2(new_n12855_), .ZN(new_n12859_));
  INV_X1     g11857(.I(\A[569] ), .ZN(new_n12860_));
  NAND2_X1   g11858(.A1(new_n12860_), .A2(\A[568] ), .ZN(new_n12861_));
  NAND2_X1   g11859(.A1(new_n12857_), .A2(new_n12861_), .ZN(new_n12862_));
  AOI22_X1   g11860(.A1(new_n12862_), .A2(new_n12855_), .B1(new_n12859_), .B2(new_n12857_), .ZN(new_n12863_));
  XNOR2_X1   g11861(.A1(new_n12863_), .A2(new_n12854_), .ZN(new_n12864_));
  NOR2_X1    g11862(.A1(new_n12860_), .A2(\A[568] ), .ZN(new_n12865_));
  NOR2_X1    g11863(.A1(new_n12865_), .A2(new_n12858_), .ZN(new_n12866_));
  NOR2_X1    g11864(.A1(new_n12856_), .A2(new_n12860_), .ZN(new_n12867_));
  INV_X1     g11865(.I(new_n12867_), .ZN(new_n12868_));
  OAI21_X1   g11866(.A1(new_n12866_), .A2(new_n12855_), .B(new_n12868_), .ZN(new_n12869_));
  NAND2_X1   g11867(.A1(new_n12851_), .A2(\A[566] ), .ZN(new_n12870_));
  NAND2_X1   g11868(.A1(new_n12870_), .A2(new_n12849_), .ZN(new_n12871_));
  NOR2_X1    g11869(.A1(new_n12851_), .A2(new_n12847_), .ZN(new_n12872_));
  AOI21_X1   g11870(.A1(new_n12871_), .A2(\A[567] ), .B(new_n12872_), .ZN(new_n12873_));
  INV_X1     g11871(.I(new_n12873_), .ZN(new_n12874_));
  INV_X1     g11872(.I(new_n12854_), .ZN(new_n12875_));
  NOR2_X1    g11873(.A1(new_n12875_), .A2(new_n12863_), .ZN(new_n12876_));
  NAND3_X1   g11874(.A1(new_n12876_), .A2(new_n12869_), .A3(new_n12874_), .ZN(new_n12877_));
  NAND2_X1   g11875(.A1(new_n12877_), .A2(new_n12864_), .ZN(new_n12878_));
  INV_X1     g11876(.I(\A[561] ), .ZN(new_n12879_));
  INV_X1     g11877(.I(\A[559] ), .ZN(new_n12880_));
  NAND2_X1   g11878(.A1(new_n12880_), .A2(\A[560] ), .ZN(new_n12881_));
  NOR2_X1    g11879(.A1(new_n12880_), .A2(\A[560] ), .ZN(new_n12882_));
  NOR2_X1    g11880(.A1(new_n12882_), .A2(new_n12879_), .ZN(new_n12883_));
  INV_X1     g11881(.I(\A[560] ), .ZN(new_n12884_));
  NAND2_X1   g11882(.A1(new_n12884_), .A2(\A[559] ), .ZN(new_n12885_));
  NAND2_X1   g11883(.A1(new_n12881_), .A2(new_n12885_), .ZN(new_n12886_));
  AOI22_X1   g11884(.A1(new_n12886_), .A2(new_n12879_), .B1(new_n12883_), .B2(new_n12881_), .ZN(new_n12887_));
  INV_X1     g11885(.I(\A[564] ), .ZN(new_n12888_));
  INV_X1     g11886(.I(\A[562] ), .ZN(new_n12889_));
  NAND2_X1   g11887(.A1(new_n12889_), .A2(\A[563] ), .ZN(new_n12890_));
  NOR2_X1    g11888(.A1(new_n12889_), .A2(\A[563] ), .ZN(new_n12891_));
  NOR2_X1    g11889(.A1(new_n12891_), .A2(new_n12888_), .ZN(new_n12892_));
  INV_X1     g11890(.I(\A[563] ), .ZN(new_n12893_));
  NAND2_X1   g11891(.A1(new_n12893_), .A2(\A[562] ), .ZN(new_n12894_));
  NAND2_X1   g11892(.A1(new_n12890_), .A2(new_n12894_), .ZN(new_n12895_));
  AOI22_X1   g11893(.A1(new_n12895_), .A2(new_n12888_), .B1(new_n12892_), .B2(new_n12890_), .ZN(new_n12896_));
  XOR2_X1    g11894(.A1(new_n12887_), .A2(new_n12896_), .Z(new_n12897_));
  NOR2_X1    g11895(.A1(new_n12893_), .A2(\A[562] ), .ZN(new_n12898_));
  NOR2_X1    g11896(.A1(new_n12898_), .A2(new_n12891_), .ZN(new_n12899_));
  NOR2_X1    g11897(.A1(new_n12889_), .A2(new_n12893_), .ZN(new_n12900_));
  INV_X1     g11898(.I(new_n12900_), .ZN(new_n12901_));
  OAI21_X1   g11899(.A1(new_n12899_), .A2(new_n12888_), .B(new_n12901_), .ZN(new_n12902_));
  NOR2_X1    g11900(.A1(new_n12880_), .A2(new_n12884_), .ZN(new_n12903_));
  AOI21_X1   g11901(.A1(new_n12886_), .A2(\A[561] ), .B(new_n12903_), .ZN(new_n12904_));
  INV_X1     g11902(.I(new_n12904_), .ZN(new_n12905_));
  NOR2_X1    g11903(.A1(new_n12887_), .A2(new_n12896_), .ZN(new_n12906_));
  NAND3_X1   g11904(.A1(new_n12906_), .A2(new_n12902_), .A3(new_n12905_), .ZN(new_n12907_));
  NAND2_X1   g11905(.A1(new_n12897_), .A2(new_n12907_), .ZN(new_n12908_));
  XOR2_X1    g11906(.A1(new_n12878_), .A2(new_n12908_), .Z(new_n12909_));
  XOR2_X1    g11907(.A1(new_n12846_), .A2(new_n12909_), .Z(new_n12910_));
  XOR2_X1    g11908(.A1(new_n12781_), .A2(new_n12910_), .Z(new_n12911_));
  XOR2_X1    g11909(.A1(new_n12652_), .A2(new_n12911_), .Z(new_n12912_));
  NAND2_X1   g11910(.A1(new_n12395_), .A2(new_n12912_), .ZN(new_n12913_));
  INV_X1     g11911(.I(new_n12913_), .ZN(new_n12914_));
  AOI21_X1   g11912(.A1(new_n12895_), .A2(\A[564] ), .B(new_n12900_), .ZN(new_n12915_));
  XOR2_X1    g11913(.A1(new_n12915_), .A2(new_n12904_), .Z(new_n12916_));
  XOR2_X1    g11914(.A1(new_n12916_), .A2(new_n12906_), .Z(new_n12917_));
  XOR2_X1    g11915(.A1(new_n12902_), .A2(new_n12904_), .Z(new_n12918_));
  INV_X1     g11916(.I(new_n12906_), .ZN(new_n12919_));
  NOR2_X1    g11917(.A1(new_n12915_), .A2(new_n12904_), .ZN(new_n12920_));
  INV_X1     g11918(.I(new_n12920_), .ZN(new_n12921_));
  OAI21_X1   g11919(.A1(new_n12918_), .A2(new_n12919_), .B(new_n12921_), .ZN(new_n12922_));
  NAND2_X1   g11920(.A1(new_n12922_), .A2(new_n12897_), .ZN(new_n12923_));
  NAND2_X1   g11921(.A1(new_n12917_), .A2(new_n12923_), .ZN(new_n12924_));
  AOI21_X1   g11922(.A1(new_n12862_), .A2(\A[570] ), .B(new_n12867_), .ZN(new_n12925_));
  XOR2_X1    g11923(.A1(new_n12925_), .A2(new_n12873_), .Z(new_n12926_));
  INV_X1     g11924(.I(new_n12863_), .ZN(new_n12927_));
  NAND2_X1   g11925(.A1(new_n12927_), .A2(new_n12854_), .ZN(new_n12928_));
  XOR2_X1    g11926(.A1(new_n12926_), .A2(new_n12928_), .Z(new_n12929_));
  INV_X1     g11927(.I(new_n12877_), .ZN(new_n12930_));
  NAND2_X1   g11928(.A1(new_n12864_), .A2(new_n12897_), .ZN(new_n12931_));
  NOR3_X1    g11929(.A1(new_n12929_), .A2(new_n12930_), .A3(new_n12931_), .ZN(new_n12932_));
  INV_X1     g11930(.I(new_n12907_), .ZN(new_n12933_));
  INV_X1     g11931(.I(new_n12864_), .ZN(new_n12934_));
  NOR2_X1    g11932(.A1(new_n12925_), .A2(new_n12873_), .ZN(new_n12935_));
  AOI21_X1   g11933(.A1(new_n12926_), .A2(new_n12876_), .B(new_n12935_), .ZN(new_n12936_));
  NOR2_X1    g11934(.A1(new_n12936_), .A2(new_n12934_), .ZN(new_n12937_));
  NOR2_X1    g11935(.A1(new_n12937_), .A2(new_n12933_), .ZN(new_n12938_));
  NAND2_X1   g11936(.A1(new_n12932_), .A2(new_n12938_), .ZN(new_n12939_));
  XNOR2_X1   g11937(.A1(new_n12887_), .A2(new_n12896_), .ZN(new_n12940_));
  NOR2_X1    g11938(.A1(new_n12934_), .A2(new_n12940_), .ZN(new_n12941_));
  NAND3_X1   g11939(.A1(new_n12941_), .A2(new_n12877_), .A3(new_n12907_), .ZN(new_n12942_));
  XOR2_X1    g11940(.A1(new_n12926_), .A2(new_n12876_), .Z(new_n12943_));
  XOR2_X1    g11941(.A1(new_n12869_), .A2(new_n12873_), .Z(new_n12944_));
  INV_X1     g11942(.I(new_n12935_), .ZN(new_n12945_));
  OAI21_X1   g11943(.A1(new_n12944_), .A2(new_n12928_), .B(new_n12945_), .ZN(new_n12946_));
  NAND2_X1   g11944(.A1(new_n12946_), .A2(new_n12864_), .ZN(new_n12947_));
  NAND2_X1   g11945(.A1(new_n12943_), .A2(new_n12947_), .ZN(new_n12948_));
  NAND2_X1   g11946(.A1(new_n12948_), .A2(new_n12942_), .ZN(new_n12949_));
  AOI21_X1   g11947(.A1(new_n12939_), .A2(new_n12949_), .B(new_n12924_), .ZN(new_n12950_));
  XOR2_X1    g11948(.A1(new_n12948_), .A2(new_n12942_), .Z(new_n12951_));
  AOI21_X1   g11949(.A1(new_n12951_), .A2(new_n12924_), .B(new_n12950_), .ZN(new_n12952_));
  XOR2_X1    g11950(.A1(new_n12836_), .A2(new_n12840_), .Z(new_n12953_));
  INV_X1     g11951(.I(new_n12830_), .ZN(new_n12954_));
  NAND2_X1   g11952(.A1(new_n12954_), .A2(new_n12821_), .ZN(new_n12955_));
  AOI21_X1   g11953(.A1(new_n12829_), .A2(\A[576] ), .B(new_n12834_), .ZN(new_n12956_));
  NOR2_X1    g11954(.A1(new_n12956_), .A2(new_n12840_), .ZN(new_n12957_));
  INV_X1     g11955(.I(new_n12957_), .ZN(new_n12958_));
  OAI21_X1   g11956(.A1(new_n12953_), .A2(new_n12955_), .B(new_n12958_), .ZN(new_n12959_));
  NAND2_X1   g11957(.A1(new_n12953_), .A2(new_n12843_), .ZN(new_n12960_));
  XOR2_X1    g11958(.A1(new_n12956_), .A2(new_n12840_), .Z(new_n12961_));
  NAND2_X1   g11959(.A1(new_n12961_), .A2(new_n12955_), .ZN(new_n12962_));
  AOI22_X1   g11960(.A1(new_n12959_), .A2(new_n12831_), .B1(new_n12960_), .B2(new_n12962_), .ZN(new_n12963_));
  XOR2_X1    g11961(.A1(new_n12804_), .A2(new_n12808_), .Z(new_n12964_));
  NAND2_X1   g11962(.A1(new_n12964_), .A2(new_n12811_), .ZN(new_n12965_));
  XNOR2_X1   g11963(.A1(new_n12804_), .A2(new_n12808_), .ZN(new_n12966_));
  INV_X1     g11964(.I(new_n12798_), .ZN(new_n12967_));
  NAND2_X1   g11965(.A1(new_n12967_), .A2(new_n12789_), .ZN(new_n12968_));
  NAND2_X1   g11966(.A1(new_n12966_), .A2(new_n12968_), .ZN(new_n12969_));
  NAND2_X1   g11967(.A1(new_n12969_), .A2(new_n12965_), .ZN(new_n12970_));
  XOR2_X1    g11968(.A1(new_n12798_), .A2(new_n12789_), .Z(new_n12971_));
  XOR2_X1    g11969(.A1(new_n12830_), .A2(new_n12821_), .Z(new_n12972_));
  NOR2_X1    g11970(.A1(new_n12971_), .A2(new_n12972_), .ZN(new_n12973_));
  NAND3_X1   g11971(.A1(new_n12970_), .A2(new_n12812_), .A3(new_n12973_), .ZN(new_n12974_));
  NAND2_X1   g11972(.A1(new_n12809_), .A2(new_n12804_), .ZN(new_n12975_));
  OAI21_X1   g11973(.A1(new_n12964_), .A2(new_n12968_), .B(new_n12975_), .ZN(new_n12976_));
  NAND2_X1   g11974(.A1(new_n12976_), .A2(new_n12799_), .ZN(new_n12977_));
  NAND2_X1   g11975(.A1(new_n12977_), .A2(new_n12844_), .ZN(new_n12978_));
  NOR2_X1    g11976(.A1(new_n12974_), .A2(new_n12978_), .ZN(new_n12979_));
  AND4_X2    g11977(.A1(new_n12799_), .A2(new_n12812_), .A3(new_n12844_), .A4(new_n12831_), .Z(new_n12980_));
  AOI22_X1   g11978(.A1(new_n12976_), .A2(new_n12799_), .B1(new_n12969_), .B2(new_n12965_), .ZN(new_n12981_));
  NOR2_X1    g11979(.A1(new_n12981_), .A2(new_n12980_), .ZN(new_n12982_));
  OAI21_X1   g11980(.A1(new_n12979_), .A2(new_n12982_), .B(new_n12963_), .ZN(new_n12983_));
  AOI21_X1   g11981(.A1(new_n12961_), .A2(new_n12843_), .B(new_n12957_), .ZN(new_n12984_));
  NOR2_X1    g11982(.A1(new_n12961_), .A2(new_n12955_), .ZN(new_n12985_));
  NOR2_X1    g11983(.A1(new_n12953_), .A2(new_n12843_), .ZN(new_n12986_));
  OAI22_X1   g11984(.A1(new_n12972_), .A2(new_n12984_), .B1(new_n12985_), .B2(new_n12986_), .ZN(new_n12987_));
  NAND3_X1   g11985(.A1(new_n12973_), .A2(new_n12812_), .A3(new_n12844_), .ZN(new_n12988_));
  NOR2_X1    g11986(.A1(new_n12981_), .A2(new_n12988_), .ZN(new_n12989_));
  NAND2_X1   g11987(.A1(new_n12977_), .A2(new_n12970_), .ZN(new_n12990_));
  NOR2_X1    g11988(.A1(new_n12990_), .A2(new_n12980_), .ZN(new_n12991_));
  OAI21_X1   g11989(.A1(new_n12991_), .A2(new_n12989_), .B(new_n12987_), .ZN(new_n12992_));
  XNOR2_X1   g11990(.A1(new_n12813_), .A2(new_n12845_), .ZN(new_n12993_));
  XNOR2_X1   g11991(.A1(new_n12878_), .A2(new_n12908_), .ZN(new_n12994_));
  NOR2_X1    g11992(.A1(new_n12993_), .A2(new_n12994_), .ZN(new_n12995_));
  NAND3_X1   g11993(.A1(new_n12983_), .A2(new_n12992_), .A3(new_n12995_), .ZN(new_n12996_));
  INV_X1     g11994(.I(new_n12996_), .ZN(new_n12997_));
  AOI21_X1   g11995(.A1(new_n12983_), .A2(new_n12992_), .B(new_n12995_), .ZN(new_n12998_));
  OAI21_X1   g11996(.A1(new_n12997_), .A2(new_n12998_), .B(new_n12952_), .ZN(new_n12999_));
  XOR2_X1    g11997(.A1(new_n12916_), .A2(new_n12919_), .Z(new_n13000_));
  AOI21_X1   g11998(.A1(new_n12916_), .A2(new_n12906_), .B(new_n12920_), .ZN(new_n13001_));
  NOR2_X1    g11999(.A1(new_n13001_), .A2(new_n12940_), .ZN(new_n13002_));
  NOR2_X1    g12000(.A1(new_n13000_), .A2(new_n13002_), .ZN(new_n13003_));
  NAND3_X1   g12001(.A1(new_n12943_), .A2(new_n12877_), .A3(new_n12941_), .ZN(new_n13004_));
  NAND2_X1   g12002(.A1(new_n12947_), .A2(new_n12907_), .ZN(new_n13005_));
  NOR2_X1    g12003(.A1(new_n13004_), .A2(new_n13005_), .ZN(new_n13006_));
  NOR3_X1    g12004(.A1(new_n12931_), .A2(new_n12930_), .A3(new_n12933_), .ZN(new_n13007_));
  NOR2_X1    g12005(.A1(new_n12929_), .A2(new_n12937_), .ZN(new_n13008_));
  NOR2_X1    g12006(.A1(new_n13008_), .A2(new_n13007_), .ZN(new_n13009_));
  OAI21_X1   g12007(.A1(new_n13006_), .A2(new_n13009_), .B(new_n13003_), .ZN(new_n13010_));
  NOR2_X1    g12008(.A1(new_n12948_), .A2(new_n13007_), .ZN(new_n13011_));
  NOR2_X1    g12009(.A1(new_n13008_), .A2(new_n12942_), .ZN(new_n13012_));
  OAI21_X1   g12010(.A1(new_n13012_), .A2(new_n13011_), .B(new_n12924_), .ZN(new_n13013_));
  NAND2_X1   g12011(.A1(new_n13010_), .A2(new_n13013_), .ZN(new_n13014_));
  NOR2_X1    g12012(.A1(new_n12966_), .A2(new_n12968_), .ZN(new_n13015_));
  NOR2_X1    g12013(.A1(new_n12964_), .A2(new_n12811_), .ZN(new_n13016_));
  NOR2_X1    g12014(.A1(new_n13015_), .A2(new_n13016_), .ZN(new_n13017_));
  NOR3_X1    g12015(.A1(new_n13017_), .A2(new_n12971_), .A3(new_n12972_), .ZN(new_n13018_));
  NAND4_X1   g12016(.A1(new_n13018_), .A2(new_n12812_), .A3(new_n12844_), .A4(new_n12977_), .ZN(new_n13019_));
  NAND2_X1   g12017(.A1(new_n12990_), .A2(new_n12988_), .ZN(new_n13020_));
  AOI21_X1   g12018(.A1(new_n13019_), .A2(new_n13020_), .B(new_n12987_), .ZN(new_n13021_));
  INV_X1     g12019(.I(new_n12989_), .ZN(new_n13022_));
  NAND2_X1   g12020(.A1(new_n12981_), .A2(new_n12988_), .ZN(new_n13023_));
  AOI21_X1   g12021(.A1(new_n13022_), .A2(new_n13023_), .B(new_n12963_), .ZN(new_n13024_));
  NOR3_X1    g12022(.A1(new_n13021_), .A2(new_n13024_), .A3(new_n12995_), .ZN(new_n13025_));
  NAND2_X1   g12023(.A1(new_n12846_), .A2(new_n12909_), .ZN(new_n13026_));
  AOI21_X1   g12024(.A1(new_n12983_), .A2(new_n12992_), .B(new_n13026_), .ZN(new_n13027_));
  OAI21_X1   g12025(.A1(new_n13025_), .A2(new_n13027_), .B(new_n13014_), .ZN(new_n13028_));
  NAND2_X1   g12026(.A1(new_n12999_), .A2(new_n13028_), .ZN(new_n13029_));
  XOR2_X1    g12027(.A1(new_n12773_), .A2(new_n12775_), .Z(new_n13030_));
  INV_X1     g12028(.I(new_n12777_), .ZN(new_n13031_));
  AOI21_X1   g12029(.A1(new_n12766_), .A2(\A[588] ), .B(new_n12771_), .ZN(new_n13032_));
  NOR2_X1    g12030(.A1(new_n13032_), .A2(new_n12775_), .ZN(new_n13033_));
  INV_X1     g12031(.I(new_n13033_), .ZN(new_n13034_));
  OAI21_X1   g12032(.A1(new_n13030_), .A2(new_n13031_), .B(new_n13034_), .ZN(new_n13035_));
  NAND2_X1   g12033(.A1(new_n13030_), .A2(new_n12777_), .ZN(new_n13036_));
  XOR2_X1    g12034(.A1(new_n13032_), .A2(new_n12775_), .Z(new_n13037_));
  NAND2_X1   g12035(.A1(new_n13037_), .A2(new_n13031_), .ZN(new_n13038_));
  AOI22_X1   g12036(.A1(new_n13035_), .A2(new_n12768_), .B1(new_n13036_), .B2(new_n13038_), .ZN(new_n13039_));
  XOR2_X1    g12037(.A1(new_n12740_), .A2(new_n12744_), .Z(new_n13040_));
  INV_X1     g12038(.I(new_n12734_), .ZN(new_n13041_));
  NAND2_X1   g12039(.A1(new_n13041_), .A2(new_n12725_), .ZN(new_n13042_));
  AOI21_X1   g12040(.A1(new_n12733_), .A2(\A[594] ), .B(new_n12738_), .ZN(new_n13043_));
  NOR2_X1    g12041(.A1(new_n13043_), .A2(new_n12744_), .ZN(new_n13044_));
  INV_X1     g12042(.I(new_n13044_), .ZN(new_n13045_));
  OAI21_X1   g12043(.A1(new_n13040_), .A2(new_n13042_), .B(new_n13045_), .ZN(new_n13046_));
  XOR2_X1    g12044(.A1(new_n13043_), .A2(new_n12744_), .Z(new_n13047_));
  NOR2_X1    g12045(.A1(new_n13047_), .A2(new_n13042_), .ZN(new_n13048_));
  NOR2_X1    g12046(.A1(new_n13040_), .A2(new_n12747_), .ZN(new_n13049_));
  NOR2_X1    g12047(.A1(new_n13049_), .A2(new_n13048_), .ZN(new_n13050_));
  NAND2_X1   g12048(.A1(new_n12735_), .A2(new_n12768_), .ZN(new_n13051_));
  NAND2_X1   g12049(.A1(new_n13046_), .A2(new_n12735_), .ZN(new_n13052_));
  NAND2_X1   g12050(.A1(new_n13052_), .A2(new_n12778_), .ZN(new_n13053_));
  NOR4_X1    g12051(.A1(new_n13053_), .A2(new_n13046_), .A3(new_n13050_), .A4(new_n13051_), .ZN(new_n13054_));
  NAND4_X1   g12052(.A1(new_n12748_), .A2(new_n12735_), .A3(new_n12768_), .A4(new_n12778_), .ZN(new_n13055_));
  INV_X1     g12053(.I(new_n13055_), .ZN(new_n13056_));
  NAND2_X1   g12054(.A1(new_n13040_), .A2(new_n12747_), .ZN(new_n13057_));
  NAND2_X1   g12055(.A1(new_n13047_), .A2(new_n13042_), .ZN(new_n13058_));
  AOI22_X1   g12056(.A1(new_n13046_), .A2(new_n12735_), .B1(new_n13057_), .B2(new_n13058_), .ZN(new_n13059_));
  NOR2_X1    g12057(.A1(new_n13059_), .A2(new_n13056_), .ZN(new_n13060_));
  OAI21_X1   g12058(.A1(new_n13054_), .A2(new_n13060_), .B(new_n13039_), .ZN(new_n13061_));
  INV_X1     g12059(.I(new_n13039_), .ZN(new_n13062_));
  NAND2_X1   g12060(.A1(new_n13057_), .A2(new_n13058_), .ZN(new_n13063_));
  NAND2_X1   g12061(.A1(new_n13052_), .A2(new_n13063_), .ZN(new_n13064_));
  NOR2_X1    g12062(.A1(new_n13064_), .A2(new_n13056_), .ZN(new_n13065_));
  NOR2_X1    g12063(.A1(new_n13059_), .A2(new_n13055_), .ZN(new_n13066_));
  OAI21_X1   g12064(.A1(new_n13065_), .A2(new_n13066_), .B(new_n13062_), .ZN(new_n13067_));
  NAND2_X1   g12065(.A1(new_n13061_), .A2(new_n13067_), .ZN(new_n13068_));
  NAND2_X1   g12066(.A1(new_n12717_), .A2(new_n12780_), .ZN(new_n13069_));
  XOR2_X1    g12067(.A1(new_n12701_), .A2(new_n12692_), .Z(new_n13070_));
  AOI21_X1   g12068(.A1(new_n12700_), .A2(\A[600] ), .B(new_n12705_), .ZN(new_n13071_));
  XOR2_X1    g12069(.A1(new_n13071_), .A2(new_n12711_), .Z(new_n13072_));
  NOR2_X1    g12070(.A1(new_n13071_), .A2(new_n12711_), .ZN(new_n13073_));
  AOI21_X1   g12071(.A1(new_n13072_), .A2(new_n12714_), .B(new_n13073_), .ZN(new_n13074_));
  INV_X1     g12072(.I(new_n12701_), .ZN(new_n13075_));
  NAND2_X1   g12073(.A1(new_n13075_), .A2(new_n12692_), .ZN(new_n13076_));
  NOR2_X1    g12074(.A1(new_n13072_), .A2(new_n13076_), .ZN(new_n13077_));
  XOR2_X1    g12075(.A1(new_n12707_), .A2(new_n12711_), .Z(new_n13078_));
  NOR2_X1    g12076(.A1(new_n13078_), .A2(new_n12714_), .ZN(new_n13079_));
  OAI22_X1   g12077(.A1(new_n13070_), .A2(new_n13074_), .B1(new_n13077_), .B2(new_n13079_), .ZN(new_n13080_));
  INV_X1     g12078(.I(new_n13080_), .ZN(new_n13081_));
  INV_X1     g12079(.I(new_n12683_), .ZN(new_n13082_));
  INV_X1     g12080(.I(new_n12715_), .ZN(new_n13083_));
  XOR2_X1    g12081(.A1(new_n12675_), .A2(new_n12679_), .Z(new_n13084_));
  NAND2_X1   g12082(.A1(new_n13084_), .A2(new_n12682_), .ZN(new_n13085_));
  AOI21_X1   g12083(.A1(new_n12668_), .A2(\A[606] ), .B(new_n12673_), .ZN(new_n13086_));
  XOR2_X1    g12084(.A1(new_n13086_), .A2(new_n12679_), .Z(new_n13087_));
  INV_X1     g12085(.I(new_n12669_), .ZN(new_n13088_));
  NAND2_X1   g12086(.A1(new_n13088_), .A2(new_n12660_), .ZN(new_n13089_));
  NAND2_X1   g12087(.A1(new_n13087_), .A2(new_n13089_), .ZN(new_n13090_));
  NAND2_X1   g12088(.A1(new_n13085_), .A2(new_n13090_), .ZN(new_n13091_));
  XOR2_X1    g12089(.A1(new_n12669_), .A2(new_n12660_), .Z(new_n13092_));
  NOR2_X1    g12090(.A1(new_n13092_), .A2(new_n13070_), .ZN(new_n13093_));
  NAND2_X1   g12091(.A1(new_n13091_), .A2(new_n13093_), .ZN(new_n13094_));
  NOR2_X1    g12092(.A1(new_n13086_), .A2(new_n12679_), .ZN(new_n13095_));
  AOI21_X1   g12093(.A1(new_n13087_), .A2(new_n12682_), .B(new_n13095_), .ZN(new_n13096_));
  NOR2_X1    g12094(.A1(new_n13096_), .A2(new_n13092_), .ZN(new_n13097_));
  NOR4_X1    g12095(.A1(new_n13094_), .A2(new_n13082_), .A3(new_n13083_), .A4(new_n13097_), .ZN(new_n13098_));
  NOR4_X1    g12096(.A1(new_n13082_), .A2(new_n13083_), .A3(new_n13092_), .A4(new_n13070_), .ZN(new_n13099_));
  NOR2_X1    g12097(.A1(new_n13087_), .A2(new_n13089_), .ZN(new_n13100_));
  NOR2_X1    g12098(.A1(new_n13084_), .A2(new_n12682_), .ZN(new_n13101_));
  NOR2_X1    g12099(.A1(new_n13101_), .A2(new_n13100_), .ZN(new_n13102_));
  NOR2_X1    g12100(.A1(new_n13097_), .A2(new_n13102_), .ZN(new_n13103_));
  NOR2_X1    g12101(.A1(new_n13103_), .A2(new_n13099_), .ZN(new_n13104_));
  OAI21_X1   g12102(.A1(new_n13098_), .A2(new_n13104_), .B(new_n13081_), .ZN(new_n13105_));
  NAND3_X1   g12103(.A1(new_n13093_), .A2(new_n12683_), .A3(new_n12715_), .ZN(new_n13106_));
  NOR2_X1    g12104(.A1(new_n13103_), .A2(new_n13106_), .ZN(new_n13107_));
  OAI22_X1   g12105(.A1(new_n13092_), .A2(new_n13096_), .B1(new_n13100_), .B2(new_n13101_), .ZN(new_n13108_));
  NOR2_X1    g12106(.A1(new_n13099_), .A2(new_n13108_), .ZN(new_n13109_));
  OAI21_X1   g12107(.A1(new_n13107_), .A2(new_n13109_), .B(new_n13080_), .ZN(new_n13110_));
  AOI21_X1   g12108(.A1(new_n13105_), .A2(new_n13110_), .B(new_n13069_), .ZN(new_n13111_));
  XNOR2_X1   g12109(.A1(new_n12684_), .A2(new_n12716_), .ZN(new_n13112_));
  XNOR2_X1   g12110(.A1(new_n12749_), .A2(new_n12779_), .ZN(new_n13113_));
  NOR2_X1    g12111(.A1(new_n13112_), .A2(new_n13113_), .ZN(new_n13114_));
  NOR2_X1    g12112(.A1(new_n13097_), .A2(new_n13083_), .ZN(new_n13115_));
  NAND4_X1   g12113(.A1(new_n13115_), .A2(new_n13096_), .A3(new_n13091_), .A4(new_n13093_), .ZN(new_n13116_));
  NAND2_X1   g12114(.A1(new_n13108_), .A2(new_n13106_), .ZN(new_n13117_));
  AOI21_X1   g12115(.A1(new_n13116_), .A2(new_n13117_), .B(new_n13080_), .ZN(new_n13118_));
  NAND2_X1   g12116(.A1(new_n13099_), .A2(new_n13108_), .ZN(new_n13119_));
  NAND2_X1   g12117(.A1(new_n13103_), .A2(new_n13106_), .ZN(new_n13120_));
  AOI21_X1   g12118(.A1(new_n13120_), .A2(new_n13119_), .B(new_n13081_), .ZN(new_n13121_));
  NOR3_X1    g12119(.A1(new_n13118_), .A2(new_n13121_), .A3(new_n13114_), .ZN(new_n13122_));
  OAI21_X1   g12120(.A1(new_n13111_), .A2(new_n13122_), .B(new_n13068_), .ZN(new_n13123_));
  NOR2_X1    g12121(.A1(new_n13050_), .A2(new_n13051_), .ZN(new_n13124_));
  NAND4_X1   g12122(.A1(new_n13124_), .A2(new_n12748_), .A3(new_n12778_), .A4(new_n13052_), .ZN(new_n13125_));
  INV_X1     g12123(.I(new_n13060_), .ZN(new_n13126_));
  AOI21_X1   g12124(.A1(new_n13126_), .A2(new_n13125_), .B(new_n13062_), .ZN(new_n13127_));
  NAND2_X1   g12125(.A1(new_n13059_), .A2(new_n13055_), .ZN(new_n13128_));
  NAND2_X1   g12126(.A1(new_n13064_), .A2(new_n13056_), .ZN(new_n13129_));
  AOI21_X1   g12127(.A1(new_n13129_), .A2(new_n13128_), .B(new_n13039_), .ZN(new_n13130_));
  NOR2_X1    g12128(.A1(new_n13127_), .A2(new_n13130_), .ZN(new_n13131_));
  AOI21_X1   g12129(.A1(new_n13105_), .A2(new_n13110_), .B(new_n13114_), .ZN(new_n13132_));
  NOR3_X1    g12130(.A1(new_n13118_), .A2(new_n13121_), .A3(new_n13069_), .ZN(new_n13133_));
  OAI21_X1   g12131(.A1(new_n13132_), .A2(new_n13133_), .B(new_n13131_), .ZN(new_n13134_));
  XOR2_X1    g12132(.A1(new_n13112_), .A2(new_n12780_), .Z(new_n13135_));
  XOR2_X1    g12133(.A1(new_n12993_), .A2(new_n12909_), .Z(new_n13136_));
  NOR2_X1    g12134(.A1(new_n13135_), .A2(new_n13136_), .ZN(new_n13137_));
  NAND3_X1   g12135(.A1(new_n13134_), .A2(new_n13123_), .A3(new_n13137_), .ZN(new_n13138_));
  NAND2_X1   g12136(.A1(new_n12781_), .A2(new_n12910_), .ZN(new_n13139_));
  NAND2_X1   g12137(.A1(new_n13134_), .A2(new_n13123_), .ZN(new_n13140_));
  NAND2_X1   g12138(.A1(new_n13140_), .A2(new_n13139_), .ZN(new_n13141_));
  AOI21_X1   g12139(.A1(new_n13141_), .A2(new_n13138_), .B(new_n13029_), .ZN(new_n13142_));
  INV_X1     g12140(.I(new_n12998_), .ZN(new_n13143_));
  AOI21_X1   g12141(.A1(new_n13143_), .A2(new_n12996_), .B(new_n13014_), .ZN(new_n13144_));
  NAND3_X1   g12142(.A1(new_n12983_), .A2(new_n12992_), .A3(new_n13026_), .ZN(new_n13145_));
  OAI21_X1   g12143(.A1(new_n13021_), .A2(new_n13024_), .B(new_n12995_), .ZN(new_n13146_));
  AOI21_X1   g12144(.A1(new_n13145_), .A2(new_n13146_), .B(new_n12952_), .ZN(new_n13147_));
  NOR2_X1    g12145(.A1(new_n13144_), .A2(new_n13147_), .ZN(new_n13148_));
  NAND3_X1   g12146(.A1(new_n13134_), .A2(new_n13123_), .A3(new_n13139_), .ZN(new_n13149_));
  OAI21_X1   g12147(.A1(new_n13118_), .A2(new_n13121_), .B(new_n13114_), .ZN(new_n13150_));
  NAND3_X1   g12148(.A1(new_n13105_), .A2(new_n13110_), .A3(new_n13069_), .ZN(new_n13151_));
  AOI21_X1   g12149(.A1(new_n13150_), .A2(new_n13151_), .B(new_n13131_), .ZN(new_n13152_));
  OAI21_X1   g12150(.A1(new_n13118_), .A2(new_n13121_), .B(new_n13069_), .ZN(new_n13153_));
  NAND3_X1   g12151(.A1(new_n13105_), .A2(new_n13110_), .A3(new_n13114_), .ZN(new_n13154_));
  AOI21_X1   g12152(.A1(new_n13153_), .A2(new_n13154_), .B(new_n13068_), .ZN(new_n13155_));
  OAI21_X1   g12153(.A1(new_n13152_), .A2(new_n13155_), .B(new_n13137_), .ZN(new_n13156_));
  AOI21_X1   g12154(.A1(new_n13149_), .A2(new_n13156_), .B(new_n13148_), .ZN(new_n13157_));
  NOR2_X1    g12155(.A1(new_n13142_), .A2(new_n13157_), .ZN(new_n13158_));
  INV_X1     g12156(.I(new_n13158_), .ZN(new_n13159_));
  XOR2_X1    g12157(.A1(new_n12634_), .A2(new_n12625_), .Z(new_n13160_));
  AOI21_X1   g12158(.A1(new_n12633_), .A2(\A[612] ), .B(new_n12638_), .ZN(new_n13161_));
  XOR2_X1    g12159(.A1(new_n13161_), .A2(new_n12644_), .Z(new_n13162_));
  NOR2_X1    g12160(.A1(new_n13161_), .A2(new_n12644_), .ZN(new_n13163_));
  AOI21_X1   g12161(.A1(new_n13162_), .A2(new_n12647_), .B(new_n13163_), .ZN(new_n13164_));
  XOR2_X1    g12162(.A1(new_n12640_), .A2(new_n12644_), .Z(new_n13165_));
  NAND2_X1   g12163(.A1(new_n13165_), .A2(new_n12647_), .ZN(new_n13166_));
  INV_X1     g12164(.I(new_n12634_), .ZN(new_n13167_));
  NAND2_X1   g12165(.A1(new_n13167_), .A2(new_n12625_), .ZN(new_n13168_));
  NAND2_X1   g12166(.A1(new_n13162_), .A2(new_n13168_), .ZN(new_n13169_));
  NAND2_X1   g12167(.A1(new_n13166_), .A2(new_n13169_), .ZN(new_n13170_));
  OAI21_X1   g12168(.A1(new_n13160_), .A2(new_n13164_), .B(new_n13170_), .ZN(new_n13171_));
  AOI21_X1   g12169(.A1(new_n12601_), .A2(\A[618] ), .B(new_n12606_), .ZN(new_n13172_));
  XOR2_X1    g12170(.A1(new_n13172_), .A2(new_n12612_), .Z(new_n13173_));
  INV_X1     g12171(.I(new_n12602_), .ZN(new_n13174_));
  NAND2_X1   g12172(.A1(new_n13174_), .A2(new_n12593_), .ZN(new_n13175_));
  NOR2_X1    g12173(.A1(new_n13173_), .A2(new_n13175_), .ZN(new_n13176_));
  XOR2_X1    g12174(.A1(new_n12608_), .A2(new_n12612_), .Z(new_n13177_));
  NOR2_X1    g12175(.A1(new_n13177_), .A2(new_n12615_), .ZN(new_n13178_));
  NOR2_X1    g12176(.A1(new_n13178_), .A2(new_n13176_), .ZN(new_n13179_));
  INV_X1     g12177(.I(new_n12616_), .ZN(new_n13180_));
  NAND2_X1   g12178(.A1(new_n12603_), .A2(new_n12635_), .ZN(new_n13181_));
  NOR3_X1    g12179(.A1(new_n13179_), .A2(new_n13180_), .A3(new_n13181_), .ZN(new_n13182_));
  INV_X1     g12180(.I(new_n12648_), .ZN(new_n13183_));
  XOR2_X1    g12181(.A1(new_n12602_), .A2(new_n12593_), .Z(new_n13184_));
  NOR2_X1    g12182(.A1(new_n13172_), .A2(new_n12612_), .ZN(new_n13185_));
  AOI21_X1   g12183(.A1(new_n13173_), .A2(new_n12615_), .B(new_n13185_), .ZN(new_n13186_));
  NOR2_X1    g12184(.A1(new_n13186_), .A2(new_n13184_), .ZN(new_n13187_));
  NOR2_X1    g12185(.A1(new_n13187_), .A2(new_n13183_), .ZN(new_n13188_));
  NAND2_X1   g12186(.A1(new_n13182_), .A2(new_n13188_), .ZN(new_n13189_));
  NOR2_X1    g12187(.A1(new_n13184_), .A2(new_n13160_), .ZN(new_n13190_));
  NAND3_X1   g12188(.A1(new_n13190_), .A2(new_n12616_), .A3(new_n12648_), .ZN(new_n13191_));
  OAI22_X1   g12189(.A1(new_n13184_), .A2(new_n13186_), .B1(new_n13176_), .B2(new_n13178_), .ZN(new_n13192_));
  NAND2_X1   g12190(.A1(new_n13192_), .A2(new_n13191_), .ZN(new_n13193_));
  AOI21_X1   g12191(.A1(new_n13189_), .A2(new_n13193_), .B(new_n13171_), .ZN(new_n13194_));
  XOR2_X1    g12192(.A1(new_n13192_), .A2(new_n13191_), .Z(new_n13195_));
  AOI21_X1   g12193(.A1(new_n13195_), .A2(new_n13171_), .B(new_n13194_), .ZN(new_n13196_));
  XOR2_X1    g12194(.A1(new_n12569_), .A2(new_n12560_), .Z(new_n13197_));
  AOI21_X1   g12195(.A1(new_n12568_), .A2(\A[624] ), .B(new_n12573_), .ZN(new_n13198_));
  XOR2_X1    g12196(.A1(new_n13198_), .A2(new_n12579_), .Z(new_n13199_));
  NOR2_X1    g12197(.A1(new_n13198_), .A2(new_n12579_), .ZN(new_n13200_));
  AOI21_X1   g12198(.A1(new_n13199_), .A2(new_n12582_), .B(new_n13200_), .ZN(new_n13201_));
  INV_X1     g12199(.I(new_n12569_), .ZN(new_n13202_));
  NAND2_X1   g12200(.A1(new_n13202_), .A2(new_n12560_), .ZN(new_n13203_));
  NOR2_X1    g12201(.A1(new_n13199_), .A2(new_n13203_), .ZN(new_n13204_));
  XOR2_X1    g12202(.A1(new_n12575_), .A2(new_n12579_), .Z(new_n13205_));
  NOR2_X1    g12203(.A1(new_n13205_), .A2(new_n12582_), .ZN(new_n13206_));
  OAI22_X1   g12204(.A1(new_n13197_), .A2(new_n13201_), .B1(new_n13204_), .B2(new_n13206_), .ZN(new_n13207_));
  XOR2_X1    g12205(.A1(new_n12537_), .A2(new_n12528_), .Z(new_n13208_));
  AOI21_X1   g12206(.A1(new_n12536_), .A2(\A[630] ), .B(new_n12541_), .ZN(new_n13209_));
  XOR2_X1    g12207(.A1(new_n13209_), .A2(new_n12547_), .Z(new_n13210_));
  INV_X1     g12208(.I(new_n12537_), .ZN(new_n13211_));
  NAND2_X1   g12209(.A1(new_n13211_), .A2(new_n12528_), .ZN(new_n13212_));
  NOR2_X1    g12210(.A1(new_n13210_), .A2(new_n13212_), .ZN(new_n13213_));
  XOR2_X1    g12211(.A1(new_n12543_), .A2(new_n12547_), .Z(new_n13214_));
  NOR2_X1    g12212(.A1(new_n13214_), .A2(new_n12550_), .ZN(new_n13215_));
  NOR2_X1    g12213(.A1(new_n13215_), .A2(new_n13213_), .ZN(new_n13216_));
  NOR3_X1    g12214(.A1(new_n13216_), .A2(new_n13208_), .A3(new_n13197_), .ZN(new_n13217_));
  NOR2_X1    g12215(.A1(new_n13209_), .A2(new_n12547_), .ZN(new_n13218_));
  INV_X1     g12216(.I(new_n13218_), .ZN(new_n13219_));
  OAI21_X1   g12217(.A1(new_n13214_), .A2(new_n13212_), .B(new_n13219_), .ZN(new_n13220_));
  NAND2_X1   g12218(.A1(new_n13220_), .A2(new_n12538_), .ZN(new_n13221_));
  NAND4_X1   g12219(.A1(new_n13217_), .A2(new_n12551_), .A3(new_n12583_), .A4(new_n13221_), .ZN(new_n13222_));
  NOR2_X1    g12220(.A1(new_n13208_), .A2(new_n13197_), .ZN(new_n13223_));
  NAND3_X1   g12221(.A1(new_n13223_), .A2(new_n12551_), .A3(new_n12583_), .ZN(new_n13224_));
  NAND2_X1   g12222(.A1(new_n13214_), .A2(new_n12550_), .ZN(new_n13225_));
  NAND2_X1   g12223(.A1(new_n13210_), .A2(new_n13212_), .ZN(new_n13226_));
  NAND2_X1   g12224(.A1(new_n13225_), .A2(new_n13226_), .ZN(new_n13227_));
  NAND2_X1   g12225(.A1(new_n13221_), .A2(new_n13227_), .ZN(new_n13228_));
  NAND2_X1   g12226(.A1(new_n13228_), .A2(new_n13224_), .ZN(new_n13229_));
  AOI21_X1   g12227(.A1(new_n13222_), .A2(new_n13229_), .B(new_n13207_), .ZN(new_n13230_));
  INV_X1     g12228(.I(new_n13201_), .ZN(new_n13231_));
  NAND2_X1   g12229(.A1(new_n13205_), .A2(new_n12582_), .ZN(new_n13232_));
  NAND2_X1   g12230(.A1(new_n13199_), .A2(new_n13203_), .ZN(new_n13233_));
  AOI22_X1   g12231(.A1(new_n13231_), .A2(new_n12570_), .B1(new_n13232_), .B2(new_n13233_), .ZN(new_n13234_));
  AND4_X2    g12232(.A1(new_n12538_), .A2(new_n12551_), .A3(new_n12583_), .A4(new_n12570_), .Z(new_n13235_));
  NAND2_X1   g12233(.A1(new_n13228_), .A2(new_n13235_), .ZN(new_n13236_));
  AOI22_X1   g12234(.A1(new_n13220_), .A2(new_n12538_), .B1(new_n13225_), .B2(new_n13226_), .ZN(new_n13237_));
  NAND2_X1   g12235(.A1(new_n13237_), .A2(new_n13224_), .ZN(new_n13238_));
  AOI21_X1   g12236(.A1(new_n13236_), .A2(new_n13238_), .B(new_n13234_), .ZN(new_n13239_));
  NAND2_X1   g12237(.A1(new_n12585_), .A2(new_n12650_), .ZN(new_n13240_));
  NOR3_X1    g12238(.A1(new_n13230_), .A2(new_n13239_), .A3(new_n13240_), .ZN(new_n13241_));
  NAND3_X1   g12239(.A1(new_n13227_), .A2(new_n12551_), .A3(new_n13223_), .ZN(new_n13242_));
  NAND2_X1   g12240(.A1(new_n13221_), .A2(new_n12583_), .ZN(new_n13243_));
  NOR2_X1    g12241(.A1(new_n13242_), .A2(new_n13243_), .ZN(new_n13244_));
  NOR2_X1    g12242(.A1(new_n13237_), .A2(new_n13235_), .ZN(new_n13245_));
  OAI21_X1   g12243(.A1(new_n13244_), .A2(new_n13245_), .B(new_n13234_), .ZN(new_n13246_));
  NOR2_X1    g12244(.A1(new_n13237_), .A2(new_n13224_), .ZN(new_n13247_));
  NOR2_X1    g12245(.A1(new_n13228_), .A2(new_n13235_), .ZN(new_n13248_));
  OAI21_X1   g12246(.A1(new_n13248_), .A2(new_n13247_), .B(new_n13207_), .ZN(new_n13249_));
  XNOR2_X1   g12247(.A1(new_n12552_), .A2(new_n12584_), .ZN(new_n13250_));
  XNOR2_X1   g12248(.A1(new_n12617_), .A2(new_n12649_), .ZN(new_n13251_));
  NOR2_X1    g12249(.A1(new_n13250_), .A2(new_n13251_), .ZN(new_n13252_));
  AOI21_X1   g12250(.A1(new_n13246_), .A2(new_n13249_), .B(new_n13252_), .ZN(new_n13253_));
  OAI21_X1   g12251(.A1(new_n13241_), .A2(new_n13253_), .B(new_n13196_), .ZN(new_n13254_));
  INV_X1     g12252(.I(new_n13164_), .ZN(new_n13255_));
  AOI22_X1   g12253(.A1(new_n13255_), .A2(new_n12635_), .B1(new_n13166_), .B2(new_n13169_), .ZN(new_n13256_));
  NAND2_X1   g12254(.A1(new_n13177_), .A2(new_n12615_), .ZN(new_n13257_));
  NAND2_X1   g12255(.A1(new_n13173_), .A2(new_n13175_), .ZN(new_n13258_));
  NAND2_X1   g12256(.A1(new_n13257_), .A2(new_n13258_), .ZN(new_n13259_));
  NAND2_X1   g12257(.A1(new_n13259_), .A2(new_n13190_), .ZN(new_n13260_));
  NOR4_X1    g12258(.A1(new_n13260_), .A2(new_n13180_), .A3(new_n13183_), .A4(new_n13187_), .ZN(new_n13261_));
  INV_X1     g12259(.I(new_n13193_), .ZN(new_n13262_));
  OAI21_X1   g12260(.A1(new_n13262_), .A2(new_n13261_), .B(new_n13256_), .ZN(new_n13263_));
  NOR3_X1    g12261(.A1(new_n13181_), .A2(new_n13180_), .A3(new_n13183_), .ZN(new_n13264_));
  NOR2_X1    g12262(.A1(new_n13264_), .A2(new_n13192_), .ZN(new_n13265_));
  INV_X1     g12263(.I(new_n13192_), .ZN(new_n13266_));
  NOR2_X1    g12264(.A1(new_n13266_), .A2(new_n13191_), .ZN(new_n13267_));
  OAI21_X1   g12265(.A1(new_n13267_), .A2(new_n13265_), .B(new_n13171_), .ZN(new_n13268_));
  NAND2_X1   g12266(.A1(new_n13263_), .A2(new_n13268_), .ZN(new_n13269_));
  NOR3_X1    g12267(.A1(new_n13230_), .A2(new_n13239_), .A3(new_n13252_), .ZN(new_n13270_));
  AOI21_X1   g12268(.A1(new_n13246_), .A2(new_n13249_), .B(new_n13240_), .ZN(new_n13271_));
  OAI21_X1   g12269(.A1(new_n13270_), .A2(new_n13271_), .B(new_n13269_), .ZN(new_n13272_));
  NAND2_X1   g12270(.A1(new_n13254_), .A2(new_n13272_), .ZN(new_n13273_));
  XOR2_X1    g12271(.A1(new_n12512_), .A2(new_n12514_), .Z(new_n13274_));
  INV_X1     g12272(.I(new_n12516_), .ZN(new_n13275_));
  AOI21_X1   g12273(.A1(new_n12505_), .A2(\A[636] ), .B(new_n12510_), .ZN(new_n13276_));
  NOR2_X1    g12274(.A1(new_n13276_), .A2(new_n12514_), .ZN(new_n13277_));
  INV_X1     g12275(.I(new_n13277_), .ZN(new_n13278_));
  OAI21_X1   g12276(.A1(new_n13274_), .A2(new_n13275_), .B(new_n13278_), .ZN(new_n13279_));
  NAND2_X1   g12277(.A1(new_n13274_), .A2(new_n12516_), .ZN(new_n13280_));
  XOR2_X1    g12278(.A1(new_n13276_), .A2(new_n12514_), .Z(new_n13281_));
  NAND2_X1   g12279(.A1(new_n13281_), .A2(new_n13275_), .ZN(new_n13282_));
  AOI22_X1   g12280(.A1(new_n13279_), .A2(new_n12507_), .B1(new_n13280_), .B2(new_n13282_), .ZN(new_n13283_));
  INV_X1     g12281(.I(new_n12487_), .ZN(new_n13284_));
  INV_X1     g12282(.I(new_n12517_), .ZN(new_n13285_));
  XOR2_X1    g12283(.A1(new_n12479_), .A2(new_n12483_), .Z(new_n13286_));
  NAND2_X1   g12284(.A1(new_n13286_), .A2(new_n12486_), .ZN(new_n13287_));
  AOI21_X1   g12285(.A1(new_n12472_), .A2(\A[642] ), .B(new_n12477_), .ZN(new_n13288_));
  XOR2_X1    g12286(.A1(new_n13288_), .A2(new_n12483_), .Z(new_n13289_));
  INV_X1     g12287(.I(new_n12473_), .ZN(new_n13290_));
  NAND2_X1   g12288(.A1(new_n13290_), .A2(new_n12464_), .ZN(new_n13291_));
  NAND2_X1   g12289(.A1(new_n13289_), .A2(new_n13291_), .ZN(new_n13292_));
  NAND2_X1   g12290(.A1(new_n13287_), .A2(new_n13292_), .ZN(new_n13293_));
  XOR2_X1    g12291(.A1(new_n12473_), .A2(new_n12464_), .Z(new_n13294_));
  XNOR2_X1   g12292(.A1(new_n12497_), .A2(new_n12506_), .ZN(new_n13295_));
  NOR2_X1    g12293(.A1(new_n13295_), .A2(new_n13294_), .ZN(new_n13296_));
  NAND2_X1   g12294(.A1(new_n13293_), .A2(new_n13296_), .ZN(new_n13297_));
  NOR2_X1    g12295(.A1(new_n13288_), .A2(new_n12483_), .ZN(new_n13298_));
  AOI21_X1   g12296(.A1(new_n13289_), .A2(new_n12486_), .B(new_n13298_), .ZN(new_n13299_));
  NOR2_X1    g12297(.A1(new_n13299_), .A2(new_n13294_), .ZN(new_n13300_));
  NOR4_X1    g12298(.A1(new_n13297_), .A2(new_n13284_), .A3(new_n13285_), .A4(new_n13300_), .ZN(new_n13301_));
  NAND2_X1   g12299(.A1(new_n12474_), .A2(new_n12507_), .ZN(new_n13302_));
  NOR3_X1    g12300(.A1(new_n13302_), .A2(new_n13284_), .A3(new_n13285_), .ZN(new_n13303_));
  NOR2_X1    g12301(.A1(new_n13289_), .A2(new_n13291_), .ZN(new_n13304_));
  NOR2_X1    g12302(.A1(new_n13286_), .A2(new_n12486_), .ZN(new_n13305_));
  NOR2_X1    g12303(.A1(new_n13305_), .A2(new_n13304_), .ZN(new_n13306_));
  NOR2_X1    g12304(.A1(new_n13300_), .A2(new_n13306_), .ZN(new_n13307_));
  NOR2_X1    g12305(.A1(new_n13307_), .A2(new_n13303_), .ZN(new_n13308_));
  OAI21_X1   g12306(.A1(new_n13301_), .A2(new_n13308_), .B(new_n13283_), .ZN(new_n13309_));
  INV_X1     g12307(.I(new_n13283_), .ZN(new_n13310_));
  INV_X1     g12308(.I(new_n13298_), .ZN(new_n13311_));
  OAI21_X1   g12309(.A1(new_n13286_), .A2(new_n13291_), .B(new_n13311_), .ZN(new_n13312_));
  NAND2_X1   g12310(.A1(new_n13312_), .A2(new_n12474_), .ZN(new_n13313_));
  NAND2_X1   g12311(.A1(new_n13313_), .A2(new_n13293_), .ZN(new_n13314_));
  NOR2_X1    g12312(.A1(new_n13314_), .A2(new_n13303_), .ZN(new_n13315_));
  NAND3_X1   g12313(.A1(new_n13296_), .A2(new_n12487_), .A3(new_n12517_), .ZN(new_n13316_));
  NOR2_X1    g12314(.A1(new_n13307_), .A2(new_n13316_), .ZN(new_n13317_));
  OAI21_X1   g12315(.A1(new_n13317_), .A2(new_n13315_), .B(new_n13310_), .ZN(new_n13318_));
  NAND2_X1   g12316(.A1(new_n13309_), .A2(new_n13318_), .ZN(new_n13319_));
  NAND2_X1   g12317(.A1(new_n12456_), .A2(new_n12519_), .ZN(new_n13320_));
  AOI21_X1   g12318(.A1(new_n12441_), .A2(\A[648] ), .B(new_n12444_), .ZN(new_n13321_));
  XOR2_X1    g12319(.A1(new_n12451_), .A2(new_n13321_), .Z(new_n13322_));
  INV_X1     g12320(.I(new_n12442_), .ZN(new_n13323_));
  NAND2_X1   g12321(.A1(new_n13323_), .A2(new_n12434_), .ZN(new_n13324_));
  NAND2_X1   g12322(.A1(new_n12431_), .A2(\A[644] ), .ZN(new_n13325_));
  NAND2_X1   g12323(.A1(new_n13325_), .A2(new_n12429_), .ZN(new_n13326_));
  AOI21_X1   g12324(.A1(new_n13326_), .A2(\A[645] ), .B(new_n12449_), .ZN(new_n13327_));
  NOR2_X1    g12325(.A1(new_n13321_), .A2(new_n13327_), .ZN(new_n13328_));
  INV_X1     g12326(.I(new_n13328_), .ZN(new_n13329_));
  OAI21_X1   g12327(.A1(new_n13322_), .A2(new_n13324_), .B(new_n13329_), .ZN(new_n13330_));
  NAND2_X1   g12328(.A1(new_n13322_), .A2(new_n12453_), .ZN(new_n13331_));
  XOR2_X1    g12329(.A1(new_n13321_), .A2(new_n13327_), .Z(new_n13332_));
  NAND2_X1   g12330(.A1(new_n13332_), .A2(new_n13324_), .ZN(new_n13333_));
  AOI22_X1   g12331(.A1(new_n13330_), .A2(new_n12443_), .B1(new_n13331_), .B2(new_n13333_), .ZN(new_n13334_));
  NAND2_X1   g12332(.A1(new_n12400_), .A2(\A[650] ), .ZN(new_n13335_));
  NAND2_X1   g12333(.A1(new_n13335_), .A2(new_n12398_), .ZN(new_n13336_));
  AOI21_X1   g12334(.A1(new_n13336_), .A2(\A[651] ), .B(new_n12420_), .ZN(new_n13337_));
  XOR2_X1    g12335(.A1(new_n12418_), .A2(new_n13337_), .Z(new_n13338_));
  INV_X1     g12336(.I(new_n12412_), .ZN(new_n13339_));
  NAND2_X1   g12337(.A1(new_n13339_), .A2(new_n12403_), .ZN(new_n13340_));
  AOI21_X1   g12338(.A1(new_n12411_), .A2(\A[654] ), .B(new_n12416_), .ZN(new_n13341_));
  NOR2_X1    g12339(.A1(new_n13341_), .A2(new_n13337_), .ZN(new_n13342_));
  INV_X1     g12340(.I(new_n13342_), .ZN(new_n13343_));
  OAI21_X1   g12341(.A1(new_n13338_), .A2(new_n13340_), .B(new_n13343_), .ZN(new_n13344_));
  NAND2_X1   g12342(.A1(new_n12418_), .A2(new_n13337_), .ZN(new_n13345_));
  NAND2_X1   g12343(.A1(new_n12422_), .A2(new_n13341_), .ZN(new_n13346_));
  NAND2_X1   g12344(.A1(new_n13345_), .A2(new_n13346_), .ZN(new_n13347_));
  XOR2_X1    g12345(.A1(new_n13347_), .A2(new_n13340_), .Z(new_n13348_));
  NAND2_X1   g12346(.A1(new_n12413_), .A2(new_n12443_), .ZN(new_n13349_));
  XOR2_X1    g12347(.A1(new_n12412_), .A2(new_n12403_), .Z(new_n13350_));
  AOI21_X1   g12348(.A1(new_n13347_), .A2(new_n12424_), .B(new_n13342_), .ZN(new_n13351_));
  OAI21_X1   g12349(.A1(new_n13351_), .A2(new_n13350_), .B(new_n12454_), .ZN(new_n13352_));
  NOR4_X1    g12350(.A1(new_n13348_), .A2(new_n13352_), .A3(new_n13344_), .A4(new_n13349_), .ZN(new_n13353_));
  NAND4_X1   g12351(.A1(new_n12425_), .A2(new_n12454_), .A3(new_n12413_), .A4(new_n12443_), .ZN(new_n13354_));
  INV_X1     g12352(.I(new_n13354_), .ZN(new_n13355_));
  NOR2_X1    g12353(.A1(new_n13351_), .A2(new_n13350_), .ZN(new_n13356_));
  NOR2_X1    g12354(.A1(new_n13348_), .A2(new_n13356_), .ZN(new_n13357_));
  NOR2_X1    g12355(.A1(new_n13357_), .A2(new_n13355_), .ZN(new_n13358_));
  OAI21_X1   g12356(.A1(new_n13358_), .A2(new_n13353_), .B(new_n13334_), .ZN(new_n13359_));
  INV_X1     g12357(.I(new_n12443_), .ZN(new_n13360_));
  AOI21_X1   g12358(.A1(new_n13332_), .A2(new_n12453_), .B(new_n13328_), .ZN(new_n13361_));
  NOR2_X1    g12359(.A1(new_n13332_), .A2(new_n13324_), .ZN(new_n13362_));
  NOR2_X1    g12360(.A1(new_n13322_), .A2(new_n12453_), .ZN(new_n13363_));
  OAI22_X1   g12361(.A1(new_n13360_), .A2(new_n13361_), .B1(new_n13363_), .B2(new_n13362_), .ZN(new_n13364_));
  NOR2_X1    g12362(.A1(new_n13357_), .A2(new_n13354_), .ZN(new_n13365_));
  NOR3_X1    g12363(.A1(new_n13355_), .A2(new_n13348_), .A3(new_n13356_), .ZN(new_n13366_));
  OAI21_X1   g12364(.A1(new_n13365_), .A2(new_n13366_), .B(new_n13364_), .ZN(new_n13367_));
  AOI21_X1   g12365(.A1(new_n13367_), .A2(new_n13359_), .B(new_n13320_), .ZN(new_n13368_));
  XNOR2_X1   g12366(.A1(new_n12426_), .A2(new_n12455_), .ZN(new_n13369_));
  XNOR2_X1   g12367(.A1(new_n12488_), .A2(new_n12518_), .ZN(new_n13370_));
  NOR2_X1    g12368(.A1(new_n13369_), .A2(new_n13370_), .ZN(new_n13371_));
  INV_X1     g12369(.I(new_n13353_), .ZN(new_n13372_));
  NAND3_X1   g12370(.A1(new_n12424_), .A2(new_n13345_), .A3(new_n13346_), .ZN(new_n13373_));
  NAND2_X1   g12371(.A1(new_n13347_), .A2(new_n13340_), .ZN(new_n13374_));
  NAND2_X1   g12372(.A1(new_n13374_), .A2(new_n13373_), .ZN(new_n13375_));
  OAI21_X1   g12373(.A1(new_n13350_), .A2(new_n13351_), .B(new_n13375_), .ZN(new_n13376_));
  NAND2_X1   g12374(.A1(new_n13376_), .A2(new_n13354_), .ZN(new_n13377_));
  AOI21_X1   g12375(.A1(new_n13372_), .A2(new_n13377_), .B(new_n13364_), .ZN(new_n13378_));
  NAND2_X1   g12376(.A1(new_n13376_), .A2(new_n13355_), .ZN(new_n13379_));
  NAND2_X1   g12377(.A1(new_n13357_), .A2(new_n13354_), .ZN(new_n13380_));
  AOI21_X1   g12378(.A1(new_n13379_), .A2(new_n13380_), .B(new_n13334_), .ZN(new_n13381_));
  NOR3_X1    g12379(.A1(new_n13378_), .A2(new_n13381_), .A3(new_n13371_), .ZN(new_n13382_));
  OAI21_X1   g12380(.A1(new_n13382_), .A2(new_n13368_), .B(new_n13319_), .ZN(new_n13383_));
  NOR2_X1    g12381(.A1(new_n13306_), .A2(new_n13302_), .ZN(new_n13384_));
  NAND4_X1   g12382(.A1(new_n13384_), .A2(new_n12487_), .A3(new_n12517_), .A4(new_n13313_), .ZN(new_n13385_));
  NAND2_X1   g12383(.A1(new_n13314_), .A2(new_n13316_), .ZN(new_n13386_));
  AOI21_X1   g12384(.A1(new_n13385_), .A2(new_n13386_), .B(new_n13310_), .ZN(new_n13387_));
  XOR2_X1    g12385(.A1(new_n13314_), .A2(new_n13316_), .Z(new_n13388_));
  AOI21_X1   g12386(.A1(new_n13388_), .A2(new_n13310_), .B(new_n13387_), .ZN(new_n13389_));
  AOI21_X1   g12387(.A1(new_n13359_), .A2(new_n13367_), .B(new_n13371_), .ZN(new_n13390_));
  NOR3_X1    g12388(.A1(new_n13378_), .A2(new_n13381_), .A3(new_n13320_), .ZN(new_n13391_));
  OAI21_X1   g12389(.A1(new_n13390_), .A2(new_n13391_), .B(new_n13389_), .ZN(new_n13392_));
  NAND2_X1   g12390(.A1(new_n12651_), .A2(new_n12520_), .ZN(new_n13393_));
  NAND3_X1   g12391(.A1(new_n13392_), .A2(new_n13383_), .A3(new_n13393_), .ZN(new_n13394_));
  OAI21_X1   g12392(.A1(new_n13378_), .A2(new_n13381_), .B(new_n13371_), .ZN(new_n13395_));
  NAND3_X1   g12393(.A1(new_n13367_), .A2(new_n13359_), .A3(new_n13320_), .ZN(new_n13396_));
  AOI21_X1   g12394(.A1(new_n13395_), .A2(new_n13396_), .B(new_n13389_), .ZN(new_n13397_));
  INV_X1     g12395(.I(new_n13390_), .ZN(new_n13398_));
  NAND3_X1   g12396(.A1(new_n13371_), .A2(new_n13367_), .A3(new_n13359_), .ZN(new_n13399_));
  AOI21_X1   g12397(.A1(new_n13398_), .A2(new_n13399_), .B(new_n13319_), .ZN(new_n13400_));
  INV_X1     g12398(.I(new_n13393_), .ZN(new_n13401_));
  OAI21_X1   g12399(.A1(new_n13400_), .A2(new_n13397_), .B(new_n13401_), .ZN(new_n13402_));
  NAND2_X1   g12400(.A1(new_n13402_), .A2(new_n13394_), .ZN(new_n13403_));
  NAND2_X1   g12401(.A1(new_n13403_), .A2(new_n13273_), .ZN(new_n13404_));
  INV_X1     g12402(.I(new_n13273_), .ZN(new_n13405_));
  NOR3_X1    g12403(.A1(new_n13400_), .A2(new_n13397_), .A3(new_n13393_), .ZN(new_n13406_));
  AOI21_X1   g12404(.A1(new_n13383_), .A2(new_n13392_), .B(new_n13401_), .ZN(new_n13407_));
  OAI21_X1   g12405(.A1(new_n13407_), .A2(new_n13406_), .B(new_n13405_), .ZN(new_n13408_));
  NAND2_X1   g12406(.A1(new_n12652_), .A2(new_n12911_), .ZN(new_n13409_));
  INV_X1     g12407(.I(new_n13409_), .ZN(new_n13410_));
  NAND3_X1   g12408(.A1(new_n13404_), .A2(new_n13408_), .A3(new_n13410_), .ZN(new_n13411_));
  AOI21_X1   g12409(.A1(new_n13394_), .A2(new_n13402_), .B(new_n13405_), .ZN(new_n13412_));
  NAND3_X1   g12410(.A1(new_n13401_), .A2(new_n13392_), .A3(new_n13383_), .ZN(new_n13413_));
  NAND2_X1   g12411(.A1(new_n13392_), .A2(new_n13383_), .ZN(new_n13414_));
  NAND2_X1   g12412(.A1(new_n13414_), .A2(new_n13393_), .ZN(new_n13415_));
  AOI21_X1   g12413(.A1(new_n13415_), .A2(new_n13413_), .B(new_n13273_), .ZN(new_n13416_));
  OAI21_X1   g12414(.A1(new_n13412_), .A2(new_n13416_), .B(new_n13409_), .ZN(new_n13417_));
  AOI21_X1   g12415(.A1(new_n13417_), .A2(new_n13411_), .B(new_n13159_), .ZN(new_n13418_));
  NAND3_X1   g12416(.A1(new_n13404_), .A2(new_n13408_), .A3(new_n13409_), .ZN(new_n13419_));
  OAI21_X1   g12417(.A1(new_n13412_), .A2(new_n13416_), .B(new_n13410_), .ZN(new_n13420_));
  AOI21_X1   g12418(.A1(new_n13419_), .A2(new_n13420_), .B(new_n13158_), .ZN(new_n13421_));
  OAI21_X1   g12419(.A1(new_n13418_), .A2(new_n13421_), .B(new_n12914_), .ZN(new_n13422_));
  NAND2_X1   g12420(.A1(new_n11914_), .A2(\A[467] ), .ZN(new_n13423_));
  NAND2_X1   g12421(.A1(new_n13423_), .A2(new_n11912_), .ZN(new_n13424_));
  AOI21_X1   g12422(.A1(new_n13424_), .A2(\A[468] ), .B(new_n11929_), .ZN(new_n13425_));
  XOR2_X1    g12423(.A1(new_n13425_), .A2(new_n11933_), .Z(new_n13426_));
  XOR2_X1    g12424(.A1(new_n13426_), .A2(new_n11936_), .Z(new_n13427_));
  XOR2_X1    g12425(.A1(new_n11931_), .A2(new_n11933_), .Z(new_n13428_));
  INV_X1     g12426(.I(new_n11936_), .ZN(new_n13429_));
  NOR2_X1    g12427(.A1(new_n13425_), .A2(new_n11933_), .ZN(new_n13430_));
  INV_X1     g12428(.I(new_n13430_), .ZN(new_n13431_));
  OAI21_X1   g12429(.A1(new_n13429_), .A2(new_n13428_), .B(new_n13431_), .ZN(new_n13432_));
  NAND2_X1   g12430(.A1(new_n13432_), .A2(new_n11927_), .ZN(new_n13433_));
  NAND2_X1   g12431(.A1(new_n13427_), .A2(new_n13433_), .ZN(new_n13434_));
  AOI21_X1   g12432(.A1(new_n11896_), .A2(\A[474] ), .B(new_n11901_), .ZN(new_n13435_));
  XOR2_X1    g12433(.A1(new_n13435_), .A2(new_n11905_), .Z(new_n13436_));
  INV_X1     g12434(.I(new_n11907_), .ZN(new_n13437_));
  XOR2_X1    g12435(.A1(new_n13436_), .A2(new_n13437_), .Z(new_n13438_));
  INV_X1     g12436(.I(new_n11908_), .ZN(new_n13439_));
  NAND2_X1   g12437(.A1(new_n11927_), .A2(new_n11898_), .ZN(new_n13440_));
  NOR3_X1    g12438(.A1(new_n13438_), .A2(new_n13439_), .A3(new_n13440_), .ZN(new_n13441_));
  INV_X1     g12439(.I(new_n11937_), .ZN(new_n13442_));
  INV_X1     g12440(.I(new_n11898_), .ZN(new_n13443_));
  NOR2_X1    g12441(.A1(new_n13435_), .A2(new_n11905_), .ZN(new_n13444_));
  AOI21_X1   g12442(.A1(new_n13436_), .A2(new_n11907_), .B(new_n13444_), .ZN(new_n13445_));
  NOR2_X1    g12443(.A1(new_n13445_), .A2(new_n13443_), .ZN(new_n13446_));
  NOR2_X1    g12444(.A1(new_n13446_), .A2(new_n13442_), .ZN(new_n13447_));
  NAND2_X1   g12445(.A1(new_n13441_), .A2(new_n13447_), .ZN(new_n13448_));
  NOR3_X1    g12446(.A1(new_n13440_), .A2(new_n13442_), .A3(new_n13439_), .ZN(new_n13449_));
  INV_X1     g12447(.I(new_n13449_), .ZN(new_n13450_));
  XOR2_X1    g12448(.A1(new_n13436_), .A2(new_n11907_), .Z(new_n13451_));
  XOR2_X1    g12449(.A1(new_n11903_), .A2(new_n11905_), .Z(new_n13452_));
  INV_X1     g12450(.I(new_n13444_), .ZN(new_n13453_));
  OAI21_X1   g12451(.A1(new_n13452_), .A2(new_n13437_), .B(new_n13453_), .ZN(new_n13454_));
  NAND2_X1   g12452(.A1(new_n13454_), .A2(new_n11898_), .ZN(new_n13455_));
  NAND2_X1   g12453(.A1(new_n13451_), .A2(new_n13455_), .ZN(new_n13456_));
  NAND2_X1   g12454(.A1(new_n13450_), .A2(new_n13456_), .ZN(new_n13457_));
  AOI21_X1   g12455(.A1(new_n13448_), .A2(new_n13457_), .B(new_n13434_), .ZN(new_n13458_));
  XOR2_X1    g12456(.A1(new_n13428_), .A2(new_n11936_), .Z(new_n13459_));
  INV_X1     g12457(.I(new_n11927_), .ZN(new_n13460_));
  AOI21_X1   g12458(.A1(new_n13426_), .A2(new_n11936_), .B(new_n13430_), .ZN(new_n13461_));
  NOR2_X1    g12459(.A1(new_n13461_), .A2(new_n13460_), .ZN(new_n13462_));
  NOR2_X1    g12460(.A1(new_n13459_), .A2(new_n13462_), .ZN(new_n13463_));
  NOR2_X1    g12461(.A1(new_n13438_), .A2(new_n13446_), .ZN(new_n13464_));
  NAND2_X1   g12462(.A1(new_n13464_), .A2(new_n13450_), .ZN(new_n13465_));
  NAND2_X1   g12463(.A1(new_n13456_), .A2(new_n13449_), .ZN(new_n13466_));
  AOI21_X1   g12464(.A1(new_n13465_), .A2(new_n13466_), .B(new_n13463_), .ZN(new_n13467_));
  NOR2_X1    g12465(.A1(new_n13458_), .A2(new_n13467_), .ZN(new_n13468_));
  AOI21_X1   g12466(.A1(new_n11987_), .A2(\A[480] ), .B(new_n11992_), .ZN(new_n13469_));
  XNOR2_X1   g12467(.A1(new_n13469_), .A2(new_n11998_), .ZN(new_n13470_));
  INV_X1     g12468(.I(new_n11988_), .ZN(new_n13471_));
  NAND2_X1   g12469(.A1(new_n13471_), .A2(new_n11979_), .ZN(new_n13472_));
  NOR2_X1    g12470(.A1(new_n13469_), .A2(new_n11998_), .ZN(new_n13473_));
  INV_X1     g12471(.I(new_n13473_), .ZN(new_n13474_));
  OAI21_X1   g12472(.A1(new_n13470_), .A2(new_n13472_), .B(new_n13474_), .ZN(new_n13475_));
  NAND2_X1   g12473(.A1(new_n13470_), .A2(new_n12001_), .ZN(new_n13476_));
  XOR2_X1    g12474(.A1(new_n13469_), .A2(new_n11998_), .Z(new_n13477_));
  NAND2_X1   g12475(.A1(new_n13477_), .A2(new_n13472_), .ZN(new_n13478_));
  AOI22_X1   g12476(.A1(new_n13475_), .A2(new_n11989_), .B1(new_n13476_), .B2(new_n13478_), .ZN(new_n13479_));
  INV_X1     g12477(.I(new_n13479_), .ZN(new_n13480_));
  XOR2_X1    g12478(.A1(new_n11956_), .A2(new_n11947_), .Z(new_n13481_));
  XNOR2_X1   g12479(.A1(new_n11962_), .A2(new_n11966_), .ZN(new_n13482_));
  INV_X1     g12480(.I(new_n11956_), .ZN(new_n13483_));
  NAND2_X1   g12481(.A1(new_n13483_), .A2(new_n11947_), .ZN(new_n13484_));
  NOR2_X1    g12482(.A1(new_n13482_), .A2(new_n13484_), .ZN(new_n13485_));
  XOR2_X1    g12483(.A1(new_n11962_), .A2(new_n11966_), .Z(new_n13486_));
  NOR2_X1    g12484(.A1(new_n13486_), .A2(new_n11969_), .ZN(new_n13487_));
  NOR2_X1    g12485(.A1(new_n13485_), .A2(new_n13487_), .ZN(new_n13488_));
  XOR2_X1    g12486(.A1(new_n11988_), .A2(new_n11979_), .Z(new_n13489_));
  NOR3_X1    g12487(.A1(new_n13488_), .A2(new_n13481_), .A3(new_n13489_), .ZN(new_n13490_));
  NAND2_X1   g12488(.A1(new_n11967_), .A2(new_n11962_), .ZN(new_n13491_));
  OAI21_X1   g12489(.A1(new_n13486_), .A2(new_n13484_), .B(new_n13491_), .ZN(new_n13492_));
  NAND2_X1   g12490(.A1(new_n13492_), .A2(new_n11957_), .ZN(new_n13493_));
  NAND4_X1   g12491(.A1(new_n13490_), .A2(new_n11970_), .A3(new_n12002_), .A4(new_n13493_), .ZN(new_n13494_));
  NOR2_X1    g12492(.A1(new_n13481_), .A2(new_n13489_), .ZN(new_n13495_));
  NAND3_X1   g12493(.A1(new_n13495_), .A2(new_n11970_), .A3(new_n12002_), .ZN(new_n13496_));
  NAND2_X1   g12494(.A1(new_n13486_), .A2(new_n11969_), .ZN(new_n13497_));
  NAND2_X1   g12495(.A1(new_n13482_), .A2(new_n13484_), .ZN(new_n13498_));
  NAND2_X1   g12496(.A1(new_n13498_), .A2(new_n13497_), .ZN(new_n13499_));
  NAND2_X1   g12497(.A1(new_n13493_), .A2(new_n13499_), .ZN(new_n13500_));
  NAND2_X1   g12498(.A1(new_n13500_), .A2(new_n13496_), .ZN(new_n13501_));
  AOI21_X1   g12499(.A1(new_n13494_), .A2(new_n13501_), .B(new_n13480_), .ZN(new_n13502_));
  XNOR2_X1   g12500(.A1(new_n11938_), .A2(new_n11909_), .ZN(new_n13503_));
  XNOR2_X1   g12501(.A1(new_n11971_), .A2(new_n12003_), .ZN(new_n13504_));
  NOR2_X1    g12502(.A1(new_n13504_), .A2(new_n13503_), .ZN(new_n13505_));
  AOI22_X1   g12503(.A1(new_n13492_), .A2(new_n11957_), .B1(new_n13498_), .B2(new_n13497_), .ZN(new_n13506_));
  NOR2_X1    g12504(.A1(new_n13506_), .A2(new_n13496_), .ZN(new_n13507_));
  AND4_X2    g12505(.A1(new_n11957_), .A2(new_n11970_), .A3(new_n12002_), .A4(new_n11989_), .Z(new_n13508_));
  NOR2_X1    g12506(.A1(new_n13500_), .A2(new_n13508_), .ZN(new_n13509_));
  OAI21_X1   g12507(.A1(new_n13509_), .A2(new_n13507_), .B(new_n13480_), .ZN(new_n13510_));
  NAND2_X1   g12508(.A1(new_n13510_), .A2(new_n13505_), .ZN(new_n13511_));
  INV_X1     g12509(.I(new_n13507_), .ZN(new_n13512_));
  NAND2_X1   g12510(.A1(new_n13506_), .A2(new_n13496_), .ZN(new_n13513_));
  AOI21_X1   g12511(.A1(new_n13512_), .A2(new_n13513_), .B(new_n13479_), .ZN(new_n13514_));
  NOR2_X1    g12512(.A1(new_n13502_), .A2(new_n13514_), .ZN(new_n13515_));
  OAI22_X1   g12513(.A1(new_n13515_), .A2(new_n13505_), .B1(new_n13511_), .B2(new_n13502_), .ZN(new_n13516_));
  NAND2_X1   g12514(.A1(new_n13516_), .A2(new_n13468_), .ZN(new_n13517_));
  INV_X1     g12515(.I(new_n13440_), .ZN(new_n13518_));
  NAND3_X1   g12516(.A1(new_n13451_), .A2(new_n13518_), .A3(new_n11908_), .ZN(new_n13519_));
  NAND2_X1   g12517(.A1(new_n13455_), .A2(new_n11937_), .ZN(new_n13520_));
  NOR2_X1    g12518(.A1(new_n13519_), .A2(new_n13520_), .ZN(new_n13521_));
  NOR2_X1    g12519(.A1(new_n13464_), .A2(new_n13449_), .ZN(new_n13522_));
  OAI21_X1   g12520(.A1(new_n13521_), .A2(new_n13522_), .B(new_n13463_), .ZN(new_n13523_));
  NOR2_X1    g12521(.A1(new_n13456_), .A2(new_n13449_), .ZN(new_n13524_));
  NOR2_X1    g12522(.A1(new_n13464_), .A2(new_n13450_), .ZN(new_n13525_));
  OAI21_X1   g12523(.A1(new_n13525_), .A2(new_n13524_), .B(new_n13434_), .ZN(new_n13526_));
  NAND2_X1   g12524(.A1(new_n13526_), .A2(new_n13523_), .ZN(new_n13527_));
  NOR3_X1    g12525(.A1(new_n13502_), .A2(new_n13514_), .A3(new_n13505_), .ZN(new_n13528_));
  NAND3_X1   g12526(.A1(new_n13499_), .A2(new_n11970_), .A3(new_n13495_), .ZN(new_n13529_));
  NAND2_X1   g12527(.A1(new_n13493_), .A2(new_n12002_), .ZN(new_n13530_));
  NOR2_X1    g12528(.A1(new_n13529_), .A2(new_n13530_), .ZN(new_n13531_));
  NOR2_X1    g12529(.A1(new_n13506_), .A2(new_n13508_), .ZN(new_n13532_));
  OAI21_X1   g12530(.A1(new_n13531_), .A2(new_n13532_), .B(new_n13479_), .ZN(new_n13533_));
  NAND2_X1   g12531(.A1(new_n12004_), .A2(new_n11939_), .ZN(new_n13534_));
  AOI21_X1   g12532(.A1(new_n13533_), .A2(new_n13510_), .B(new_n13534_), .ZN(new_n13535_));
  OAI21_X1   g12533(.A1(new_n13528_), .A2(new_n13535_), .B(new_n13527_), .ZN(new_n13536_));
  NAND2_X1   g12534(.A1(new_n13517_), .A2(new_n13536_), .ZN(new_n13537_));
  AOI21_X1   g12535(.A1(new_n12117_), .A2(\A[492] ), .B(new_n12122_), .ZN(new_n13538_));
  XOR2_X1    g12536(.A1(new_n13538_), .A2(new_n12126_), .Z(new_n13539_));
  INV_X1     g12537(.I(new_n12128_), .ZN(new_n13540_));
  XOR2_X1    g12538(.A1(new_n13539_), .A2(new_n13540_), .Z(new_n13541_));
  XNOR2_X1   g12539(.A1(new_n12109_), .A2(new_n12118_), .ZN(new_n13542_));
  NOR2_X1    g12540(.A1(new_n13538_), .A2(new_n12126_), .ZN(new_n13543_));
  AOI21_X1   g12541(.A1(new_n13539_), .A2(new_n12128_), .B(new_n13543_), .ZN(new_n13544_));
  NOR2_X1    g12542(.A1(new_n13544_), .A2(new_n13542_), .ZN(new_n13545_));
  NOR2_X1    g12543(.A1(new_n13541_), .A2(new_n13545_), .ZN(new_n13546_));
  AOI21_X1   g12544(.A1(new_n12087_), .A2(\A[498] ), .B(new_n12092_), .ZN(new_n13547_));
  XOR2_X1    g12545(.A1(new_n13547_), .A2(new_n12096_), .Z(new_n13548_));
  XOR2_X1    g12546(.A1(new_n13548_), .A2(new_n12098_), .Z(new_n13549_));
  INV_X1     g12547(.I(new_n12089_), .ZN(new_n13550_));
  NOR2_X1    g12548(.A1(new_n13550_), .A2(new_n13542_), .ZN(new_n13551_));
  NAND3_X1   g12549(.A1(new_n13549_), .A2(new_n12099_), .A3(new_n13551_), .ZN(new_n13552_));
  XOR2_X1    g12550(.A1(new_n12094_), .A2(new_n12096_), .Z(new_n13553_));
  INV_X1     g12551(.I(new_n12098_), .ZN(new_n13554_));
  NOR2_X1    g12552(.A1(new_n13547_), .A2(new_n12096_), .ZN(new_n13555_));
  INV_X1     g12553(.I(new_n13555_), .ZN(new_n13556_));
  OAI21_X1   g12554(.A1(new_n13553_), .A2(new_n13554_), .B(new_n13556_), .ZN(new_n13557_));
  NAND2_X1   g12555(.A1(new_n13557_), .A2(new_n12089_), .ZN(new_n13558_));
  NAND2_X1   g12556(.A1(new_n13558_), .A2(new_n12129_), .ZN(new_n13559_));
  NOR2_X1    g12557(.A1(new_n13552_), .A2(new_n13559_), .ZN(new_n13560_));
  INV_X1     g12558(.I(new_n12099_), .ZN(new_n13561_));
  INV_X1     g12559(.I(new_n12129_), .ZN(new_n13562_));
  NAND2_X1   g12560(.A1(new_n12089_), .A2(new_n12119_), .ZN(new_n13563_));
  NOR3_X1    g12561(.A1(new_n13563_), .A2(new_n13561_), .A3(new_n13562_), .ZN(new_n13564_));
  XOR2_X1    g12562(.A1(new_n13548_), .A2(new_n13554_), .Z(new_n13565_));
  AOI21_X1   g12563(.A1(new_n13548_), .A2(new_n12098_), .B(new_n13555_), .ZN(new_n13566_));
  NOR2_X1    g12564(.A1(new_n13566_), .A2(new_n13550_), .ZN(new_n13567_));
  NOR2_X1    g12565(.A1(new_n13565_), .A2(new_n13567_), .ZN(new_n13568_));
  NOR2_X1    g12566(.A1(new_n13568_), .A2(new_n13564_), .ZN(new_n13569_));
  OAI21_X1   g12567(.A1(new_n13560_), .A2(new_n13569_), .B(new_n13546_), .ZN(new_n13570_));
  XOR2_X1    g12568(.A1(new_n13539_), .A2(new_n12128_), .Z(new_n13571_));
  XOR2_X1    g12569(.A1(new_n12124_), .A2(new_n12126_), .Z(new_n13572_));
  INV_X1     g12570(.I(new_n13543_), .ZN(new_n13573_));
  OAI21_X1   g12571(.A1(new_n13572_), .A2(new_n13540_), .B(new_n13573_), .ZN(new_n13574_));
  NAND2_X1   g12572(.A1(new_n13574_), .A2(new_n12119_), .ZN(new_n13575_));
  NAND2_X1   g12573(.A1(new_n13571_), .A2(new_n13575_), .ZN(new_n13576_));
  NOR3_X1    g12574(.A1(new_n13564_), .A2(new_n13565_), .A3(new_n13567_), .ZN(new_n13577_));
  NAND3_X1   g12575(.A1(new_n13551_), .A2(new_n12099_), .A3(new_n12129_), .ZN(new_n13578_));
  NOR2_X1    g12576(.A1(new_n13568_), .A2(new_n13578_), .ZN(new_n13579_));
  OAI21_X1   g12577(.A1(new_n13579_), .A2(new_n13577_), .B(new_n13576_), .ZN(new_n13580_));
  NAND2_X1   g12578(.A1(new_n13570_), .A2(new_n13580_), .ZN(new_n13581_));
  NAND2_X1   g12579(.A1(new_n12070_), .A2(new_n12131_), .ZN(new_n13582_));
  XOR2_X1    g12580(.A1(new_n12054_), .A2(new_n12045_), .Z(new_n13583_));
  AOI21_X1   g12581(.A1(new_n12053_), .A2(\A[504] ), .B(new_n12058_), .ZN(new_n13584_));
  XOR2_X1    g12582(.A1(new_n13584_), .A2(new_n12064_), .Z(new_n13585_));
  NOR2_X1    g12583(.A1(new_n13584_), .A2(new_n12064_), .ZN(new_n13586_));
  AOI21_X1   g12584(.A1(new_n13585_), .A2(new_n12067_), .B(new_n13586_), .ZN(new_n13587_));
  INV_X1     g12585(.I(new_n12054_), .ZN(new_n13588_));
  NAND2_X1   g12586(.A1(new_n13588_), .A2(new_n12045_), .ZN(new_n13589_));
  NOR2_X1    g12587(.A1(new_n13585_), .A2(new_n13589_), .ZN(new_n13590_));
  XOR2_X1    g12588(.A1(new_n12060_), .A2(new_n12064_), .Z(new_n13591_));
  NOR2_X1    g12589(.A1(new_n13591_), .A2(new_n12067_), .ZN(new_n13592_));
  OAI22_X1   g12590(.A1(new_n13583_), .A2(new_n13587_), .B1(new_n13590_), .B2(new_n13592_), .ZN(new_n13593_));
  INV_X1     g12591(.I(new_n13593_), .ZN(new_n13594_));
  INV_X1     g12592(.I(new_n12036_), .ZN(new_n13595_));
  INV_X1     g12593(.I(new_n12068_), .ZN(new_n13596_));
  XOR2_X1    g12594(.A1(new_n12028_), .A2(new_n12032_), .Z(new_n13597_));
  NAND2_X1   g12595(.A1(new_n13597_), .A2(new_n12035_), .ZN(new_n13598_));
  AOI21_X1   g12596(.A1(new_n12021_), .A2(\A[510] ), .B(new_n12026_), .ZN(new_n13599_));
  XOR2_X1    g12597(.A1(new_n13599_), .A2(new_n12032_), .Z(new_n13600_));
  INV_X1     g12598(.I(new_n12022_), .ZN(new_n13601_));
  NAND2_X1   g12599(.A1(new_n13601_), .A2(new_n12013_), .ZN(new_n13602_));
  NAND2_X1   g12600(.A1(new_n13600_), .A2(new_n13602_), .ZN(new_n13603_));
  NAND2_X1   g12601(.A1(new_n13598_), .A2(new_n13603_), .ZN(new_n13604_));
  XOR2_X1    g12602(.A1(new_n12022_), .A2(new_n12013_), .Z(new_n13605_));
  NOR2_X1    g12603(.A1(new_n13605_), .A2(new_n13583_), .ZN(new_n13606_));
  NAND2_X1   g12604(.A1(new_n13604_), .A2(new_n13606_), .ZN(new_n13607_));
  NOR2_X1    g12605(.A1(new_n13599_), .A2(new_n12032_), .ZN(new_n13608_));
  AOI21_X1   g12606(.A1(new_n13600_), .A2(new_n12035_), .B(new_n13608_), .ZN(new_n13609_));
  NOR2_X1    g12607(.A1(new_n13609_), .A2(new_n13605_), .ZN(new_n13610_));
  NOR4_X1    g12608(.A1(new_n13607_), .A2(new_n13595_), .A3(new_n13596_), .A4(new_n13610_), .ZN(new_n13611_));
  NAND2_X1   g12609(.A1(new_n12023_), .A2(new_n12055_), .ZN(new_n13612_));
  NOR3_X1    g12610(.A1(new_n13612_), .A2(new_n13595_), .A3(new_n13596_), .ZN(new_n13613_));
  NOR2_X1    g12611(.A1(new_n13600_), .A2(new_n13602_), .ZN(new_n13614_));
  NOR2_X1    g12612(.A1(new_n13597_), .A2(new_n12035_), .ZN(new_n13615_));
  NOR2_X1    g12613(.A1(new_n13615_), .A2(new_n13614_), .ZN(new_n13616_));
  NOR2_X1    g12614(.A1(new_n13610_), .A2(new_n13616_), .ZN(new_n13617_));
  NOR2_X1    g12615(.A1(new_n13617_), .A2(new_n13613_), .ZN(new_n13618_));
  OAI21_X1   g12616(.A1(new_n13611_), .A2(new_n13618_), .B(new_n13594_), .ZN(new_n13619_));
  NAND3_X1   g12617(.A1(new_n13606_), .A2(new_n12036_), .A3(new_n12068_), .ZN(new_n13620_));
  NOR2_X1    g12618(.A1(new_n13617_), .A2(new_n13620_), .ZN(new_n13621_));
  OAI22_X1   g12619(.A1(new_n13605_), .A2(new_n13609_), .B1(new_n13614_), .B2(new_n13615_), .ZN(new_n13622_));
  NOR2_X1    g12620(.A1(new_n13613_), .A2(new_n13622_), .ZN(new_n13623_));
  OAI21_X1   g12621(.A1(new_n13621_), .A2(new_n13623_), .B(new_n13593_), .ZN(new_n13624_));
  AOI21_X1   g12622(.A1(new_n13619_), .A2(new_n13624_), .B(new_n13582_), .ZN(new_n13625_));
  XNOR2_X1   g12623(.A1(new_n12037_), .A2(new_n12069_), .ZN(new_n13626_));
  XNOR2_X1   g12624(.A1(new_n12100_), .A2(new_n12130_), .ZN(new_n13627_));
  NOR2_X1    g12625(.A1(new_n13626_), .A2(new_n13627_), .ZN(new_n13628_));
  NOR3_X1    g12626(.A1(new_n13616_), .A2(new_n13595_), .A3(new_n13612_), .ZN(new_n13629_));
  NOR2_X1    g12627(.A1(new_n13610_), .A2(new_n13596_), .ZN(new_n13630_));
  NAND2_X1   g12628(.A1(new_n13629_), .A2(new_n13630_), .ZN(new_n13631_));
  NAND2_X1   g12629(.A1(new_n13622_), .A2(new_n13620_), .ZN(new_n13632_));
  AOI21_X1   g12630(.A1(new_n13631_), .A2(new_n13632_), .B(new_n13593_), .ZN(new_n13633_));
  NAND2_X1   g12631(.A1(new_n13613_), .A2(new_n13622_), .ZN(new_n13634_));
  NAND2_X1   g12632(.A1(new_n13617_), .A2(new_n13620_), .ZN(new_n13635_));
  AOI21_X1   g12633(.A1(new_n13635_), .A2(new_n13634_), .B(new_n13594_), .ZN(new_n13636_));
  NOR3_X1    g12634(.A1(new_n13633_), .A2(new_n13636_), .A3(new_n13628_), .ZN(new_n13637_));
  OAI21_X1   g12635(.A1(new_n13637_), .A2(new_n13625_), .B(new_n13581_), .ZN(new_n13638_));
  NOR3_X1    g12636(.A1(new_n13565_), .A2(new_n13561_), .A3(new_n13563_), .ZN(new_n13639_));
  NOR2_X1    g12637(.A1(new_n13567_), .A2(new_n13562_), .ZN(new_n13640_));
  NAND2_X1   g12638(.A1(new_n13639_), .A2(new_n13640_), .ZN(new_n13641_));
  NAND2_X1   g12639(.A1(new_n13549_), .A2(new_n13558_), .ZN(new_n13642_));
  NAND2_X1   g12640(.A1(new_n13642_), .A2(new_n13578_), .ZN(new_n13643_));
  AOI21_X1   g12641(.A1(new_n13641_), .A2(new_n13643_), .B(new_n13576_), .ZN(new_n13644_));
  INV_X1     g12642(.I(new_n13577_), .ZN(new_n13645_));
  NAND2_X1   g12643(.A1(new_n13642_), .A2(new_n13564_), .ZN(new_n13646_));
  AOI21_X1   g12644(.A1(new_n13645_), .A2(new_n13646_), .B(new_n13546_), .ZN(new_n13647_));
  NOR2_X1    g12645(.A1(new_n13647_), .A2(new_n13644_), .ZN(new_n13648_));
  AOI21_X1   g12646(.A1(new_n13619_), .A2(new_n13624_), .B(new_n13628_), .ZN(new_n13649_));
  NAND3_X1   g12647(.A1(new_n13619_), .A2(new_n13624_), .A3(new_n13628_), .ZN(new_n13650_));
  INV_X1     g12648(.I(new_n13650_), .ZN(new_n13651_));
  OAI21_X1   g12649(.A1(new_n13651_), .A2(new_n13649_), .B(new_n13648_), .ZN(new_n13652_));
  XOR2_X1    g12650(.A1(new_n13504_), .A2(new_n11939_), .Z(new_n13653_));
  XOR2_X1    g12651(.A1(new_n12070_), .A2(new_n13627_), .Z(new_n13654_));
  NOR2_X1    g12652(.A1(new_n13653_), .A2(new_n13654_), .ZN(new_n13655_));
  NAND3_X1   g12653(.A1(new_n13652_), .A2(new_n13638_), .A3(new_n13655_), .ZN(new_n13656_));
  OAI21_X1   g12654(.A1(new_n13633_), .A2(new_n13636_), .B(new_n13628_), .ZN(new_n13657_));
  NAND3_X1   g12655(.A1(new_n13619_), .A2(new_n13624_), .A3(new_n13582_), .ZN(new_n13658_));
  AOI21_X1   g12656(.A1(new_n13657_), .A2(new_n13658_), .B(new_n13648_), .ZN(new_n13659_));
  OAI21_X1   g12657(.A1(new_n13633_), .A2(new_n13636_), .B(new_n13582_), .ZN(new_n13660_));
  AOI21_X1   g12658(.A1(new_n13660_), .A2(new_n13650_), .B(new_n13581_), .ZN(new_n13661_));
  NAND2_X1   g12659(.A1(new_n12005_), .A2(new_n12132_), .ZN(new_n13662_));
  OAI21_X1   g12660(.A1(new_n13659_), .A2(new_n13661_), .B(new_n13662_), .ZN(new_n13663_));
  AOI21_X1   g12661(.A1(new_n13663_), .A2(new_n13656_), .B(new_n13537_), .ZN(new_n13664_));
  NAND3_X1   g12662(.A1(new_n13533_), .A2(new_n13510_), .A3(new_n13534_), .ZN(new_n13665_));
  OAI21_X1   g12663(.A1(new_n13502_), .A2(new_n13514_), .B(new_n13505_), .ZN(new_n13666_));
  AOI21_X1   g12664(.A1(new_n13666_), .A2(new_n13665_), .B(new_n13468_), .ZN(new_n13667_));
  AOI21_X1   g12665(.A1(new_n13468_), .A2(new_n13516_), .B(new_n13667_), .ZN(new_n13668_));
  NAND3_X1   g12666(.A1(new_n13652_), .A2(new_n13638_), .A3(new_n13662_), .ZN(new_n13669_));
  OAI21_X1   g12667(.A1(new_n13659_), .A2(new_n13661_), .B(new_n13655_), .ZN(new_n13670_));
  AOI21_X1   g12668(.A1(new_n13669_), .A2(new_n13670_), .B(new_n13668_), .ZN(new_n13671_));
  NOR2_X1    g12669(.A1(new_n13664_), .A2(new_n13671_), .ZN(new_n13672_));
  AOI21_X1   g12670(.A1(new_n12375_), .A2(\A[516] ), .B(new_n12380_), .ZN(new_n13673_));
  XOR2_X1    g12671(.A1(new_n13673_), .A2(new_n12386_), .Z(new_n13674_));
  XOR2_X1    g12672(.A1(new_n13674_), .A2(new_n12389_), .Z(new_n13675_));
  XOR2_X1    g12673(.A1(new_n12382_), .A2(new_n12386_), .Z(new_n13676_));
  INV_X1     g12674(.I(new_n12376_), .ZN(new_n13677_));
  NAND2_X1   g12675(.A1(new_n13677_), .A2(new_n12367_), .ZN(new_n13678_));
  NOR2_X1    g12676(.A1(new_n13673_), .A2(new_n12386_), .ZN(new_n13679_));
  INV_X1     g12677(.I(new_n13679_), .ZN(new_n13680_));
  OAI21_X1   g12678(.A1(new_n13676_), .A2(new_n13678_), .B(new_n13680_), .ZN(new_n13681_));
  NAND2_X1   g12679(.A1(new_n13681_), .A2(new_n12377_), .ZN(new_n13682_));
  NAND2_X1   g12680(.A1(new_n13675_), .A2(new_n13682_), .ZN(new_n13683_));
  AOI21_X1   g12681(.A1(new_n12343_), .A2(\A[522] ), .B(new_n12348_), .ZN(new_n13684_));
  XOR2_X1    g12682(.A1(new_n13684_), .A2(new_n12354_), .Z(new_n13685_));
  INV_X1     g12683(.I(new_n12344_), .ZN(new_n13686_));
  NAND2_X1   g12684(.A1(new_n13686_), .A2(new_n12335_), .ZN(new_n13687_));
  XOR2_X1    g12685(.A1(new_n13685_), .A2(new_n13687_), .Z(new_n13688_));
  INV_X1     g12686(.I(new_n12358_), .ZN(new_n13689_));
  NAND2_X1   g12687(.A1(new_n12345_), .A2(new_n12377_), .ZN(new_n13690_));
  NOR3_X1    g12688(.A1(new_n13688_), .A2(new_n13689_), .A3(new_n13690_), .ZN(new_n13691_));
  INV_X1     g12689(.I(new_n12390_), .ZN(new_n13692_));
  INV_X1     g12690(.I(new_n12345_), .ZN(new_n13693_));
  NOR2_X1    g12691(.A1(new_n13684_), .A2(new_n12354_), .ZN(new_n13694_));
  AOI21_X1   g12692(.A1(new_n13685_), .A2(new_n12357_), .B(new_n13694_), .ZN(new_n13695_));
  NOR2_X1    g12693(.A1(new_n13695_), .A2(new_n13693_), .ZN(new_n13696_));
  NOR2_X1    g12694(.A1(new_n13696_), .A2(new_n13692_), .ZN(new_n13697_));
  NAND2_X1   g12695(.A1(new_n13691_), .A2(new_n13697_), .ZN(new_n13698_));
  XOR2_X1    g12696(.A1(new_n12376_), .A2(new_n12367_), .Z(new_n13699_));
  NOR2_X1    g12697(.A1(new_n13693_), .A2(new_n13699_), .ZN(new_n13700_));
  NAND3_X1   g12698(.A1(new_n13700_), .A2(new_n12358_), .A3(new_n12390_), .ZN(new_n13701_));
  XOR2_X1    g12699(.A1(new_n13685_), .A2(new_n12357_), .Z(new_n13702_));
  XOR2_X1    g12700(.A1(new_n12350_), .A2(new_n12354_), .Z(new_n13703_));
  INV_X1     g12701(.I(new_n13694_), .ZN(new_n13704_));
  OAI21_X1   g12702(.A1(new_n13703_), .A2(new_n13687_), .B(new_n13704_), .ZN(new_n13705_));
  NAND2_X1   g12703(.A1(new_n13705_), .A2(new_n12345_), .ZN(new_n13706_));
  NAND2_X1   g12704(.A1(new_n13702_), .A2(new_n13706_), .ZN(new_n13707_));
  NAND2_X1   g12705(.A1(new_n13707_), .A2(new_n13701_), .ZN(new_n13708_));
  AOI21_X1   g12706(.A1(new_n13698_), .A2(new_n13708_), .B(new_n13683_), .ZN(new_n13709_));
  XOR2_X1    g12707(.A1(new_n13707_), .A2(new_n13701_), .Z(new_n13710_));
  AOI21_X1   g12708(.A1(new_n13710_), .A2(new_n13683_), .B(new_n13709_), .ZN(new_n13711_));
  XOR2_X1    g12709(.A1(new_n12311_), .A2(new_n12302_), .Z(new_n13712_));
  AOI21_X1   g12710(.A1(new_n12310_), .A2(\A[528] ), .B(new_n12315_), .ZN(new_n13713_));
  XOR2_X1    g12711(.A1(new_n13713_), .A2(new_n12321_), .Z(new_n13714_));
  NOR2_X1    g12712(.A1(new_n13713_), .A2(new_n12321_), .ZN(new_n13715_));
  AOI21_X1   g12713(.A1(new_n13714_), .A2(new_n12324_), .B(new_n13715_), .ZN(new_n13716_));
  XOR2_X1    g12714(.A1(new_n12317_), .A2(new_n12321_), .Z(new_n13717_));
  NAND2_X1   g12715(.A1(new_n13717_), .A2(new_n12324_), .ZN(new_n13718_));
  INV_X1     g12716(.I(new_n12311_), .ZN(new_n13719_));
  NAND2_X1   g12717(.A1(new_n13719_), .A2(new_n12302_), .ZN(new_n13720_));
  NAND2_X1   g12718(.A1(new_n13714_), .A2(new_n13720_), .ZN(new_n13721_));
  NAND2_X1   g12719(.A1(new_n13718_), .A2(new_n13721_), .ZN(new_n13722_));
  OAI21_X1   g12720(.A1(new_n13712_), .A2(new_n13716_), .B(new_n13722_), .ZN(new_n13723_));
  AOI21_X1   g12721(.A1(new_n12278_), .A2(\A[534] ), .B(new_n12283_), .ZN(new_n13724_));
  XOR2_X1    g12722(.A1(new_n13724_), .A2(new_n12289_), .Z(new_n13725_));
  INV_X1     g12723(.I(new_n12279_), .ZN(new_n13726_));
  NAND2_X1   g12724(.A1(new_n13726_), .A2(new_n12270_), .ZN(new_n13727_));
  NOR2_X1    g12725(.A1(new_n13725_), .A2(new_n13727_), .ZN(new_n13728_));
  XOR2_X1    g12726(.A1(new_n12285_), .A2(new_n12289_), .Z(new_n13729_));
  NOR2_X1    g12727(.A1(new_n13729_), .A2(new_n12292_), .ZN(new_n13730_));
  NOR2_X1    g12728(.A1(new_n13730_), .A2(new_n13728_), .ZN(new_n13731_));
  NAND2_X1   g12729(.A1(new_n12280_), .A2(new_n12312_), .ZN(new_n13732_));
  NOR2_X1    g12730(.A1(new_n13731_), .A2(new_n13732_), .ZN(new_n13733_));
  NAND2_X1   g12731(.A1(new_n12290_), .A2(new_n12285_), .ZN(new_n13734_));
  OAI21_X1   g12732(.A1(new_n13729_), .A2(new_n13727_), .B(new_n13734_), .ZN(new_n13735_));
  NAND2_X1   g12733(.A1(new_n13735_), .A2(new_n12280_), .ZN(new_n13736_));
  NAND4_X1   g12734(.A1(new_n13733_), .A2(new_n12293_), .A3(new_n12325_), .A4(new_n13736_), .ZN(new_n13737_));
  XOR2_X1    g12735(.A1(new_n12279_), .A2(new_n12270_), .Z(new_n13738_));
  NOR2_X1    g12736(.A1(new_n13738_), .A2(new_n13712_), .ZN(new_n13739_));
  NAND3_X1   g12737(.A1(new_n13739_), .A2(new_n12293_), .A3(new_n12325_), .ZN(new_n13740_));
  NAND2_X1   g12738(.A1(new_n13729_), .A2(new_n12292_), .ZN(new_n13741_));
  NAND2_X1   g12739(.A1(new_n13725_), .A2(new_n13727_), .ZN(new_n13742_));
  NAND2_X1   g12740(.A1(new_n13741_), .A2(new_n13742_), .ZN(new_n13743_));
  NAND2_X1   g12741(.A1(new_n13736_), .A2(new_n13743_), .ZN(new_n13744_));
  NAND2_X1   g12742(.A1(new_n13744_), .A2(new_n13740_), .ZN(new_n13745_));
  AOI21_X1   g12743(.A1(new_n13737_), .A2(new_n13745_), .B(new_n13723_), .ZN(new_n13746_));
  INV_X1     g12744(.I(new_n13716_), .ZN(new_n13747_));
  NOR2_X1    g12745(.A1(new_n13714_), .A2(new_n13720_), .ZN(new_n13748_));
  NOR2_X1    g12746(.A1(new_n13717_), .A2(new_n12324_), .ZN(new_n13749_));
  NOR2_X1    g12747(.A1(new_n13749_), .A2(new_n13748_), .ZN(new_n13750_));
  AOI21_X1   g12748(.A1(new_n12312_), .A2(new_n13747_), .B(new_n13750_), .ZN(new_n13751_));
  AND4_X2    g12749(.A1(new_n12280_), .A2(new_n12293_), .A3(new_n12325_), .A4(new_n12312_), .Z(new_n13752_));
  NAND2_X1   g12750(.A1(new_n13744_), .A2(new_n13752_), .ZN(new_n13753_));
  AOI22_X1   g12751(.A1(new_n13735_), .A2(new_n12280_), .B1(new_n13741_), .B2(new_n13742_), .ZN(new_n13754_));
  NAND2_X1   g12752(.A1(new_n13754_), .A2(new_n13740_), .ZN(new_n13755_));
  AOI21_X1   g12753(.A1(new_n13753_), .A2(new_n13755_), .B(new_n13751_), .ZN(new_n13756_));
  NAND2_X1   g12754(.A1(new_n12327_), .A2(new_n12392_), .ZN(new_n13757_));
  NOR3_X1    g12755(.A1(new_n13746_), .A2(new_n13756_), .A3(new_n13757_), .ZN(new_n13758_));
  NAND3_X1   g12756(.A1(new_n13743_), .A2(new_n12293_), .A3(new_n13739_), .ZN(new_n13759_));
  NAND2_X1   g12757(.A1(new_n13736_), .A2(new_n12325_), .ZN(new_n13760_));
  NOR2_X1    g12758(.A1(new_n13759_), .A2(new_n13760_), .ZN(new_n13761_));
  NOR2_X1    g12759(.A1(new_n13754_), .A2(new_n13752_), .ZN(new_n13762_));
  OAI21_X1   g12760(.A1(new_n13761_), .A2(new_n13762_), .B(new_n13751_), .ZN(new_n13763_));
  NOR2_X1    g12761(.A1(new_n13754_), .A2(new_n13740_), .ZN(new_n13764_));
  NOR2_X1    g12762(.A1(new_n13744_), .A2(new_n13752_), .ZN(new_n13765_));
  OAI21_X1   g12763(.A1(new_n13765_), .A2(new_n13764_), .B(new_n13723_), .ZN(new_n13766_));
  XNOR2_X1   g12764(.A1(new_n12294_), .A2(new_n12326_), .ZN(new_n13767_));
  XNOR2_X1   g12765(.A1(new_n12359_), .A2(new_n12391_), .ZN(new_n13768_));
  NOR2_X1    g12766(.A1(new_n13767_), .A2(new_n13768_), .ZN(new_n13769_));
  AOI21_X1   g12767(.A1(new_n13763_), .A2(new_n13766_), .B(new_n13769_), .ZN(new_n13770_));
  NOR2_X1    g12768(.A1(new_n13770_), .A2(new_n13758_), .ZN(new_n13771_));
  NOR3_X1    g12769(.A1(new_n13746_), .A2(new_n13769_), .A3(new_n13756_), .ZN(new_n13772_));
  AOI21_X1   g12770(.A1(new_n13763_), .A2(new_n13766_), .B(new_n13757_), .ZN(new_n13773_));
  NOR2_X1    g12771(.A1(new_n13772_), .A2(new_n13773_), .ZN(new_n13774_));
  MUX2_X1    g12772(.I0(new_n13774_), .I1(new_n13771_), .S(new_n13711_), .Z(new_n13775_));
  XOR2_X1    g12773(.A1(new_n12254_), .A2(new_n12256_), .Z(new_n13776_));
  INV_X1     g12774(.I(new_n12258_), .ZN(new_n13777_));
  AOI21_X1   g12775(.A1(new_n12247_), .A2(\A[540] ), .B(new_n12252_), .ZN(new_n13778_));
  NOR2_X1    g12776(.A1(new_n13778_), .A2(new_n12256_), .ZN(new_n13779_));
  INV_X1     g12777(.I(new_n13779_), .ZN(new_n13780_));
  OAI21_X1   g12778(.A1(new_n13776_), .A2(new_n13777_), .B(new_n13780_), .ZN(new_n13781_));
  NAND2_X1   g12779(.A1(new_n13776_), .A2(new_n12258_), .ZN(new_n13782_));
  XOR2_X1    g12780(.A1(new_n13778_), .A2(new_n12256_), .Z(new_n13783_));
  NAND2_X1   g12781(.A1(new_n13783_), .A2(new_n13777_), .ZN(new_n13784_));
  AOI22_X1   g12782(.A1(new_n13781_), .A2(new_n12249_), .B1(new_n13782_), .B2(new_n13784_), .ZN(new_n13785_));
  INV_X1     g12783(.I(new_n12229_), .ZN(new_n13786_));
  INV_X1     g12784(.I(new_n12259_), .ZN(new_n13787_));
  XOR2_X1    g12785(.A1(new_n12221_), .A2(new_n12225_), .Z(new_n13788_));
  NAND2_X1   g12786(.A1(new_n13788_), .A2(new_n12228_), .ZN(new_n13789_));
  AOI21_X1   g12787(.A1(new_n12214_), .A2(\A[546] ), .B(new_n12219_), .ZN(new_n13790_));
  XOR2_X1    g12788(.A1(new_n13790_), .A2(new_n12225_), .Z(new_n13791_));
  INV_X1     g12789(.I(new_n12215_), .ZN(new_n13792_));
  NAND2_X1   g12790(.A1(new_n13792_), .A2(new_n12206_), .ZN(new_n13793_));
  NAND2_X1   g12791(.A1(new_n13791_), .A2(new_n13793_), .ZN(new_n13794_));
  NAND2_X1   g12792(.A1(new_n13789_), .A2(new_n13794_), .ZN(new_n13795_));
  XOR2_X1    g12793(.A1(new_n12215_), .A2(new_n12206_), .Z(new_n13796_));
  XNOR2_X1   g12794(.A1(new_n12239_), .A2(new_n12248_), .ZN(new_n13797_));
  NOR2_X1    g12795(.A1(new_n13797_), .A2(new_n13796_), .ZN(new_n13798_));
  NAND2_X1   g12796(.A1(new_n13795_), .A2(new_n13798_), .ZN(new_n13799_));
  NOR2_X1    g12797(.A1(new_n13790_), .A2(new_n12225_), .ZN(new_n13800_));
  AOI21_X1   g12798(.A1(new_n13791_), .A2(new_n12228_), .B(new_n13800_), .ZN(new_n13801_));
  NOR2_X1    g12799(.A1(new_n13801_), .A2(new_n13796_), .ZN(new_n13802_));
  NOR4_X1    g12800(.A1(new_n13799_), .A2(new_n13786_), .A3(new_n13787_), .A4(new_n13802_), .ZN(new_n13803_));
  NAND2_X1   g12801(.A1(new_n12216_), .A2(new_n12249_), .ZN(new_n13804_));
  NOR3_X1    g12802(.A1(new_n13804_), .A2(new_n13786_), .A3(new_n13787_), .ZN(new_n13805_));
  NOR2_X1    g12803(.A1(new_n13791_), .A2(new_n13793_), .ZN(new_n13806_));
  NOR2_X1    g12804(.A1(new_n13788_), .A2(new_n12228_), .ZN(new_n13807_));
  NOR2_X1    g12805(.A1(new_n13807_), .A2(new_n13806_), .ZN(new_n13808_));
  NOR2_X1    g12806(.A1(new_n13802_), .A2(new_n13808_), .ZN(new_n13809_));
  NOR2_X1    g12807(.A1(new_n13809_), .A2(new_n13805_), .ZN(new_n13810_));
  OAI21_X1   g12808(.A1(new_n13803_), .A2(new_n13810_), .B(new_n13785_), .ZN(new_n13811_));
  INV_X1     g12809(.I(new_n13785_), .ZN(new_n13812_));
  INV_X1     g12810(.I(new_n13800_), .ZN(new_n13813_));
  OAI21_X1   g12811(.A1(new_n13788_), .A2(new_n13793_), .B(new_n13813_), .ZN(new_n13814_));
  NAND2_X1   g12812(.A1(new_n13814_), .A2(new_n12216_), .ZN(new_n13815_));
  NAND2_X1   g12813(.A1(new_n13815_), .A2(new_n13795_), .ZN(new_n13816_));
  NOR2_X1    g12814(.A1(new_n13816_), .A2(new_n13805_), .ZN(new_n13817_));
  NAND3_X1   g12815(.A1(new_n13798_), .A2(new_n12229_), .A3(new_n12259_), .ZN(new_n13818_));
  NOR2_X1    g12816(.A1(new_n13809_), .A2(new_n13818_), .ZN(new_n13819_));
  OAI21_X1   g12817(.A1(new_n13819_), .A2(new_n13817_), .B(new_n13812_), .ZN(new_n13820_));
  NAND2_X1   g12818(.A1(new_n13811_), .A2(new_n13820_), .ZN(new_n13821_));
  NAND2_X1   g12819(.A1(new_n12198_), .A2(new_n12261_), .ZN(new_n13822_));
  XOR2_X1    g12820(.A1(new_n12182_), .A2(new_n12173_), .Z(new_n13823_));
  AOI21_X1   g12821(.A1(new_n12181_), .A2(\A[552] ), .B(new_n12186_), .ZN(new_n13824_));
  XOR2_X1    g12822(.A1(new_n13824_), .A2(new_n12192_), .Z(new_n13825_));
  NOR2_X1    g12823(.A1(new_n13824_), .A2(new_n12192_), .ZN(new_n13826_));
  AOI21_X1   g12824(.A1(new_n13825_), .A2(new_n12195_), .B(new_n13826_), .ZN(new_n13827_));
  INV_X1     g12825(.I(new_n12182_), .ZN(new_n13828_));
  NAND2_X1   g12826(.A1(new_n13828_), .A2(new_n12173_), .ZN(new_n13829_));
  NOR2_X1    g12827(.A1(new_n13825_), .A2(new_n13829_), .ZN(new_n13830_));
  XOR2_X1    g12828(.A1(new_n12188_), .A2(new_n12192_), .Z(new_n13831_));
  NOR2_X1    g12829(.A1(new_n13831_), .A2(new_n12195_), .ZN(new_n13832_));
  OAI22_X1   g12830(.A1(new_n13823_), .A2(new_n13827_), .B1(new_n13830_), .B2(new_n13832_), .ZN(new_n13833_));
  INV_X1     g12831(.I(new_n13833_), .ZN(new_n13834_));
  INV_X1     g12832(.I(new_n12164_), .ZN(new_n13835_));
  INV_X1     g12833(.I(new_n12196_), .ZN(new_n13836_));
  XOR2_X1    g12834(.A1(new_n12156_), .A2(new_n12160_), .Z(new_n13837_));
  NAND2_X1   g12835(.A1(new_n13837_), .A2(new_n12163_), .ZN(new_n13838_));
  AOI21_X1   g12836(.A1(new_n12149_), .A2(\A[558] ), .B(new_n12154_), .ZN(new_n13839_));
  XOR2_X1    g12837(.A1(new_n13839_), .A2(new_n12160_), .Z(new_n13840_));
  INV_X1     g12838(.I(new_n12150_), .ZN(new_n13841_));
  NAND2_X1   g12839(.A1(new_n13841_), .A2(new_n12141_), .ZN(new_n13842_));
  NAND2_X1   g12840(.A1(new_n13840_), .A2(new_n13842_), .ZN(new_n13843_));
  NAND2_X1   g12841(.A1(new_n13838_), .A2(new_n13843_), .ZN(new_n13844_));
  XOR2_X1    g12842(.A1(new_n12150_), .A2(new_n12141_), .Z(new_n13845_));
  NOR2_X1    g12843(.A1(new_n13845_), .A2(new_n13823_), .ZN(new_n13846_));
  NAND2_X1   g12844(.A1(new_n13844_), .A2(new_n13846_), .ZN(new_n13847_));
  NOR2_X1    g12845(.A1(new_n13839_), .A2(new_n12160_), .ZN(new_n13848_));
  AOI21_X1   g12846(.A1(new_n13840_), .A2(new_n12163_), .B(new_n13848_), .ZN(new_n13849_));
  NOR2_X1    g12847(.A1(new_n13849_), .A2(new_n13845_), .ZN(new_n13850_));
  NOR4_X1    g12848(.A1(new_n13847_), .A2(new_n13835_), .A3(new_n13836_), .A4(new_n13850_), .ZN(new_n13851_));
  NAND2_X1   g12849(.A1(new_n12151_), .A2(new_n12183_), .ZN(new_n13852_));
  NOR3_X1    g12850(.A1(new_n13852_), .A2(new_n13835_), .A3(new_n13836_), .ZN(new_n13853_));
  NOR2_X1    g12851(.A1(new_n13840_), .A2(new_n13842_), .ZN(new_n13854_));
  NOR2_X1    g12852(.A1(new_n13837_), .A2(new_n12163_), .ZN(new_n13855_));
  NOR2_X1    g12853(.A1(new_n13855_), .A2(new_n13854_), .ZN(new_n13856_));
  NOR2_X1    g12854(.A1(new_n13850_), .A2(new_n13856_), .ZN(new_n13857_));
  NOR2_X1    g12855(.A1(new_n13857_), .A2(new_n13853_), .ZN(new_n13858_));
  OAI21_X1   g12856(.A1(new_n13851_), .A2(new_n13858_), .B(new_n13834_), .ZN(new_n13859_));
  NAND3_X1   g12857(.A1(new_n13846_), .A2(new_n12164_), .A3(new_n12196_), .ZN(new_n13860_));
  NOR2_X1    g12858(.A1(new_n13857_), .A2(new_n13860_), .ZN(new_n13861_));
  OAI22_X1   g12859(.A1(new_n13845_), .A2(new_n13849_), .B1(new_n13854_), .B2(new_n13855_), .ZN(new_n13862_));
  NOR2_X1    g12860(.A1(new_n13853_), .A2(new_n13862_), .ZN(new_n13863_));
  OAI21_X1   g12861(.A1(new_n13861_), .A2(new_n13863_), .B(new_n13833_), .ZN(new_n13864_));
  AOI21_X1   g12862(.A1(new_n13859_), .A2(new_n13864_), .B(new_n13822_), .ZN(new_n13865_));
  XNOR2_X1   g12863(.A1(new_n12165_), .A2(new_n12197_), .ZN(new_n13866_));
  XNOR2_X1   g12864(.A1(new_n12230_), .A2(new_n12260_), .ZN(new_n13867_));
  NOR2_X1    g12865(.A1(new_n13866_), .A2(new_n13867_), .ZN(new_n13868_));
  NOR3_X1    g12866(.A1(new_n13856_), .A2(new_n13835_), .A3(new_n13852_), .ZN(new_n13869_));
  NOR2_X1    g12867(.A1(new_n13850_), .A2(new_n13836_), .ZN(new_n13870_));
  NAND2_X1   g12868(.A1(new_n13869_), .A2(new_n13870_), .ZN(new_n13871_));
  NAND2_X1   g12869(.A1(new_n13862_), .A2(new_n13860_), .ZN(new_n13872_));
  AOI21_X1   g12870(.A1(new_n13871_), .A2(new_n13872_), .B(new_n13833_), .ZN(new_n13873_));
  NAND2_X1   g12871(.A1(new_n13853_), .A2(new_n13862_), .ZN(new_n13874_));
  NAND2_X1   g12872(.A1(new_n13857_), .A2(new_n13860_), .ZN(new_n13875_));
  AOI21_X1   g12873(.A1(new_n13875_), .A2(new_n13874_), .B(new_n13834_), .ZN(new_n13876_));
  NOR3_X1    g12874(.A1(new_n13873_), .A2(new_n13876_), .A3(new_n13868_), .ZN(new_n13877_));
  OAI21_X1   g12875(.A1(new_n13865_), .A2(new_n13877_), .B(new_n13821_), .ZN(new_n13878_));
  NOR2_X1    g12876(.A1(new_n13808_), .A2(new_n13804_), .ZN(new_n13879_));
  NAND4_X1   g12877(.A1(new_n13879_), .A2(new_n12229_), .A3(new_n12259_), .A4(new_n13815_), .ZN(new_n13880_));
  NAND2_X1   g12878(.A1(new_n13816_), .A2(new_n13818_), .ZN(new_n13881_));
  AOI21_X1   g12879(.A1(new_n13880_), .A2(new_n13881_), .B(new_n13812_), .ZN(new_n13882_));
  NAND2_X1   g12880(.A1(new_n13809_), .A2(new_n13818_), .ZN(new_n13883_));
  NAND2_X1   g12881(.A1(new_n13816_), .A2(new_n13805_), .ZN(new_n13884_));
  AOI21_X1   g12882(.A1(new_n13883_), .A2(new_n13884_), .B(new_n13785_), .ZN(new_n13885_));
  NOR2_X1    g12883(.A1(new_n13882_), .A2(new_n13885_), .ZN(new_n13886_));
  AOI21_X1   g12884(.A1(new_n13859_), .A2(new_n13864_), .B(new_n13868_), .ZN(new_n13887_));
  NOR3_X1    g12885(.A1(new_n13873_), .A2(new_n13876_), .A3(new_n13822_), .ZN(new_n13888_));
  OAI21_X1   g12886(.A1(new_n13887_), .A2(new_n13888_), .B(new_n13886_), .ZN(new_n13889_));
  NAND2_X1   g12887(.A1(new_n12393_), .A2(new_n12262_), .ZN(new_n13890_));
  NAND3_X1   g12888(.A1(new_n13889_), .A2(new_n13878_), .A3(new_n13890_), .ZN(new_n13891_));
  OAI21_X1   g12889(.A1(new_n13873_), .A2(new_n13876_), .B(new_n13868_), .ZN(new_n13892_));
  NAND3_X1   g12890(.A1(new_n13859_), .A2(new_n13864_), .A3(new_n13822_), .ZN(new_n13893_));
  AOI21_X1   g12891(.A1(new_n13892_), .A2(new_n13893_), .B(new_n13886_), .ZN(new_n13894_));
  OAI21_X1   g12892(.A1(new_n13873_), .A2(new_n13876_), .B(new_n13822_), .ZN(new_n13895_));
  NAND3_X1   g12893(.A1(new_n13859_), .A2(new_n13864_), .A3(new_n13868_), .ZN(new_n13896_));
  AOI21_X1   g12894(.A1(new_n13895_), .A2(new_n13896_), .B(new_n13821_), .ZN(new_n13897_));
  XOR2_X1    g12895(.A1(new_n13866_), .A2(new_n12261_), .Z(new_n13898_));
  XOR2_X1    g12896(.A1(new_n13767_), .A2(new_n12392_), .Z(new_n13899_));
  NOR2_X1    g12897(.A1(new_n13899_), .A2(new_n13898_), .ZN(new_n13900_));
  OAI21_X1   g12898(.A1(new_n13894_), .A2(new_n13897_), .B(new_n13900_), .ZN(new_n13901_));
  AOI21_X1   g12899(.A1(new_n13891_), .A2(new_n13901_), .B(new_n13775_), .ZN(new_n13902_));
  XOR2_X1    g12900(.A1(new_n13674_), .A2(new_n13678_), .Z(new_n13903_));
  AOI21_X1   g12901(.A1(new_n13674_), .A2(new_n12389_), .B(new_n13679_), .ZN(new_n13904_));
  NOR2_X1    g12902(.A1(new_n13904_), .A2(new_n13699_), .ZN(new_n13905_));
  NOR2_X1    g12903(.A1(new_n13903_), .A2(new_n13905_), .ZN(new_n13906_));
  NAND3_X1   g12904(.A1(new_n13702_), .A2(new_n12358_), .A3(new_n13700_), .ZN(new_n13907_));
  NAND2_X1   g12905(.A1(new_n13706_), .A2(new_n12390_), .ZN(new_n13908_));
  NOR2_X1    g12906(.A1(new_n13907_), .A2(new_n13908_), .ZN(new_n13909_));
  NOR3_X1    g12907(.A1(new_n13690_), .A2(new_n13689_), .A3(new_n13692_), .ZN(new_n13910_));
  NOR2_X1    g12908(.A1(new_n13688_), .A2(new_n13696_), .ZN(new_n13911_));
  NOR2_X1    g12909(.A1(new_n13911_), .A2(new_n13910_), .ZN(new_n13912_));
  OAI21_X1   g12910(.A1(new_n13909_), .A2(new_n13912_), .B(new_n13906_), .ZN(new_n13913_));
  NOR2_X1    g12911(.A1(new_n13707_), .A2(new_n13910_), .ZN(new_n13914_));
  NOR2_X1    g12912(.A1(new_n13911_), .A2(new_n13701_), .ZN(new_n13915_));
  OAI21_X1   g12913(.A1(new_n13915_), .A2(new_n13914_), .B(new_n13683_), .ZN(new_n13916_));
  NAND2_X1   g12914(.A1(new_n13913_), .A2(new_n13916_), .ZN(new_n13917_));
  OAI21_X1   g12915(.A1(new_n13773_), .A2(new_n13772_), .B(new_n13917_), .ZN(new_n13918_));
  OAI21_X1   g12916(.A1(new_n13917_), .A2(new_n13771_), .B(new_n13918_), .ZN(new_n13919_));
  NAND3_X1   g12917(.A1(new_n13889_), .A2(new_n13878_), .A3(new_n13900_), .ZN(new_n13920_));
  NAND2_X1   g12918(.A1(new_n13889_), .A2(new_n13878_), .ZN(new_n13921_));
  NAND2_X1   g12919(.A1(new_n13921_), .A2(new_n13890_), .ZN(new_n13922_));
  AOI21_X1   g12920(.A1(new_n13922_), .A2(new_n13920_), .B(new_n13919_), .ZN(new_n13923_));
  NAND2_X1   g12921(.A1(new_n12133_), .A2(new_n12394_), .ZN(new_n13924_));
  NOR3_X1    g12922(.A1(new_n13923_), .A2(new_n13902_), .A3(new_n13924_), .ZN(new_n13925_));
  INV_X1     g12923(.I(new_n13924_), .ZN(new_n13926_));
  NOR2_X1    g12924(.A1(new_n13923_), .A2(new_n13902_), .ZN(new_n13927_));
  NOR2_X1    g12925(.A1(new_n13927_), .A2(new_n13926_), .ZN(new_n13928_));
  OAI21_X1   g12926(.A1(new_n13928_), .A2(new_n13925_), .B(new_n13672_), .ZN(new_n13929_));
  NOR3_X1    g12927(.A1(new_n13923_), .A2(new_n13902_), .A3(new_n13926_), .ZN(new_n13930_));
  NOR2_X1    g12928(.A1(new_n13927_), .A2(new_n13924_), .ZN(new_n13931_));
  OAI22_X1   g12929(.A1(new_n13931_), .A2(new_n13930_), .B1(new_n13664_), .B2(new_n13671_), .ZN(new_n13932_));
  NAND2_X1   g12930(.A1(new_n13932_), .A2(new_n13929_), .ZN(new_n13933_));
  INV_X1     g12931(.I(new_n13933_), .ZN(new_n13934_));
  NOR3_X1    g12932(.A1(new_n13418_), .A2(new_n12914_), .A3(new_n13421_), .ZN(new_n13935_));
  OAI21_X1   g12933(.A1(new_n13934_), .A2(new_n13935_), .B(new_n13422_), .ZN(new_n13936_));
  NOR2_X1    g12934(.A1(new_n13930_), .A2(new_n13672_), .ZN(new_n13937_));
  NOR2_X1    g12935(.A1(new_n13937_), .A2(new_n13931_), .ZN(new_n13938_));
  NOR3_X1    g12936(.A1(new_n13659_), .A2(new_n13661_), .A3(new_n13655_), .ZN(new_n13939_));
  OAI21_X1   g12937(.A1(new_n13668_), .A2(new_n13939_), .B(new_n13670_), .ZN(new_n13940_));
  AOI21_X1   g12938(.A1(new_n13527_), .A2(new_n13665_), .B(new_n13535_), .ZN(new_n13941_));
  AOI21_X1   g12939(.A1(new_n13451_), .A2(new_n11898_), .B(new_n13445_), .ZN(new_n13942_));
  OAI21_X1   g12940(.A1(new_n13459_), .A2(new_n13460_), .B(new_n13432_), .ZN(new_n13943_));
  NOR2_X1    g12941(.A1(new_n13942_), .A2(new_n13943_), .ZN(new_n13944_));
  OAI21_X1   g12942(.A1(new_n13438_), .A2(new_n13443_), .B(new_n13454_), .ZN(new_n13945_));
  AOI21_X1   g12943(.A1(new_n13427_), .A2(new_n11927_), .B(new_n13461_), .ZN(new_n13946_));
  NOR2_X1    g12944(.A1(new_n13946_), .A2(new_n13945_), .ZN(new_n13947_));
  AOI21_X1   g12945(.A1(new_n13450_), .A2(new_n13456_), .B(new_n13434_), .ZN(new_n13948_));
  OAI22_X1   g12946(.A1(new_n13521_), .A2(new_n13948_), .B1(new_n13944_), .B2(new_n13947_), .ZN(new_n13949_));
  NAND2_X1   g12947(.A1(new_n13946_), .A2(new_n13945_), .ZN(new_n13950_));
  NAND2_X1   g12948(.A1(new_n13942_), .A2(new_n13943_), .ZN(new_n13951_));
  OAI21_X1   g12949(.A1(new_n13449_), .A2(new_n13464_), .B(new_n13463_), .ZN(new_n13952_));
  NAND4_X1   g12950(.A1(new_n13952_), .A2(new_n13951_), .A3(new_n13950_), .A4(new_n13448_), .ZN(new_n13953_));
  NAND2_X1   g12951(.A1(new_n13949_), .A2(new_n13953_), .ZN(new_n13954_));
  OAI21_X1   g12952(.A1(new_n13488_), .A2(new_n13481_), .B(new_n13492_), .ZN(new_n13955_));
  INV_X1     g12953(.I(new_n13475_), .ZN(new_n13956_));
  NAND2_X1   g12954(.A1(new_n13476_), .A2(new_n13478_), .ZN(new_n13957_));
  AOI21_X1   g12955(.A1(new_n13957_), .A2(new_n11989_), .B(new_n13956_), .ZN(new_n13958_));
  NAND2_X1   g12956(.A1(new_n13958_), .A2(new_n13955_), .ZN(new_n13959_));
  NAND2_X1   g12957(.A1(new_n13482_), .A2(new_n11969_), .ZN(new_n13960_));
  AOI22_X1   g12958(.A1(new_n13499_), .A2(new_n11957_), .B1(new_n13960_), .B2(new_n13491_), .ZN(new_n13961_));
  XOR2_X1    g12959(.A1(new_n13477_), .A2(new_n13472_), .Z(new_n13962_));
  OAI21_X1   g12960(.A1(new_n13962_), .A2(new_n13489_), .B(new_n13475_), .ZN(new_n13963_));
  NAND2_X1   g12961(.A1(new_n13963_), .A2(new_n13961_), .ZN(new_n13964_));
  OAI21_X1   g12962(.A1(new_n13508_), .A2(new_n13506_), .B(new_n13479_), .ZN(new_n13965_));
  AOI22_X1   g12963(.A1(new_n13964_), .A2(new_n13959_), .B1(new_n13494_), .B2(new_n13965_), .ZN(new_n13966_));
  NOR2_X1    g12964(.A1(new_n13963_), .A2(new_n13961_), .ZN(new_n13967_));
  NOR2_X1    g12965(.A1(new_n13958_), .A2(new_n13955_), .ZN(new_n13968_));
  INV_X1     g12966(.I(new_n13965_), .ZN(new_n13969_));
  NOR4_X1    g12967(.A1(new_n13969_), .A2(new_n13967_), .A3(new_n13531_), .A4(new_n13968_), .ZN(new_n13970_));
  NOR2_X1    g12968(.A1(new_n13970_), .A2(new_n13966_), .ZN(new_n13971_));
  NAND2_X1   g12969(.A1(new_n13954_), .A2(new_n13971_), .ZN(new_n13972_));
  AOI22_X1   g12970(.A1(new_n13448_), .A2(new_n13952_), .B1(new_n13950_), .B2(new_n13951_), .ZN(new_n13973_));
  NOR4_X1    g12971(.A1(new_n13948_), .A2(new_n13944_), .A3(new_n13947_), .A4(new_n13521_), .ZN(new_n13974_));
  NOR2_X1    g12972(.A1(new_n13973_), .A2(new_n13974_), .ZN(new_n13975_));
  OAI22_X1   g12973(.A1(new_n13969_), .A2(new_n13531_), .B1(new_n13967_), .B2(new_n13968_), .ZN(new_n13976_));
  NAND4_X1   g12974(.A1(new_n13964_), .A2(new_n13494_), .A3(new_n13959_), .A4(new_n13965_), .ZN(new_n13977_));
  NAND2_X1   g12975(.A1(new_n13976_), .A2(new_n13977_), .ZN(new_n13978_));
  NAND2_X1   g12976(.A1(new_n13975_), .A2(new_n13978_), .ZN(new_n13979_));
  AOI21_X1   g12977(.A1(new_n13972_), .A2(new_n13979_), .B(new_n13941_), .ZN(new_n13980_));
  OAI21_X1   g12978(.A1(new_n13468_), .A2(new_n13528_), .B(new_n13666_), .ZN(new_n13981_));
  NOR2_X1    g12979(.A1(new_n13975_), .A2(new_n13978_), .ZN(new_n13982_));
  NOR2_X1    g12980(.A1(new_n13954_), .A2(new_n13971_), .ZN(new_n13983_));
  NOR3_X1    g12981(.A1(new_n13982_), .A2(new_n13983_), .A3(new_n13981_), .ZN(new_n13984_));
  NOR2_X1    g12982(.A1(new_n13984_), .A2(new_n13980_), .ZN(new_n13985_));
  OAI21_X1   g12983(.A1(new_n13648_), .A2(new_n13637_), .B(new_n13657_), .ZN(new_n13986_));
  OAI21_X1   g12984(.A1(new_n13565_), .A2(new_n13550_), .B(new_n13557_), .ZN(new_n13987_));
  AOI21_X1   g12985(.A1(new_n13571_), .A2(new_n12119_), .B(new_n13544_), .ZN(new_n13988_));
  NAND2_X1   g12986(.A1(new_n13988_), .A2(new_n13987_), .ZN(new_n13989_));
  AOI21_X1   g12987(.A1(new_n13549_), .A2(new_n12089_), .B(new_n13566_), .ZN(new_n13990_));
  OAI21_X1   g12988(.A1(new_n13541_), .A2(new_n13542_), .B(new_n13574_), .ZN(new_n13991_));
  NAND2_X1   g12989(.A1(new_n13990_), .A2(new_n13991_), .ZN(new_n13992_));
  OAI21_X1   g12990(.A1(new_n13564_), .A2(new_n13568_), .B(new_n13546_), .ZN(new_n13993_));
  AOI22_X1   g12991(.A1(new_n13989_), .A2(new_n13992_), .B1(new_n13993_), .B2(new_n13641_), .ZN(new_n13994_));
  NOR2_X1    g12992(.A1(new_n13990_), .A2(new_n13991_), .ZN(new_n13995_));
  NOR2_X1    g12993(.A1(new_n13988_), .A2(new_n13987_), .ZN(new_n13996_));
  AOI21_X1   g12994(.A1(new_n13578_), .A2(new_n13642_), .B(new_n13576_), .ZN(new_n13997_));
  NOR4_X1    g12995(.A1(new_n13995_), .A2(new_n13997_), .A3(new_n13996_), .A4(new_n13560_), .ZN(new_n13998_));
  NOR2_X1    g12996(.A1(new_n13994_), .A2(new_n13998_), .ZN(new_n13999_));
  AOI21_X1   g12997(.A1(new_n13604_), .A2(new_n12023_), .B(new_n13609_), .ZN(new_n14000_));
  INV_X1     g12998(.I(new_n13587_), .ZN(new_n14001_));
  NOR2_X1    g12999(.A1(new_n13592_), .A2(new_n13590_), .ZN(new_n14002_));
  OAI21_X1   g13000(.A1(new_n14002_), .A2(new_n13583_), .B(new_n14001_), .ZN(new_n14003_));
  NOR2_X1    g13001(.A1(new_n14003_), .A2(new_n14000_), .ZN(new_n14004_));
  NOR2_X1    g13002(.A1(new_n13597_), .A2(new_n13602_), .ZN(new_n14005_));
  OAI22_X1   g13003(.A1(new_n13616_), .A2(new_n13605_), .B1(new_n14005_), .B2(new_n13608_), .ZN(new_n14006_));
  NAND2_X1   g13004(.A1(new_n13591_), .A2(new_n12067_), .ZN(new_n14007_));
  NAND2_X1   g13005(.A1(new_n13585_), .A2(new_n13589_), .ZN(new_n14008_));
  NAND2_X1   g13006(.A1(new_n14007_), .A2(new_n14008_), .ZN(new_n14009_));
  AOI21_X1   g13007(.A1(new_n14009_), .A2(new_n12055_), .B(new_n13587_), .ZN(new_n14010_));
  NOR2_X1    g13008(.A1(new_n14006_), .A2(new_n14010_), .ZN(new_n14011_));
  AOI21_X1   g13009(.A1(new_n13620_), .A2(new_n13622_), .B(new_n13593_), .ZN(new_n14012_));
  OAI22_X1   g13010(.A1(new_n14004_), .A2(new_n14011_), .B1(new_n13611_), .B2(new_n14012_), .ZN(new_n14013_));
  NAND2_X1   g13011(.A1(new_n14006_), .A2(new_n14010_), .ZN(new_n14014_));
  NAND2_X1   g13012(.A1(new_n14003_), .A2(new_n14000_), .ZN(new_n14015_));
  NAND2_X1   g13013(.A1(new_n13632_), .A2(new_n13594_), .ZN(new_n14016_));
  NAND4_X1   g13014(.A1(new_n14016_), .A2(new_n14014_), .A3(new_n14015_), .A4(new_n13631_), .ZN(new_n14017_));
  NAND2_X1   g13015(.A1(new_n14013_), .A2(new_n14017_), .ZN(new_n14018_));
  NOR2_X1    g13016(.A1(new_n13999_), .A2(new_n14018_), .ZN(new_n14019_));
  OAI22_X1   g13017(.A1(new_n13995_), .A2(new_n13996_), .B1(new_n13997_), .B2(new_n13560_), .ZN(new_n14020_));
  NAND4_X1   g13018(.A1(new_n13989_), .A2(new_n13993_), .A3(new_n13992_), .A4(new_n13641_), .ZN(new_n14021_));
  NAND2_X1   g13019(.A1(new_n14020_), .A2(new_n14021_), .ZN(new_n14022_));
  AOI22_X1   g13020(.A1(new_n14016_), .A2(new_n13631_), .B1(new_n14014_), .B2(new_n14015_), .ZN(new_n14023_));
  NOR4_X1    g13021(.A1(new_n13611_), .A2(new_n14011_), .A3(new_n14004_), .A4(new_n14012_), .ZN(new_n14024_));
  NOR2_X1    g13022(.A1(new_n14023_), .A2(new_n14024_), .ZN(new_n14025_));
  NOR2_X1    g13023(.A1(new_n14022_), .A2(new_n14025_), .ZN(new_n14026_));
  OAI21_X1   g13024(.A1(new_n14019_), .A2(new_n14026_), .B(new_n13986_), .ZN(new_n14027_));
  AOI21_X1   g13025(.A1(new_n13581_), .A2(new_n13658_), .B(new_n13625_), .ZN(new_n14028_));
  NAND2_X1   g13026(.A1(new_n14022_), .A2(new_n14025_), .ZN(new_n14029_));
  NAND2_X1   g13027(.A1(new_n13999_), .A2(new_n14018_), .ZN(new_n14030_));
  NAND3_X1   g13028(.A1(new_n14030_), .A2(new_n14029_), .A3(new_n14028_), .ZN(new_n14031_));
  NAND2_X1   g13029(.A1(new_n14027_), .A2(new_n14031_), .ZN(new_n14032_));
  NOR2_X1    g13030(.A1(new_n13985_), .A2(new_n14032_), .ZN(new_n14033_));
  OAI21_X1   g13031(.A1(new_n13983_), .A2(new_n13982_), .B(new_n13981_), .ZN(new_n14034_));
  NAND3_X1   g13032(.A1(new_n13972_), .A2(new_n13979_), .A3(new_n13941_), .ZN(new_n14035_));
  NAND2_X1   g13033(.A1(new_n14034_), .A2(new_n14035_), .ZN(new_n14036_));
  AOI21_X1   g13034(.A1(new_n14030_), .A2(new_n14029_), .B(new_n14028_), .ZN(new_n14037_));
  NOR3_X1    g13035(.A1(new_n14019_), .A2(new_n14026_), .A3(new_n13986_), .ZN(new_n14038_));
  NOR2_X1    g13036(.A1(new_n14037_), .A2(new_n14038_), .ZN(new_n14039_));
  NOR2_X1    g13037(.A1(new_n14036_), .A2(new_n14039_), .ZN(new_n14040_));
  OAI21_X1   g13038(.A1(new_n14040_), .A2(new_n14033_), .B(new_n13940_), .ZN(new_n14041_));
  AOI21_X1   g13039(.A1(new_n13652_), .A2(new_n13638_), .B(new_n13662_), .ZN(new_n14042_));
  AOI21_X1   g13040(.A1(new_n13537_), .A2(new_n13669_), .B(new_n14042_), .ZN(new_n14043_));
  NAND2_X1   g13041(.A1(new_n14036_), .A2(new_n14039_), .ZN(new_n14044_));
  NAND2_X1   g13042(.A1(new_n13985_), .A2(new_n14032_), .ZN(new_n14045_));
  NAND3_X1   g13043(.A1(new_n14044_), .A2(new_n14045_), .A3(new_n14043_), .ZN(new_n14046_));
  NAND2_X1   g13044(.A1(new_n14041_), .A2(new_n14046_), .ZN(new_n14047_));
  AOI22_X1   g13045(.A1(new_n13919_), .A2(new_n13891_), .B1(new_n13921_), .B2(new_n13900_), .ZN(new_n14048_));
  OAI21_X1   g13046(.A1(new_n13746_), .A2(new_n13756_), .B(new_n13769_), .ZN(new_n14049_));
  OAI21_X1   g13047(.A1(new_n13711_), .A2(new_n13772_), .B(new_n14049_), .ZN(new_n14050_));
  OAI21_X1   g13048(.A1(new_n13688_), .A2(new_n13693_), .B(new_n13705_), .ZN(new_n14051_));
  AOI21_X1   g13049(.A1(new_n13675_), .A2(new_n12377_), .B(new_n13904_), .ZN(new_n14052_));
  NAND2_X1   g13050(.A1(new_n14052_), .A2(new_n14051_), .ZN(new_n14053_));
  AOI21_X1   g13051(.A1(new_n13702_), .A2(new_n12345_), .B(new_n13695_), .ZN(new_n14054_));
  OAI21_X1   g13052(.A1(new_n13903_), .A2(new_n13699_), .B(new_n13681_), .ZN(new_n14055_));
  NAND2_X1   g13053(.A1(new_n14054_), .A2(new_n14055_), .ZN(new_n14056_));
  OAI21_X1   g13054(.A1(new_n13910_), .A2(new_n13911_), .B(new_n13906_), .ZN(new_n14057_));
  AOI22_X1   g13055(.A1(new_n14053_), .A2(new_n14056_), .B1(new_n14057_), .B2(new_n13698_), .ZN(new_n14058_));
  NOR2_X1    g13056(.A1(new_n14054_), .A2(new_n14055_), .ZN(new_n14059_));
  NOR2_X1    g13057(.A1(new_n14052_), .A2(new_n14051_), .ZN(new_n14060_));
  AOI21_X1   g13058(.A1(new_n13701_), .A2(new_n13707_), .B(new_n13683_), .ZN(new_n14061_));
  NOR4_X1    g13059(.A1(new_n14059_), .A2(new_n14061_), .A3(new_n14060_), .A4(new_n13909_), .ZN(new_n14062_));
  NOR2_X1    g13060(.A1(new_n14058_), .A2(new_n14062_), .ZN(new_n14063_));
  NAND2_X1   g13061(.A1(new_n13725_), .A2(new_n12292_), .ZN(new_n14064_));
  AOI22_X1   g13062(.A1(new_n13743_), .A2(new_n12280_), .B1(new_n14064_), .B2(new_n13734_), .ZN(new_n14065_));
  OAI21_X1   g13063(.A1(new_n13750_), .A2(new_n13712_), .B(new_n13747_), .ZN(new_n14066_));
  NOR2_X1    g13064(.A1(new_n14065_), .A2(new_n14066_), .ZN(new_n14067_));
  OAI21_X1   g13065(.A1(new_n13731_), .A2(new_n13738_), .B(new_n13735_), .ZN(new_n14068_));
  AOI21_X1   g13066(.A1(new_n13722_), .A2(new_n12312_), .B(new_n13716_), .ZN(new_n14069_));
  NOR2_X1    g13067(.A1(new_n14068_), .A2(new_n14069_), .ZN(new_n14070_));
  NOR2_X1    g13068(.A1(new_n13762_), .A2(new_n13723_), .ZN(new_n14071_));
  OAI22_X1   g13069(.A1(new_n14071_), .A2(new_n13761_), .B1(new_n14067_), .B2(new_n14070_), .ZN(new_n14072_));
  NAND2_X1   g13070(.A1(new_n14068_), .A2(new_n14069_), .ZN(new_n14073_));
  NAND2_X1   g13071(.A1(new_n14065_), .A2(new_n14066_), .ZN(new_n14074_));
  NAND2_X1   g13072(.A1(new_n13745_), .A2(new_n13751_), .ZN(new_n14075_));
  NAND4_X1   g13073(.A1(new_n14075_), .A2(new_n14073_), .A3(new_n14074_), .A4(new_n13737_), .ZN(new_n14076_));
  NAND2_X1   g13074(.A1(new_n14076_), .A2(new_n14072_), .ZN(new_n14077_));
  NOR2_X1    g13075(.A1(new_n14063_), .A2(new_n14077_), .ZN(new_n14078_));
  OAI22_X1   g13076(.A1(new_n14059_), .A2(new_n14060_), .B1(new_n14061_), .B2(new_n13909_), .ZN(new_n14079_));
  NAND4_X1   g13077(.A1(new_n14053_), .A2(new_n14057_), .A3(new_n14056_), .A4(new_n13698_), .ZN(new_n14080_));
  NAND2_X1   g13078(.A1(new_n14079_), .A2(new_n14080_), .ZN(new_n14081_));
  AOI22_X1   g13079(.A1(new_n14075_), .A2(new_n13737_), .B1(new_n14073_), .B2(new_n14074_), .ZN(new_n14082_));
  NOR4_X1    g13080(.A1(new_n14071_), .A2(new_n14067_), .A3(new_n14070_), .A4(new_n13761_), .ZN(new_n14083_));
  NOR2_X1    g13081(.A1(new_n14082_), .A2(new_n14083_), .ZN(new_n14084_));
  NOR2_X1    g13082(.A1(new_n14084_), .A2(new_n14081_), .ZN(new_n14085_));
  OAI21_X1   g13083(.A1(new_n14085_), .A2(new_n14078_), .B(new_n14050_), .ZN(new_n14086_));
  NAND3_X1   g13084(.A1(new_n13763_), .A2(new_n13766_), .A3(new_n13757_), .ZN(new_n14087_));
  AOI21_X1   g13085(.A1(new_n13917_), .A2(new_n14087_), .B(new_n13773_), .ZN(new_n14088_));
  NAND2_X1   g13086(.A1(new_n14084_), .A2(new_n14081_), .ZN(new_n14089_));
  NAND2_X1   g13087(.A1(new_n14063_), .A2(new_n14077_), .ZN(new_n14090_));
  NAND3_X1   g13088(.A1(new_n14089_), .A2(new_n14090_), .A3(new_n14088_), .ZN(new_n14091_));
  NAND2_X1   g13089(.A1(new_n14086_), .A2(new_n14091_), .ZN(new_n14092_));
  AOI21_X1   g13090(.A1(new_n13821_), .A2(new_n13893_), .B(new_n13865_), .ZN(new_n14093_));
  AOI21_X1   g13091(.A1(new_n13795_), .A2(new_n12216_), .B(new_n13801_), .ZN(new_n14094_));
  XOR2_X1    g13092(.A1(new_n13783_), .A2(new_n13777_), .Z(new_n14095_));
  OAI21_X1   g13093(.A1(new_n14095_), .A2(new_n13797_), .B(new_n13781_), .ZN(new_n14096_));
  NOR2_X1    g13094(.A1(new_n14096_), .A2(new_n14094_), .ZN(new_n14097_));
  OAI21_X1   g13095(.A1(new_n13808_), .A2(new_n13796_), .B(new_n13814_), .ZN(new_n14098_));
  INV_X1     g13096(.I(new_n13781_), .ZN(new_n14099_));
  NAND2_X1   g13097(.A1(new_n13782_), .A2(new_n13784_), .ZN(new_n14100_));
  AOI21_X1   g13098(.A1(new_n14100_), .A2(new_n12249_), .B(new_n14099_), .ZN(new_n14101_));
  NOR2_X1    g13099(.A1(new_n14101_), .A2(new_n14098_), .ZN(new_n14102_));
  AOI21_X1   g13100(.A1(new_n13818_), .A2(new_n13816_), .B(new_n13812_), .ZN(new_n14103_));
  OAI22_X1   g13101(.A1(new_n14103_), .A2(new_n13803_), .B1(new_n14097_), .B2(new_n14102_), .ZN(new_n14104_));
  NAND2_X1   g13102(.A1(new_n14101_), .A2(new_n14098_), .ZN(new_n14105_));
  NAND2_X1   g13103(.A1(new_n14096_), .A2(new_n14094_), .ZN(new_n14106_));
  OAI21_X1   g13104(.A1(new_n13809_), .A2(new_n13805_), .B(new_n13785_), .ZN(new_n14107_));
  NAND4_X1   g13105(.A1(new_n14105_), .A2(new_n14106_), .A3(new_n14107_), .A4(new_n13880_), .ZN(new_n14108_));
  NAND2_X1   g13106(.A1(new_n14104_), .A2(new_n14108_), .ZN(new_n14109_));
  NOR2_X1    g13107(.A1(new_n13837_), .A2(new_n13842_), .ZN(new_n14110_));
  OAI22_X1   g13108(.A1(new_n13856_), .A2(new_n13845_), .B1(new_n14110_), .B2(new_n13848_), .ZN(new_n14111_));
  NAND2_X1   g13109(.A1(new_n13831_), .A2(new_n12195_), .ZN(new_n14112_));
  NAND2_X1   g13110(.A1(new_n13825_), .A2(new_n13829_), .ZN(new_n14113_));
  NAND2_X1   g13111(.A1(new_n14112_), .A2(new_n14113_), .ZN(new_n14114_));
  AOI21_X1   g13112(.A1(new_n14114_), .A2(new_n12183_), .B(new_n13827_), .ZN(new_n14115_));
  NAND2_X1   g13113(.A1(new_n14111_), .A2(new_n14115_), .ZN(new_n14116_));
  AOI21_X1   g13114(.A1(new_n13844_), .A2(new_n12151_), .B(new_n13849_), .ZN(new_n14117_));
  INV_X1     g13115(.I(new_n13827_), .ZN(new_n14118_));
  NOR2_X1    g13116(.A1(new_n13832_), .A2(new_n13830_), .ZN(new_n14119_));
  OAI21_X1   g13117(.A1(new_n14119_), .A2(new_n13823_), .B(new_n14118_), .ZN(new_n14120_));
  NAND2_X1   g13118(.A1(new_n14120_), .A2(new_n14117_), .ZN(new_n14121_));
  NAND2_X1   g13119(.A1(new_n13872_), .A2(new_n13834_), .ZN(new_n14122_));
  AOI22_X1   g13120(.A1(new_n14122_), .A2(new_n13871_), .B1(new_n14116_), .B2(new_n14121_), .ZN(new_n14123_));
  NOR2_X1    g13121(.A1(new_n14120_), .A2(new_n14117_), .ZN(new_n14124_));
  NOR2_X1    g13122(.A1(new_n14111_), .A2(new_n14115_), .ZN(new_n14125_));
  AOI21_X1   g13123(.A1(new_n13860_), .A2(new_n13862_), .B(new_n13833_), .ZN(new_n14126_));
  NOR4_X1    g13124(.A1(new_n13851_), .A2(new_n14125_), .A3(new_n14124_), .A4(new_n14126_), .ZN(new_n14127_));
  NOR2_X1    g13125(.A1(new_n14123_), .A2(new_n14127_), .ZN(new_n14128_));
  NAND2_X1   g13126(.A1(new_n14109_), .A2(new_n14128_), .ZN(new_n14129_));
  AOI22_X1   g13127(.A1(new_n14105_), .A2(new_n14106_), .B1(new_n14107_), .B2(new_n13880_), .ZN(new_n14130_));
  NOR4_X1    g13128(.A1(new_n14103_), .A2(new_n14097_), .A3(new_n14102_), .A4(new_n13803_), .ZN(new_n14131_));
  NOR2_X1    g13129(.A1(new_n14131_), .A2(new_n14130_), .ZN(new_n14132_));
  OAI22_X1   g13130(.A1(new_n14124_), .A2(new_n14125_), .B1(new_n13851_), .B2(new_n14126_), .ZN(new_n14133_));
  NAND4_X1   g13131(.A1(new_n14122_), .A2(new_n14116_), .A3(new_n14121_), .A4(new_n13871_), .ZN(new_n14134_));
  NAND2_X1   g13132(.A1(new_n14133_), .A2(new_n14134_), .ZN(new_n14135_));
  NAND2_X1   g13133(.A1(new_n14132_), .A2(new_n14135_), .ZN(new_n14136_));
  AOI21_X1   g13134(.A1(new_n14129_), .A2(new_n14136_), .B(new_n14093_), .ZN(new_n14137_));
  OAI21_X1   g13135(.A1(new_n13886_), .A2(new_n13877_), .B(new_n13892_), .ZN(new_n14138_));
  NOR2_X1    g13136(.A1(new_n14132_), .A2(new_n14135_), .ZN(new_n14139_));
  NOR2_X1    g13137(.A1(new_n14109_), .A2(new_n14128_), .ZN(new_n14140_));
  NOR3_X1    g13138(.A1(new_n14140_), .A2(new_n14139_), .A3(new_n14138_), .ZN(new_n14141_));
  NOR2_X1    g13139(.A1(new_n14137_), .A2(new_n14141_), .ZN(new_n14142_));
  NAND2_X1   g13140(.A1(new_n14092_), .A2(new_n14142_), .ZN(new_n14143_));
  AOI21_X1   g13141(.A1(new_n14089_), .A2(new_n14090_), .B(new_n14088_), .ZN(new_n14144_));
  NOR3_X1    g13142(.A1(new_n14085_), .A2(new_n14078_), .A3(new_n14050_), .ZN(new_n14145_));
  NOR2_X1    g13143(.A1(new_n14144_), .A2(new_n14145_), .ZN(new_n14146_));
  OAI21_X1   g13144(.A1(new_n14140_), .A2(new_n14139_), .B(new_n14138_), .ZN(new_n14147_));
  NAND3_X1   g13145(.A1(new_n14129_), .A2(new_n14136_), .A3(new_n14093_), .ZN(new_n14148_));
  NAND2_X1   g13146(.A1(new_n14147_), .A2(new_n14148_), .ZN(new_n14149_));
  NAND2_X1   g13147(.A1(new_n14146_), .A2(new_n14149_), .ZN(new_n14150_));
  AOI21_X1   g13148(.A1(new_n14150_), .A2(new_n14143_), .B(new_n14048_), .ZN(new_n14151_));
  NOR3_X1    g13149(.A1(new_n13894_), .A2(new_n13897_), .A3(new_n13900_), .ZN(new_n14152_));
  OAI21_X1   g13150(.A1(new_n13775_), .A2(new_n14152_), .B(new_n13901_), .ZN(new_n14153_));
  NOR2_X1    g13151(.A1(new_n14146_), .A2(new_n14149_), .ZN(new_n14154_));
  NOR2_X1    g13152(.A1(new_n14092_), .A2(new_n14142_), .ZN(new_n14155_));
  NOR3_X1    g13153(.A1(new_n14154_), .A2(new_n14155_), .A3(new_n14153_), .ZN(new_n14156_));
  NOR2_X1    g13154(.A1(new_n14151_), .A2(new_n14156_), .ZN(new_n14157_));
  NAND2_X1   g13155(.A1(new_n14157_), .A2(new_n14047_), .ZN(new_n14158_));
  AOI21_X1   g13156(.A1(new_n14044_), .A2(new_n14045_), .B(new_n14043_), .ZN(new_n14159_));
  NOR3_X1    g13157(.A1(new_n14040_), .A2(new_n14033_), .A3(new_n13940_), .ZN(new_n14160_));
  NOR2_X1    g13158(.A1(new_n14159_), .A2(new_n14160_), .ZN(new_n14161_));
  OAI21_X1   g13159(.A1(new_n14154_), .A2(new_n14155_), .B(new_n14153_), .ZN(new_n14162_));
  NAND3_X1   g13160(.A1(new_n14150_), .A2(new_n14143_), .A3(new_n14048_), .ZN(new_n14163_));
  NAND2_X1   g13161(.A1(new_n14162_), .A2(new_n14163_), .ZN(new_n14164_));
  NAND2_X1   g13162(.A1(new_n14161_), .A2(new_n14164_), .ZN(new_n14165_));
  AOI21_X1   g13163(.A1(new_n14158_), .A2(new_n14165_), .B(new_n13938_), .ZN(new_n14166_));
  OAI22_X1   g13164(.A1(new_n13930_), .A2(new_n13672_), .B1(new_n13927_), .B2(new_n13924_), .ZN(new_n14167_));
  NOR2_X1    g13165(.A1(new_n14161_), .A2(new_n14164_), .ZN(new_n14168_));
  NOR2_X1    g13166(.A1(new_n14157_), .A2(new_n14047_), .ZN(new_n14169_));
  NOR3_X1    g13167(.A1(new_n14169_), .A2(new_n14168_), .A3(new_n14167_), .ZN(new_n14170_));
  NOR2_X1    g13168(.A1(new_n14166_), .A2(new_n14170_), .ZN(new_n14171_));
  NOR3_X1    g13169(.A1(new_n13412_), .A2(new_n13416_), .A3(new_n13410_), .ZN(new_n14172_));
  OAI21_X1   g13170(.A1(new_n13158_), .A2(new_n14172_), .B(new_n13420_), .ZN(new_n14173_));
  AOI22_X1   g13171(.A1(new_n13029_), .A2(new_n13149_), .B1(new_n13140_), .B2(new_n13137_), .ZN(new_n14174_));
  OAI21_X1   g13172(.A1(new_n12952_), .A2(new_n13025_), .B(new_n13146_), .ZN(new_n14175_));
  OAI21_X1   g13173(.A1(new_n12929_), .A2(new_n12934_), .B(new_n12946_), .ZN(new_n14176_));
  AOI21_X1   g13174(.A1(new_n12917_), .A2(new_n12897_), .B(new_n13001_), .ZN(new_n14177_));
  NAND2_X1   g13175(.A1(new_n14177_), .A2(new_n14176_), .ZN(new_n14178_));
  AOI21_X1   g13176(.A1(new_n12943_), .A2(new_n12864_), .B(new_n12936_), .ZN(new_n14179_));
  OAI21_X1   g13177(.A1(new_n13000_), .A2(new_n12940_), .B(new_n12922_), .ZN(new_n14180_));
  NAND2_X1   g13178(.A1(new_n14179_), .A2(new_n14180_), .ZN(new_n14181_));
  OAI21_X1   g13179(.A1(new_n13007_), .A2(new_n13008_), .B(new_n13003_), .ZN(new_n14182_));
  AOI22_X1   g13180(.A1(new_n14178_), .A2(new_n14181_), .B1(new_n14182_), .B2(new_n12939_), .ZN(new_n14183_));
  NOR2_X1    g13181(.A1(new_n14179_), .A2(new_n14180_), .ZN(new_n14184_));
  NOR2_X1    g13182(.A1(new_n14177_), .A2(new_n14176_), .ZN(new_n14185_));
  AOI21_X1   g13183(.A1(new_n12942_), .A2(new_n12948_), .B(new_n12924_), .ZN(new_n14186_));
  NOR4_X1    g13184(.A1(new_n14184_), .A2(new_n14186_), .A3(new_n14185_), .A4(new_n13006_), .ZN(new_n14187_));
  NOR2_X1    g13185(.A1(new_n14183_), .A2(new_n14187_), .ZN(new_n14188_));
  NAND2_X1   g13186(.A1(new_n12966_), .A2(new_n12811_), .ZN(new_n14189_));
  AOI22_X1   g13187(.A1(new_n12970_), .A2(new_n12799_), .B1(new_n14189_), .B2(new_n12975_), .ZN(new_n14190_));
  NOR2_X1    g13188(.A1(new_n12986_), .A2(new_n12985_), .ZN(new_n14191_));
  OAI21_X1   g13189(.A1(new_n14191_), .A2(new_n12972_), .B(new_n12959_), .ZN(new_n14192_));
  NOR2_X1    g13190(.A1(new_n14190_), .A2(new_n14192_), .ZN(new_n14193_));
  OAI21_X1   g13191(.A1(new_n13017_), .A2(new_n12971_), .B(new_n12976_), .ZN(new_n14194_));
  NAND2_X1   g13192(.A1(new_n12960_), .A2(new_n12962_), .ZN(new_n14195_));
  AOI21_X1   g13193(.A1(new_n14195_), .A2(new_n12831_), .B(new_n12984_), .ZN(new_n14196_));
  NOR2_X1    g13194(.A1(new_n14194_), .A2(new_n14196_), .ZN(new_n14197_));
  AOI21_X1   g13195(.A1(new_n12990_), .A2(new_n12988_), .B(new_n12987_), .ZN(new_n14198_));
  OAI22_X1   g13196(.A1(new_n14193_), .A2(new_n14197_), .B1(new_n14198_), .B2(new_n12979_), .ZN(new_n14199_));
  NAND2_X1   g13197(.A1(new_n14194_), .A2(new_n14196_), .ZN(new_n14200_));
  NAND2_X1   g13198(.A1(new_n14190_), .A2(new_n14192_), .ZN(new_n14201_));
  OAI21_X1   g13199(.A1(new_n12980_), .A2(new_n12981_), .B(new_n12963_), .ZN(new_n14202_));
  NAND4_X1   g13200(.A1(new_n13019_), .A2(new_n14201_), .A3(new_n14200_), .A4(new_n14202_), .ZN(new_n14203_));
  NAND2_X1   g13201(.A1(new_n14199_), .A2(new_n14203_), .ZN(new_n14204_));
  NOR2_X1    g13202(.A1(new_n14188_), .A2(new_n14204_), .ZN(new_n14205_));
  OAI22_X1   g13203(.A1(new_n14184_), .A2(new_n14185_), .B1(new_n14186_), .B2(new_n13006_), .ZN(new_n14206_));
  NAND4_X1   g13204(.A1(new_n14178_), .A2(new_n14182_), .A3(new_n14181_), .A4(new_n12939_), .ZN(new_n14207_));
  NAND2_X1   g13205(.A1(new_n14206_), .A2(new_n14207_), .ZN(new_n14208_));
  AOI22_X1   g13206(.A1(new_n13019_), .A2(new_n14202_), .B1(new_n14201_), .B2(new_n14200_), .ZN(new_n14209_));
  NOR4_X1    g13207(.A1(new_n14193_), .A2(new_n14197_), .A3(new_n14198_), .A4(new_n12979_), .ZN(new_n14210_));
  NOR2_X1    g13208(.A1(new_n14209_), .A2(new_n14210_), .ZN(new_n14211_));
  NOR2_X1    g13209(.A1(new_n14208_), .A2(new_n14211_), .ZN(new_n14212_));
  OAI21_X1   g13210(.A1(new_n14205_), .A2(new_n14212_), .B(new_n14175_), .ZN(new_n14213_));
  AOI21_X1   g13211(.A1(new_n13014_), .A2(new_n13145_), .B(new_n13027_), .ZN(new_n14214_));
  NAND2_X1   g13212(.A1(new_n14208_), .A2(new_n14211_), .ZN(new_n14215_));
  NAND2_X1   g13213(.A1(new_n14188_), .A2(new_n14204_), .ZN(new_n14216_));
  NAND3_X1   g13214(.A1(new_n14216_), .A2(new_n14215_), .A3(new_n14214_), .ZN(new_n14217_));
  NAND2_X1   g13215(.A1(new_n14213_), .A2(new_n14217_), .ZN(new_n14218_));
  AOI21_X1   g13216(.A1(new_n13068_), .A2(new_n13151_), .B(new_n13111_), .ZN(new_n14219_));
  NAND2_X1   g13217(.A1(new_n13047_), .A2(new_n12747_), .ZN(new_n14220_));
  AOI22_X1   g13218(.A1(new_n13063_), .A2(new_n12735_), .B1(new_n14220_), .B2(new_n13045_), .ZN(new_n14221_));
  XNOR2_X1   g13219(.A1(new_n12758_), .A2(new_n12767_), .ZN(new_n14222_));
  XOR2_X1    g13220(.A1(new_n13037_), .A2(new_n13031_), .Z(new_n14223_));
  OAI21_X1   g13221(.A1(new_n14223_), .A2(new_n14222_), .B(new_n13035_), .ZN(new_n14224_));
  NOR2_X1    g13222(.A1(new_n14224_), .A2(new_n14221_), .ZN(new_n14225_));
  INV_X1     g13223(.I(new_n12735_), .ZN(new_n14226_));
  OAI21_X1   g13224(.A1(new_n13050_), .A2(new_n14226_), .B(new_n13046_), .ZN(new_n14227_));
  INV_X1     g13225(.I(new_n13035_), .ZN(new_n14228_));
  NAND2_X1   g13226(.A1(new_n13036_), .A2(new_n13038_), .ZN(new_n14229_));
  AOI21_X1   g13227(.A1(new_n14229_), .A2(new_n12768_), .B(new_n14228_), .ZN(new_n14230_));
  NOR2_X1    g13228(.A1(new_n14230_), .A2(new_n14227_), .ZN(new_n14231_));
  OAI21_X1   g13229(.A1(new_n13059_), .A2(new_n13056_), .B(new_n13039_), .ZN(new_n14232_));
  INV_X1     g13230(.I(new_n14232_), .ZN(new_n14233_));
  OAI22_X1   g13231(.A1(new_n14233_), .A2(new_n13054_), .B1(new_n14225_), .B2(new_n14231_), .ZN(new_n14234_));
  NAND2_X1   g13232(.A1(new_n14230_), .A2(new_n14227_), .ZN(new_n14235_));
  NAND2_X1   g13233(.A1(new_n14224_), .A2(new_n14221_), .ZN(new_n14236_));
  NAND4_X1   g13234(.A1(new_n14236_), .A2(new_n14235_), .A3(new_n13125_), .A4(new_n14232_), .ZN(new_n14237_));
  NAND2_X1   g13235(.A1(new_n14234_), .A2(new_n14237_), .ZN(new_n14238_));
  NOR2_X1    g13236(.A1(new_n13084_), .A2(new_n13089_), .ZN(new_n14239_));
  OAI22_X1   g13237(.A1(new_n13102_), .A2(new_n13092_), .B1(new_n14239_), .B2(new_n13095_), .ZN(new_n14240_));
  NAND2_X1   g13238(.A1(new_n13078_), .A2(new_n12714_), .ZN(new_n14241_));
  NAND2_X1   g13239(.A1(new_n13072_), .A2(new_n13076_), .ZN(new_n14242_));
  NAND2_X1   g13240(.A1(new_n14241_), .A2(new_n14242_), .ZN(new_n14243_));
  AOI21_X1   g13241(.A1(new_n14243_), .A2(new_n12702_), .B(new_n13074_), .ZN(new_n14244_));
  NAND2_X1   g13242(.A1(new_n14240_), .A2(new_n14244_), .ZN(new_n14245_));
  AOI21_X1   g13243(.A1(new_n13091_), .A2(new_n12670_), .B(new_n13096_), .ZN(new_n14246_));
  INV_X1     g13244(.I(new_n13074_), .ZN(new_n14247_));
  NOR2_X1    g13245(.A1(new_n13079_), .A2(new_n13077_), .ZN(new_n14248_));
  OAI21_X1   g13246(.A1(new_n14248_), .A2(new_n13070_), .B(new_n14247_), .ZN(new_n14249_));
  NAND2_X1   g13247(.A1(new_n14249_), .A2(new_n14246_), .ZN(new_n14250_));
  NAND2_X1   g13248(.A1(new_n13117_), .A2(new_n13081_), .ZN(new_n14251_));
  AOI22_X1   g13249(.A1(new_n14251_), .A2(new_n13116_), .B1(new_n14245_), .B2(new_n14250_), .ZN(new_n14252_));
  NOR2_X1    g13250(.A1(new_n14249_), .A2(new_n14246_), .ZN(new_n14253_));
  NOR2_X1    g13251(.A1(new_n14240_), .A2(new_n14244_), .ZN(new_n14254_));
  AOI21_X1   g13252(.A1(new_n13106_), .A2(new_n13108_), .B(new_n13080_), .ZN(new_n14255_));
  NOR4_X1    g13253(.A1(new_n13098_), .A2(new_n14254_), .A3(new_n14253_), .A4(new_n14255_), .ZN(new_n14256_));
  NOR2_X1    g13254(.A1(new_n14252_), .A2(new_n14256_), .ZN(new_n14257_));
  NAND2_X1   g13255(.A1(new_n14238_), .A2(new_n14257_), .ZN(new_n14258_));
  AOI22_X1   g13256(.A1(new_n14236_), .A2(new_n14235_), .B1(new_n13125_), .B2(new_n14232_), .ZN(new_n14259_));
  NOR4_X1    g13257(.A1(new_n14233_), .A2(new_n14225_), .A3(new_n14231_), .A4(new_n13054_), .ZN(new_n14260_));
  NOR2_X1    g13258(.A1(new_n14260_), .A2(new_n14259_), .ZN(new_n14261_));
  OAI22_X1   g13259(.A1(new_n14253_), .A2(new_n14254_), .B1(new_n13098_), .B2(new_n14255_), .ZN(new_n14262_));
  NAND4_X1   g13260(.A1(new_n13116_), .A2(new_n14251_), .A3(new_n14245_), .A4(new_n14250_), .ZN(new_n14263_));
  NAND2_X1   g13261(.A1(new_n14263_), .A2(new_n14262_), .ZN(new_n14264_));
  NAND2_X1   g13262(.A1(new_n14261_), .A2(new_n14264_), .ZN(new_n14265_));
  AOI21_X1   g13263(.A1(new_n14258_), .A2(new_n14265_), .B(new_n14219_), .ZN(new_n14266_));
  OAI21_X1   g13264(.A1(new_n13131_), .A2(new_n13122_), .B(new_n13150_), .ZN(new_n14267_));
  NOR2_X1    g13265(.A1(new_n14261_), .A2(new_n14264_), .ZN(new_n14268_));
  NOR2_X1    g13266(.A1(new_n14238_), .A2(new_n14257_), .ZN(new_n14269_));
  NOR3_X1    g13267(.A1(new_n14269_), .A2(new_n14268_), .A3(new_n14267_), .ZN(new_n14270_));
  NOR2_X1    g13268(.A1(new_n14266_), .A2(new_n14270_), .ZN(new_n14271_));
  NAND2_X1   g13269(.A1(new_n14271_), .A2(new_n14218_), .ZN(new_n14272_));
  AOI21_X1   g13270(.A1(new_n14216_), .A2(new_n14215_), .B(new_n14214_), .ZN(new_n14273_));
  NOR3_X1    g13271(.A1(new_n14175_), .A2(new_n14205_), .A3(new_n14212_), .ZN(new_n14274_));
  NOR2_X1    g13272(.A1(new_n14274_), .A2(new_n14273_), .ZN(new_n14275_));
  OAI21_X1   g13273(.A1(new_n14269_), .A2(new_n14268_), .B(new_n14267_), .ZN(new_n14276_));
  NAND3_X1   g13274(.A1(new_n14258_), .A2(new_n14265_), .A3(new_n14219_), .ZN(new_n14277_));
  NAND2_X1   g13275(.A1(new_n14276_), .A2(new_n14277_), .ZN(new_n14278_));
  NAND2_X1   g13276(.A1(new_n14275_), .A2(new_n14278_), .ZN(new_n14279_));
  AOI21_X1   g13277(.A1(new_n14272_), .A2(new_n14279_), .B(new_n14174_), .ZN(new_n14280_));
  NOR3_X1    g13278(.A1(new_n13152_), .A2(new_n13155_), .A3(new_n13137_), .ZN(new_n14281_));
  OAI21_X1   g13279(.A1(new_n13148_), .A2(new_n14281_), .B(new_n13156_), .ZN(new_n14282_));
  NOR2_X1    g13280(.A1(new_n14275_), .A2(new_n14278_), .ZN(new_n14283_));
  NOR2_X1    g13281(.A1(new_n14271_), .A2(new_n14218_), .ZN(new_n14284_));
  NOR3_X1    g13282(.A1(new_n14284_), .A2(new_n14283_), .A3(new_n14282_), .ZN(new_n14285_));
  NOR2_X1    g13283(.A1(new_n14280_), .A2(new_n14285_), .ZN(new_n14286_));
  NAND2_X1   g13284(.A1(new_n13394_), .A2(new_n13273_), .ZN(new_n14287_));
  NAND2_X1   g13285(.A1(new_n14287_), .A2(new_n13402_), .ZN(new_n14288_));
  NAND3_X1   g13286(.A1(new_n13246_), .A2(new_n13249_), .A3(new_n13240_), .ZN(new_n14289_));
  AOI21_X1   g13287(.A1(new_n13269_), .A2(new_n14289_), .B(new_n13271_), .ZN(new_n14290_));
  AOI21_X1   g13288(.A1(new_n13259_), .A2(new_n12603_), .B(new_n13186_), .ZN(new_n14291_));
  XOR2_X1    g13289(.A1(new_n13162_), .A2(new_n13168_), .Z(new_n14292_));
  OAI21_X1   g13290(.A1(new_n14292_), .A2(new_n13160_), .B(new_n13255_), .ZN(new_n14293_));
  NOR2_X1    g13291(.A1(new_n14293_), .A2(new_n14291_), .ZN(new_n14294_));
  NOR2_X1    g13292(.A1(new_n13177_), .A2(new_n13175_), .ZN(new_n14295_));
  OAI22_X1   g13293(.A1(new_n13179_), .A2(new_n13184_), .B1(new_n14295_), .B2(new_n13185_), .ZN(new_n14296_));
  AOI21_X1   g13294(.A1(new_n13170_), .A2(new_n12635_), .B(new_n13164_), .ZN(new_n14297_));
  NOR2_X1    g13295(.A1(new_n14296_), .A2(new_n14297_), .ZN(new_n14298_));
  AOI21_X1   g13296(.A1(new_n13191_), .A2(new_n13192_), .B(new_n13171_), .ZN(new_n14299_));
  OAI22_X1   g13297(.A1(new_n14299_), .A2(new_n13261_), .B1(new_n14294_), .B2(new_n14298_), .ZN(new_n14300_));
  NAND2_X1   g13298(.A1(new_n14296_), .A2(new_n14297_), .ZN(new_n14301_));
  NAND2_X1   g13299(.A1(new_n14293_), .A2(new_n14291_), .ZN(new_n14302_));
  NAND2_X1   g13300(.A1(new_n13193_), .A2(new_n13256_), .ZN(new_n14303_));
  NAND4_X1   g13301(.A1(new_n14303_), .A2(new_n14302_), .A3(new_n14301_), .A4(new_n13189_), .ZN(new_n14304_));
  NAND2_X1   g13302(.A1(new_n14300_), .A2(new_n14304_), .ZN(new_n14305_));
  OAI21_X1   g13303(.A1(new_n13216_), .A2(new_n13208_), .B(new_n13220_), .ZN(new_n14306_));
  NAND2_X1   g13304(.A1(new_n13232_), .A2(new_n13233_), .ZN(new_n14307_));
  AOI21_X1   g13305(.A1(new_n14307_), .A2(new_n12570_), .B(new_n13201_), .ZN(new_n14308_));
  NAND2_X1   g13306(.A1(new_n14306_), .A2(new_n14308_), .ZN(new_n14309_));
  AOI21_X1   g13307(.A1(new_n13210_), .A2(new_n12550_), .B(new_n13218_), .ZN(new_n14310_));
  AOI21_X1   g13308(.A1(new_n13227_), .A2(new_n12538_), .B(new_n14310_), .ZN(new_n14311_));
  NOR2_X1    g13309(.A1(new_n13206_), .A2(new_n13204_), .ZN(new_n14312_));
  OAI21_X1   g13310(.A1(new_n14312_), .A2(new_n13197_), .B(new_n13231_), .ZN(new_n14313_));
  NAND2_X1   g13311(.A1(new_n14313_), .A2(new_n14311_), .ZN(new_n14314_));
  OAI21_X1   g13312(.A1(new_n13237_), .A2(new_n13235_), .B(new_n13234_), .ZN(new_n14315_));
  AOI22_X1   g13313(.A1(new_n14315_), .A2(new_n13222_), .B1(new_n14309_), .B2(new_n14314_), .ZN(new_n14316_));
  NOR2_X1    g13314(.A1(new_n14313_), .A2(new_n14311_), .ZN(new_n14317_));
  NOR2_X1    g13315(.A1(new_n14306_), .A2(new_n14308_), .ZN(new_n14318_));
  AOI21_X1   g13316(.A1(new_n13228_), .A2(new_n13224_), .B(new_n13207_), .ZN(new_n14319_));
  NOR4_X1    g13317(.A1(new_n14317_), .A2(new_n14318_), .A3(new_n14319_), .A4(new_n13244_), .ZN(new_n14320_));
  NOR2_X1    g13318(.A1(new_n14316_), .A2(new_n14320_), .ZN(new_n14321_));
  NAND2_X1   g13319(.A1(new_n14305_), .A2(new_n14321_), .ZN(new_n14322_));
  AOI22_X1   g13320(.A1(new_n14303_), .A2(new_n13189_), .B1(new_n14302_), .B2(new_n14301_), .ZN(new_n14323_));
  NOR4_X1    g13321(.A1(new_n14299_), .A2(new_n14294_), .A3(new_n14298_), .A4(new_n13261_), .ZN(new_n14324_));
  NOR2_X1    g13322(.A1(new_n14324_), .A2(new_n14323_), .ZN(new_n14325_));
  OAI22_X1   g13323(.A1(new_n14317_), .A2(new_n14318_), .B1(new_n14319_), .B2(new_n13244_), .ZN(new_n14326_));
  NAND4_X1   g13324(.A1(new_n14315_), .A2(new_n13222_), .A3(new_n14309_), .A4(new_n14314_), .ZN(new_n14327_));
  NAND2_X1   g13325(.A1(new_n14327_), .A2(new_n14326_), .ZN(new_n14328_));
  NAND2_X1   g13326(.A1(new_n14325_), .A2(new_n14328_), .ZN(new_n14329_));
  AOI21_X1   g13327(.A1(new_n14329_), .A2(new_n14322_), .B(new_n14290_), .ZN(new_n14330_));
  NOR2_X1    g13328(.A1(new_n13230_), .A2(new_n13239_), .ZN(new_n14331_));
  OAI22_X1   g13329(.A1(new_n13270_), .A2(new_n13196_), .B1(new_n14331_), .B2(new_n13240_), .ZN(new_n14332_));
  NOR2_X1    g13330(.A1(new_n14325_), .A2(new_n14328_), .ZN(new_n14333_));
  NOR2_X1    g13331(.A1(new_n14305_), .A2(new_n14321_), .ZN(new_n14334_));
  NOR3_X1    g13332(.A1(new_n14332_), .A2(new_n14333_), .A3(new_n14334_), .ZN(new_n14335_));
  NOR2_X1    g13333(.A1(new_n14335_), .A2(new_n14330_), .ZN(new_n14336_));
  OAI21_X1   g13334(.A1(new_n13389_), .A2(new_n13382_), .B(new_n13395_), .ZN(new_n14337_));
  OAI21_X1   g13335(.A1(new_n13306_), .A2(new_n13294_), .B(new_n13312_), .ZN(new_n14338_));
  INV_X1     g13336(.I(new_n13279_), .ZN(new_n14339_));
  NAND2_X1   g13337(.A1(new_n13280_), .A2(new_n13282_), .ZN(new_n14340_));
  AOI21_X1   g13338(.A1(new_n14340_), .A2(new_n12507_), .B(new_n14339_), .ZN(new_n14341_));
  NAND2_X1   g13339(.A1(new_n14341_), .A2(new_n14338_), .ZN(new_n14342_));
  AOI21_X1   g13340(.A1(new_n13293_), .A2(new_n12474_), .B(new_n13299_), .ZN(new_n14343_));
  NOR2_X1    g13341(.A1(new_n13281_), .A2(new_n13275_), .ZN(new_n14344_));
  NOR2_X1    g13342(.A1(new_n13274_), .A2(new_n12516_), .ZN(new_n14345_));
  NOR2_X1    g13343(.A1(new_n14345_), .A2(new_n14344_), .ZN(new_n14346_));
  OAI21_X1   g13344(.A1(new_n14346_), .A2(new_n13295_), .B(new_n13279_), .ZN(new_n14347_));
  NAND2_X1   g13345(.A1(new_n14347_), .A2(new_n14343_), .ZN(new_n14348_));
  OAI21_X1   g13346(.A1(new_n13307_), .A2(new_n13303_), .B(new_n13283_), .ZN(new_n14349_));
  AOI22_X1   g13347(.A1(new_n14349_), .A2(new_n13385_), .B1(new_n14342_), .B2(new_n14348_), .ZN(new_n14350_));
  NOR2_X1    g13348(.A1(new_n14347_), .A2(new_n14343_), .ZN(new_n14351_));
  NOR2_X1    g13349(.A1(new_n14341_), .A2(new_n14338_), .ZN(new_n14352_));
  AOI21_X1   g13350(.A1(new_n13316_), .A2(new_n13314_), .B(new_n13310_), .ZN(new_n14353_));
  NOR4_X1    g13351(.A1(new_n14353_), .A2(new_n14351_), .A3(new_n14352_), .A4(new_n13301_), .ZN(new_n14354_));
  NOR2_X1    g13352(.A1(new_n14354_), .A2(new_n14350_), .ZN(new_n14355_));
  AOI21_X1   g13353(.A1(new_n13375_), .A2(new_n12413_), .B(new_n13351_), .ZN(new_n14356_));
  NOR2_X1    g13354(.A1(new_n13363_), .A2(new_n13362_), .ZN(new_n14357_));
  OAI21_X1   g13355(.A1(new_n14357_), .A2(new_n13360_), .B(new_n13330_), .ZN(new_n14358_));
  NOR2_X1    g13356(.A1(new_n14358_), .A2(new_n14356_), .ZN(new_n14359_));
  OAI21_X1   g13357(.A1(new_n13348_), .A2(new_n13350_), .B(new_n13344_), .ZN(new_n14360_));
  NAND2_X1   g13358(.A1(new_n13331_), .A2(new_n13333_), .ZN(new_n14361_));
  AOI21_X1   g13359(.A1(new_n14361_), .A2(new_n12443_), .B(new_n13361_), .ZN(new_n14362_));
  NOR2_X1    g13360(.A1(new_n14360_), .A2(new_n14362_), .ZN(new_n14363_));
  AOI21_X1   g13361(.A1(new_n13376_), .A2(new_n13354_), .B(new_n13364_), .ZN(new_n14364_));
  OAI22_X1   g13362(.A1(new_n14363_), .A2(new_n14359_), .B1(new_n14364_), .B2(new_n13353_), .ZN(new_n14365_));
  NAND2_X1   g13363(.A1(new_n14360_), .A2(new_n14362_), .ZN(new_n14366_));
  NAND2_X1   g13364(.A1(new_n14358_), .A2(new_n14356_), .ZN(new_n14367_));
  OAI21_X1   g13365(.A1(new_n13357_), .A2(new_n13355_), .B(new_n13334_), .ZN(new_n14368_));
  NAND4_X1   g13366(.A1(new_n13372_), .A2(new_n14366_), .A3(new_n14367_), .A4(new_n14368_), .ZN(new_n14369_));
  NAND2_X1   g13367(.A1(new_n14369_), .A2(new_n14365_), .ZN(new_n14370_));
  NOR2_X1    g13368(.A1(new_n14355_), .A2(new_n14370_), .ZN(new_n14371_));
  OAI22_X1   g13369(.A1(new_n14353_), .A2(new_n13301_), .B1(new_n14351_), .B2(new_n14352_), .ZN(new_n14372_));
  NAND4_X1   g13370(.A1(new_n13385_), .A2(new_n14342_), .A3(new_n14349_), .A4(new_n14348_), .ZN(new_n14373_));
  NAND2_X1   g13371(.A1(new_n14372_), .A2(new_n14373_), .ZN(new_n14374_));
  AOI22_X1   g13372(.A1(new_n14366_), .A2(new_n14367_), .B1(new_n13372_), .B2(new_n14368_), .ZN(new_n14375_));
  NOR4_X1    g13373(.A1(new_n14363_), .A2(new_n14364_), .A3(new_n14359_), .A4(new_n13353_), .ZN(new_n14376_));
  NOR2_X1    g13374(.A1(new_n14375_), .A2(new_n14376_), .ZN(new_n14377_));
  NOR2_X1    g13375(.A1(new_n14374_), .A2(new_n14377_), .ZN(new_n14378_));
  OAI21_X1   g13376(.A1(new_n14371_), .A2(new_n14378_), .B(new_n14337_), .ZN(new_n14379_));
  AOI21_X1   g13377(.A1(new_n13319_), .A2(new_n13396_), .B(new_n13368_), .ZN(new_n14380_));
  NAND2_X1   g13378(.A1(new_n14374_), .A2(new_n14377_), .ZN(new_n14381_));
  NAND2_X1   g13379(.A1(new_n14355_), .A2(new_n14370_), .ZN(new_n14382_));
  NAND3_X1   g13380(.A1(new_n14382_), .A2(new_n14381_), .A3(new_n14380_), .ZN(new_n14383_));
  NAND2_X1   g13381(.A1(new_n14379_), .A2(new_n14383_), .ZN(new_n14384_));
  NOR2_X1    g13382(.A1(new_n14336_), .A2(new_n14384_), .ZN(new_n14385_));
  OAI21_X1   g13383(.A1(new_n14334_), .A2(new_n14333_), .B(new_n14332_), .ZN(new_n14386_));
  NAND3_X1   g13384(.A1(new_n14329_), .A2(new_n14322_), .A3(new_n14290_), .ZN(new_n14387_));
  NAND2_X1   g13385(.A1(new_n14386_), .A2(new_n14387_), .ZN(new_n14388_));
  AOI21_X1   g13386(.A1(new_n14382_), .A2(new_n14381_), .B(new_n14380_), .ZN(new_n14389_));
  NOR3_X1    g13387(.A1(new_n14371_), .A2(new_n14378_), .A3(new_n14337_), .ZN(new_n14390_));
  NOR2_X1    g13388(.A1(new_n14390_), .A2(new_n14389_), .ZN(new_n14391_));
  NOR2_X1    g13389(.A1(new_n14388_), .A2(new_n14391_), .ZN(new_n14392_));
  OAI21_X1   g13390(.A1(new_n14392_), .A2(new_n14385_), .B(new_n14288_), .ZN(new_n14393_));
  AOI22_X1   g13391(.A1(new_n13394_), .A2(new_n13273_), .B1(new_n13414_), .B2(new_n13401_), .ZN(new_n14394_));
  NAND2_X1   g13392(.A1(new_n14388_), .A2(new_n14391_), .ZN(new_n14395_));
  NAND2_X1   g13393(.A1(new_n14336_), .A2(new_n14384_), .ZN(new_n14396_));
  NAND3_X1   g13394(.A1(new_n14395_), .A2(new_n14396_), .A3(new_n14394_), .ZN(new_n14397_));
  NAND2_X1   g13395(.A1(new_n14393_), .A2(new_n14397_), .ZN(new_n14398_));
  NOR2_X1    g13396(.A1(new_n14286_), .A2(new_n14398_), .ZN(new_n14399_));
  OAI21_X1   g13397(.A1(new_n14284_), .A2(new_n14283_), .B(new_n14282_), .ZN(new_n14400_));
  NAND3_X1   g13398(.A1(new_n14272_), .A2(new_n14279_), .A3(new_n14174_), .ZN(new_n14401_));
  NAND2_X1   g13399(.A1(new_n14400_), .A2(new_n14401_), .ZN(new_n14402_));
  AOI21_X1   g13400(.A1(new_n14395_), .A2(new_n14396_), .B(new_n14394_), .ZN(new_n14403_));
  NOR3_X1    g13401(.A1(new_n14392_), .A2(new_n14385_), .A3(new_n14288_), .ZN(new_n14404_));
  NOR2_X1    g13402(.A1(new_n14403_), .A2(new_n14404_), .ZN(new_n14405_));
  NOR2_X1    g13403(.A1(new_n14402_), .A2(new_n14405_), .ZN(new_n14406_));
  OAI21_X1   g13404(.A1(new_n14406_), .A2(new_n14399_), .B(new_n14173_), .ZN(new_n14407_));
  AOI21_X1   g13405(.A1(new_n13404_), .A2(new_n13408_), .B(new_n13409_), .ZN(new_n14408_));
  AOI21_X1   g13406(.A1(new_n13159_), .A2(new_n13419_), .B(new_n14408_), .ZN(new_n14409_));
  NAND2_X1   g13407(.A1(new_n14402_), .A2(new_n14405_), .ZN(new_n14410_));
  NAND2_X1   g13408(.A1(new_n14286_), .A2(new_n14398_), .ZN(new_n14411_));
  NAND3_X1   g13409(.A1(new_n14410_), .A2(new_n14411_), .A3(new_n14409_), .ZN(new_n14412_));
  NAND2_X1   g13410(.A1(new_n14407_), .A2(new_n14412_), .ZN(new_n14413_));
  NOR2_X1    g13411(.A1(new_n14171_), .A2(new_n14413_), .ZN(new_n14414_));
  OAI21_X1   g13412(.A1(new_n14169_), .A2(new_n14168_), .B(new_n14167_), .ZN(new_n14415_));
  NAND3_X1   g13413(.A1(new_n14158_), .A2(new_n14165_), .A3(new_n13938_), .ZN(new_n14416_));
  NAND2_X1   g13414(.A1(new_n14415_), .A2(new_n14416_), .ZN(new_n14417_));
  AOI21_X1   g13415(.A1(new_n14410_), .A2(new_n14411_), .B(new_n14409_), .ZN(new_n14418_));
  NOR3_X1    g13416(.A1(new_n14406_), .A2(new_n14399_), .A3(new_n14173_), .ZN(new_n14419_));
  NOR2_X1    g13417(.A1(new_n14418_), .A2(new_n14419_), .ZN(new_n14420_));
  NOR2_X1    g13418(.A1(new_n14420_), .A2(new_n14417_), .ZN(new_n14421_));
  OAI21_X1   g13419(.A1(new_n14421_), .A2(new_n14414_), .B(new_n13936_), .ZN(new_n14422_));
  NAND2_X1   g13420(.A1(new_n13411_), .A2(new_n13417_), .ZN(new_n14423_));
  NAND2_X1   g13421(.A1(new_n14423_), .A2(new_n13158_), .ZN(new_n14424_));
  INV_X1     g13422(.I(new_n13421_), .ZN(new_n14425_));
  NAND2_X1   g13423(.A1(new_n14425_), .A2(new_n14424_), .ZN(new_n14426_));
  NAND3_X1   g13424(.A1(new_n14425_), .A2(new_n14424_), .A3(new_n12913_), .ZN(new_n14427_));
  AOI22_X1   g13425(.A1(new_n13933_), .A2(new_n14427_), .B1(new_n14426_), .B2(new_n12914_), .ZN(new_n14428_));
  NAND2_X1   g13426(.A1(new_n14420_), .A2(new_n14417_), .ZN(new_n14429_));
  NAND2_X1   g13427(.A1(new_n14171_), .A2(new_n14413_), .ZN(new_n14430_));
  NAND3_X1   g13428(.A1(new_n14429_), .A2(new_n14430_), .A3(new_n14428_), .ZN(new_n14431_));
  INV_X1     g13429(.I(\A[798] ), .ZN(new_n14432_));
  INV_X1     g13430(.I(\A[796] ), .ZN(new_n14433_));
  INV_X1     g13431(.I(\A[797] ), .ZN(new_n14434_));
  NOR2_X1    g13432(.A1(new_n14433_), .A2(new_n14434_), .ZN(new_n14435_));
  INV_X1     g13433(.I(new_n14435_), .ZN(new_n14436_));
  NOR2_X1    g13434(.A1(new_n14433_), .A2(\A[797] ), .ZN(new_n14437_));
  NOR2_X1    g13435(.A1(new_n14434_), .A2(\A[796] ), .ZN(new_n14438_));
  NOR2_X1    g13436(.A1(new_n14437_), .A2(new_n14438_), .ZN(new_n14439_));
  OAI21_X1   g13437(.A1(new_n14439_), .A2(new_n14432_), .B(new_n14436_), .ZN(new_n14440_));
  INV_X1     g13438(.I(\A[795] ), .ZN(new_n14441_));
  INV_X1     g13439(.I(\A[793] ), .ZN(new_n14442_));
  INV_X1     g13440(.I(\A[794] ), .ZN(new_n14443_));
  NOR2_X1    g13441(.A1(new_n14442_), .A2(new_n14443_), .ZN(new_n14444_));
  INV_X1     g13442(.I(new_n14444_), .ZN(new_n14445_));
  NOR2_X1    g13443(.A1(new_n14442_), .A2(\A[794] ), .ZN(new_n14446_));
  NOR2_X1    g13444(.A1(new_n14443_), .A2(\A[793] ), .ZN(new_n14447_));
  NOR2_X1    g13445(.A1(new_n14446_), .A2(new_n14447_), .ZN(new_n14448_));
  OAI21_X1   g13446(.A1(new_n14448_), .A2(new_n14441_), .B(new_n14445_), .ZN(new_n14449_));
  NAND2_X1   g13447(.A1(new_n14443_), .A2(\A[793] ), .ZN(new_n14450_));
  NAND2_X1   g13448(.A1(new_n14450_), .A2(\A[795] ), .ZN(new_n14451_));
  OAI22_X1   g13449(.A1(new_n14448_), .A2(\A[795] ), .B1(new_n14451_), .B2(new_n14447_), .ZN(new_n14452_));
  NAND2_X1   g13450(.A1(new_n14434_), .A2(\A[796] ), .ZN(new_n14453_));
  NAND2_X1   g13451(.A1(new_n14453_), .A2(\A[798] ), .ZN(new_n14454_));
  OAI22_X1   g13452(.A1(new_n14439_), .A2(\A[798] ), .B1(new_n14454_), .B2(new_n14438_), .ZN(new_n14455_));
  AND2_X2    g13453(.A1(new_n14452_), .A2(new_n14455_), .Z(new_n14456_));
  NAND3_X1   g13454(.A1(new_n14456_), .A2(new_n14440_), .A3(new_n14449_), .ZN(new_n14457_));
  XOR2_X1    g13455(.A1(new_n14452_), .A2(new_n14455_), .Z(new_n14458_));
  NAND2_X1   g13456(.A1(new_n14457_), .A2(new_n14458_), .ZN(new_n14459_));
  INV_X1     g13457(.I(\A[788] ), .ZN(new_n14460_));
  NOR2_X1    g13458(.A1(new_n14460_), .A2(\A[787] ), .ZN(new_n14461_));
  INV_X1     g13459(.I(\A[787] ), .ZN(new_n14462_));
  NOR2_X1    g13460(.A1(new_n14462_), .A2(\A[788] ), .ZN(new_n14463_));
  NOR2_X1    g13461(.A1(new_n14463_), .A2(new_n14461_), .ZN(new_n14464_));
  NAND2_X1   g13462(.A1(new_n14460_), .A2(\A[787] ), .ZN(new_n14465_));
  NAND2_X1   g13463(.A1(new_n14465_), .A2(\A[789] ), .ZN(new_n14466_));
  OAI22_X1   g13464(.A1(new_n14464_), .A2(\A[789] ), .B1(new_n14466_), .B2(new_n14461_), .ZN(new_n14467_));
  INV_X1     g13465(.I(\A[792] ), .ZN(new_n14468_));
  INV_X1     g13466(.I(\A[790] ), .ZN(new_n14469_));
  NAND2_X1   g13467(.A1(new_n14469_), .A2(\A[791] ), .ZN(new_n14470_));
  INV_X1     g13468(.I(\A[791] ), .ZN(new_n14471_));
  NAND2_X1   g13469(.A1(new_n14471_), .A2(\A[790] ), .ZN(new_n14472_));
  NAND2_X1   g13470(.A1(new_n14472_), .A2(new_n14470_), .ZN(new_n14473_));
  AOI21_X1   g13471(.A1(\A[790] ), .A2(new_n14471_), .B(new_n14468_), .ZN(new_n14474_));
  AOI22_X1   g13472(.A1(new_n14473_), .A2(new_n14468_), .B1(new_n14470_), .B2(new_n14474_), .ZN(new_n14475_));
  XNOR2_X1   g13473(.A1(new_n14467_), .A2(new_n14475_), .ZN(new_n14476_));
  NOR2_X1    g13474(.A1(new_n14469_), .A2(new_n14471_), .ZN(new_n14477_));
  INV_X1     g13475(.I(new_n14477_), .ZN(new_n14478_));
  NAND2_X1   g13476(.A1(new_n14473_), .A2(\A[792] ), .ZN(new_n14479_));
  NAND2_X1   g13477(.A1(new_n14479_), .A2(new_n14478_), .ZN(new_n14480_));
  INV_X1     g13478(.I(\A[789] ), .ZN(new_n14481_));
  NOR2_X1    g13479(.A1(new_n14462_), .A2(new_n14460_), .ZN(new_n14482_));
  INV_X1     g13480(.I(new_n14482_), .ZN(new_n14483_));
  OAI21_X1   g13481(.A1(new_n14464_), .A2(new_n14481_), .B(new_n14483_), .ZN(new_n14484_));
  INV_X1     g13482(.I(new_n14467_), .ZN(new_n14485_));
  NOR2_X1    g13483(.A1(new_n14485_), .A2(new_n14475_), .ZN(new_n14486_));
  NAND3_X1   g13484(.A1(new_n14486_), .A2(new_n14480_), .A3(new_n14484_), .ZN(new_n14487_));
  NAND2_X1   g13485(.A1(new_n14487_), .A2(new_n14476_), .ZN(new_n14488_));
  XOR2_X1    g13486(.A1(new_n14459_), .A2(new_n14488_), .Z(new_n14489_));
  INV_X1     g13487(.I(\A[784] ), .ZN(new_n14490_));
  INV_X1     g13488(.I(\A[785] ), .ZN(new_n14491_));
  NOR2_X1    g13489(.A1(new_n14490_), .A2(new_n14491_), .ZN(new_n14492_));
  NAND2_X1   g13490(.A1(new_n14491_), .A2(\A[784] ), .ZN(new_n14493_));
  NAND2_X1   g13491(.A1(new_n14490_), .A2(\A[785] ), .ZN(new_n14494_));
  NAND2_X1   g13492(.A1(new_n14493_), .A2(new_n14494_), .ZN(new_n14495_));
  AOI21_X1   g13493(.A1(new_n14495_), .A2(\A[786] ), .B(new_n14492_), .ZN(new_n14496_));
  INV_X1     g13494(.I(new_n14496_), .ZN(new_n14497_));
  INV_X1     g13495(.I(\A[781] ), .ZN(new_n14498_));
  INV_X1     g13496(.I(\A[782] ), .ZN(new_n14499_));
  NOR2_X1    g13497(.A1(new_n14498_), .A2(new_n14499_), .ZN(new_n14500_));
  NAND2_X1   g13498(.A1(new_n14499_), .A2(\A[781] ), .ZN(new_n14501_));
  NAND2_X1   g13499(.A1(new_n14498_), .A2(\A[782] ), .ZN(new_n14502_));
  NAND2_X1   g13500(.A1(new_n14501_), .A2(new_n14502_), .ZN(new_n14503_));
  AOI21_X1   g13501(.A1(new_n14503_), .A2(\A[783] ), .B(new_n14500_), .ZN(new_n14504_));
  INV_X1     g13502(.I(new_n14504_), .ZN(new_n14505_));
  INV_X1     g13503(.I(\A[783] ), .ZN(new_n14506_));
  AOI21_X1   g13504(.A1(\A[781] ), .A2(new_n14499_), .B(new_n14506_), .ZN(new_n14507_));
  AOI22_X1   g13505(.A1(new_n14503_), .A2(new_n14506_), .B1(new_n14502_), .B2(new_n14507_), .ZN(new_n14508_));
  INV_X1     g13506(.I(\A[786] ), .ZN(new_n14509_));
  AOI21_X1   g13507(.A1(\A[784] ), .A2(new_n14491_), .B(new_n14509_), .ZN(new_n14510_));
  AOI22_X1   g13508(.A1(new_n14495_), .A2(new_n14509_), .B1(new_n14494_), .B2(new_n14510_), .ZN(new_n14511_));
  NOR2_X1    g13509(.A1(new_n14508_), .A2(new_n14511_), .ZN(new_n14512_));
  NAND3_X1   g13510(.A1(new_n14512_), .A2(new_n14497_), .A3(new_n14505_), .ZN(new_n14513_));
  XOR2_X1    g13511(.A1(new_n14508_), .A2(new_n14511_), .Z(new_n14514_));
  NAND2_X1   g13512(.A1(new_n14514_), .A2(new_n14513_), .ZN(new_n14515_));
  INV_X1     g13513(.I(\A[776] ), .ZN(new_n14516_));
  NOR2_X1    g13514(.A1(new_n14516_), .A2(\A[775] ), .ZN(new_n14517_));
  INV_X1     g13515(.I(\A[775] ), .ZN(new_n14518_));
  NOR2_X1    g13516(.A1(new_n14518_), .A2(\A[776] ), .ZN(new_n14519_));
  NOR2_X1    g13517(.A1(new_n14519_), .A2(new_n14517_), .ZN(new_n14520_));
  NAND2_X1   g13518(.A1(new_n14516_), .A2(\A[775] ), .ZN(new_n14521_));
  NAND2_X1   g13519(.A1(new_n14521_), .A2(\A[777] ), .ZN(new_n14522_));
  OAI22_X1   g13520(.A1(new_n14520_), .A2(\A[777] ), .B1(new_n14522_), .B2(new_n14517_), .ZN(new_n14523_));
  INV_X1     g13521(.I(\A[780] ), .ZN(new_n14524_));
  INV_X1     g13522(.I(\A[778] ), .ZN(new_n14525_));
  NAND2_X1   g13523(.A1(new_n14525_), .A2(\A[779] ), .ZN(new_n14526_));
  INV_X1     g13524(.I(\A[779] ), .ZN(new_n14527_));
  NAND2_X1   g13525(.A1(new_n14527_), .A2(\A[778] ), .ZN(new_n14528_));
  NAND2_X1   g13526(.A1(new_n14528_), .A2(new_n14526_), .ZN(new_n14529_));
  AOI21_X1   g13527(.A1(\A[778] ), .A2(new_n14527_), .B(new_n14524_), .ZN(new_n14530_));
  AOI22_X1   g13528(.A1(new_n14529_), .A2(new_n14524_), .B1(new_n14526_), .B2(new_n14530_), .ZN(new_n14531_));
  XNOR2_X1   g13529(.A1(new_n14523_), .A2(new_n14531_), .ZN(new_n14532_));
  NOR2_X1    g13530(.A1(new_n14525_), .A2(new_n14527_), .ZN(new_n14533_));
  AOI21_X1   g13531(.A1(new_n14529_), .A2(\A[780] ), .B(new_n14533_), .ZN(new_n14534_));
  INV_X1     g13532(.I(new_n14534_), .ZN(new_n14535_));
  INV_X1     g13533(.I(\A[777] ), .ZN(new_n14536_));
  NOR2_X1    g13534(.A1(new_n14518_), .A2(new_n14516_), .ZN(new_n14537_));
  INV_X1     g13535(.I(new_n14537_), .ZN(new_n14538_));
  OAI21_X1   g13536(.A1(new_n14520_), .A2(new_n14536_), .B(new_n14538_), .ZN(new_n14539_));
  INV_X1     g13537(.I(new_n14523_), .ZN(new_n14540_));
  NOR2_X1    g13538(.A1(new_n14540_), .A2(new_n14531_), .ZN(new_n14541_));
  NAND3_X1   g13539(.A1(new_n14541_), .A2(new_n14535_), .A3(new_n14539_), .ZN(new_n14542_));
  NAND2_X1   g13540(.A1(new_n14542_), .A2(new_n14532_), .ZN(new_n14543_));
  XOR2_X1    g13541(.A1(new_n14543_), .A2(new_n14515_), .Z(new_n14544_));
  XOR2_X1    g13542(.A1(new_n14489_), .A2(new_n14544_), .Z(new_n14545_));
  INV_X1     g13543(.I(\A[770] ), .ZN(new_n14546_));
  NOR2_X1    g13544(.A1(new_n14546_), .A2(\A[769] ), .ZN(new_n14547_));
  NAND2_X1   g13545(.A1(new_n14546_), .A2(\A[769] ), .ZN(new_n14548_));
  NAND2_X1   g13546(.A1(new_n14548_), .A2(\A[771] ), .ZN(new_n14549_));
  INV_X1     g13547(.I(\A[769] ), .ZN(new_n14550_));
  NOR2_X1    g13548(.A1(new_n14550_), .A2(\A[770] ), .ZN(new_n14551_));
  NOR2_X1    g13549(.A1(new_n14547_), .A2(new_n14551_), .ZN(new_n14552_));
  OAI22_X1   g13550(.A1(new_n14552_), .A2(\A[771] ), .B1(new_n14549_), .B2(new_n14547_), .ZN(new_n14553_));
  INV_X1     g13551(.I(\A[774] ), .ZN(new_n14554_));
  INV_X1     g13552(.I(\A[772] ), .ZN(new_n14555_));
  NAND2_X1   g13553(.A1(new_n14555_), .A2(\A[773] ), .ZN(new_n14556_));
  NOR2_X1    g13554(.A1(new_n14555_), .A2(\A[773] ), .ZN(new_n14557_));
  NOR2_X1    g13555(.A1(new_n14557_), .A2(new_n14554_), .ZN(new_n14558_));
  INV_X1     g13556(.I(\A[773] ), .ZN(new_n14559_));
  NAND2_X1   g13557(.A1(new_n14559_), .A2(\A[772] ), .ZN(new_n14560_));
  NAND2_X1   g13558(.A1(new_n14556_), .A2(new_n14560_), .ZN(new_n14561_));
  AOI22_X1   g13559(.A1(new_n14561_), .A2(new_n14554_), .B1(new_n14558_), .B2(new_n14556_), .ZN(new_n14562_));
  XNOR2_X1   g13560(.A1(new_n14562_), .A2(new_n14553_), .ZN(new_n14563_));
  NOR2_X1    g13561(.A1(new_n14559_), .A2(\A[772] ), .ZN(new_n14564_));
  NOR2_X1    g13562(.A1(new_n14564_), .A2(new_n14557_), .ZN(new_n14565_));
  NOR2_X1    g13563(.A1(new_n14555_), .A2(new_n14559_), .ZN(new_n14566_));
  INV_X1     g13564(.I(new_n14566_), .ZN(new_n14567_));
  OAI21_X1   g13565(.A1(new_n14565_), .A2(new_n14554_), .B(new_n14567_), .ZN(new_n14568_));
  NAND2_X1   g13566(.A1(new_n14550_), .A2(\A[770] ), .ZN(new_n14569_));
  NAND2_X1   g13567(.A1(new_n14569_), .A2(new_n14548_), .ZN(new_n14570_));
  NOR2_X1    g13568(.A1(new_n14550_), .A2(new_n14546_), .ZN(new_n14571_));
  AOI21_X1   g13569(.A1(new_n14570_), .A2(\A[771] ), .B(new_n14571_), .ZN(new_n14572_));
  INV_X1     g13570(.I(new_n14572_), .ZN(new_n14573_));
  INV_X1     g13571(.I(new_n14553_), .ZN(new_n14574_));
  NOR2_X1    g13572(.A1(new_n14574_), .A2(new_n14562_), .ZN(new_n14575_));
  NAND3_X1   g13573(.A1(new_n14575_), .A2(new_n14568_), .A3(new_n14573_), .ZN(new_n14576_));
  NAND2_X1   g13574(.A1(new_n14576_), .A2(new_n14563_), .ZN(new_n14577_));
  INV_X1     g13575(.I(\A[764] ), .ZN(new_n14578_));
  NOR2_X1    g13576(.A1(new_n14578_), .A2(\A[763] ), .ZN(new_n14579_));
  NAND2_X1   g13577(.A1(new_n14578_), .A2(\A[763] ), .ZN(new_n14580_));
  NAND2_X1   g13578(.A1(new_n14580_), .A2(\A[765] ), .ZN(new_n14581_));
  INV_X1     g13579(.I(\A[763] ), .ZN(new_n14582_));
  NOR2_X1    g13580(.A1(new_n14582_), .A2(\A[764] ), .ZN(new_n14583_));
  NOR2_X1    g13581(.A1(new_n14579_), .A2(new_n14583_), .ZN(new_n14584_));
  OAI22_X1   g13582(.A1(new_n14584_), .A2(\A[765] ), .B1(new_n14581_), .B2(new_n14579_), .ZN(new_n14585_));
  INV_X1     g13583(.I(\A[768] ), .ZN(new_n14586_));
  INV_X1     g13584(.I(\A[766] ), .ZN(new_n14587_));
  NAND2_X1   g13585(.A1(new_n14587_), .A2(\A[767] ), .ZN(new_n14588_));
  NOR2_X1    g13586(.A1(new_n14587_), .A2(\A[767] ), .ZN(new_n14589_));
  NOR2_X1    g13587(.A1(new_n14589_), .A2(new_n14586_), .ZN(new_n14590_));
  INV_X1     g13588(.I(\A[767] ), .ZN(new_n14591_));
  NAND2_X1   g13589(.A1(new_n14591_), .A2(\A[766] ), .ZN(new_n14592_));
  NAND2_X1   g13590(.A1(new_n14588_), .A2(new_n14592_), .ZN(new_n14593_));
  AOI22_X1   g13591(.A1(new_n14593_), .A2(new_n14586_), .B1(new_n14590_), .B2(new_n14588_), .ZN(new_n14594_));
  XNOR2_X1   g13592(.A1(new_n14594_), .A2(new_n14585_), .ZN(new_n14595_));
  NOR2_X1    g13593(.A1(new_n14591_), .A2(\A[766] ), .ZN(new_n14596_));
  NOR2_X1    g13594(.A1(new_n14596_), .A2(new_n14589_), .ZN(new_n14597_));
  NOR2_X1    g13595(.A1(new_n14587_), .A2(new_n14591_), .ZN(new_n14598_));
  INV_X1     g13596(.I(new_n14598_), .ZN(new_n14599_));
  OAI21_X1   g13597(.A1(new_n14597_), .A2(new_n14586_), .B(new_n14599_), .ZN(new_n14600_));
  NAND2_X1   g13598(.A1(new_n14582_), .A2(\A[764] ), .ZN(new_n14601_));
  NAND2_X1   g13599(.A1(new_n14601_), .A2(new_n14580_), .ZN(new_n14602_));
  NOR2_X1    g13600(.A1(new_n14582_), .A2(new_n14578_), .ZN(new_n14603_));
  AOI21_X1   g13601(.A1(new_n14602_), .A2(\A[765] ), .B(new_n14603_), .ZN(new_n14604_));
  INV_X1     g13602(.I(new_n14604_), .ZN(new_n14605_));
  INV_X1     g13603(.I(new_n14585_), .ZN(new_n14606_));
  NOR2_X1    g13604(.A1(new_n14606_), .A2(new_n14594_), .ZN(new_n14607_));
  NAND3_X1   g13605(.A1(new_n14607_), .A2(new_n14600_), .A3(new_n14605_), .ZN(new_n14608_));
  NAND2_X1   g13606(.A1(new_n14608_), .A2(new_n14595_), .ZN(new_n14609_));
  XOR2_X1    g13607(.A1(new_n14577_), .A2(new_n14609_), .Z(new_n14610_));
  INV_X1     g13608(.I(\A[758] ), .ZN(new_n14611_));
  NOR2_X1    g13609(.A1(new_n14611_), .A2(\A[757] ), .ZN(new_n14612_));
  NAND2_X1   g13610(.A1(new_n14611_), .A2(\A[757] ), .ZN(new_n14613_));
  NAND2_X1   g13611(.A1(new_n14613_), .A2(\A[759] ), .ZN(new_n14614_));
  INV_X1     g13612(.I(\A[757] ), .ZN(new_n14615_));
  NOR2_X1    g13613(.A1(new_n14615_), .A2(\A[758] ), .ZN(new_n14616_));
  NOR2_X1    g13614(.A1(new_n14612_), .A2(new_n14616_), .ZN(new_n14617_));
  OAI22_X1   g13615(.A1(new_n14617_), .A2(\A[759] ), .B1(new_n14614_), .B2(new_n14612_), .ZN(new_n14618_));
  INV_X1     g13616(.I(\A[762] ), .ZN(new_n14619_));
  INV_X1     g13617(.I(\A[760] ), .ZN(new_n14620_));
  NAND2_X1   g13618(.A1(new_n14620_), .A2(\A[761] ), .ZN(new_n14621_));
  NOR2_X1    g13619(.A1(new_n14620_), .A2(\A[761] ), .ZN(new_n14622_));
  NOR2_X1    g13620(.A1(new_n14622_), .A2(new_n14619_), .ZN(new_n14623_));
  INV_X1     g13621(.I(\A[761] ), .ZN(new_n14624_));
  NAND2_X1   g13622(.A1(new_n14624_), .A2(\A[760] ), .ZN(new_n14625_));
  NAND2_X1   g13623(.A1(new_n14621_), .A2(new_n14625_), .ZN(new_n14626_));
  AOI22_X1   g13624(.A1(new_n14626_), .A2(new_n14619_), .B1(new_n14623_), .B2(new_n14621_), .ZN(new_n14627_));
  XNOR2_X1   g13625(.A1(new_n14627_), .A2(new_n14618_), .ZN(new_n14628_));
  NOR2_X1    g13626(.A1(new_n14624_), .A2(\A[760] ), .ZN(new_n14629_));
  NOR2_X1    g13627(.A1(new_n14629_), .A2(new_n14622_), .ZN(new_n14630_));
  NOR2_X1    g13628(.A1(new_n14620_), .A2(new_n14624_), .ZN(new_n14631_));
  INV_X1     g13629(.I(new_n14631_), .ZN(new_n14632_));
  OAI21_X1   g13630(.A1(new_n14630_), .A2(new_n14619_), .B(new_n14632_), .ZN(new_n14633_));
  NAND2_X1   g13631(.A1(new_n14615_), .A2(\A[758] ), .ZN(new_n14634_));
  NAND2_X1   g13632(.A1(new_n14634_), .A2(new_n14613_), .ZN(new_n14635_));
  NOR2_X1    g13633(.A1(new_n14615_), .A2(new_n14611_), .ZN(new_n14636_));
  AOI21_X1   g13634(.A1(new_n14635_), .A2(\A[759] ), .B(new_n14636_), .ZN(new_n14637_));
  INV_X1     g13635(.I(new_n14637_), .ZN(new_n14638_));
  INV_X1     g13636(.I(new_n14618_), .ZN(new_n14639_));
  NOR2_X1    g13637(.A1(new_n14639_), .A2(new_n14627_), .ZN(new_n14640_));
  NAND3_X1   g13638(.A1(new_n14640_), .A2(new_n14633_), .A3(new_n14638_), .ZN(new_n14641_));
  NAND2_X1   g13639(.A1(new_n14641_), .A2(new_n14628_), .ZN(new_n14642_));
  INV_X1     g13640(.I(\A[752] ), .ZN(new_n14643_));
  NOR2_X1    g13641(.A1(new_n14643_), .A2(\A[751] ), .ZN(new_n14644_));
  NAND2_X1   g13642(.A1(new_n14643_), .A2(\A[751] ), .ZN(new_n14645_));
  NAND2_X1   g13643(.A1(new_n14645_), .A2(\A[753] ), .ZN(new_n14646_));
  INV_X1     g13644(.I(\A[751] ), .ZN(new_n14647_));
  NOR2_X1    g13645(.A1(new_n14647_), .A2(\A[752] ), .ZN(new_n14648_));
  NOR2_X1    g13646(.A1(new_n14644_), .A2(new_n14648_), .ZN(new_n14649_));
  OAI22_X1   g13647(.A1(new_n14649_), .A2(\A[753] ), .B1(new_n14646_), .B2(new_n14644_), .ZN(new_n14650_));
  INV_X1     g13648(.I(\A[756] ), .ZN(new_n14651_));
  INV_X1     g13649(.I(\A[754] ), .ZN(new_n14652_));
  NAND2_X1   g13650(.A1(new_n14652_), .A2(\A[755] ), .ZN(new_n14653_));
  NOR2_X1    g13651(.A1(new_n14652_), .A2(\A[755] ), .ZN(new_n14654_));
  NOR2_X1    g13652(.A1(new_n14654_), .A2(new_n14651_), .ZN(new_n14655_));
  INV_X1     g13653(.I(\A[755] ), .ZN(new_n14656_));
  NAND2_X1   g13654(.A1(new_n14656_), .A2(\A[754] ), .ZN(new_n14657_));
  NAND2_X1   g13655(.A1(new_n14653_), .A2(new_n14657_), .ZN(new_n14658_));
  AOI22_X1   g13656(.A1(new_n14658_), .A2(new_n14651_), .B1(new_n14655_), .B2(new_n14653_), .ZN(new_n14659_));
  XNOR2_X1   g13657(.A1(new_n14659_), .A2(new_n14650_), .ZN(new_n14660_));
  NOR2_X1    g13658(.A1(new_n14656_), .A2(\A[754] ), .ZN(new_n14661_));
  NOR2_X1    g13659(.A1(new_n14661_), .A2(new_n14654_), .ZN(new_n14662_));
  NOR2_X1    g13660(.A1(new_n14652_), .A2(new_n14656_), .ZN(new_n14663_));
  INV_X1     g13661(.I(new_n14663_), .ZN(new_n14664_));
  OAI21_X1   g13662(.A1(new_n14662_), .A2(new_n14651_), .B(new_n14664_), .ZN(new_n14665_));
  NAND2_X1   g13663(.A1(new_n14647_), .A2(\A[752] ), .ZN(new_n14666_));
  NAND2_X1   g13664(.A1(new_n14666_), .A2(new_n14645_), .ZN(new_n14667_));
  NOR2_X1    g13665(.A1(new_n14647_), .A2(new_n14643_), .ZN(new_n14668_));
  AOI21_X1   g13666(.A1(new_n14667_), .A2(\A[753] ), .B(new_n14668_), .ZN(new_n14669_));
  INV_X1     g13667(.I(new_n14669_), .ZN(new_n14670_));
  INV_X1     g13668(.I(new_n14650_), .ZN(new_n14671_));
  NOR2_X1    g13669(.A1(new_n14671_), .A2(new_n14659_), .ZN(new_n14672_));
  NAND3_X1   g13670(.A1(new_n14672_), .A2(new_n14665_), .A3(new_n14670_), .ZN(new_n14673_));
  NAND2_X1   g13671(.A1(new_n14673_), .A2(new_n14660_), .ZN(new_n14674_));
  XOR2_X1    g13672(.A1(new_n14642_), .A2(new_n14674_), .Z(new_n14675_));
  XOR2_X1    g13673(.A1(new_n14610_), .A2(new_n14675_), .Z(new_n14676_));
  XNOR2_X1   g13674(.A1(new_n14676_), .A2(new_n14545_), .ZN(new_n14677_));
  INV_X1     g13675(.I(\A[836] ), .ZN(new_n14678_));
  NOR2_X1    g13676(.A1(new_n14678_), .A2(\A[835] ), .ZN(new_n14679_));
  INV_X1     g13677(.I(\A[835] ), .ZN(new_n14680_));
  NOR2_X1    g13678(.A1(new_n14680_), .A2(\A[836] ), .ZN(new_n14681_));
  NOR2_X1    g13679(.A1(new_n14681_), .A2(new_n14679_), .ZN(new_n14682_));
  NAND2_X1   g13680(.A1(new_n14678_), .A2(\A[835] ), .ZN(new_n14683_));
  NAND2_X1   g13681(.A1(new_n14683_), .A2(\A[837] ), .ZN(new_n14684_));
  OAI22_X1   g13682(.A1(new_n14682_), .A2(\A[837] ), .B1(new_n14684_), .B2(new_n14679_), .ZN(new_n14685_));
  INV_X1     g13683(.I(\A[840] ), .ZN(new_n14686_));
  INV_X1     g13684(.I(\A[838] ), .ZN(new_n14687_));
  NAND2_X1   g13685(.A1(new_n14687_), .A2(\A[839] ), .ZN(new_n14688_));
  INV_X1     g13686(.I(\A[839] ), .ZN(new_n14689_));
  NAND2_X1   g13687(.A1(new_n14689_), .A2(\A[838] ), .ZN(new_n14690_));
  NAND2_X1   g13688(.A1(new_n14690_), .A2(new_n14688_), .ZN(new_n14691_));
  AOI21_X1   g13689(.A1(\A[838] ), .A2(new_n14689_), .B(new_n14686_), .ZN(new_n14692_));
  AOI22_X1   g13690(.A1(new_n14691_), .A2(new_n14686_), .B1(new_n14688_), .B2(new_n14692_), .ZN(new_n14693_));
  XNOR2_X1   g13691(.A1(new_n14685_), .A2(new_n14693_), .ZN(new_n14694_));
  AND2_X2    g13692(.A1(new_n14690_), .A2(new_n14688_), .Z(new_n14695_));
  NOR2_X1    g13693(.A1(new_n14687_), .A2(new_n14689_), .ZN(new_n14696_));
  INV_X1     g13694(.I(new_n14696_), .ZN(new_n14697_));
  OAI21_X1   g13695(.A1(new_n14695_), .A2(new_n14686_), .B(new_n14697_), .ZN(new_n14698_));
  INV_X1     g13696(.I(\A[837] ), .ZN(new_n14699_));
  NOR2_X1    g13697(.A1(new_n14680_), .A2(new_n14678_), .ZN(new_n14700_));
  INV_X1     g13698(.I(new_n14700_), .ZN(new_n14701_));
  OAI21_X1   g13699(.A1(new_n14682_), .A2(new_n14699_), .B(new_n14701_), .ZN(new_n14702_));
  INV_X1     g13700(.I(new_n14685_), .ZN(new_n14703_));
  NOR2_X1    g13701(.A1(new_n14703_), .A2(new_n14693_), .ZN(new_n14704_));
  NAND3_X1   g13702(.A1(new_n14704_), .A2(new_n14698_), .A3(new_n14702_), .ZN(new_n14705_));
  NAND2_X1   g13703(.A1(new_n14705_), .A2(new_n14694_), .ZN(new_n14706_));
  INV_X1     g13704(.I(\A[843] ), .ZN(new_n14707_));
  INV_X1     g13705(.I(\A[841] ), .ZN(new_n14708_));
  NAND2_X1   g13706(.A1(new_n14708_), .A2(\A[842] ), .ZN(new_n14709_));
  INV_X1     g13707(.I(\A[842] ), .ZN(new_n14710_));
  NAND2_X1   g13708(.A1(new_n14710_), .A2(\A[841] ), .ZN(new_n14711_));
  NAND2_X1   g13709(.A1(new_n14711_), .A2(new_n14709_), .ZN(new_n14712_));
  NOR2_X1    g13710(.A1(new_n14708_), .A2(\A[842] ), .ZN(new_n14713_));
  NOR2_X1    g13711(.A1(new_n14713_), .A2(new_n14707_), .ZN(new_n14714_));
  AOI22_X1   g13712(.A1(new_n14712_), .A2(new_n14707_), .B1(new_n14714_), .B2(new_n14709_), .ZN(new_n14715_));
  INV_X1     g13713(.I(\A[846] ), .ZN(new_n14716_));
  INV_X1     g13714(.I(\A[844] ), .ZN(new_n14717_));
  NAND2_X1   g13715(.A1(new_n14717_), .A2(\A[845] ), .ZN(new_n14718_));
  INV_X1     g13716(.I(\A[845] ), .ZN(new_n14719_));
  NAND2_X1   g13717(.A1(new_n14719_), .A2(\A[844] ), .ZN(new_n14720_));
  NAND2_X1   g13718(.A1(new_n14720_), .A2(new_n14718_), .ZN(new_n14721_));
  AOI21_X1   g13719(.A1(\A[844] ), .A2(new_n14719_), .B(new_n14716_), .ZN(new_n14722_));
  AOI22_X1   g13720(.A1(new_n14721_), .A2(new_n14716_), .B1(new_n14718_), .B2(new_n14722_), .ZN(new_n14723_));
  XOR2_X1    g13721(.A1(new_n14715_), .A2(new_n14723_), .Z(new_n14724_));
  AND2_X2    g13722(.A1(new_n14720_), .A2(new_n14718_), .Z(new_n14725_));
  NOR2_X1    g13723(.A1(new_n14717_), .A2(new_n14719_), .ZN(new_n14726_));
  INV_X1     g13724(.I(new_n14726_), .ZN(new_n14727_));
  OAI21_X1   g13725(.A1(new_n14725_), .A2(new_n14716_), .B(new_n14727_), .ZN(new_n14728_));
  NOR2_X1    g13726(.A1(new_n14710_), .A2(\A[841] ), .ZN(new_n14729_));
  NOR2_X1    g13727(.A1(new_n14713_), .A2(new_n14729_), .ZN(new_n14730_));
  NOR2_X1    g13728(.A1(new_n14708_), .A2(new_n14710_), .ZN(new_n14731_));
  INV_X1     g13729(.I(new_n14731_), .ZN(new_n14732_));
  OAI21_X1   g13730(.A1(new_n14730_), .A2(new_n14707_), .B(new_n14732_), .ZN(new_n14733_));
  NOR2_X1    g13731(.A1(new_n14715_), .A2(new_n14723_), .ZN(new_n14734_));
  NAND3_X1   g13732(.A1(new_n14734_), .A2(new_n14728_), .A3(new_n14733_), .ZN(new_n14735_));
  NAND2_X1   g13733(.A1(new_n14724_), .A2(new_n14735_), .ZN(new_n14736_));
  XOR2_X1    g13734(.A1(new_n14706_), .A2(new_n14736_), .Z(new_n14737_));
  INV_X1     g13735(.I(\A[825] ), .ZN(new_n14738_));
  INV_X1     g13736(.I(\A[823] ), .ZN(new_n14739_));
  NAND2_X1   g13737(.A1(new_n14739_), .A2(\A[824] ), .ZN(new_n14740_));
  INV_X1     g13738(.I(\A[824] ), .ZN(new_n14741_));
  NAND2_X1   g13739(.A1(new_n14741_), .A2(\A[823] ), .ZN(new_n14742_));
  NAND2_X1   g13740(.A1(new_n14742_), .A2(new_n14740_), .ZN(new_n14743_));
  NOR2_X1    g13741(.A1(new_n14739_), .A2(\A[824] ), .ZN(new_n14744_));
  NOR2_X1    g13742(.A1(new_n14744_), .A2(new_n14738_), .ZN(new_n14745_));
  AOI22_X1   g13743(.A1(new_n14743_), .A2(new_n14738_), .B1(new_n14745_), .B2(new_n14740_), .ZN(new_n14746_));
  INV_X1     g13744(.I(\A[828] ), .ZN(new_n14747_));
  INV_X1     g13745(.I(\A[826] ), .ZN(new_n14748_));
  NAND2_X1   g13746(.A1(new_n14748_), .A2(\A[827] ), .ZN(new_n14749_));
  INV_X1     g13747(.I(\A[827] ), .ZN(new_n14750_));
  NAND2_X1   g13748(.A1(new_n14750_), .A2(\A[826] ), .ZN(new_n14751_));
  NAND2_X1   g13749(.A1(new_n14751_), .A2(new_n14749_), .ZN(new_n14752_));
  AOI21_X1   g13750(.A1(\A[826] ), .A2(new_n14750_), .B(new_n14747_), .ZN(new_n14753_));
  AOI22_X1   g13751(.A1(new_n14752_), .A2(new_n14747_), .B1(new_n14749_), .B2(new_n14753_), .ZN(new_n14754_));
  XOR2_X1    g13752(.A1(new_n14746_), .A2(new_n14754_), .Z(new_n14755_));
  NOR2_X1    g13753(.A1(new_n14748_), .A2(new_n14750_), .ZN(new_n14756_));
  AOI21_X1   g13754(.A1(new_n14752_), .A2(\A[828] ), .B(new_n14756_), .ZN(new_n14757_));
  INV_X1     g13755(.I(new_n14757_), .ZN(new_n14758_));
  NOR2_X1    g13756(.A1(new_n14741_), .A2(\A[823] ), .ZN(new_n14759_));
  NOR2_X1    g13757(.A1(new_n14744_), .A2(new_n14759_), .ZN(new_n14760_));
  NOR2_X1    g13758(.A1(new_n14739_), .A2(new_n14741_), .ZN(new_n14761_));
  INV_X1     g13759(.I(new_n14761_), .ZN(new_n14762_));
  OAI21_X1   g13760(.A1(new_n14760_), .A2(new_n14738_), .B(new_n14762_), .ZN(new_n14763_));
  NOR2_X1    g13761(.A1(new_n14746_), .A2(new_n14754_), .ZN(new_n14764_));
  NAND3_X1   g13762(.A1(new_n14764_), .A2(new_n14758_), .A3(new_n14763_), .ZN(new_n14765_));
  NAND2_X1   g13763(.A1(new_n14755_), .A2(new_n14765_), .ZN(new_n14766_));
  INV_X1     g13764(.I(\A[831] ), .ZN(new_n14767_));
  INV_X1     g13765(.I(\A[829] ), .ZN(new_n14768_));
  NAND2_X1   g13766(.A1(new_n14768_), .A2(\A[830] ), .ZN(new_n14769_));
  INV_X1     g13767(.I(\A[830] ), .ZN(new_n14770_));
  NAND2_X1   g13768(.A1(new_n14770_), .A2(\A[829] ), .ZN(new_n14771_));
  NAND2_X1   g13769(.A1(new_n14771_), .A2(new_n14769_), .ZN(new_n14772_));
  NOR2_X1    g13770(.A1(new_n14768_), .A2(\A[830] ), .ZN(new_n14773_));
  NOR2_X1    g13771(.A1(new_n14773_), .A2(new_n14767_), .ZN(new_n14774_));
  AOI22_X1   g13772(.A1(new_n14772_), .A2(new_n14767_), .B1(new_n14774_), .B2(new_n14769_), .ZN(new_n14775_));
  INV_X1     g13773(.I(\A[834] ), .ZN(new_n14776_));
  INV_X1     g13774(.I(\A[832] ), .ZN(new_n14777_));
  NAND2_X1   g13775(.A1(new_n14777_), .A2(\A[833] ), .ZN(new_n14778_));
  INV_X1     g13776(.I(\A[833] ), .ZN(new_n14779_));
  NAND2_X1   g13777(.A1(new_n14779_), .A2(\A[832] ), .ZN(new_n14780_));
  NAND2_X1   g13778(.A1(new_n14780_), .A2(new_n14778_), .ZN(new_n14781_));
  AOI21_X1   g13779(.A1(\A[832] ), .A2(new_n14779_), .B(new_n14776_), .ZN(new_n14782_));
  AOI22_X1   g13780(.A1(new_n14781_), .A2(new_n14776_), .B1(new_n14778_), .B2(new_n14782_), .ZN(new_n14783_));
  XOR2_X1    g13781(.A1(new_n14775_), .A2(new_n14783_), .Z(new_n14784_));
  NOR2_X1    g13782(.A1(new_n14777_), .A2(new_n14779_), .ZN(new_n14785_));
  AOI21_X1   g13783(.A1(new_n14781_), .A2(\A[834] ), .B(new_n14785_), .ZN(new_n14786_));
  INV_X1     g13784(.I(new_n14786_), .ZN(new_n14787_));
  NOR2_X1    g13785(.A1(new_n14770_), .A2(\A[829] ), .ZN(new_n14788_));
  NOR2_X1    g13786(.A1(new_n14773_), .A2(new_n14788_), .ZN(new_n14789_));
  NOR2_X1    g13787(.A1(new_n14768_), .A2(new_n14770_), .ZN(new_n14790_));
  INV_X1     g13788(.I(new_n14790_), .ZN(new_n14791_));
  OAI21_X1   g13789(.A1(new_n14789_), .A2(new_n14767_), .B(new_n14791_), .ZN(new_n14792_));
  NOR2_X1    g13790(.A1(new_n14775_), .A2(new_n14783_), .ZN(new_n14793_));
  NAND3_X1   g13791(.A1(new_n14793_), .A2(new_n14787_), .A3(new_n14792_), .ZN(new_n14794_));
  NAND2_X1   g13792(.A1(new_n14784_), .A2(new_n14794_), .ZN(new_n14795_));
  XOR2_X1    g13793(.A1(new_n14766_), .A2(new_n14795_), .Z(new_n14796_));
  XOR2_X1    g13794(.A1(new_n14737_), .A2(new_n14796_), .Z(new_n14797_));
  INV_X1     g13795(.I(\A[813] ), .ZN(new_n14798_));
  INV_X1     g13796(.I(\A[811] ), .ZN(new_n14799_));
  NAND2_X1   g13797(.A1(new_n14799_), .A2(\A[812] ), .ZN(new_n14800_));
  INV_X1     g13798(.I(\A[812] ), .ZN(new_n14801_));
  NAND2_X1   g13799(.A1(new_n14801_), .A2(\A[811] ), .ZN(new_n14802_));
  NAND2_X1   g13800(.A1(new_n14802_), .A2(new_n14800_), .ZN(new_n14803_));
  AOI21_X1   g13801(.A1(\A[811] ), .A2(new_n14801_), .B(new_n14798_), .ZN(new_n14804_));
  AOI22_X1   g13802(.A1(new_n14803_), .A2(new_n14798_), .B1(new_n14800_), .B2(new_n14804_), .ZN(new_n14805_));
  INV_X1     g13803(.I(\A[816] ), .ZN(new_n14806_));
  INV_X1     g13804(.I(\A[814] ), .ZN(new_n14807_));
  NAND2_X1   g13805(.A1(new_n14807_), .A2(\A[815] ), .ZN(new_n14808_));
  INV_X1     g13806(.I(\A[815] ), .ZN(new_n14809_));
  NAND2_X1   g13807(.A1(new_n14809_), .A2(\A[814] ), .ZN(new_n14810_));
  NAND2_X1   g13808(.A1(new_n14810_), .A2(new_n14808_), .ZN(new_n14811_));
  AOI21_X1   g13809(.A1(\A[814] ), .A2(new_n14809_), .B(new_n14806_), .ZN(new_n14812_));
  AOI22_X1   g13810(.A1(new_n14811_), .A2(new_n14806_), .B1(new_n14808_), .B2(new_n14812_), .ZN(new_n14813_));
  XOR2_X1    g13811(.A1(new_n14805_), .A2(new_n14813_), .Z(new_n14814_));
  NOR2_X1    g13812(.A1(new_n14807_), .A2(new_n14809_), .ZN(new_n14815_));
  AOI21_X1   g13813(.A1(new_n14811_), .A2(\A[816] ), .B(new_n14815_), .ZN(new_n14816_));
  INV_X1     g13814(.I(new_n14816_), .ZN(new_n14817_));
  NOR2_X1    g13815(.A1(new_n14799_), .A2(new_n14801_), .ZN(new_n14818_));
  AOI21_X1   g13816(.A1(new_n14803_), .A2(\A[813] ), .B(new_n14818_), .ZN(new_n14819_));
  INV_X1     g13817(.I(new_n14819_), .ZN(new_n14820_));
  NOR2_X1    g13818(.A1(new_n14805_), .A2(new_n14813_), .ZN(new_n14821_));
  NAND3_X1   g13819(.A1(new_n14821_), .A2(new_n14817_), .A3(new_n14820_), .ZN(new_n14822_));
  NAND2_X1   g13820(.A1(new_n14814_), .A2(new_n14822_), .ZN(new_n14823_));
  INV_X1     g13821(.I(\A[818] ), .ZN(new_n14824_));
  NOR2_X1    g13822(.A1(new_n14824_), .A2(\A[817] ), .ZN(new_n14825_));
  INV_X1     g13823(.I(\A[817] ), .ZN(new_n14826_));
  NOR2_X1    g13824(.A1(new_n14826_), .A2(\A[818] ), .ZN(new_n14827_));
  NOR2_X1    g13825(.A1(new_n14827_), .A2(new_n14825_), .ZN(new_n14828_));
  NAND2_X1   g13826(.A1(new_n14824_), .A2(\A[817] ), .ZN(new_n14829_));
  NAND2_X1   g13827(.A1(new_n14829_), .A2(\A[819] ), .ZN(new_n14830_));
  OAI22_X1   g13828(.A1(new_n14828_), .A2(\A[819] ), .B1(new_n14830_), .B2(new_n14825_), .ZN(new_n14831_));
  INV_X1     g13829(.I(\A[822] ), .ZN(new_n14832_));
  INV_X1     g13830(.I(\A[820] ), .ZN(new_n14833_));
  NAND2_X1   g13831(.A1(new_n14833_), .A2(\A[821] ), .ZN(new_n14834_));
  INV_X1     g13832(.I(\A[821] ), .ZN(new_n14835_));
  NAND2_X1   g13833(.A1(new_n14835_), .A2(\A[820] ), .ZN(new_n14836_));
  NAND2_X1   g13834(.A1(new_n14836_), .A2(new_n14834_), .ZN(new_n14837_));
  AOI21_X1   g13835(.A1(\A[820] ), .A2(new_n14835_), .B(new_n14832_), .ZN(new_n14838_));
  AOI22_X1   g13836(.A1(new_n14837_), .A2(new_n14832_), .B1(new_n14834_), .B2(new_n14838_), .ZN(new_n14839_));
  XNOR2_X1   g13837(.A1(new_n14831_), .A2(new_n14839_), .ZN(new_n14840_));
  NOR2_X1    g13838(.A1(new_n14833_), .A2(new_n14835_), .ZN(new_n14841_));
  INV_X1     g13839(.I(new_n14841_), .ZN(new_n14842_));
  NAND2_X1   g13840(.A1(new_n14837_), .A2(\A[822] ), .ZN(new_n14843_));
  NAND2_X1   g13841(.A1(new_n14843_), .A2(new_n14842_), .ZN(new_n14844_));
  INV_X1     g13842(.I(\A[819] ), .ZN(new_n14845_));
  NOR2_X1    g13843(.A1(new_n14826_), .A2(new_n14824_), .ZN(new_n14846_));
  INV_X1     g13844(.I(new_n14846_), .ZN(new_n14847_));
  OAI21_X1   g13845(.A1(new_n14828_), .A2(new_n14845_), .B(new_n14847_), .ZN(new_n14848_));
  INV_X1     g13846(.I(new_n14831_), .ZN(new_n14849_));
  NOR2_X1    g13847(.A1(new_n14849_), .A2(new_n14839_), .ZN(new_n14850_));
  NAND3_X1   g13848(.A1(new_n14850_), .A2(new_n14844_), .A3(new_n14848_), .ZN(new_n14851_));
  NAND2_X1   g13849(.A1(new_n14851_), .A2(new_n14840_), .ZN(new_n14852_));
  XOR2_X1    g13850(.A1(new_n14852_), .A2(new_n14823_), .Z(new_n14853_));
  INV_X1     g13851(.I(\A[806] ), .ZN(new_n14854_));
  NOR2_X1    g13852(.A1(new_n14854_), .A2(\A[805] ), .ZN(new_n14855_));
  NAND2_X1   g13853(.A1(new_n14854_), .A2(\A[805] ), .ZN(new_n14856_));
  NAND2_X1   g13854(.A1(new_n14856_), .A2(\A[807] ), .ZN(new_n14857_));
  INV_X1     g13855(.I(\A[805] ), .ZN(new_n14858_));
  NOR2_X1    g13856(.A1(new_n14858_), .A2(\A[806] ), .ZN(new_n14859_));
  NOR2_X1    g13857(.A1(new_n14855_), .A2(new_n14859_), .ZN(new_n14860_));
  OAI22_X1   g13858(.A1(new_n14860_), .A2(\A[807] ), .B1(new_n14857_), .B2(new_n14855_), .ZN(new_n14861_));
  INV_X1     g13859(.I(\A[810] ), .ZN(new_n14862_));
  INV_X1     g13860(.I(\A[808] ), .ZN(new_n14863_));
  NAND2_X1   g13861(.A1(new_n14863_), .A2(\A[809] ), .ZN(new_n14864_));
  NOR2_X1    g13862(.A1(new_n14863_), .A2(\A[809] ), .ZN(new_n14865_));
  NOR2_X1    g13863(.A1(new_n14865_), .A2(new_n14862_), .ZN(new_n14866_));
  INV_X1     g13864(.I(\A[809] ), .ZN(new_n14867_));
  NAND2_X1   g13865(.A1(new_n14867_), .A2(\A[808] ), .ZN(new_n14868_));
  NAND2_X1   g13866(.A1(new_n14864_), .A2(new_n14868_), .ZN(new_n14869_));
  AOI22_X1   g13867(.A1(new_n14869_), .A2(new_n14862_), .B1(new_n14866_), .B2(new_n14864_), .ZN(new_n14870_));
  XNOR2_X1   g13868(.A1(new_n14870_), .A2(new_n14861_), .ZN(new_n14871_));
  NOR2_X1    g13869(.A1(new_n14867_), .A2(\A[808] ), .ZN(new_n14872_));
  NOR2_X1    g13870(.A1(new_n14872_), .A2(new_n14865_), .ZN(new_n14873_));
  NOR2_X1    g13871(.A1(new_n14863_), .A2(new_n14867_), .ZN(new_n14874_));
  INV_X1     g13872(.I(new_n14874_), .ZN(new_n14875_));
  OAI21_X1   g13873(.A1(new_n14873_), .A2(new_n14862_), .B(new_n14875_), .ZN(new_n14876_));
  NAND2_X1   g13874(.A1(new_n14858_), .A2(\A[806] ), .ZN(new_n14877_));
  NAND2_X1   g13875(.A1(new_n14877_), .A2(new_n14856_), .ZN(new_n14878_));
  NOR2_X1    g13876(.A1(new_n14858_), .A2(new_n14854_), .ZN(new_n14879_));
  AOI21_X1   g13877(.A1(new_n14878_), .A2(\A[807] ), .B(new_n14879_), .ZN(new_n14880_));
  INV_X1     g13878(.I(new_n14880_), .ZN(new_n14881_));
  INV_X1     g13879(.I(new_n14861_), .ZN(new_n14882_));
  NOR2_X1    g13880(.A1(new_n14882_), .A2(new_n14870_), .ZN(new_n14883_));
  NAND3_X1   g13881(.A1(new_n14883_), .A2(new_n14876_), .A3(new_n14881_), .ZN(new_n14884_));
  NAND2_X1   g13882(.A1(new_n14884_), .A2(new_n14871_), .ZN(new_n14885_));
  INV_X1     g13883(.I(\A[801] ), .ZN(new_n14886_));
  INV_X1     g13884(.I(\A[799] ), .ZN(new_n14887_));
  NAND2_X1   g13885(.A1(new_n14887_), .A2(\A[800] ), .ZN(new_n14888_));
  NOR2_X1    g13886(.A1(new_n14887_), .A2(\A[800] ), .ZN(new_n14889_));
  NOR2_X1    g13887(.A1(new_n14889_), .A2(new_n14886_), .ZN(new_n14890_));
  INV_X1     g13888(.I(\A[800] ), .ZN(new_n14891_));
  NAND2_X1   g13889(.A1(new_n14891_), .A2(\A[799] ), .ZN(new_n14892_));
  NAND2_X1   g13890(.A1(new_n14888_), .A2(new_n14892_), .ZN(new_n14893_));
  AOI22_X1   g13891(.A1(new_n14893_), .A2(new_n14886_), .B1(new_n14890_), .B2(new_n14888_), .ZN(new_n14894_));
  INV_X1     g13892(.I(\A[804] ), .ZN(new_n14895_));
  INV_X1     g13893(.I(\A[802] ), .ZN(new_n14896_));
  NAND2_X1   g13894(.A1(new_n14896_), .A2(\A[803] ), .ZN(new_n14897_));
  NOR2_X1    g13895(.A1(new_n14896_), .A2(\A[803] ), .ZN(new_n14898_));
  NOR2_X1    g13896(.A1(new_n14898_), .A2(new_n14895_), .ZN(new_n14899_));
  INV_X1     g13897(.I(\A[803] ), .ZN(new_n14900_));
  NAND2_X1   g13898(.A1(new_n14900_), .A2(\A[802] ), .ZN(new_n14901_));
  NAND2_X1   g13899(.A1(new_n14897_), .A2(new_n14901_), .ZN(new_n14902_));
  AOI22_X1   g13900(.A1(new_n14902_), .A2(new_n14895_), .B1(new_n14899_), .B2(new_n14897_), .ZN(new_n14903_));
  XOR2_X1    g13901(.A1(new_n14894_), .A2(new_n14903_), .Z(new_n14904_));
  NOR2_X1    g13902(.A1(new_n14896_), .A2(new_n14900_), .ZN(new_n14905_));
  AOI21_X1   g13903(.A1(new_n14902_), .A2(\A[804] ), .B(new_n14905_), .ZN(new_n14906_));
  NOR2_X1    g13904(.A1(new_n14887_), .A2(new_n14891_), .ZN(new_n14907_));
  AOI21_X1   g13905(.A1(new_n14893_), .A2(\A[801] ), .B(new_n14907_), .ZN(new_n14908_));
  OR4_X2     g13906(.A1(new_n14894_), .A2(new_n14903_), .A3(new_n14906_), .A4(new_n14908_), .Z(new_n14909_));
  NAND2_X1   g13907(.A1(new_n14904_), .A2(new_n14909_), .ZN(new_n14910_));
  XOR2_X1    g13908(.A1(new_n14885_), .A2(new_n14910_), .Z(new_n14911_));
  XOR2_X1    g13909(.A1(new_n14911_), .A2(new_n14853_), .Z(new_n14912_));
  XNOR2_X1   g13910(.A1(new_n14912_), .A2(new_n14797_), .ZN(new_n14913_));
  XOR2_X1    g13911(.A1(new_n14677_), .A2(new_n14913_), .Z(new_n14914_));
  INV_X1     g13912(.I(\A[741] ), .ZN(new_n14915_));
  INV_X1     g13913(.I(\A[739] ), .ZN(new_n14916_));
  NAND2_X1   g13914(.A1(new_n14916_), .A2(\A[740] ), .ZN(new_n14917_));
  INV_X1     g13915(.I(\A[740] ), .ZN(new_n14918_));
  NAND2_X1   g13916(.A1(new_n14918_), .A2(\A[739] ), .ZN(new_n14919_));
  NAND2_X1   g13917(.A1(new_n14919_), .A2(new_n14917_), .ZN(new_n14920_));
  AOI21_X1   g13918(.A1(\A[739] ), .A2(new_n14918_), .B(new_n14915_), .ZN(new_n14921_));
  AOI22_X1   g13919(.A1(new_n14920_), .A2(new_n14915_), .B1(new_n14917_), .B2(new_n14921_), .ZN(new_n14922_));
  INV_X1     g13920(.I(\A[744] ), .ZN(new_n14923_));
  INV_X1     g13921(.I(\A[742] ), .ZN(new_n14924_));
  NAND2_X1   g13922(.A1(new_n14924_), .A2(\A[743] ), .ZN(new_n14925_));
  INV_X1     g13923(.I(\A[743] ), .ZN(new_n14926_));
  NAND2_X1   g13924(.A1(new_n14926_), .A2(\A[742] ), .ZN(new_n14927_));
  NAND2_X1   g13925(.A1(new_n14927_), .A2(new_n14925_), .ZN(new_n14928_));
  AOI21_X1   g13926(.A1(\A[742] ), .A2(new_n14926_), .B(new_n14923_), .ZN(new_n14929_));
  AOI22_X1   g13927(.A1(new_n14928_), .A2(new_n14923_), .B1(new_n14925_), .B2(new_n14929_), .ZN(new_n14930_));
  XOR2_X1    g13928(.A1(new_n14922_), .A2(new_n14930_), .Z(new_n14931_));
  NOR2_X1    g13929(.A1(new_n14924_), .A2(new_n14926_), .ZN(new_n14932_));
  AOI21_X1   g13930(.A1(new_n14928_), .A2(\A[744] ), .B(new_n14932_), .ZN(new_n14933_));
  INV_X1     g13931(.I(new_n14933_), .ZN(new_n14934_));
  AND2_X2    g13932(.A1(new_n14919_), .A2(new_n14917_), .Z(new_n14935_));
  NOR2_X1    g13933(.A1(new_n14916_), .A2(new_n14918_), .ZN(new_n14936_));
  INV_X1     g13934(.I(new_n14936_), .ZN(new_n14937_));
  OAI21_X1   g13935(.A1(new_n14935_), .A2(new_n14915_), .B(new_n14937_), .ZN(new_n14938_));
  NOR2_X1    g13936(.A1(new_n14922_), .A2(new_n14930_), .ZN(new_n14939_));
  NAND3_X1   g13937(.A1(new_n14939_), .A2(new_n14934_), .A3(new_n14938_), .ZN(new_n14940_));
  NAND2_X1   g13938(.A1(new_n14931_), .A2(new_n14940_), .ZN(new_n14941_));
  INV_X1     g13939(.I(\A[746] ), .ZN(new_n14942_));
  NOR2_X1    g13940(.A1(new_n14942_), .A2(\A[745] ), .ZN(new_n14943_));
  INV_X1     g13941(.I(\A[745] ), .ZN(new_n14944_));
  NOR2_X1    g13942(.A1(new_n14944_), .A2(\A[746] ), .ZN(new_n14945_));
  NOR2_X1    g13943(.A1(new_n14945_), .A2(new_n14943_), .ZN(new_n14946_));
  NAND2_X1   g13944(.A1(new_n14942_), .A2(\A[745] ), .ZN(new_n14947_));
  NAND2_X1   g13945(.A1(new_n14947_), .A2(\A[747] ), .ZN(new_n14948_));
  OAI22_X1   g13946(.A1(new_n14946_), .A2(\A[747] ), .B1(new_n14948_), .B2(new_n14943_), .ZN(new_n14949_));
  INV_X1     g13947(.I(\A[750] ), .ZN(new_n14950_));
  INV_X1     g13948(.I(\A[748] ), .ZN(new_n14951_));
  NAND2_X1   g13949(.A1(new_n14951_), .A2(\A[749] ), .ZN(new_n14952_));
  INV_X1     g13950(.I(\A[749] ), .ZN(new_n14953_));
  NAND2_X1   g13951(.A1(new_n14953_), .A2(\A[748] ), .ZN(new_n14954_));
  NAND2_X1   g13952(.A1(new_n14954_), .A2(new_n14952_), .ZN(new_n14955_));
  AOI21_X1   g13953(.A1(\A[748] ), .A2(new_n14953_), .B(new_n14950_), .ZN(new_n14956_));
  AOI22_X1   g13954(.A1(new_n14955_), .A2(new_n14950_), .B1(new_n14952_), .B2(new_n14956_), .ZN(new_n14957_));
  XNOR2_X1   g13955(.A1(new_n14949_), .A2(new_n14957_), .ZN(new_n14958_));
  AND2_X2    g13956(.A1(new_n14954_), .A2(new_n14952_), .Z(new_n14959_));
  NOR2_X1    g13957(.A1(new_n14951_), .A2(new_n14953_), .ZN(new_n14960_));
  INV_X1     g13958(.I(new_n14960_), .ZN(new_n14961_));
  OAI21_X1   g13959(.A1(new_n14959_), .A2(new_n14950_), .B(new_n14961_), .ZN(new_n14962_));
  INV_X1     g13960(.I(\A[747] ), .ZN(new_n14963_));
  NOR2_X1    g13961(.A1(new_n14944_), .A2(new_n14942_), .ZN(new_n14964_));
  INV_X1     g13962(.I(new_n14964_), .ZN(new_n14965_));
  OAI21_X1   g13963(.A1(new_n14946_), .A2(new_n14963_), .B(new_n14965_), .ZN(new_n14966_));
  INV_X1     g13964(.I(new_n14949_), .ZN(new_n14967_));
  NOR2_X1    g13965(.A1(new_n14967_), .A2(new_n14957_), .ZN(new_n14968_));
  NAND3_X1   g13966(.A1(new_n14968_), .A2(new_n14962_), .A3(new_n14966_), .ZN(new_n14969_));
  NAND2_X1   g13967(.A1(new_n14969_), .A2(new_n14958_), .ZN(new_n14970_));
  XOR2_X1    g13968(.A1(new_n14970_), .A2(new_n14941_), .Z(new_n14971_));
  INV_X1     g13969(.I(\A[728] ), .ZN(new_n14972_));
  NOR2_X1    g13970(.A1(new_n14972_), .A2(\A[727] ), .ZN(new_n14973_));
  INV_X1     g13971(.I(\A[727] ), .ZN(new_n14974_));
  NOR2_X1    g13972(.A1(new_n14974_), .A2(\A[728] ), .ZN(new_n14975_));
  NOR2_X1    g13973(.A1(new_n14975_), .A2(new_n14973_), .ZN(new_n14976_));
  NAND2_X1   g13974(.A1(new_n14972_), .A2(\A[727] ), .ZN(new_n14977_));
  NAND2_X1   g13975(.A1(new_n14977_), .A2(\A[729] ), .ZN(new_n14978_));
  OAI22_X1   g13976(.A1(new_n14976_), .A2(\A[729] ), .B1(new_n14978_), .B2(new_n14973_), .ZN(new_n14979_));
  INV_X1     g13977(.I(\A[732] ), .ZN(new_n14980_));
  INV_X1     g13978(.I(\A[730] ), .ZN(new_n14981_));
  NAND2_X1   g13979(.A1(new_n14981_), .A2(\A[731] ), .ZN(new_n14982_));
  INV_X1     g13980(.I(\A[731] ), .ZN(new_n14983_));
  NAND2_X1   g13981(.A1(new_n14983_), .A2(\A[730] ), .ZN(new_n14984_));
  NAND2_X1   g13982(.A1(new_n14984_), .A2(new_n14982_), .ZN(new_n14985_));
  AOI21_X1   g13983(.A1(\A[730] ), .A2(new_n14983_), .B(new_n14980_), .ZN(new_n14986_));
  AOI22_X1   g13984(.A1(new_n14985_), .A2(new_n14980_), .B1(new_n14982_), .B2(new_n14986_), .ZN(new_n14987_));
  XNOR2_X1   g13985(.A1(new_n14979_), .A2(new_n14987_), .ZN(new_n14988_));
  NOR2_X1    g13986(.A1(new_n14981_), .A2(new_n14983_), .ZN(new_n14989_));
  AOI21_X1   g13987(.A1(new_n14985_), .A2(\A[732] ), .B(new_n14989_), .ZN(new_n14990_));
  INV_X1     g13988(.I(new_n14990_), .ZN(new_n14991_));
  INV_X1     g13989(.I(\A[729] ), .ZN(new_n14992_));
  NOR2_X1    g13990(.A1(new_n14974_), .A2(new_n14972_), .ZN(new_n14993_));
  INV_X1     g13991(.I(new_n14993_), .ZN(new_n14994_));
  OAI21_X1   g13992(.A1(new_n14976_), .A2(new_n14992_), .B(new_n14994_), .ZN(new_n14995_));
  INV_X1     g13993(.I(new_n14979_), .ZN(new_n14996_));
  NOR2_X1    g13994(.A1(new_n14996_), .A2(new_n14987_), .ZN(new_n14997_));
  NAND3_X1   g13995(.A1(new_n14997_), .A2(new_n14991_), .A3(new_n14995_), .ZN(new_n14998_));
  NAND2_X1   g13996(.A1(new_n14998_), .A2(new_n14988_), .ZN(new_n14999_));
  INV_X1     g13997(.I(\A[735] ), .ZN(new_n15000_));
  INV_X1     g13998(.I(\A[733] ), .ZN(new_n15001_));
  NAND2_X1   g13999(.A1(new_n15001_), .A2(\A[734] ), .ZN(new_n15002_));
  INV_X1     g14000(.I(\A[734] ), .ZN(new_n15003_));
  NAND2_X1   g14001(.A1(new_n15003_), .A2(\A[733] ), .ZN(new_n15004_));
  NAND2_X1   g14002(.A1(new_n15004_), .A2(new_n15002_), .ZN(new_n15005_));
  NOR2_X1    g14003(.A1(new_n15001_), .A2(\A[734] ), .ZN(new_n15006_));
  NOR2_X1    g14004(.A1(new_n15006_), .A2(new_n15000_), .ZN(new_n15007_));
  AOI22_X1   g14005(.A1(new_n15005_), .A2(new_n15000_), .B1(new_n15007_), .B2(new_n15002_), .ZN(new_n15008_));
  INV_X1     g14006(.I(\A[738] ), .ZN(new_n15009_));
  INV_X1     g14007(.I(\A[736] ), .ZN(new_n15010_));
  NAND2_X1   g14008(.A1(new_n15010_), .A2(\A[737] ), .ZN(new_n15011_));
  INV_X1     g14009(.I(\A[737] ), .ZN(new_n15012_));
  NAND2_X1   g14010(.A1(new_n15012_), .A2(\A[736] ), .ZN(new_n15013_));
  NAND2_X1   g14011(.A1(new_n15013_), .A2(new_n15011_), .ZN(new_n15014_));
  AOI21_X1   g14012(.A1(\A[736] ), .A2(new_n15012_), .B(new_n15009_), .ZN(new_n15015_));
  AOI22_X1   g14013(.A1(new_n15014_), .A2(new_n15009_), .B1(new_n15011_), .B2(new_n15015_), .ZN(new_n15016_));
  XOR2_X1    g14014(.A1(new_n15008_), .A2(new_n15016_), .Z(new_n15017_));
  NOR2_X1    g14015(.A1(new_n15010_), .A2(new_n15012_), .ZN(new_n15018_));
  AOI21_X1   g14016(.A1(new_n15014_), .A2(\A[738] ), .B(new_n15018_), .ZN(new_n15019_));
  INV_X1     g14017(.I(new_n15019_), .ZN(new_n15020_));
  NOR2_X1    g14018(.A1(new_n15003_), .A2(\A[733] ), .ZN(new_n15021_));
  NOR2_X1    g14019(.A1(new_n15006_), .A2(new_n15021_), .ZN(new_n15022_));
  NOR2_X1    g14020(.A1(new_n15001_), .A2(new_n15003_), .ZN(new_n15023_));
  INV_X1     g14021(.I(new_n15023_), .ZN(new_n15024_));
  OAI21_X1   g14022(.A1(new_n15022_), .A2(new_n15000_), .B(new_n15024_), .ZN(new_n15025_));
  NOR2_X1    g14023(.A1(new_n15008_), .A2(new_n15016_), .ZN(new_n15026_));
  NAND3_X1   g14024(.A1(new_n15026_), .A2(new_n15020_), .A3(new_n15025_), .ZN(new_n15027_));
  NAND2_X1   g14025(.A1(new_n15017_), .A2(new_n15027_), .ZN(new_n15028_));
  XOR2_X1    g14026(.A1(new_n14999_), .A2(new_n15028_), .Z(new_n15029_));
  XOR2_X1    g14027(.A1(new_n14971_), .A2(new_n15029_), .Z(new_n15030_));
  INV_X1     g14028(.I(\A[717] ), .ZN(new_n15031_));
  INV_X1     g14029(.I(\A[715] ), .ZN(new_n15032_));
  NAND2_X1   g14030(.A1(new_n15032_), .A2(\A[716] ), .ZN(new_n15033_));
  INV_X1     g14031(.I(\A[716] ), .ZN(new_n15034_));
  NAND2_X1   g14032(.A1(new_n15034_), .A2(\A[715] ), .ZN(new_n15035_));
  NAND2_X1   g14033(.A1(new_n15035_), .A2(new_n15033_), .ZN(new_n15036_));
  AOI21_X1   g14034(.A1(\A[715] ), .A2(new_n15034_), .B(new_n15031_), .ZN(new_n15037_));
  AOI22_X1   g14035(.A1(new_n15036_), .A2(new_n15031_), .B1(new_n15033_), .B2(new_n15037_), .ZN(new_n15038_));
  INV_X1     g14036(.I(\A[720] ), .ZN(new_n15039_));
  INV_X1     g14037(.I(\A[718] ), .ZN(new_n15040_));
  NAND2_X1   g14038(.A1(new_n15040_), .A2(\A[719] ), .ZN(new_n15041_));
  INV_X1     g14039(.I(\A[719] ), .ZN(new_n15042_));
  NAND2_X1   g14040(.A1(new_n15042_), .A2(\A[718] ), .ZN(new_n15043_));
  NAND2_X1   g14041(.A1(new_n15043_), .A2(new_n15041_), .ZN(new_n15044_));
  AOI21_X1   g14042(.A1(\A[718] ), .A2(new_n15042_), .B(new_n15039_), .ZN(new_n15045_));
  AOI22_X1   g14043(.A1(new_n15044_), .A2(new_n15039_), .B1(new_n15041_), .B2(new_n15045_), .ZN(new_n15046_));
  XOR2_X1    g14044(.A1(new_n15038_), .A2(new_n15046_), .Z(new_n15047_));
  NOR2_X1    g14045(.A1(new_n15040_), .A2(new_n15042_), .ZN(new_n15048_));
  AOI21_X1   g14046(.A1(new_n15044_), .A2(\A[720] ), .B(new_n15048_), .ZN(new_n15049_));
  NOR2_X1    g14047(.A1(new_n15032_), .A2(new_n15034_), .ZN(new_n15050_));
  AOI21_X1   g14048(.A1(new_n15036_), .A2(\A[717] ), .B(new_n15050_), .ZN(new_n15051_));
  OR4_X2     g14049(.A1(new_n15038_), .A2(new_n15046_), .A3(new_n15049_), .A4(new_n15051_), .Z(new_n15052_));
  NAND2_X1   g14050(.A1(new_n15047_), .A2(new_n15052_), .ZN(new_n15053_));
  INV_X1     g14051(.I(\A[723] ), .ZN(new_n15054_));
  INV_X1     g14052(.I(\A[721] ), .ZN(new_n15055_));
  NAND2_X1   g14053(.A1(new_n15055_), .A2(\A[722] ), .ZN(new_n15056_));
  INV_X1     g14054(.I(\A[722] ), .ZN(new_n15057_));
  NAND2_X1   g14055(.A1(new_n15057_), .A2(\A[721] ), .ZN(new_n15058_));
  NAND2_X1   g14056(.A1(new_n15058_), .A2(new_n15056_), .ZN(new_n15059_));
  AOI21_X1   g14057(.A1(\A[721] ), .A2(new_n15057_), .B(new_n15054_), .ZN(new_n15060_));
  AOI22_X1   g14058(.A1(new_n15059_), .A2(new_n15054_), .B1(new_n15056_), .B2(new_n15060_), .ZN(new_n15061_));
  INV_X1     g14059(.I(\A[726] ), .ZN(new_n15062_));
  INV_X1     g14060(.I(\A[724] ), .ZN(new_n15063_));
  NAND2_X1   g14061(.A1(new_n15063_), .A2(\A[725] ), .ZN(new_n15064_));
  INV_X1     g14062(.I(\A[725] ), .ZN(new_n15065_));
  NAND2_X1   g14063(.A1(new_n15065_), .A2(\A[724] ), .ZN(new_n15066_));
  NAND2_X1   g14064(.A1(new_n15066_), .A2(new_n15064_), .ZN(new_n15067_));
  AOI21_X1   g14065(.A1(\A[724] ), .A2(new_n15065_), .B(new_n15062_), .ZN(new_n15068_));
  AOI22_X1   g14066(.A1(new_n15067_), .A2(new_n15062_), .B1(new_n15064_), .B2(new_n15068_), .ZN(new_n15069_));
  XOR2_X1    g14067(.A1(new_n15061_), .A2(new_n15069_), .Z(new_n15070_));
  NOR2_X1    g14068(.A1(new_n15063_), .A2(new_n15065_), .ZN(new_n15071_));
  AOI21_X1   g14069(.A1(new_n15067_), .A2(\A[726] ), .B(new_n15071_), .ZN(new_n15072_));
  NOR2_X1    g14070(.A1(new_n15055_), .A2(new_n15057_), .ZN(new_n15073_));
  AOI21_X1   g14071(.A1(new_n15059_), .A2(\A[723] ), .B(new_n15073_), .ZN(new_n15074_));
  OR4_X2     g14072(.A1(new_n15061_), .A2(new_n15069_), .A3(new_n15072_), .A4(new_n15074_), .Z(new_n15075_));
  NAND2_X1   g14073(.A1(new_n15070_), .A2(new_n15075_), .ZN(new_n15076_));
  XOR2_X1    g14074(.A1(new_n15053_), .A2(new_n15076_), .Z(new_n15077_));
  INV_X1     g14075(.I(\A[710] ), .ZN(new_n15078_));
  NOR2_X1    g14076(.A1(new_n15078_), .A2(\A[709] ), .ZN(new_n15079_));
  NAND2_X1   g14077(.A1(new_n15078_), .A2(\A[709] ), .ZN(new_n15080_));
  NAND2_X1   g14078(.A1(new_n15080_), .A2(\A[711] ), .ZN(new_n15081_));
  INV_X1     g14079(.I(\A[709] ), .ZN(new_n15082_));
  NOR2_X1    g14080(.A1(new_n15082_), .A2(\A[710] ), .ZN(new_n15083_));
  NOR2_X1    g14081(.A1(new_n15079_), .A2(new_n15083_), .ZN(new_n15084_));
  OAI22_X1   g14082(.A1(new_n15084_), .A2(\A[711] ), .B1(new_n15081_), .B2(new_n15079_), .ZN(new_n15085_));
  INV_X1     g14083(.I(\A[714] ), .ZN(new_n15086_));
  INV_X1     g14084(.I(\A[712] ), .ZN(new_n15087_));
  NAND2_X1   g14085(.A1(new_n15087_), .A2(\A[713] ), .ZN(new_n15088_));
  NOR2_X1    g14086(.A1(new_n15087_), .A2(\A[713] ), .ZN(new_n15089_));
  NOR2_X1    g14087(.A1(new_n15089_), .A2(new_n15086_), .ZN(new_n15090_));
  INV_X1     g14088(.I(\A[713] ), .ZN(new_n15091_));
  NAND2_X1   g14089(.A1(new_n15091_), .A2(\A[712] ), .ZN(new_n15092_));
  NAND2_X1   g14090(.A1(new_n15088_), .A2(new_n15092_), .ZN(new_n15093_));
  AOI22_X1   g14091(.A1(new_n15093_), .A2(new_n15086_), .B1(new_n15090_), .B2(new_n15088_), .ZN(new_n15094_));
  XNOR2_X1   g14092(.A1(new_n15094_), .A2(new_n15085_), .ZN(new_n15095_));
  NOR2_X1    g14093(.A1(new_n15091_), .A2(\A[712] ), .ZN(new_n15096_));
  NOR2_X1    g14094(.A1(new_n15096_), .A2(new_n15089_), .ZN(new_n15097_));
  NOR2_X1    g14095(.A1(new_n15087_), .A2(new_n15091_), .ZN(new_n15098_));
  INV_X1     g14096(.I(new_n15098_), .ZN(new_n15099_));
  OAI21_X1   g14097(.A1(new_n15097_), .A2(new_n15086_), .B(new_n15099_), .ZN(new_n15100_));
  NAND2_X1   g14098(.A1(new_n15082_), .A2(\A[710] ), .ZN(new_n15101_));
  NAND2_X1   g14099(.A1(new_n15101_), .A2(new_n15080_), .ZN(new_n15102_));
  NOR2_X1    g14100(.A1(new_n15082_), .A2(new_n15078_), .ZN(new_n15103_));
  AOI21_X1   g14101(.A1(new_n15102_), .A2(\A[711] ), .B(new_n15103_), .ZN(new_n15104_));
  INV_X1     g14102(.I(new_n15104_), .ZN(new_n15105_));
  INV_X1     g14103(.I(new_n15085_), .ZN(new_n15106_));
  NOR2_X1    g14104(.A1(new_n15106_), .A2(new_n15094_), .ZN(new_n15107_));
  NAND3_X1   g14105(.A1(new_n15107_), .A2(new_n15100_), .A3(new_n15105_), .ZN(new_n15108_));
  NAND2_X1   g14106(.A1(new_n15108_), .A2(new_n15095_), .ZN(new_n15109_));
  INV_X1     g14107(.I(\A[704] ), .ZN(new_n15110_));
  NOR2_X1    g14108(.A1(new_n15110_), .A2(\A[703] ), .ZN(new_n15111_));
  NAND2_X1   g14109(.A1(new_n15110_), .A2(\A[703] ), .ZN(new_n15112_));
  NAND2_X1   g14110(.A1(new_n15112_), .A2(\A[705] ), .ZN(new_n15113_));
  INV_X1     g14111(.I(\A[703] ), .ZN(new_n15114_));
  NOR2_X1    g14112(.A1(new_n15114_), .A2(\A[704] ), .ZN(new_n15115_));
  NOR2_X1    g14113(.A1(new_n15111_), .A2(new_n15115_), .ZN(new_n15116_));
  OAI22_X1   g14114(.A1(new_n15116_), .A2(\A[705] ), .B1(new_n15113_), .B2(new_n15111_), .ZN(new_n15117_));
  INV_X1     g14115(.I(\A[708] ), .ZN(new_n15118_));
  INV_X1     g14116(.I(\A[706] ), .ZN(new_n15119_));
  NAND2_X1   g14117(.A1(new_n15119_), .A2(\A[707] ), .ZN(new_n15120_));
  NOR2_X1    g14118(.A1(new_n15119_), .A2(\A[707] ), .ZN(new_n15121_));
  NOR2_X1    g14119(.A1(new_n15121_), .A2(new_n15118_), .ZN(new_n15122_));
  INV_X1     g14120(.I(\A[707] ), .ZN(new_n15123_));
  NAND2_X1   g14121(.A1(new_n15123_), .A2(\A[706] ), .ZN(new_n15124_));
  NAND2_X1   g14122(.A1(new_n15120_), .A2(new_n15124_), .ZN(new_n15125_));
  AOI22_X1   g14123(.A1(new_n15125_), .A2(new_n15118_), .B1(new_n15122_), .B2(new_n15120_), .ZN(new_n15126_));
  XNOR2_X1   g14124(.A1(new_n15126_), .A2(new_n15117_), .ZN(new_n15127_));
  NOR2_X1    g14125(.A1(new_n15123_), .A2(\A[706] ), .ZN(new_n15128_));
  NOR2_X1    g14126(.A1(new_n15128_), .A2(new_n15121_), .ZN(new_n15129_));
  NOR2_X1    g14127(.A1(new_n15119_), .A2(new_n15123_), .ZN(new_n15130_));
  INV_X1     g14128(.I(new_n15130_), .ZN(new_n15131_));
  OAI21_X1   g14129(.A1(new_n15129_), .A2(new_n15118_), .B(new_n15131_), .ZN(new_n15132_));
  NAND2_X1   g14130(.A1(new_n15114_), .A2(\A[704] ), .ZN(new_n15133_));
  NAND2_X1   g14131(.A1(new_n15133_), .A2(new_n15112_), .ZN(new_n15134_));
  NOR2_X1    g14132(.A1(new_n15114_), .A2(new_n15110_), .ZN(new_n15135_));
  AOI21_X1   g14133(.A1(new_n15134_), .A2(\A[705] ), .B(new_n15135_), .ZN(new_n15136_));
  INV_X1     g14134(.I(new_n15136_), .ZN(new_n15137_));
  INV_X1     g14135(.I(new_n15117_), .ZN(new_n15138_));
  NOR2_X1    g14136(.A1(new_n15138_), .A2(new_n15126_), .ZN(new_n15139_));
  NAND3_X1   g14137(.A1(new_n15139_), .A2(new_n15132_), .A3(new_n15137_), .ZN(new_n15140_));
  NAND2_X1   g14138(.A1(new_n15140_), .A2(new_n15127_), .ZN(new_n15141_));
  XOR2_X1    g14139(.A1(new_n15109_), .A2(new_n15141_), .Z(new_n15142_));
  XOR2_X1    g14140(.A1(new_n15142_), .A2(new_n15077_), .Z(new_n15143_));
  XNOR2_X1   g14141(.A1(new_n15143_), .A2(new_n15030_), .ZN(new_n15144_));
  INV_X1     g14142(.I(\A[698] ), .ZN(new_n15145_));
  NOR2_X1    g14143(.A1(new_n15145_), .A2(\A[697] ), .ZN(new_n15146_));
  NAND2_X1   g14144(.A1(new_n15145_), .A2(\A[697] ), .ZN(new_n15147_));
  NAND2_X1   g14145(.A1(new_n15147_), .A2(\A[699] ), .ZN(new_n15148_));
  INV_X1     g14146(.I(\A[697] ), .ZN(new_n15149_));
  NOR2_X1    g14147(.A1(new_n15149_), .A2(\A[698] ), .ZN(new_n15150_));
  NOR2_X1    g14148(.A1(new_n15146_), .A2(new_n15150_), .ZN(new_n15151_));
  OAI22_X1   g14149(.A1(new_n15151_), .A2(\A[699] ), .B1(new_n15148_), .B2(new_n15146_), .ZN(new_n15152_));
  INV_X1     g14150(.I(\A[702] ), .ZN(new_n15153_));
  INV_X1     g14151(.I(\A[700] ), .ZN(new_n15154_));
  NAND2_X1   g14152(.A1(new_n15154_), .A2(\A[701] ), .ZN(new_n15155_));
  NOR2_X1    g14153(.A1(new_n15154_), .A2(\A[701] ), .ZN(new_n15156_));
  NOR2_X1    g14154(.A1(new_n15156_), .A2(new_n15153_), .ZN(new_n15157_));
  INV_X1     g14155(.I(\A[701] ), .ZN(new_n15158_));
  NAND2_X1   g14156(.A1(new_n15158_), .A2(\A[700] ), .ZN(new_n15159_));
  NAND2_X1   g14157(.A1(new_n15155_), .A2(new_n15159_), .ZN(new_n15160_));
  AOI22_X1   g14158(.A1(new_n15160_), .A2(new_n15153_), .B1(new_n15157_), .B2(new_n15155_), .ZN(new_n15161_));
  XNOR2_X1   g14159(.A1(new_n15161_), .A2(new_n15152_), .ZN(new_n15162_));
  NOR2_X1    g14160(.A1(new_n15158_), .A2(\A[700] ), .ZN(new_n15163_));
  NOR2_X1    g14161(.A1(new_n15163_), .A2(new_n15156_), .ZN(new_n15164_));
  NOR2_X1    g14162(.A1(new_n15154_), .A2(new_n15158_), .ZN(new_n15165_));
  INV_X1     g14163(.I(new_n15165_), .ZN(new_n15166_));
  OAI21_X1   g14164(.A1(new_n15164_), .A2(new_n15153_), .B(new_n15166_), .ZN(new_n15167_));
  NAND2_X1   g14165(.A1(new_n15149_), .A2(\A[698] ), .ZN(new_n15168_));
  NAND2_X1   g14166(.A1(new_n15168_), .A2(new_n15147_), .ZN(new_n15169_));
  NOR2_X1    g14167(.A1(new_n15149_), .A2(new_n15145_), .ZN(new_n15170_));
  AOI21_X1   g14168(.A1(new_n15169_), .A2(\A[699] ), .B(new_n15170_), .ZN(new_n15171_));
  INV_X1     g14169(.I(new_n15171_), .ZN(new_n15172_));
  INV_X1     g14170(.I(new_n15152_), .ZN(new_n15173_));
  NOR2_X1    g14171(.A1(new_n15173_), .A2(new_n15161_), .ZN(new_n15174_));
  NAND3_X1   g14172(.A1(new_n15174_), .A2(new_n15167_), .A3(new_n15172_), .ZN(new_n15175_));
  NAND2_X1   g14173(.A1(new_n15175_), .A2(new_n15162_), .ZN(new_n15176_));
  INV_X1     g14174(.I(\A[692] ), .ZN(new_n15177_));
  NOR2_X1    g14175(.A1(new_n15177_), .A2(\A[691] ), .ZN(new_n15178_));
  NAND2_X1   g14176(.A1(new_n15177_), .A2(\A[691] ), .ZN(new_n15179_));
  NAND2_X1   g14177(.A1(new_n15179_), .A2(\A[693] ), .ZN(new_n15180_));
  INV_X1     g14178(.I(\A[691] ), .ZN(new_n15181_));
  NOR2_X1    g14179(.A1(new_n15181_), .A2(\A[692] ), .ZN(new_n15182_));
  NOR2_X1    g14180(.A1(new_n15178_), .A2(new_n15182_), .ZN(new_n15183_));
  OAI22_X1   g14181(.A1(new_n15183_), .A2(\A[693] ), .B1(new_n15180_), .B2(new_n15178_), .ZN(new_n15184_));
  INV_X1     g14182(.I(\A[696] ), .ZN(new_n15185_));
  INV_X1     g14183(.I(\A[694] ), .ZN(new_n15186_));
  NAND2_X1   g14184(.A1(new_n15186_), .A2(\A[695] ), .ZN(new_n15187_));
  NOR2_X1    g14185(.A1(new_n15186_), .A2(\A[695] ), .ZN(new_n15188_));
  NOR2_X1    g14186(.A1(new_n15188_), .A2(new_n15185_), .ZN(new_n15189_));
  INV_X1     g14187(.I(\A[695] ), .ZN(new_n15190_));
  NAND2_X1   g14188(.A1(new_n15190_), .A2(\A[694] ), .ZN(new_n15191_));
  NAND2_X1   g14189(.A1(new_n15187_), .A2(new_n15191_), .ZN(new_n15192_));
  AOI22_X1   g14190(.A1(new_n15192_), .A2(new_n15185_), .B1(new_n15189_), .B2(new_n15187_), .ZN(new_n15193_));
  XNOR2_X1   g14191(.A1(new_n15193_), .A2(new_n15184_), .ZN(new_n15194_));
  NOR2_X1    g14192(.A1(new_n15190_), .A2(\A[694] ), .ZN(new_n15195_));
  NOR2_X1    g14193(.A1(new_n15195_), .A2(new_n15188_), .ZN(new_n15196_));
  NOR2_X1    g14194(.A1(new_n15186_), .A2(new_n15190_), .ZN(new_n15197_));
  INV_X1     g14195(.I(new_n15197_), .ZN(new_n15198_));
  OAI21_X1   g14196(.A1(new_n15196_), .A2(new_n15185_), .B(new_n15198_), .ZN(new_n15199_));
  NAND2_X1   g14197(.A1(new_n15181_), .A2(\A[692] ), .ZN(new_n15200_));
  NAND2_X1   g14198(.A1(new_n15200_), .A2(new_n15179_), .ZN(new_n15201_));
  NOR2_X1    g14199(.A1(new_n15181_), .A2(new_n15177_), .ZN(new_n15202_));
  AOI21_X1   g14200(.A1(new_n15201_), .A2(\A[693] ), .B(new_n15202_), .ZN(new_n15203_));
  INV_X1     g14201(.I(new_n15203_), .ZN(new_n15204_));
  INV_X1     g14202(.I(new_n15184_), .ZN(new_n15205_));
  NOR2_X1    g14203(.A1(new_n15205_), .A2(new_n15193_), .ZN(new_n15206_));
  NAND3_X1   g14204(.A1(new_n15206_), .A2(new_n15199_), .A3(new_n15204_), .ZN(new_n15207_));
  NAND2_X1   g14205(.A1(new_n15207_), .A2(new_n15194_), .ZN(new_n15208_));
  XOR2_X1    g14206(.A1(new_n15176_), .A2(new_n15208_), .Z(new_n15209_));
  INV_X1     g14207(.I(\A[686] ), .ZN(new_n15210_));
  NOR2_X1    g14208(.A1(new_n15210_), .A2(\A[685] ), .ZN(new_n15211_));
  NAND2_X1   g14209(.A1(new_n15210_), .A2(\A[685] ), .ZN(new_n15212_));
  NAND2_X1   g14210(.A1(new_n15212_), .A2(\A[687] ), .ZN(new_n15213_));
  INV_X1     g14211(.I(\A[685] ), .ZN(new_n15214_));
  NOR2_X1    g14212(.A1(new_n15214_), .A2(\A[686] ), .ZN(new_n15215_));
  NOR2_X1    g14213(.A1(new_n15211_), .A2(new_n15215_), .ZN(new_n15216_));
  OAI22_X1   g14214(.A1(new_n15216_), .A2(\A[687] ), .B1(new_n15213_), .B2(new_n15211_), .ZN(new_n15217_));
  INV_X1     g14215(.I(\A[690] ), .ZN(new_n15218_));
  INV_X1     g14216(.I(\A[688] ), .ZN(new_n15219_));
  NAND2_X1   g14217(.A1(new_n15219_), .A2(\A[689] ), .ZN(new_n15220_));
  NOR2_X1    g14218(.A1(new_n15219_), .A2(\A[689] ), .ZN(new_n15221_));
  NOR2_X1    g14219(.A1(new_n15221_), .A2(new_n15218_), .ZN(new_n15222_));
  INV_X1     g14220(.I(\A[689] ), .ZN(new_n15223_));
  NAND2_X1   g14221(.A1(new_n15223_), .A2(\A[688] ), .ZN(new_n15224_));
  NAND2_X1   g14222(.A1(new_n15220_), .A2(new_n15224_), .ZN(new_n15225_));
  AOI22_X1   g14223(.A1(new_n15225_), .A2(new_n15218_), .B1(new_n15222_), .B2(new_n15220_), .ZN(new_n15226_));
  XNOR2_X1   g14224(.A1(new_n15226_), .A2(new_n15217_), .ZN(new_n15227_));
  NOR2_X1    g14225(.A1(new_n15223_), .A2(\A[688] ), .ZN(new_n15228_));
  NOR2_X1    g14226(.A1(new_n15228_), .A2(new_n15221_), .ZN(new_n15229_));
  NOR2_X1    g14227(.A1(new_n15219_), .A2(new_n15223_), .ZN(new_n15230_));
  INV_X1     g14228(.I(new_n15230_), .ZN(new_n15231_));
  OAI21_X1   g14229(.A1(new_n15229_), .A2(new_n15218_), .B(new_n15231_), .ZN(new_n15232_));
  NAND2_X1   g14230(.A1(new_n15214_), .A2(\A[686] ), .ZN(new_n15233_));
  NAND2_X1   g14231(.A1(new_n15233_), .A2(new_n15212_), .ZN(new_n15234_));
  NOR2_X1    g14232(.A1(new_n15214_), .A2(new_n15210_), .ZN(new_n15235_));
  AOI21_X1   g14233(.A1(new_n15234_), .A2(\A[687] ), .B(new_n15235_), .ZN(new_n15236_));
  INV_X1     g14234(.I(new_n15236_), .ZN(new_n15237_));
  INV_X1     g14235(.I(new_n15217_), .ZN(new_n15238_));
  NOR2_X1    g14236(.A1(new_n15238_), .A2(new_n15226_), .ZN(new_n15239_));
  NAND3_X1   g14237(.A1(new_n15239_), .A2(new_n15232_), .A3(new_n15237_), .ZN(new_n15240_));
  NAND2_X1   g14238(.A1(new_n15240_), .A2(new_n15227_), .ZN(new_n15241_));
  INV_X1     g14239(.I(\A[681] ), .ZN(new_n15242_));
  INV_X1     g14240(.I(\A[679] ), .ZN(new_n15243_));
  NAND2_X1   g14241(.A1(new_n15243_), .A2(\A[680] ), .ZN(new_n15244_));
  NOR2_X1    g14242(.A1(new_n15243_), .A2(\A[680] ), .ZN(new_n15245_));
  NOR2_X1    g14243(.A1(new_n15245_), .A2(new_n15242_), .ZN(new_n15246_));
  INV_X1     g14244(.I(\A[680] ), .ZN(new_n15247_));
  NAND2_X1   g14245(.A1(new_n15247_), .A2(\A[679] ), .ZN(new_n15248_));
  NAND2_X1   g14246(.A1(new_n15244_), .A2(new_n15248_), .ZN(new_n15249_));
  AOI22_X1   g14247(.A1(new_n15249_), .A2(new_n15242_), .B1(new_n15246_), .B2(new_n15244_), .ZN(new_n15250_));
  INV_X1     g14248(.I(\A[684] ), .ZN(new_n15251_));
  INV_X1     g14249(.I(\A[682] ), .ZN(new_n15252_));
  NAND2_X1   g14250(.A1(new_n15252_), .A2(\A[683] ), .ZN(new_n15253_));
  NOR2_X1    g14251(.A1(new_n15252_), .A2(\A[683] ), .ZN(new_n15254_));
  NOR2_X1    g14252(.A1(new_n15254_), .A2(new_n15251_), .ZN(new_n15255_));
  INV_X1     g14253(.I(\A[683] ), .ZN(new_n15256_));
  NAND2_X1   g14254(.A1(new_n15256_), .A2(\A[682] ), .ZN(new_n15257_));
  NAND2_X1   g14255(.A1(new_n15253_), .A2(new_n15257_), .ZN(new_n15258_));
  AOI22_X1   g14256(.A1(new_n15258_), .A2(new_n15251_), .B1(new_n15255_), .B2(new_n15253_), .ZN(new_n15259_));
  XOR2_X1    g14257(.A1(new_n15250_), .A2(new_n15259_), .Z(new_n15260_));
  NOR2_X1    g14258(.A1(new_n15256_), .A2(\A[682] ), .ZN(new_n15261_));
  NOR2_X1    g14259(.A1(new_n15261_), .A2(new_n15254_), .ZN(new_n15262_));
  NOR2_X1    g14260(.A1(new_n15252_), .A2(new_n15256_), .ZN(new_n15263_));
  INV_X1     g14261(.I(new_n15263_), .ZN(new_n15264_));
  OAI21_X1   g14262(.A1(new_n15262_), .A2(new_n15251_), .B(new_n15264_), .ZN(new_n15265_));
  NOR2_X1    g14263(.A1(new_n15243_), .A2(new_n15247_), .ZN(new_n15266_));
  AOI21_X1   g14264(.A1(new_n15249_), .A2(\A[681] ), .B(new_n15266_), .ZN(new_n15267_));
  INV_X1     g14265(.I(new_n15267_), .ZN(new_n15268_));
  NOR2_X1    g14266(.A1(new_n15250_), .A2(new_n15259_), .ZN(new_n15269_));
  NAND3_X1   g14267(.A1(new_n15269_), .A2(new_n15265_), .A3(new_n15268_), .ZN(new_n15270_));
  NAND2_X1   g14268(.A1(new_n15260_), .A2(new_n15270_), .ZN(new_n15271_));
  XOR2_X1    g14269(.A1(new_n15241_), .A2(new_n15271_), .Z(new_n15272_));
  XOR2_X1    g14270(.A1(new_n15209_), .A2(new_n15272_), .Z(new_n15273_));
  INV_X1     g14271(.I(\A[674] ), .ZN(new_n15274_));
  NOR2_X1    g14272(.A1(new_n15274_), .A2(\A[673] ), .ZN(new_n15275_));
  NAND2_X1   g14273(.A1(new_n15274_), .A2(\A[673] ), .ZN(new_n15276_));
  NAND2_X1   g14274(.A1(new_n15276_), .A2(\A[675] ), .ZN(new_n15277_));
  INV_X1     g14275(.I(\A[673] ), .ZN(new_n15278_));
  NOR2_X1    g14276(.A1(new_n15278_), .A2(\A[674] ), .ZN(new_n15279_));
  NOR2_X1    g14277(.A1(new_n15275_), .A2(new_n15279_), .ZN(new_n15280_));
  OAI22_X1   g14278(.A1(new_n15280_), .A2(\A[675] ), .B1(new_n15277_), .B2(new_n15275_), .ZN(new_n15281_));
  INV_X1     g14279(.I(\A[678] ), .ZN(new_n15282_));
  INV_X1     g14280(.I(\A[676] ), .ZN(new_n15283_));
  NAND2_X1   g14281(.A1(new_n15283_), .A2(\A[677] ), .ZN(new_n15284_));
  NOR2_X1    g14282(.A1(new_n15283_), .A2(\A[677] ), .ZN(new_n15285_));
  NOR2_X1    g14283(.A1(new_n15285_), .A2(new_n15282_), .ZN(new_n15286_));
  INV_X1     g14284(.I(\A[677] ), .ZN(new_n15287_));
  NAND2_X1   g14285(.A1(new_n15287_), .A2(\A[676] ), .ZN(new_n15288_));
  NAND2_X1   g14286(.A1(new_n15284_), .A2(new_n15288_), .ZN(new_n15289_));
  AOI22_X1   g14287(.A1(new_n15289_), .A2(new_n15282_), .B1(new_n15286_), .B2(new_n15284_), .ZN(new_n15290_));
  XNOR2_X1   g14288(.A1(new_n15290_), .A2(new_n15281_), .ZN(new_n15291_));
  NOR2_X1    g14289(.A1(new_n15287_), .A2(\A[676] ), .ZN(new_n15292_));
  NOR2_X1    g14290(.A1(new_n15292_), .A2(new_n15285_), .ZN(new_n15293_));
  NOR2_X1    g14291(.A1(new_n15283_), .A2(new_n15287_), .ZN(new_n15294_));
  INV_X1     g14292(.I(new_n15294_), .ZN(new_n15295_));
  OAI21_X1   g14293(.A1(new_n15293_), .A2(new_n15282_), .B(new_n15295_), .ZN(new_n15296_));
  NAND2_X1   g14294(.A1(new_n15278_), .A2(\A[674] ), .ZN(new_n15297_));
  NAND2_X1   g14295(.A1(new_n15297_), .A2(new_n15276_), .ZN(new_n15298_));
  NOR2_X1    g14296(.A1(new_n15278_), .A2(new_n15274_), .ZN(new_n15299_));
  AOI21_X1   g14297(.A1(new_n15298_), .A2(\A[675] ), .B(new_n15299_), .ZN(new_n15300_));
  INV_X1     g14298(.I(new_n15300_), .ZN(new_n15301_));
  INV_X1     g14299(.I(new_n15281_), .ZN(new_n15302_));
  NOR2_X1    g14300(.A1(new_n15302_), .A2(new_n15290_), .ZN(new_n15303_));
  NAND3_X1   g14301(.A1(new_n15303_), .A2(new_n15296_), .A3(new_n15301_), .ZN(new_n15304_));
  NAND2_X1   g14302(.A1(new_n15304_), .A2(new_n15291_), .ZN(new_n15305_));
  INV_X1     g14303(.I(\A[668] ), .ZN(new_n15306_));
  NOR2_X1    g14304(.A1(new_n15306_), .A2(\A[667] ), .ZN(new_n15307_));
  NAND2_X1   g14305(.A1(new_n15306_), .A2(\A[667] ), .ZN(new_n15308_));
  NAND2_X1   g14306(.A1(new_n15308_), .A2(\A[669] ), .ZN(new_n15309_));
  INV_X1     g14307(.I(\A[667] ), .ZN(new_n15310_));
  NOR2_X1    g14308(.A1(new_n15310_), .A2(\A[668] ), .ZN(new_n15311_));
  NOR2_X1    g14309(.A1(new_n15307_), .A2(new_n15311_), .ZN(new_n15312_));
  OAI22_X1   g14310(.A1(new_n15312_), .A2(\A[669] ), .B1(new_n15309_), .B2(new_n15307_), .ZN(new_n15313_));
  INV_X1     g14311(.I(\A[672] ), .ZN(new_n15314_));
  INV_X1     g14312(.I(\A[670] ), .ZN(new_n15315_));
  NAND2_X1   g14313(.A1(new_n15315_), .A2(\A[671] ), .ZN(new_n15316_));
  NOR2_X1    g14314(.A1(new_n15315_), .A2(\A[671] ), .ZN(new_n15317_));
  NOR2_X1    g14315(.A1(new_n15317_), .A2(new_n15314_), .ZN(new_n15318_));
  INV_X1     g14316(.I(\A[671] ), .ZN(new_n15319_));
  NAND2_X1   g14317(.A1(new_n15319_), .A2(\A[670] ), .ZN(new_n15320_));
  NAND2_X1   g14318(.A1(new_n15316_), .A2(new_n15320_), .ZN(new_n15321_));
  AOI22_X1   g14319(.A1(new_n15321_), .A2(new_n15314_), .B1(new_n15318_), .B2(new_n15316_), .ZN(new_n15322_));
  XNOR2_X1   g14320(.A1(new_n15322_), .A2(new_n15313_), .ZN(new_n15323_));
  NOR2_X1    g14321(.A1(new_n15319_), .A2(\A[670] ), .ZN(new_n15324_));
  NOR2_X1    g14322(.A1(new_n15324_), .A2(new_n15317_), .ZN(new_n15325_));
  NOR2_X1    g14323(.A1(new_n15315_), .A2(new_n15319_), .ZN(new_n15326_));
  INV_X1     g14324(.I(new_n15326_), .ZN(new_n15327_));
  OAI21_X1   g14325(.A1(new_n15325_), .A2(new_n15314_), .B(new_n15327_), .ZN(new_n15328_));
  NAND2_X1   g14326(.A1(new_n15310_), .A2(\A[668] ), .ZN(new_n15329_));
  NAND2_X1   g14327(.A1(new_n15329_), .A2(new_n15308_), .ZN(new_n15330_));
  NOR2_X1    g14328(.A1(new_n15310_), .A2(new_n15306_), .ZN(new_n15331_));
  AOI21_X1   g14329(.A1(new_n15330_), .A2(\A[669] ), .B(new_n15331_), .ZN(new_n15332_));
  INV_X1     g14330(.I(new_n15332_), .ZN(new_n15333_));
  INV_X1     g14331(.I(new_n15313_), .ZN(new_n15334_));
  NOR2_X1    g14332(.A1(new_n15334_), .A2(new_n15322_), .ZN(new_n15335_));
  NAND3_X1   g14333(.A1(new_n15335_), .A2(new_n15328_), .A3(new_n15333_), .ZN(new_n15336_));
  NAND2_X1   g14334(.A1(new_n15336_), .A2(new_n15323_), .ZN(new_n15337_));
  XNOR2_X1   g14335(.A1(new_n15305_), .A2(new_n15337_), .ZN(new_n15338_));
  INV_X1     g14336(.I(\A[662] ), .ZN(new_n15339_));
  NOR2_X1    g14337(.A1(new_n15339_), .A2(\A[661] ), .ZN(new_n15340_));
  NAND2_X1   g14338(.A1(new_n15339_), .A2(\A[661] ), .ZN(new_n15341_));
  NAND2_X1   g14339(.A1(new_n15341_), .A2(\A[663] ), .ZN(new_n15342_));
  INV_X1     g14340(.I(\A[661] ), .ZN(new_n15343_));
  NOR2_X1    g14341(.A1(new_n15343_), .A2(\A[662] ), .ZN(new_n15344_));
  NOR2_X1    g14342(.A1(new_n15340_), .A2(new_n15344_), .ZN(new_n15345_));
  OAI22_X1   g14343(.A1(new_n15345_), .A2(\A[663] ), .B1(new_n15342_), .B2(new_n15340_), .ZN(new_n15346_));
  INV_X1     g14344(.I(\A[666] ), .ZN(new_n15347_));
  INV_X1     g14345(.I(\A[664] ), .ZN(new_n15348_));
  NAND2_X1   g14346(.A1(new_n15348_), .A2(\A[665] ), .ZN(new_n15349_));
  NOR2_X1    g14347(.A1(new_n15348_), .A2(\A[665] ), .ZN(new_n15350_));
  NOR2_X1    g14348(.A1(new_n15350_), .A2(new_n15347_), .ZN(new_n15351_));
  INV_X1     g14349(.I(\A[665] ), .ZN(new_n15352_));
  NAND2_X1   g14350(.A1(new_n15352_), .A2(\A[664] ), .ZN(new_n15353_));
  NAND2_X1   g14351(.A1(new_n15349_), .A2(new_n15353_), .ZN(new_n15354_));
  AOI22_X1   g14352(.A1(new_n15354_), .A2(new_n15347_), .B1(new_n15351_), .B2(new_n15349_), .ZN(new_n15355_));
  XNOR2_X1   g14353(.A1(new_n15355_), .A2(new_n15346_), .ZN(new_n15356_));
  NOR2_X1    g14354(.A1(new_n15352_), .A2(\A[664] ), .ZN(new_n15357_));
  NOR2_X1    g14355(.A1(new_n15357_), .A2(new_n15350_), .ZN(new_n15358_));
  NOR2_X1    g14356(.A1(new_n15348_), .A2(new_n15352_), .ZN(new_n15359_));
  INV_X1     g14357(.I(new_n15359_), .ZN(new_n15360_));
  OAI21_X1   g14358(.A1(new_n15358_), .A2(new_n15347_), .B(new_n15360_), .ZN(new_n15361_));
  NAND2_X1   g14359(.A1(new_n15343_), .A2(\A[662] ), .ZN(new_n15362_));
  NAND2_X1   g14360(.A1(new_n15362_), .A2(new_n15341_), .ZN(new_n15363_));
  NOR2_X1    g14361(.A1(new_n15343_), .A2(new_n15339_), .ZN(new_n15364_));
  AOI21_X1   g14362(.A1(new_n15363_), .A2(\A[663] ), .B(new_n15364_), .ZN(new_n15365_));
  INV_X1     g14363(.I(new_n15365_), .ZN(new_n15366_));
  INV_X1     g14364(.I(new_n15346_), .ZN(new_n15367_));
  NOR2_X1    g14365(.A1(new_n15367_), .A2(new_n15355_), .ZN(new_n15368_));
  NAND3_X1   g14366(.A1(new_n15368_), .A2(new_n15361_), .A3(new_n15366_), .ZN(new_n15369_));
  NAND2_X1   g14367(.A1(new_n15369_), .A2(new_n15356_), .ZN(new_n15370_));
  INV_X1     g14368(.I(\A[656] ), .ZN(new_n15371_));
  NOR2_X1    g14369(.A1(new_n15371_), .A2(\A[655] ), .ZN(new_n15372_));
  NAND2_X1   g14370(.A1(new_n15371_), .A2(\A[655] ), .ZN(new_n15373_));
  NAND2_X1   g14371(.A1(new_n15373_), .A2(\A[657] ), .ZN(new_n15374_));
  INV_X1     g14372(.I(\A[655] ), .ZN(new_n15375_));
  NOR2_X1    g14373(.A1(new_n15375_), .A2(\A[656] ), .ZN(new_n15376_));
  NOR2_X1    g14374(.A1(new_n15372_), .A2(new_n15376_), .ZN(new_n15377_));
  OAI22_X1   g14375(.A1(new_n15377_), .A2(\A[657] ), .B1(new_n15374_), .B2(new_n15372_), .ZN(new_n15378_));
  INV_X1     g14376(.I(\A[660] ), .ZN(new_n15379_));
  INV_X1     g14377(.I(\A[658] ), .ZN(new_n15380_));
  NAND2_X1   g14378(.A1(new_n15380_), .A2(\A[659] ), .ZN(new_n15381_));
  NOR2_X1    g14379(.A1(new_n15380_), .A2(\A[659] ), .ZN(new_n15382_));
  NOR2_X1    g14380(.A1(new_n15382_), .A2(new_n15379_), .ZN(new_n15383_));
  INV_X1     g14381(.I(\A[659] ), .ZN(new_n15384_));
  NAND2_X1   g14382(.A1(new_n15384_), .A2(\A[658] ), .ZN(new_n15385_));
  NAND2_X1   g14383(.A1(new_n15381_), .A2(new_n15385_), .ZN(new_n15386_));
  AOI22_X1   g14384(.A1(new_n15386_), .A2(new_n15379_), .B1(new_n15383_), .B2(new_n15381_), .ZN(new_n15387_));
  XNOR2_X1   g14385(.A1(new_n15387_), .A2(new_n15378_), .ZN(new_n15388_));
  NOR2_X1    g14386(.A1(new_n15384_), .A2(\A[658] ), .ZN(new_n15389_));
  NOR2_X1    g14387(.A1(new_n15389_), .A2(new_n15382_), .ZN(new_n15390_));
  NOR2_X1    g14388(.A1(new_n15380_), .A2(new_n15384_), .ZN(new_n15391_));
  INV_X1     g14389(.I(new_n15391_), .ZN(new_n15392_));
  OAI21_X1   g14390(.A1(new_n15390_), .A2(new_n15379_), .B(new_n15392_), .ZN(new_n15393_));
  NAND2_X1   g14391(.A1(new_n15375_), .A2(\A[656] ), .ZN(new_n15394_));
  NAND2_X1   g14392(.A1(new_n15394_), .A2(new_n15373_), .ZN(new_n15395_));
  NOR2_X1    g14393(.A1(new_n15375_), .A2(new_n15371_), .ZN(new_n15396_));
  AOI21_X1   g14394(.A1(new_n15395_), .A2(\A[657] ), .B(new_n15396_), .ZN(new_n15397_));
  INV_X1     g14395(.I(new_n15397_), .ZN(new_n15398_));
  INV_X1     g14396(.I(new_n15378_), .ZN(new_n15399_));
  NOR2_X1    g14397(.A1(new_n15399_), .A2(new_n15387_), .ZN(new_n15400_));
  NAND3_X1   g14398(.A1(new_n15400_), .A2(new_n15393_), .A3(new_n15398_), .ZN(new_n15401_));
  NAND2_X1   g14399(.A1(new_n15401_), .A2(new_n15388_), .ZN(new_n15402_));
  XOR2_X1    g14400(.A1(new_n15370_), .A2(new_n15402_), .Z(new_n15403_));
  XOR2_X1    g14401(.A1(new_n15338_), .A2(new_n15403_), .Z(new_n15404_));
  XOR2_X1    g14402(.A1(new_n15404_), .A2(new_n15273_), .Z(new_n15405_));
  XOR2_X1    g14403(.A1(new_n15144_), .A2(new_n15405_), .Z(new_n15406_));
  NAND2_X1   g14404(.A1(new_n15406_), .A2(new_n14914_), .ZN(new_n15407_));
  INV_X1     g14405(.I(new_n15407_), .ZN(new_n15408_));
  XOR2_X1    g14406(.A1(new_n14665_), .A2(new_n14669_), .Z(new_n15409_));
  NAND2_X1   g14407(.A1(new_n15409_), .A2(new_n14672_), .ZN(new_n15410_));
  AOI21_X1   g14408(.A1(new_n14658_), .A2(\A[756] ), .B(new_n14663_), .ZN(new_n15411_));
  XOR2_X1    g14409(.A1(new_n15411_), .A2(new_n14669_), .Z(new_n15412_));
  INV_X1     g14410(.I(new_n14659_), .ZN(new_n15413_));
  NAND2_X1   g14411(.A1(new_n15413_), .A2(new_n14650_), .ZN(new_n15414_));
  NAND2_X1   g14412(.A1(new_n15412_), .A2(new_n15414_), .ZN(new_n15415_));
  NAND2_X1   g14413(.A1(new_n15410_), .A2(new_n15415_), .ZN(new_n15416_));
  NAND2_X1   g14414(.A1(new_n14670_), .A2(new_n14665_), .ZN(new_n15417_));
  OAI21_X1   g14415(.A1(new_n15409_), .A2(new_n15414_), .B(new_n15417_), .ZN(new_n15418_));
  NAND2_X1   g14416(.A1(new_n15418_), .A2(new_n14660_), .ZN(new_n15419_));
  NAND2_X1   g14417(.A1(new_n15419_), .A2(new_n15416_), .ZN(new_n15420_));
  INV_X1     g14418(.I(new_n15420_), .ZN(new_n15421_));
  XOR2_X1    g14419(.A1(new_n14633_), .A2(new_n14637_), .Z(new_n15422_));
  NAND2_X1   g14420(.A1(new_n15422_), .A2(new_n14640_), .ZN(new_n15423_));
  AOI21_X1   g14421(.A1(new_n14626_), .A2(\A[762] ), .B(new_n14631_), .ZN(new_n15424_));
  XOR2_X1    g14422(.A1(new_n15424_), .A2(new_n14637_), .Z(new_n15425_));
  INV_X1     g14423(.I(new_n14627_), .ZN(new_n15426_));
  NAND2_X1   g14424(.A1(new_n15426_), .A2(new_n14618_), .ZN(new_n15427_));
  NAND2_X1   g14425(.A1(new_n15425_), .A2(new_n15427_), .ZN(new_n15428_));
  NAND2_X1   g14426(.A1(new_n15423_), .A2(new_n15428_), .ZN(new_n15429_));
  XOR2_X1    g14427(.A1(new_n14627_), .A2(new_n14618_), .Z(new_n15430_));
  XOR2_X1    g14428(.A1(new_n14659_), .A2(new_n14650_), .Z(new_n15431_));
  NOR2_X1    g14429(.A1(new_n15430_), .A2(new_n15431_), .ZN(new_n15432_));
  NAND3_X1   g14430(.A1(new_n15429_), .A2(new_n14641_), .A3(new_n15432_), .ZN(new_n15433_));
  NOR2_X1    g14431(.A1(new_n15424_), .A2(new_n14637_), .ZN(new_n15434_));
  INV_X1     g14432(.I(new_n15434_), .ZN(new_n15435_));
  OAI21_X1   g14433(.A1(new_n15422_), .A2(new_n15427_), .B(new_n15435_), .ZN(new_n15436_));
  NAND2_X1   g14434(.A1(new_n15436_), .A2(new_n14628_), .ZN(new_n15437_));
  NAND2_X1   g14435(.A1(new_n15437_), .A2(new_n14673_), .ZN(new_n15438_));
  NOR2_X1    g14436(.A1(new_n15433_), .A2(new_n15438_), .ZN(new_n15439_));
  NAND3_X1   g14437(.A1(new_n15432_), .A2(new_n14641_), .A3(new_n14673_), .ZN(new_n15440_));
  NAND2_X1   g14438(.A1(new_n15437_), .A2(new_n15429_), .ZN(new_n15441_));
  NAND2_X1   g14439(.A1(new_n15441_), .A2(new_n15440_), .ZN(new_n15442_));
  INV_X1     g14440(.I(new_n15442_), .ZN(new_n15443_));
  OAI21_X1   g14441(.A1(new_n15443_), .A2(new_n15439_), .B(new_n15421_), .ZN(new_n15444_));
  INV_X1     g14442(.I(new_n14641_), .ZN(new_n15445_));
  INV_X1     g14443(.I(new_n14673_), .ZN(new_n15446_));
  NAND2_X1   g14444(.A1(new_n14628_), .A2(new_n14660_), .ZN(new_n15447_));
  NOR3_X1    g14445(.A1(new_n15447_), .A2(new_n15445_), .A3(new_n15446_), .ZN(new_n15448_));
  NOR2_X1    g14446(.A1(new_n15441_), .A2(new_n15448_), .ZN(new_n15449_));
  AOI21_X1   g14447(.A1(new_n15429_), .A2(new_n15437_), .B(new_n15440_), .ZN(new_n15450_));
  OAI21_X1   g14448(.A1(new_n15449_), .A2(new_n15450_), .B(new_n15420_), .ZN(new_n15451_));
  NAND2_X1   g14449(.A1(new_n15444_), .A2(new_n15451_), .ZN(new_n15452_));
  XOR2_X1    g14450(.A1(new_n14594_), .A2(new_n14585_), .Z(new_n15453_));
  AOI21_X1   g14451(.A1(new_n14593_), .A2(\A[768] ), .B(new_n14598_), .ZN(new_n15454_));
  XOR2_X1    g14452(.A1(new_n15454_), .A2(new_n14604_), .Z(new_n15455_));
  NOR2_X1    g14453(.A1(new_n15454_), .A2(new_n14604_), .ZN(new_n15456_));
  AOI21_X1   g14454(.A1(new_n15455_), .A2(new_n14607_), .B(new_n15456_), .ZN(new_n15457_));
  INV_X1     g14455(.I(new_n14594_), .ZN(new_n15458_));
  NAND2_X1   g14456(.A1(new_n15458_), .A2(new_n14585_), .ZN(new_n15459_));
  NOR2_X1    g14457(.A1(new_n15455_), .A2(new_n15459_), .ZN(new_n15460_));
  XOR2_X1    g14458(.A1(new_n14600_), .A2(new_n14604_), .Z(new_n15461_));
  NOR2_X1    g14459(.A1(new_n15461_), .A2(new_n14607_), .ZN(new_n15462_));
  OAI22_X1   g14460(.A1(new_n15453_), .A2(new_n15457_), .B1(new_n15460_), .B2(new_n15462_), .ZN(new_n15463_));
  XOR2_X1    g14461(.A1(new_n14562_), .A2(new_n14553_), .Z(new_n15464_));
  AOI21_X1   g14462(.A1(new_n14561_), .A2(\A[774] ), .B(new_n14566_), .ZN(new_n15465_));
  XOR2_X1    g14463(.A1(new_n15465_), .A2(new_n14572_), .Z(new_n15466_));
  INV_X1     g14464(.I(new_n14562_), .ZN(new_n15467_));
  NAND2_X1   g14465(.A1(new_n15467_), .A2(new_n14553_), .ZN(new_n15468_));
  NOR2_X1    g14466(.A1(new_n15466_), .A2(new_n15468_), .ZN(new_n15469_));
  XOR2_X1    g14467(.A1(new_n14568_), .A2(new_n14572_), .Z(new_n15470_));
  NOR2_X1    g14468(.A1(new_n15470_), .A2(new_n14575_), .ZN(new_n15471_));
  NOR2_X1    g14469(.A1(new_n15471_), .A2(new_n15469_), .ZN(new_n15472_));
  NOR3_X1    g14470(.A1(new_n15472_), .A2(new_n15464_), .A3(new_n15453_), .ZN(new_n15473_));
  NOR2_X1    g14471(.A1(new_n15465_), .A2(new_n14572_), .ZN(new_n15474_));
  INV_X1     g14472(.I(new_n15474_), .ZN(new_n15475_));
  OAI21_X1   g14473(.A1(new_n15470_), .A2(new_n15468_), .B(new_n15475_), .ZN(new_n15476_));
  NAND2_X1   g14474(.A1(new_n15476_), .A2(new_n14563_), .ZN(new_n15477_));
  NAND4_X1   g14475(.A1(new_n15473_), .A2(new_n14576_), .A3(new_n14608_), .A4(new_n15477_), .ZN(new_n15478_));
  NOR2_X1    g14476(.A1(new_n15464_), .A2(new_n15453_), .ZN(new_n15479_));
  NAND3_X1   g14477(.A1(new_n15479_), .A2(new_n14576_), .A3(new_n14608_), .ZN(new_n15480_));
  NAND2_X1   g14478(.A1(new_n15470_), .A2(new_n14575_), .ZN(new_n15481_));
  NAND2_X1   g14479(.A1(new_n15466_), .A2(new_n15468_), .ZN(new_n15482_));
  NAND2_X1   g14480(.A1(new_n15481_), .A2(new_n15482_), .ZN(new_n15483_));
  NAND2_X1   g14481(.A1(new_n15477_), .A2(new_n15483_), .ZN(new_n15484_));
  NAND2_X1   g14482(.A1(new_n15484_), .A2(new_n15480_), .ZN(new_n15485_));
  AOI21_X1   g14483(.A1(new_n15478_), .A2(new_n15485_), .B(new_n15463_), .ZN(new_n15486_));
  INV_X1     g14484(.I(new_n15457_), .ZN(new_n15487_));
  NAND2_X1   g14485(.A1(new_n15461_), .A2(new_n14607_), .ZN(new_n15488_));
  NAND2_X1   g14486(.A1(new_n15455_), .A2(new_n15459_), .ZN(new_n15489_));
  AOI22_X1   g14487(.A1(new_n15487_), .A2(new_n14595_), .B1(new_n15488_), .B2(new_n15489_), .ZN(new_n15490_));
  AND4_X2    g14488(.A1(new_n14563_), .A2(new_n14576_), .A3(new_n14608_), .A4(new_n14595_), .Z(new_n15491_));
  NAND2_X1   g14489(.A1(new_n15484_), .A2(new_n15491_), .ZN(new_n15492_));
  AOI22_X1   g14490(.A1(new_n15476_), .A2(new_n14563_), .B1(new_n15481_), .B2(new_n15482_), .ZN(new_n15493_));
  NAND2_X1   g14491(.A1(new_n15493_), .A2(new_n15480_), .ZN(new_n15494_));
  AOI21_X1   g14492(.A1(new_n15492_), .A2(new_n15494_), .B(new_n15490_), .ZN(new_n15495_));
  NAND2_X1   g14493(.A1(new_n14610_), .A2(new_n14675_), .ZN(new_n15496_));
  NOR3_X1    g14494(.A1(new_n15486_), .A2(new_n15495_), .A3(new_n15496_), .ZN(new_n15497_));
  NAND3_X1   g14495(.A1(new_n15483_), .A2(new_n14576_), .A3(new_n15479_), .ZN(new_n15498_));
  NAND2_X1   g14496(.A1(new_n15477_), .A2(new_n14608_), .ZN(new_n15499_));
  NOR2_X1    g14497(.A1(new_n15498_), .A2(new_n15499_), .ZN(new_n15500_));
  NOR2_X1    g14498(.A1(new_n15493_), .A2(new_n15491_), .ZN(new_n15501_));
  OAI21_X1   g14499(.A1(new_n15500_), .A2(new_n15501_), .B(new_n15490_), .ZN(new_n15502_));
  NOR2_X1    g14500(.A1(new_n15493_), .A2(new_n15480_), .ZN(new_n15503_));
  NOR2_X1    g14501(.A1(new_n15484_), .A2(new_n15491_), .ZN(new_n15504_));
  OAI21_X1   g14502(.A1(new_n15504_), .A2(new_n15503_), .B(new_n15463_), .ZN(new_n15505_));
  XNOR2_X1   g14503(.A1(new_n14577_), .A2(new_n14609_), .ZN(new_n15506_));
  XNOR2_X1   g14504(.A1(new_n14642_), .A2(new_n14674_), .ZN(new_n15507_));
  NOR2_X1    g14505(.A1(new_n15506_), .A2(new_n15507_), .ZN(new_n15508_));
  AOI21_X1   g14506(.A1(new_n15502_), .A2(new_n15505_), .B(new_n15508_), .ZN(new_n15509_));
  NOR2_X1    g14507(.A1(new_n15497_), .A2(new_n15509_), .ZN(new_n15510_));
  NOR2_X1    g14508(.A1(new_n15510_), .A2(new_n15452_), .ZN(new_n15511_));
  NOR2_X1    g14509(.A1(new_n15425_), .A2(new_n15427_), .ZN(new_n15512_));
  NOR2_X1    g14510(.A1(new_n15422_), .A2(new_n14640_), .ZN(new_n15513_));
  NOR2_X1    g14511(.A1(new_n15513_), .A2(new_n15512_), .ZN(new_n15514_));
  NOR3_X1    g14512(.A1(new_n15514_), .A2(new_n15445_), .A3(new_n15447_), .ZN(new_n15515_));
  AOI21_X1   g14513(.A1(new_n15425_), .A2(new_n14640_), .B(new_n15434_), .ZN(new_n15516_));
  NOR2_X1    g14514(.A1(new_n15516_), .A2(new_n15430_), .ZN(new_n15517_));
  NOR2_X1    g14515(.A1(new_n15517_), .A2(new_n15446_), .ZN(new_n15518_));
  NAND2_X1   g14516(.A1(new_n15515_), .A2(new_n15518_), .ZN(new_n15519_));
  AOI21_X1   g14517(.A1(new_n15519_), .A2(new_n15442_), .B(new_n15420_), .ZN(new_n15520_));
  OR2_X2     g14518(.A1(new_n15449_), .A2(new_n15450_), .Z(new_n15521_));
  AOI21_X1   g14519(.A1(new_n15521_), .A2(new_n15420_), .B(new_n15520_), .ZN(new_n15522_));
  NAND3_X1   g14520(.A1(new_n15502_), .A2(new_n15505_), .A3(new_n15496_), .ZN(new_n15523_));
  OAI21_X1   g14521(.A1(new_n15486_), .A2(new_n15495_), .B(new_n15508_), .ZN(new_n15524_));
  AOI21_X1   g14522(.A1(new_n15523_), .A2(new_n15524_), .B(new_n15522_), .ZN(new_n15525_));
  NOR2_X1    g14523(.A1(new_n15511_), .A2(new_n15525_), .ZN(new_n15526_));
  NAND2_X1   g14524(.A1(new_n14676_), .A2(new_n14545_), .ZN(new_n15527_));
  INV_X1     g14525(.I(new_n15527_), .ZN(new_n15528_));
  XOR2_X1    g14526(.A1(new_n14523_), .A2(new_n14531_), .Z(new_n15529_));
  NAND2_X1   g14527(.A1(new_n14518_), .A2(\A[776] ), .ZN(new_n15530_));
  NAND2_X1   g14528(.A1(new_n14521_), .A2(new_n15530_), .ZN(new_n15531_));
  AOI21_X1   g14529(.A1(new_n15531_), .A2(\A[777] ), .B(new_n14537_), .ZN(new_n15532_));
  XOR2_X1    g14530(.A1(new_n14534_), .A2(new_n15532_), .Z(new_n15533_));
  NOR2_X1    g14531(.A1(new_n14534_), .A2(new_n15532_), .ZN(new_n15534_));
  AOI21_X1   g14532(.A1(new_n15533_), .A2(new_n14541_), .B(new_n15534_), .ZN(new_n15535_));
  XOR2_X1    g14533(.A1(new_n14539_), .A2(new_n14534_), .Z(new_n15536_));
  NAND2_X1   g14534(.A1(new_n15536_), .A2(new_n14541_), .ZN(new_n15537_));
  INV_X1     g14535(.I(new_n14531_), .ZN(new_n15538_));
  NAND2_X1   g14536(.A1(new_n15538_), .A2(new_n14523_), .ZN(new_n15539_));
  NAND2_X1   g14537(.A1(new_n15533_), .A2(new_n15539_), .ZN(new_n15540_));
  NAND2_X1   g14538(.A1(new_n15537_), .A2(new_n15540_), .ZN(new_n15541_));
  OAI21_X1   g14539(.A1(new_n15529_), .A2(new_n15535_), .B(new_n15541_), .ZN(new_n15542_));
  XNOR2_X1   g14540(.A1(new_n14508_), .A2(new_n14511_), .ZN(new_n15543_));
  NOR2_X1    g14541(.A1(new_n15543_), .A2(new_n15529_), .ZN(new_n15544_));
  NAND3_X1   g14542(.A1(new_n15544_), .A2(new_n14513_), .A3(new_n14542_), .ZN(new_n15545_));
  INV_X1     g14543(.I(new_n15545_), .ZN(new_n15546_));
  NOR2_X1    g14544(.A1(new_n14496_), .A2(new_n14504_), .ZN(new_n15547_));
  XOR2_X1    g14545(.A1(new_n14496_), .A2(new_n14504_), .Z(new_n15548_));
  AOI21_X1   g14546(.A1(new_n15548_), .A2(new_n14512_), .B(new_n15547_), .ZN(new_n15549_));
  XNOR2_X1   g14547(.A1(new_n14496_), .A2(new_n14504_), .ZN(new_n15550_));
  NOR2_X1    g14548(.A1(new_n15550_), .A2(new_n14512_), .ZN(new_n15551_));
  INV_X1     g14549(.I(new_n14512_), .ZN(new_n15552_));
  NOR2_X1    g14550(.A1(new_n15548_), .A2(new_n15552_), .ZN(new_n15553_));
  OAI22_X1   g14551(.A1(new_n15549_), .A2(new_n15543_), .B1(new_n15551_), .B2(new_n15553_), .ZN(new_n15554_));
  NOR2_X1    g14552(.A1(new_n15546_), .A2(new_n15554_), .ZN(new_n15555_));
  INV_X1     g14553(.I(new_n15554_), .ZN(new_n15556_));
  NOR2_X1    g14554(.A1(new_n15556_), .A2(new_n15545_), .ZN(new_n15557_));
  OAI21_X1   g14555(.A1(new_n15557_), .A2(new_n15555_), .B(new_n15542_), .ZN(new_n15558_));
  INV_X1     g14556(.I(new_n15535_), .ZN(new_n15559_));
  NOR2_X1    g14557(.A1(new_n15533_), .A2(new_n15539_), .ZN(new_n15560_));
  NOR2_X1    g14558(.A1(new_n15536_), .A2(new_n14541_), .ZN(new_n15561_));
  NOR2_X1    g14559(.A1(new_n15561_), .A2(new_n15560_), .ZN(new_n15562_));
  AOI21_X1   g14560(.A1(new_n14532_), .A2(new_n15559_), .B(new_n15562_), .ZN(new_n15563_));
  INV_X1     g14561(.I(new_n14542_), .ZN(new_n15564_));
  NOR2_X1    g14562(.A1(new_n15549_), .A2(new_n15543_), .ZN(new_n15565_));
  NAND2_X1   g14563(.A1(new_n15548_), .A2(new_n15552_), .ZN(new_n15566_));
  NAND2_X1   g14564(.A1(new_n15550_), .A2(new_n14512_), .ZN(new_n15567_));
  NAND2_X1   g14565(.A1(new_n15567_), .A2(new_n15566_), .ZN(new_n15568_));
  NAND3_X1   g14566(.A1(new_n15568_), .A2(new_n14513_), .A3(new_n15544_), .ZN(new_n15569_));
  NOR3_X1    g14567(.A1(new_n15569_), .A2(new_n15564_), .A3(new_n15565_), .ZN(new_n15570_));
  NAND2_X1   g14568(.A1(new_n15554_), .A2(new_n15545_), .ZN(new_n15571_));
  INV_X1     g14569(.I(new_n15571_), .ZN(new_n15572_));
  OAI21_X1   g14570(.A1(new_n15572_), .A2(new_n15570_), .B(new_n15563_), .ZN(new_n15573_));
  NAND2_X1   g14571(.A1(new_n15573_), .A2(new_n15558_), .ZN(new_n15574_));
  AOI21_X1   g14572(.A1(new_n14473_), .A2(\A[792] ), .B(new_n14477_), .ZN(new_n15575_));
  XOR2_X1    g14573(.A1(new_n14484_), .A2(new_n15575_), .Z(new_n15576_));
  INV_X1     g14574(.I(new_n14475_), .ZN(new_n15577_));
  NAND2_X1   g14575(.A1(new_n15577_), .A2(new_n14467_), .ZN(new_n15578_));
  NAND2_X1   g14576(.A1(new_n14462_), .A2(\A[788] ), .ZN(new_n15579_));
  NAND2_X1   g14577(.A1(new_n14465_), .A2(new_n15579_), .ZN(new_n15580_));
  AOI21_X1   g14578(.A1(new_n15580_), .A2(\A[789] ), .B(new_n14482_), .ZN(new_n15581_));
  NOR2_X1    g14579(.A1(new_n15575_), .A2(new_n15581_), .ZN(new_n15582_));
  INV_X1     g14580(.I(new_n15582_), .ZN(new_n15583_));
  OAI21_X1   g14581(.A1(new_n15576_), .A2(new_n15578_), .B(new_n15583_), .ZN(new_n15584_));
  NAND2_X1   g14582(.A1(new_n15576_), .A2(new_n14486_), .ZN(new_n15585_));
  XOR2_X1    g14583(.A1(new_n15575_), .A2(new_n15581_), .Z(new_n15586_));
  NAND2_X1   g14584(.A1(new_n15586_), .A2(new_n15578_), .ZN(new_n15587_));
  AOI22_X1   g14585(.A1(new_n15584_), .A2(new_n14476_), .B1(new_n15585_), .B2(new_n15587_), .ZN(new_n15588_));
  NAND2_X1   g14586(.A1(new_n14433_), .A2(\A[797] ), .ZN(new_n15589_));
  NAND2_X1   g14587(.A1(new_n14453_), .A2(new_n15589_), .ZN(new_n15590_));
  AOI21_X1   g14588(.A1(new_n15590_), .A2(\A[798] ), .B(new_n14435_), .ZN(new_n15591_));
  NAND2_X1   g14589(.A1(new_n14442_), .A2(\A[794] ), .ZN(new_n15592_));
  NAND2_X1   g14590(.A1(new_n14450_), .A2(new_n15592_), .ZN(new_n15593_));
  AOI21_X1   g14591(.A1(new_n15593_), .A2(\A[795] ), .B(new_n14444_), .ZN(new_n15594_));
  NAND2_X1   g14592(.A1(new_n14452_), .A2(new_n14455_), .ZN(new_n15595_));
  NOR3_X1    g14593(.A1(new_n15595_), .A2(new_n15591_), .A3(new_n15594_), .ZN(new_n15596_));
  INV_X1     g14594(.I(new_n14487_), .ZN(new_n15597_));
  NAND2_X1   g14595(.A1(new_n14440_), .A2(new_n15594_), .ZN(new_n15598_));
  NAND2_X1   g14596(.A1(new_n14449_), .A2(new_n15591_), .ZN(new_n15599_));
  NAND2_X1   g14597(.A1(new_n15598_), .A2(new_n15599_), .ZN(new_n15600_));
  NAND2_X1   g14598(.A1(new_n15600_), .A2(new_n15595_), .ZN(new_n15601_));
  NAND3_X1   g14599(.A1(new_n14456_), .A2(new_n15598_), .A3(new_n15599_), .ZN(new_n15602_));
  NAND2_X1   g14600(.A1(new_n15601_), .A2(new_n15602_), .ZN(new_n15603_));
  XNOR2_X1   g14601(.A1(new_n14452_), .A2(new_n14455_), .ZN(new_n15604_));
  XOR2_X1    g14602(.A1(new_n14467_), .A2(new_n14475_), .Z(new_n15605_));
  NOR2_X1    g14603(.A1(new_n15604_), .A2(new_n15605_), .ZN(new_n15606_));
  NAND2_X1   g14604(.A1(new_n15603_), .A2(new_n15606_), .ZN(new_n15607_));
  NOR2_X1    g14605(.A1(new_n15591_), .A2(new_n15594_), .ZN(new_n15608_));
  AOI21_X1   g14606(.A1(new_n15600_), .A2(new_n14456_), .B(new_n15608_), .ZN(new_n15609_));
  NOR2_X1    g14607(.A1(new_n15609_), .A2(new_n15604_), .ZN(new_n15610_));
  NOR4_X1    g14608(.A1(new_n15607_), .A2(new_n15596_), .A3(new_n15597_), .A4(new_n15610_), .ZN(new_n15611_));
  NOR4_X1    g14609(.A1(new_n15597_), .A2(new_n15596_), .A3(new_n15604_), .A4(new_n15605_), .ZN(new_n15612_));
  XOR2_X1    g14610(.A1(new_n15600_), .A2(new_n15595_), .Z(new_n15613_));
  NOR2_X1    g14611(.A1(new_n15613_), .A2(new_n15610_), .ZN(new_n15614_));
  NOR2_X1    g14612(.A1(new_n15614_), .A2(new_n15612_), .ZN(new_n15615_));
  OAI21_X1   g14613(.A1(new_n15615_), .A2(new_n15611_), .B(new_n15588_), .ZN(new_n15616_));
  AOI21_X1   g14614(.A1(new_n15586_), .A2(new_n14486_), .B(new_n15582_), .ZN(new_n15617_));
  NOR2_X1    g14615(.A1(new_n15586_), .A2(new_n15578_), .ZN(new_n15618_));
  NOR2_X1    g14616(.A1(new_n15576_), .A2(new_n14486_), .ZN(new_n15619_));
  OAI22_X1   g14617(.A1(new_n15605_), .A2(new_n15617_), .B1(new_n15619_), .B2(new_n15618_), .ZN(new_n15620_));
  OAI21_X1   g14618(.A1(new_n15609_), .A2(new_n15604_), .B(new_n15603_), .ZN(new_n15621_));
  NOR2_X1    g14619(.A1(new_n15621_), .A2(new_n15612_), .ZN(new_n15622_));
  NAND3_X1   g14620(.A1(new_n15606_), .A2(new_n14457_), .A3(new_n14487_), .ZN(new_n15623_));
  NOR2_X1    g14621(.A1(new_n15614_), .A2(new_n15623_), .ZN(new_n15624_));
  OAI21_X1   g14622(.A1(new_n15622_), .A2(new_n15624_), .B(new_n15620_), .ZN(new_n15625_));
  XNOR2_X1   g14623(.A1(new_n14459_), .A2(new_n14488_), .ZN(new_n15626_));
  XNOR2_X1   g14624(.A1(new_n14543_), .A2(new_n14515_), .ZN(new_n15627_));
  NOR2_X1    g14625(.A1(new_n15626_), .A2(new_n15627_), .ZN(new_n15628_));
  NAND3_X1   g14626(.A1(new_n15616_), .A2(new_n15625_), .A3(new_n15628_), .ZN(new_n15629_));
  NOR2_X1    g14627(.A1(new_n15610_), .A2(new_n15597_), .ZN(new_n15630_));
  NAND4_X1   g14628(.A1(new_n15630_), .A2(new_n15609_), .A3(new_n15603_), .A4(new_n15606_), .ZN(new_n15631_));
  NAND2_X1   g14629(.A1(new_n15621_), .A2(new_n15623_), .ZN(new_n15632_));
  AOI21_X1   g14630(.A1(new_n15631_), .A2(new_n15632_), .B(new_n15620_), .ZN(new_n15633_));
  NAND2_X1   g14631(.A1(new_n15614_), .A2(new_n15623_), .ZN(new_n15634_));
  NAND2_X1   g14632(.A1(new_n15621_), .A2(new_n15612_), .ZN(new_n15635_));
  AOI21_X1   g14633(.A1(new_n15635_), .A2(new_n15634_), .B(new_n15588_), .ZN(new_n15636_));
  NAND2_X1   g14634(.A1(new_n14489_), .A2(new_n14544_), .ZN(new_n15637_));
  OAI21_X1   g14635(.A1(new_n15633_), .A2(new_n15636_), .B(new_n15637_), .ZN(new_n15638_));
  AOI21_X1   g14636(.A1(new_n15638_), .A2(new_n15629_), .B(new_n15574_), .ZN(new_n15639_));
  XOR2_X1    g14637(.A1(new_n15554_), .A2(new_n15545_), .Z(new_n15640_));
  NOR2_X1    g14638(.A1(new_n15565_), .A2(new_n15564_), .ZN(new_n15641_));
  NAND4_X1   g14639(.A1(new_n15641_), .A2(new_n15549_), .A3(new_n15568_), .A4(new_n15544_), .ZN(new_n15642_));
  AOI21_X1   g14640(.A1(new_n15642_), .A2(new_n15571_), .B(new_n15542_), .ZN(new_n15643_));
  AOI21_X1   g14641(.A1(new_n15640_), .A2(new_n15542_), .B(new_n15643_), .ZN(new_n15644_));
  NAND3_X1   g14642(.A1(new_n15625_), .A2(new_n15616_), .A3(new_n15637_), .ZN(new_n15645_));
  OAI21_X1   g14643(.A1(new_n15633_), .A2(new_n15636_), .B(new_n15628_), .ZN(new_n15646_));
  AOI21_X1   g14644(.A1(new_n15645_), .A2(new_n15646_), .B(new_n15644_), .ZN(new_n15647_));
  NOR2_X1    g14645(.A1(new_n15647_), .A2(new_n15639_), .ZN(new_n15648_));
  NOR2_X1    g14646(.A1(new_n15648_), .A2(new_n15528_), .ZN(new_n15649_));
  NOR3_X1    g14647(.A1(new_n15647_), .A2(new_n15639_), .A3(new_n15527_), .ZN(new_n15650_));
  OAI21_X1   g14648(.A1(new_n15649_), .A2(new_n15650_), .B(new_n15526_), .ZN(new_n15651_));
  OAI21_X1   g14649(.A1(new_n15497_), .A2(new_n15509_), .B(new_n15522_), .ZN(new_n15652_));
  NOR3_X1    g14650(.A1(new_n15486_), .A2(new_n15495_), .A3(new_n15508_), .ZN(new_n15653_));
  AOI21_X1   g14651(.A1(new_n15502_), .A2(new_n15505_), .B(new_n15496_), .ZN(new_n15654_));
  OAI21_X1   g14652(.A1(new_n15654_), .A2(new_n15653_), .B(new_n15452_), .ZN(new_n15655_));
  NAND2_X1   g14653(.A1(new_n15652_), .A2(new_n15655_), .ZN(new_n15656_));
  NOR2_X1    g14654(.A1(new_n15648_), .A2(new_n15527_), .ZN(new_n15657_));
  NOR3_X1    g14655(.A1(new_n15528_), .A2(new_n15647_), .A3(new_n15639_), .ZN(new_n15658_));
  OAI21_X1   g14656(.A1(new_n15657_), .A2(new_n15658_), .B(new_n15656_), .ZN(new_n15659_));
  NAND2_X1   g14657(.A1(new_n15651_), .A2(new_n15659_), .ZN(new_n15660_));
  XNOR2_X1   g14658(.A1(new_n14894_), .A2(new_n14903_), .ZN(new_n15661_));
  XOR2_X1    g14659(.A1(new_n14906_), .A2(new_n14908_), .Z(new_n15662_));
  NOR2_X1    g14660(.A1(new_n14894_), .A2(new_n14903_), .ZN(new_n15663_));
  NOR2_X1    g14661(.A1(new_n14906_), .A2(new_n14908_), .ZN(new_n15664_));
  AOI21_X1   g14662(.A1(new_n15662_), .A2(new_n15663_), .B(new_n15664_), .ZN(new_n15665_));
  INV_X1     g14663(.I(new_n15663_), .ZN(new_n15666_));
  NOR2_X1    g14664(.A1(new_n15662_), .A2(new_n15666_), .ZN(new_n15667_));
  XNOR2_X1   g14665(.A1(new_n14906_), .A2(new_n14908_), .ZN(new_n15668_));
  NOR2_X1    g14666(.A1(new_n15668_), .A2(new_n15663_), .ZN(new_n15669_));
  OAI22_X1   g14667(.A1(new_n15661_), .A2(new_n15665_), .B1(new_n15669_), .B2(new_n15667_), .ZN(new_n15670_));
  AOI21_X1   g14668(.A1(new_n14869_), .A2(\A[810] ), .B(new_n14874_), .ZN(new_n15671_));
  XOR2_X1    g14669(.A1(new_n15671_), .A2(new_n14880_), .Z(new_n15672_));
  INV_X1     g14670(.I(new_n14870_), .ZN(new_n15673_));
  NAND2_X1   g14671(.A1(new_n15673_), .A2(new_n14861_), .ZN(new_n15674_));
  NOR2_X1    g14672(.A1(new_n15672_), .A2(new_n15674_), .ZN(new_n15675_));
  XOR2_X1    g14673(.A1(new_n14876_), .A2(new_n14880_), .Z(new_n15676_));
  NOR2_X1    g14674(.A1(new_n15676_), .A2(new_n14883_), .ZN(new_n15677_));
  NOR2_X1    g14675(.A1(new_n15677_), .A2(new_n15675_), .ZN(new_n15678_));
  NAND2_X1   g14676(.A1(new_n14871_), .A2(new_n14904_), .ZN(new_n15679_));
  NOR2_X1    g14677(.A1(new_n15678_), .A2(new_n15679_), .ZN(new_n15680_));
  NOR2_X1    g14678(.A1(new_n15671_), .A2(new_n14880_), .ZN(new_n15681_));
  INV_X1     g14679(.I(new_n15681_), .ZN(new_n15682_));
  OAI21_X1   g14680(.A1(new_n15676_), .A2(new_n15674_), .B(new_n15682_), .ZN(new_n15683_));
  NAND2_X1   g14681(.A1(new_n15683_), .A2(new_n14871_), .ZN(new_n15684_));
  NAND4_X1   g14682(.A1(new_n15680_), .A2(new_n14884_), .A3(new_n14909_), .A4(new_n15684_), .ZN(new_n15685_));
  INV_X1     g14683(.I(new_n14871_), .ZN(new_n15686_));
  NOR2_X1    g14684(.A1(new_n15686_), .A2(new_n15661_), .ZN(new_n15687_));
  NAND3_X1   g14685(.A1(new_n15687_), .A2(new_n14884_), .A3(new_n14909_), .ZN(new_n15688_));
  NAND2_X1   g14686(.A1(new_n15676_), .A2(new_n14883_), .ZN(new_n15689_));
  NAND2_X1   g14687(.A1(new_n15672_), .A2(new_n15674_), .ZN(new_n15690_));
  NAND2_X1   g14688(.A1(new_n15689_), .A2(new_n15690_), .ZN(new_n15691_));
  NAND2_X1   g14689(.A1(new_n15684_), .A2(new_n15691_), .ZN(new_n15692_));
  NAND2_X1   g14690(.A1(new_n15688_), .A2(new_n15692_), .ZN(new_n15693_));
  AOI21_X1   g14691(.A1(new_n15685_), .A2(new_n15693_), .B(new_n15670_), .ZN(new_n15694_));
  INV_X1     g14692(.I(new_n15665_), .ZN(new_n15695_));
  NAND2_X1   g14693(.A1(new_n15668_), .A2(new_n15663_), .ZN(new_n15696_));
  NAND2_X1   g14694(.A1(new_n15662_), .A2(new_n15666_), .ZN(new_n15697_));
  AOI22_X1   g14695(.A1(new_n15695_), .A2(new_n14904_), .B1(new_n15696_), .B2(new_n15697_), .ZN(new_n15698_));
  AOI21_X1   g14696(.A1(new_n14871_), .A2(new_n15683_), .B(new_n15678_), .ZN(new_n15699_));
  NAND2_X1   g14697(.A1(new_n15699_), .A2(new_n15688_), .ZN(new_n15700_));
  INV_X1     g14698(.I(new_n14884_), .ZN(new_n15701_));
  INV_X1     g14699(.I(new_n14909_), .ZN(new_n15702_));
  NOR3_X1    g14700(.A1(new_n15679_), .A2(new_n15701_), .A3(new_n15702_), .ZN(new_n15703_));
  NAND2_X1   g14701(.A1(new_n15692_), .A2(new_n15703_), .ZN(new_n15704_));
  AOI21_X1   g14702(.A1(new_n15700_), .A2(new_n15704_), .B(new_n15698_), .ZN(new_n15705_));
  NOR2_X1    g14703(.A1(new_n15694_), .A2(new_n15705_), .ZN(new_n15706_));
  XNOR2_X1   g14704(.A1(new_n14805_), .A2(new_n14813_), .ZN(new_n15707_));
  XOR2_X1    g14705(.A1(new_n14816_), .A2(new_n14819_), .Z(new_n15708_));
  NOR2_X1    g14706(.A1(new_n14816_), .A2(new_n14819_), .ZN(new_n15709_));
  AOI21_X1   g14707(.A1(new_n15708_), .A2(new_n14821_), .B(new_n15709_), .ZN(new_n15710_));
  NAND2_X1   g14708(.A1(new_n14817_), .A2(new_n14819_), .ZN(new_n15711_));
  NAND2_X1   g14709(.A1(new_n14820_), .A2(new_n14816_), .ZN(new_n15712_));
  NAND3_X1   g14710(.A1(new_n15711_), .A2(new_n15712_), .A3(new_n14821_), .ZN(new_n15713_));
  INV_X1     g14711(.I(new_n15713_), .ZN(new_n15714_));
  XNOR2_X1   g14712(.A1(new_n14816_), .A2(new_n14819_), .ZN(new_n15715_));
  NOR2_X1    g14713(.A1(new_n15715_), .A2(new_n14821_), .ZN(new_n15716_));
  OAI22_X1   g14714(.A1(new_n15714_), .A2(new_n15716_), .B1(new_n15710_), .B2(new_n15707_), .ZN(new_n15717_));
  XOR2_X1    g14715(.A1(new_n14831_), .A2(new_n14839_), .Z(new_n15718_));
  AOI21_X1   g14716(.A1(new_n14837_), .A2(\A[822] ), .B(new_n14841_), .ZN(new_n15719_));
  NAND2_X1   g14717(.A1(new_n14848_), .A2(new_n15719_), .ZN(new_n15720_));
  NAND2_X1   g14718(.A1(new_n14826_), .A2(\A[818] ), .ZN(new_n15721_));
  NAND2_X1   g14719(.A1(new_n14829_), .A2(new_n15721_), .ZN(new_n15722_));
  AOI21_X1   g14720(.A1(new_n15722_), .A2(\A[819] ), .B(new_n14846_), .ZN(new_n15723_));
  NAND2_X1   g14721(.A1(new_n14844_), .A2(new_n15723_), .ZN(new_n15724_));
  NAND2_X1   g14722(.A1(new_n15724_), .A2(new_n15720_), .ZN(new_n15725_));
  INV_X1     g14723(.I(new_n14839_), .ZN(new_n15726_));
  NAND2_X1   g14724(.A1(new_n15726_), .A2(new_n14831_), .ZN(new_n15727_));
  NOR2_X1    g14725(.A1(new_n15725_), .A2(new_n15727_), .ZN(new_n15728_));
  AOI21_X1   g14726(.A1(new_n15720_), .A2(new_n15724_), .B(new_n14850_), .ZN(new_n15729_));
  NOR2_X1    g14727(.A1(new_n15728_), .A2(new_n15729_), .ZN(new_n15730_));
  NOR3_X1    g14728(.A1(new_n15730_), .A2(new_n15707_), .A3(new_n15718_), .ZN(new_n15731_));
  NOR2_X1    g14729(.A1(new_n15719_), .A2(new_n15723_), .ZN(new_n15732_));
  AOI21_X1   g14730(.A1(new_n15725_), .A2(new_n14850_), .B(new_n15732_), .ZN(new_n15733_));
  NOR2_X1    g14731(.A1(new_n15733_), .A2(new_n15718_), .ZN(new_n15734_));
  INV_X1     g14732(.I(new_n15734_), .ZN(new_n15735_));
  NAND4_X1   g14733(.A1(new_n15731_), .A2(new_n14822_), .A3(new_n15735_), .A4(new_n14851_), .ZN(new_n15736_));
  NOR2_X1    g14734(.A1(new_n15707_), .A2(new_n15718_), .ZN(new_n15737_));
  NAND3_X1   g14735(.A1(new_n15737_), .A2(new_n14822_), .A3(new_n14851_), .ZN(new_n15738_));
  NAND3_X1   g14736(.A1(new_n14850_), .A2(new_n15720_), .A3(new_n15724_), .ZN(new_n15739_));
  NAND2_X1   g14737(.A1(new_n15725_), .A2(new_n15727_), .ZN(new_n15740_));
  NAND2_X1   g14738(.A1(new_n15740_), .A2(new_n15739_), .ZN(new_n15741_));
  OAI21_X1   g14739(.A1(new_n15718_), .A2(new_n15733_), .B(new_n15741_), .ZN(new_n15742_));
  NAND2_X1   g14740(.A1(new_n15742_), .A2(new_n15738_), .ZN(new_n15743_));
  AOI21_X1   g14741(.A1(new_n15736_), .A2(new_n15743_), .B(new_n15717_), .ZN(new_n15744_));
  INV_X1     g14742(.I(new_n14821_), .ZN(new_n15745_));
  INV_X1     g14743(.I(new_n15709_), .ZN(new_n15746_));
  OAI21_X1   g14744(.A1(new_n15715_), .A2(new_n15745_), .B(new_n15746_), .ZN(new_n15747_));
  NAND2_X1   g14745(.A1(new_n15708_), .A2(new_n15745_), .ZN(new_n15748_));
  AOI22_X1   g14746(.A1(new_n15747_), .A2(new_n14814_), .B1(new_n15748_), .B2(new_n15713_), .ZN(new_n15749_));
  NOR2_X1    g14747(.A1(new_n15734_), .A2(new_n15730_), .ZN(new_n15750_));
  NAND2_X1   g14748(.A1(new_n15750_), .A2(new_n15738_), .ZN(new_n15751_));
  AND4_X2    g14749(.A1(new_n14814_), .A2(new_n14851_), .A3(new_n14822_), .A4(new_n14840_), .Z(new_n15752_));
  NAND2_X1   g14750(.A1(new_n15742_), .A2(new_n15752_), .ZN(new_n15753_));
  AOI21_X1   g14751(.A1(new_n15753_), .A2(new_n15751_), .B(new_n15749_), .ZN(new_n15754_));
  NAND2_X1   g14752(.A1(new_n14911_), .A2(new_n14853_), .ZN(new_n15755_));
  NOR3_X1    g14753(.A1(new_n15744_), .A2(new_n15754_), .A3(new_n15755_), .ZN(new_n15756_));
  NAND3_X1   g14754(.A1(new_n15741_), .A2(new_n14822_), .A3(new_n15737_), .ZN(new_n15757_));
  OAI21_X1   g14755(.A1(new_n15733_), .A2(new_n15718_), .B(new_n14851_), .ZN(new_n15758_));
  NOR2_X1    g14756(.A1(new_n15757_), .A2(new_n15758_), .ZN(new_n15759_));
  NOR2_X1    g14757(.A1(new_n15750_), .A2(new_n15752_), .ZN(new_n15760_));
  OAI21_X1   g14758(.A1(new_n15760_), .A2(new_n15759_), .B(new_n15749_), .ZN(new_n15761_));
  NOR2_X1    g14759(.A1(new_n15742_), .A2(new_n15752_), .ZN(new_n15762_));
  NOR2_X1    g14760(.A1(new_n15750_), .A2(new_n15738_), .ZN(new_n15763_));
  OAI21_X1   g14761(.A1(new_n15762_), .A2(new_n15763_), .B(new_n15717_), .ZN(new_n15764_));
  AND2_X2    g14762(.A1(new_n14911_), .A2(new_n14853_), .Z(new_n15765_));
  AOI21_X1   g14763(.A1(new_n15764_), .A2(new_n15761_), .B(new_n15765_), .ZN(new_n15766_));
  OAI21_X1   g14764(.A1(new_n15766_), .A2(new_n15756_), .B(new_n15706_), .ZN(new_n15767_));
  NAND3_X1   g14765(.A1(new_n15687_), .A2(new_n15691_), .A3(new_n14884_), .ZN(new_n15768_));
  NAND2_X1   g14766(.A1(new_n15684_), .A2(new_n14909_), .ZN(new_n15769_));
  NOR2_X1    g14767(.A1(new_n15768_), .A2(new_n15769_), .ZN(new_n15770_));
  NOR2_X1    g14768(.A1(new_n15699_), .A2(new_n15703_), .ZN(new_n15771_));
  OAI21_X1   g14769(.A1(new_n15771_), .A2(new_n15770_), .B(new_n15698_), .ZN(new_n15772_));
  NOR2_X1    g14770(.A1(new_n15692_), .A2(new_n15703_), .ZN(new_n15773_));
  NOR2_X1    g14771(.A1(new_n15699_), .A2(new_n15688_), .ZN(new_n15774_));
  OAI21_X1   g14772(.A1(new_n15774_), .A2(new_n15773_), .B(new_n15670_), .ZN(new_n15775_));
  NAND2_X1   g14773(.A1(new_n15772_), .A2(new_n15775_), .ZN(new_n15776_));
  NOR3_X1    g14774(.A1(new_n15765_), .A2(new_n15744_), .A3(new_n15754_), .ZN(new_n15777_));
  AOI21_X1   g14775(.A1(new_n15764_), .A2(new_n15761_), .B(new_n15755_), .ZN(new_n15778_));
  OAI21_X1   g14776(.A1(new_n15777_), .A2(new_n15778_), .B(new_n15776_), .ZN(new_n15779_));
  NAND2_X1   g14777(.A1(new_n15767_), .A2(new_n15779_), .ZN(new_n15780_));
  INV_X1     g14778(.I(new_n15780_), .ZN(new_n15781_));
  AOI21_X1   g14779(.A1(new_n14743_), .A2(\A[825] ), .B(new_n14761_), .ZN(new_n15782_));
  XOR2_X1    g14780(.A1(new_n14757_), .A2(new_n15782_), .Z(new_n15783_));
  NOR2_X1    g14781(.A1(new_n14757_), .A2(new_n15782_), .ZN(new_n15784_));
  AOI21_X1   g14782(.A1(new_n15783_), .A2(new_n14764_), .B(new_n15784_), .ZN(new_n15785_));
  INV_X1     g14783(.I(new_n15785_), .ZN(new_n15786_));
  XOR2_X1    g14784(.A1(new_n14763_), .A2(new_n14757_), .Z(new_n15787_));
  NAND2_X1   g14785(.A1(new_n15787_), .A2(new_n14764_), .ZN(new_n15788_));
  INV_X1     g14786(.I(new_n14764_), .ZN(new_n15789_));
  NAND2_X1   g14787(.A1(new_n15783_), .A2(new_n15789_), .ZN(new_n15790_));
  AOI22_X1   g14788(.A1(new_n15786_), .A2(new_n14755_), .B1(new_n15788_), .B2(new_n15790_), .ZN(new_n15791_));
  XOR2_X1    g14789(.A1(new_n14792_), .A2(new_n14786_), .Z(new_n15792_));
  NAND2_X1   g14790(.A1(new_n15792_), .A2(new_n14793_), .ZN(new_n15793_));
  AOI21_X1   g14791(.A1(new_n14772_), .A2(\A[831] ), .B(new_n14790_), .ZN(new_n15794_));
  XOR2_X1    g14792(.A1(new_n14786_), .A2(new_n15794_), .Z(new_n15795_));
  INV_X1     g14793(.I(new_n14793_), .ZN(new_n15796_));
  NAND2_X1   g14794(.A1(new_n15795_), .A2(new_n15796_), .ZN(new_n15797_));
  NAND2_X1   g14795(.A1(new_n15793_), .A2(new_n15797_), .ZN(new_n15798_));
  XNOR2_X1   g14796(.A1(new_n14746_), .A2(new_n14754_), .ZN(new_n15799_));
  XNOR2_X1   g14797(.A1(new_n14775_), .A2(new_n14783_), .ZN(new_n15800_));
  NOR2_X1    g14798(.A1(new_n15799_), .A2(new_n15800_), .ZN(new_n15801_));
  NAND3_X1   g14799(.A1(new_n15798_), .A2(new_n14765_), .A3(new_n15801_), .ZN(new_n15802_));
  NOR2_X1    g14800(.A1(new_n14786_), .A2(new_n15794_), .ZN(new_n15803_));
  INV_X1     g14801(.I(new_n15803_), .ZN(new_n15804_));
  OAI21_X1   g14802(.A1(new_n15792_), .A2(new_n15796_), .B(new_n15804_), .ZN(new_n15805_));
  NAND2_X1   g14803(.A1(new_n15805_), .A2(new_n14784_), .ZN(new_n15806_));
  NAND2_X1   g14804(.A1(new_n15806_), .A2(new_n14794_), .ZN(new_n15807_));
  NOR2_X1    g14805(.A1(new_n15802_), .A2(new_n15807_), .ZN(new_n15808_));
  AND4_X2    g14806(.A1(new_n14755_), .A2(new_n14784_), .A3(new_n14765_), .A4(new_n14794_), .Z(new_n15809_));
  AOI22_X1   g14807(.A1(new_n15805_), .A2(new_n14784_), .B1(new_n15793_), .B2(new_n15797_), .ZN(new_n15810_));
  NOR2_X1    g14808(.A1(new_n15810_), .A2(new_n15809_), .ZN(new_n15811_));
  OAI21_X1   g14809(.A1(new_n15808_), .A2(new_n15811_), .B(new_n15791_), .ZN(new_n15812_));
  NOR2_X1    g14810(.A1(new_n15783_), .A2(new_n15789_), .ZN(new_n15813_));
  NOR2_X1    g14811(.A1(new_n15787_), .A2(new_n14764_), .ZN(new_n15814_));
  OAI22_X1   g14812(.A1(new_n15799_), .A2(new_n15785_), .B1(new_n15813_), .B2(new_n15814_), .ZN(new_n15815_));
  NAND3_X1   g14813(.A1(new_n15801_), .A2(new_n14765_), .A3(new_n14794_), .ZN(new_n15816_));
  NOR2_X1    g14814(.A1(new_n15810_), .A2(new_n15816_), .ZN(new_n15817_));
  NAND2_X1   g14815(.A1(new_n15806_), .A2(new_n15798_), .ZN(new_n15818_));
  NOR2_X1    g14816(.A1(new_n15818_), .A2(new_n15809_), .ZN(new_n15819_));
  OAI21_X1   g14817(.A1(new_n15819_), .A2(new_n15817_), .B(new_n15815_), .ZN(new_n15820_));
  NAND2_X1   g14818(.A1(new_n15812_), .A2(new_n15820_), .ZN(new_n15821_));
  NAND2_X1   g14819(.A1(new_n14737_), .A2(new_n14796_), .ZN(new_n15822_));
  AOI21_X1   g14820(.A1(new_n14691_), .A2(\A[840] ), .B(new_n14696_), .ZN(new_n15823_));
  XOR2_X1    g14821(.A1(new_n14702_), .A2(new_n15823_), .Z(new_n15824_));
  INV_X1     g14822(.I(new_n14693_), .ZN(new_n15825_));
  NAND2_X1   g14823(.A1(new_n15825_), .A2(new_n14685_), .ZN(new_n15826_));
  NAND2_X1   g14824(.A1(new_n14680_), .A2(\A[836] ), .ZN(new_n15827_));
  NAND2_X1   g14825(.A1(new_n14683_), .A2(new_n15827_), .ZN(new_n15828_));
  AOI21_X1   g14826(.A1(new_n15828_), .A2(\A[837] ), .B(new_n14700_), .ZN(new_n15829_));
  NOR2_X1    g14827(.A1(new_n15823_), .A2(new_n15829_), .ZN(new_n15830_));
  INV_X1     g14828(.I(new_n15830_), .ZN(new_n15831_));
  OAI21_X1   g14829(.A1(new_n15824_), .A2(new_n15826_), .B(new_n15831_), .ZN(new_n15832_));
  NAND2_X1   g14830(.A1(new_n14698_), .A2(new_n15829_), .ZN(new_n15833_));
  NAND2_X1   g14831(.A1(new_n14702_), .A2(new_n15823_), .ZN(new_n15834_));
  NAND3_X1   g14832(.A1(new_n14704_), .A2(new_n15833_), .A3(new_n15834_), .ZN(new_n15835_));
  NAND2_X1   g14833(.A1(new_n15833_), .A2(new_n15834_), .ZN(new_n15836_));
  NAND2_X1   g14834(.A1(new_n15836_), .A2(new_n15826_), .ZN(new_n15837_));
  AOI22_X1   g14835(.A1(new_n15832_), .A2(new_n14694_), .B1(new_n15837_), .B2(new_n15835_), .ZN(new_n15838_));
  AOI21_X1   g14836(.A1(new_n14721_), .A2(\A[846] ), .B(new_n14726_), .ZN(new_n15839_));
  NAND2_X1   g14837(.A1(new_n14733_), .A2(new_n15839_), .ZN(new_n15840_));
  AOI21_X1   g14838(.A1(new_n14712_), .A2(\A[843] ), .B(new_n14731_), .ZN(new_n15841_));
  NAND2_X1   g14839(.A1(new_n14728_), .A2(new_n15841_), .ZN(new_n15842_));
  NAND3_X1   g14840(.A1(new_n15842_), .A2(new_n14734_), .A3(new_n15840_), .ZN(new_n15843_));
  NAND2_X1   g14841(.A1(new_n15842_), .A2(new_n15840_), .ZN(new_n15844_));
  INV_X1     g14842(.I(new_n14734_), .ZN(new_n15845_));
  NAND2_X1   g14843(.A1(new_n15844_), .A2(new_n15845_), .ZN(new_n15846_));
  NAND2_X1   g14844(.A1(new_n15846_), .A2(new_n15843_), .ZN(new_n15847_));
  XOR2_X1    g14845(.A1(new_n14685_), .A2(new_n14693_), .Z(new_n15848_));
  XNOR2_X1   g14846(.A1(new_n14715_), .A2(new_n14723_), .ZN(new_n15849_));
  NOR2_X1    g14847(.A1(new_n15849_), .A2(new_n15848_), .ZN(new_n15850_));
  NAND3_X1   g14848(.A1(new_n15847_), .A2(new_n14705_), .A3(new_n15850_), .ZN(new_n15851_));
  NOR2_X1    g14849(.A1(new_n15839_), .A2(new_n15841_), .ZN(new_n15852_));
  AOI21_X1   g14850(.A1(new_n15844_), .A2(new_n14734_), .B(new_n15852_), .ZN(new_n15853_));
  OAI21_X1   g14851(.A1(new_n15853_), .A2(new_n15849_), .B(new_n14735_), .ZN(new_n15854_));
  NOR2_X1    g14852(.A1(new_n15851_), .A2(new_n15854_), .ZN(new_n15855_));
  AND4_X2    g14853(.A1(new_n14694_), .A2(new_n14705_), .A3(new_n14724_), .A4(new_n14735_), .Z(new_n15856_));
  XOR2_X1    g14854(.A1(new_n14733_), .A2(new_n15839_), .Z(new_n15857_));
  INV_X1     g14855(.I(new_n15852_), .ZN(new_n15858_));
  OAI21_X1   g14856(.A1(new_n15857_), .A2(new_n15845_), .B(new_n15858_), .ZN(new_n15859_));
  AOI22_X1   g14857(.A1(new_n15859_), .A2(new_n14724_), .B1(new_n15846_), .B2(new_n15843_), .ZN(new_n15860_));
  NOR2_X1    g14858(.A1(new_n15856_), .A2(new_n15860_), .ZN(new_n15861_));
  OAI21_X1   g14859(.A1(new_n15855_), .A2(new_n15861_), .B(new_n15838_), .ZN(new_n15862_));
  AOI21_X1   g14860(.A1(new_n15836_), .A2(new_n14704_), .B(new_n15830_), .ZN(new_n15863_));
  NAND2_X1   g14861(.A1(new_n15837_), .A2(new_n15835_), .ZN(new_n15864_));
  OAI21_X1   g14862(.A1(new_n15848_), .A2(new_n15863_), .B(new_n15864_), .ZN(new_n15865_));
  INV_X1     g14863(.I(new_n15843_), .ZN(new_n15866_));
  NOR2_X1    g14864(.A1(new_n15857_), .A2(new_n14734_), .ZN(new_n15867_));
  OAI22_X1   g14865(.A1(new_n15849_), .A2(new_n15853_), .B1(new_n15867_), .B2(new_n15866_), .ZN(new_n15868_));
  NOR2_X1    g14866(.A1(new_n15856_), .A2(new_n15868_), .ZN(new_n15869_));
  NAND3_X1   g14867(.A1(new_n15850_), .A2(new_n14705_), .A3(new_n14735_), .ZN(new_n15870_));
  NOR2_X1    g14868(.A1(new_n15860_), .A2(new_n15870_), .ZN(new_n15871_));
  OAI21_X1   g14869(.A1(new_n15869_), .A2(new_n15871_), .B(new_n15865_), .ZN(new_n15872_));
  AOI21_X1   g14870(.A1(new_n15862_), .A2(new_n15872_), .B(new_n15822_), .ZN(new_n15873_));
  XNOR2_X1   g14871(.A1(new_n14706_), .A2(new_n14736_), .ZN(new_n15874_));
  XNOR2_X1   g14872(.A1(new_n14766_), .A2(new_n14795_), .ZN(new_n15875_));
  NOR2_X1    g14873(.A1(new_n15874_), .A2(new_n15875_), .ZN(new_n15876_));
  OAI21_X1   g14874(.A1(new_n15847_), .A2(new_n14724_), .B(new_n15859_), .ZN(new_n15877_));
  NAND4_X1   g14875(.A1(new_n15877_), .A2(new_n14705_), .A3(new_n15847_), .A4(new_n15850_), .ZN(new_n15878_));
  NAND2_X1   g14876(.A1(new_n15868_), .A2(new_n15870_), .ZN(new_n15879_));
  AOI21_X1   g14877(.A1(new_n15878_), .A2(new_n15879_), .B(new_n15865_), .ZN(new_n15880_));
  NAND2_X1   g14878(.A1(new_n15860_), .A2(new_n15870_), .ZN(new_n15881_));
  NAND2_X1   g14879(.A1(new_n15856_), .A2(new_n15868_), .ZN(new_n15882_));
  AOI21_X1   g14880(.A1(new_n15882_), .A2(new_n15881_), .B(new_n15838_), .ZN(new_n15883_));
  NOR3_X1    g14881(.A1(new_n15880_), .A2(new_n15883_), .A3(new_n15876_), .ZN(new_n15884_));
  OAI21_X1   g14882(.A1(new_n15884_), .A2(new_n15873_), .B(new_n15821_), .ZN(new_n15885_));
  OAI21_X1   g14883(.A1(new_n15798_), .A2(new_n14784_), .B(new_n15805_), .ZN(new_n15886_));
  NAND4_X1   g14884(.A1(new_n15886_), .A2(new_n14765_), .A3(new_n15798_), .A4(new_n15801_), .ZN(new_n15887_));
  NAND2_X1   g14885(.A1(new_n15818_), .A2(new_n15816_), .ZN(new_n15888_));
  AOI21_X1   g14886(.A1(new_n15887_), .A2(new_n15888_), .B(new_n15815_), .ZN(new_n15889_));
  NAND2_X1   g14887(.A1(new_n15818_), .A2(new_n15809_), .ZN(new_n15890_));
  NAND2_X1   g14888(.A1(new_n15810_), .A2(new_n15816_), .ZN(new_n15891_));
  AOI21_X1   g14889(.A1(new_n15890_), .A2(new_n15891_), .B(new_n15791_), .ZN(new_n15892_));
  NOR2_X1    g14890(.A1(new_n15889_), .A2(new_n15892_), .ZN(new_n15893_));
  AOI21_X1   g14891(.A1(new_n15862_), .A2(new_n15872_), .B(new_n15876_), .ZN(new_n15894_));
  NOR3_X1    g14892(.A1(new_n15880_), .A2(new_n15883_), .A3(new_n15822_), .ZN(new_n15895_));
  OAI21_X1   g14893(.A1(new_n15895_), .A2(new_n15894_), .B(new_n15893_), .ZN(new_n15896_));
  NAND2_X1   g14894(.A1(new_n14912_), .A2(new_n14797_), .ZN(new_n15897_));
  NAND3_X1   g14895(.A1(new_n15896_), .A2(new_n15885_), .A3(new_n15897_), .ZN(new_n15898_));
  INV_X1     g14896(.I(new_n15897_), .ZN(new_n15899_));
  NAND2_X1   g14897(.A1(new_n15896_), .A2(new_n15885_), .ZN(new_n15900_));
  NAND2_X1   g14898(.A1(new_n15900_), .A2(new_n15899_), .ZN(new_n15901_));
  AOI21_X1   g14899(.A1(new_n15901_), .A2(new_n15898_), .B(new_n15781_), .ZN(new_n15902_));
  NAND3_X1   g14900(.A1(new_n15899_), .A2(new_n15896_), .A3(new_n15885_), .ZN(new_n15903_));
  NAND2_X1   g14901(.A1(new_n15900_), .A2(new_n15897_), .ZN(new_n15904_));
  AOI21_X1   g14902(.A1(new_n15904_), .A2(new_n15903_), .B(new_n15780_), .ZN(new_n15905_));
  NOR2_X1    g14903(.A1(new_n14677_), .A2(new_n14913_), .ZN(new_n15906_));
  INV_X1     g14904(.I(new_n15906_), .ZN(new_n15907_));
  NOR3_X1    g14905(.A1(new_n15902_), .A2(new_n15905_), .A3(new_n15907_), .ZN(new_n15908_));
  NAND2_X1   g14906(.A1(new_n15901_), .A2(new_n15898_), .ZN(new_n15909_));
  NAND2_X1   g14907(.A1(new_n15909_), .A2(new_n15780_), .ZN(new_n15910_));
  INV_X1     g14908(.I(new_n15905_), .ZN(new_n15911_));
  AOI21_X1   g14909(.A1(new_n15911_), .A2(new_n15910_), .B(new_n15906_), .ZN(new_n15912_));
  NOR2_X1    g14910(.A1(new_n15912_), .A2(new_n15908_), .ZN(new_n15913_));
  NOR2_X1    g14911(.A1(new_n15913_), .A2(new_n15660_), .ZN(new_n15914_));
  AND2_X2    g14912(.A1(new_n15651_), .A2(new_n15659_), .Z(new_n15915_));
  NAND3_X1   g14913(.A1(new_n15911_), .A2(new_n15910_), .A3(new_n15907_), .ZN(new_n15916_));
  OAI21_X1   g14914(.A1(new_n15902_), .A2(new_n15905_), .B(new_n15906_), .ZN(new_n15917_));
  AOI21_X1   g14915(.A1(new_n15916_), .A2(new_n15917_), .B(new_n15915_), .ZN(new_n15918_));
  OAI21_X1   g14916(.A1(new_n15914_), .A2(new_n15918_), .B(new_n15408_), .ZN(new_n15919_));
  XOR2_X1    g14917(.A1(new_n15387_), .A2(new_n15378_), .Z(new_n15920_));
  AOI21_X1   g14918(.A1(new_n15386_), .A2(\A[660] ), .B(new_n15391_), .ZN(new_n15921_));
  XOR2_X1    g14919(.A1(new_n15921_), .A2(new_n15397_), .Z(new_n15922_));
  NOR2_X1    g14920(.A1(new_n15921_), .A2(new_n15397_), .ZN(new_n15923_));
  AOI21_X1   g14921(.A1(new_n15922_), .A2(new_n15400_), .B(new_n15923_), .ZN(new_n15924_));
  XOR2_X1    g14922(.A1(new_n15393_), .A2(new_n15397_), .Z(new_n15925_));
  NAND2_X1   g14923(.A1(new_n15925_), .A2(new_n15400_), .ZN(new_n15926_));
  INV_X1     g14924(.I(new_n15387_), .ZN(new_n15927_));
  NAND2_X1   g14925(.A1(new_n15927_), .A2(new_n15378_), .ZN(new_n15928_));
  NAND2_X1   g14926(.A1(new_n15922_), .A2(new_n15928_), .ZN(new_n15929_));
  NAND2_X1   g14927(.A1(new_n15926_), .A2(new_n15929_), .ZN(new_n15930_));
  OAI21_X1   g14928(.A1(new_n15920_), .A2(new_n15924_), .B(new_n15930_), .ZN(new_n15931_));
  AOI21_X1   g14929(.A1(new_n15354_), .A2(\A[666] ), .B(new_n15359_), .ZN(new_n15932_));
  XOR2_X1    g14930(.A1(new_n15932_), .A2(new_n15365_), .Z(new_n15933_));
  INV_X1     g14931(.I(new_n15355_), .ZN(new_n15934_));
  NAND2_X1   g14932(.A1(new_n15934_), .A2(new_n15346_), .ZN(new_n15935_));
  XOR2_X1    g14933(.A1(new_n15933_), .A2(new_n15935_), .Z(new_n15936_));
  INV_X1     g14934(.I(new_n15369_), .ZN(new_n15937_));
  NAND2_X1   g14935(.A1(new_n15356_), .A2(new_n15388_), .ZN(new_n15938_));
  NOR3_X1    g14936(.A1(new_n15936_), .A2(new_n15937_), .A3(new_n15938_), .ZN(new_n15939_));
  INV_X1     g14937(.I(new_n15401_), .ZN(new_n15940_));
  INV_X1     g14938(.I(new_n15356_), .ZN(new_n15941_));
  NOR2_X1    g14939(.A1(new_n15932_), .A2(new_n15365_), .ZN(new_n15942_));
  AOI21_X1   g14940(.A1(new_n15933_), .A2(new_n15368_), .B(new_n15942_), .ZN(new_n15943_));
  NOR2_X1    g14941(.A1(new_n15943_), .A2(new_n15941_), .ZN(new_n15944_));
  NOR2_X1    g14942(.A1(new_n15944_), .A2(new_n15940_), .ZN(new_n15945_));
  NAND2_X1   g14943(.A1(new_n15939_), .A2(new_n15945_), .ZN(new_n15946_));
  NOR3_X1    g14944(.A1(new_n15938_), .A2(new_n15937_), .A3(new_n15940_), .ZN(new_n15947_));
  INV_X1     g14945(.I(new_n15947_), .ZN(new_n15948_));
  XOR2_X1    g14946(.A1(new_n15933_), .A2(new_n15368_), .Z(new_n15949_));
  XOR2_X1    g14947(.A1(new_n15361_), .A2(new_n15365_), .Z(new_n15950_));
  INV_X1     g14948(.I(new_n15942_), .ZN(new_n15951_));
  OAI21_X1   g14949(.A1(new_n15950_), .A2(new_n15935_), .B(new_n15951_), .ZN(new_n15952_));
  NAND2_X1   g14950(.A1(new_n15952_), .A2(new_n15356_), .ZN(new_n15953_));
  NAND2_X1   g14951(.A1(new_n15949_), .A2(new_n15953_), .ZN(new_n15954_));
  NAND2_X1   g14952(.A1(new_n15948_), .A2(new_n15954_), .ZN(new_n15955_));
  AOI21_X1   g14953(.A1(new_n15946_), .A2(new_n15955_), .B(new_n15931_), .ZN(new_n15956_));
  INV_X1     g14954(.I(new_n15924_), .ZN(new_n15957_));
  AOI22_X1   g14955(.A1(new_n15957_), .A2(new_n15388_), .B1(new_n15926_), .B2(new_n15929_), .ZN(new_n15958_));
  NOR2_X1    g14956(.A1(new_n15936_), .A2(new_n15944_), .ZN(new_n15959_));
  NAND2_X1   g14957(.A1(new_n15948_), .A2(new_n15959_), .ZN(new_n15960_));
  NAND2_X1   g14958(.A1(new_n15954_), .A2(new_n15947_), .ZN(new_n15961_));
  AOI21_X1   g14959(.A1(new_n15960_), .A2(new_n15961_), .B(new_n15958_), .ZN(new_n15962_));
  NOR2_X1    g14960(.A1(new_n15956_), .A2(new_n15962_), .ZN(new_n15963_));
  XOR2_X1    g14961(.A1(new_n15322_), .A2(new_n15313_), .Z(new_n15964_));
  AOI21_X1   g14962(.A1(new_n15321_), .A2(\A[672] ), .B(new_n15326_), .ZN(new_n15965_));
  XOR2_X1    g14963(.A1(new_n15965_), .A2(new_n15332_), .Z(new_n15966_));
  NOR2_X1    g14964(.A1(new_n15965_), .A2(new_n15332_), .ZN(new_n15967_));
  AOI21_X1   g14965(.A1(new_n15966_), .A2(new_n15335_), .B(new_n15967_), .ZN(new_n15968_));
  XOR2_X1    g14966(.A1(new_n15328_), .A2(new_n15332_), .Z(new_n15969_));
  NAND2_X1   g14967(.A1(new_n15969_), .A2(new_n15335_), .ZN(new_n15970_));
  INV_X1     g14968(.I(new_n15322_), .ZN(new_n15971_));
  NAND2_X1   g14969(.A1(new_n15971_), .A2(new_n15313_), .ZN(new_n15972_));
  NAND2_X1   g14970(.A1(new_n15966_), .A2(new_n15972_), .ZN(new_n15973_));
  NAND2_X1   g14971(.A1(new_n15970_), .A2(new_n15973_), .ZN(new_n15974_));
  OAI21_X1   g14972(.A1(new_n15964_), .A2(new_n15968_), .B(new_n15974_), .ZN(new_n15975_));
  XOR2_X1    g14973(.A1(new_n15290_), .A2(new_n15281_), .Z(new_n15976_));
  XNOR2_X1   g14974(.A1(new_n15296_), .A2(new_n15300_), .ZN(new_n15977_));
  INV_X1     g14975(.I(new_n15290_), .ZN(new_n15978_));
  NAND2_X1   g14976(.A1(new_n15978_), .A2(new_n15281_), .ZN(new_n15979_));
  NOR2_X1    g14977(.A1(new_n15977_), .A2(new_n15979_), .ZN(new_n15980_));
  XOR2_X1    g14978(.A1(new_n15296_), .A2(new_n15300_), .Z(new_n15981_));
  NOR2_X1    g14979(.A1(new_n15981_), .A2(new_n15303_), .ZN(new_n15982_));
  NOR2_X1    g14980(.A1(new_n15980_), .A2(new_n15982_), .ZN(new_n15983_));
  NOR3_X1    g14981(.A1(new_n15983_), .A2(new_n15976_), .A3(new_n15964_), .ZN(new_n15984_));
  NAND2_X1   g14982(.A1(new_n15301_), .A2(new_n15296_), .ZN(new_n15985_));
  OAI21_X1   g14983(.A1(new_n15981_), .A2(new_n15979_), .B(new_n15985_), .ZN(new_n15986_));
  NAND2_X1   g14984(.A1(new_n15986_), .A2(new_n15291_), .ZN(new_n15987_));
  NAND4_X1   g14985(.A1(new_n15984_), .A2(new_n15304_), .A3(new_n15336_), .A4(new_n15987_), .ZN(new_n15988_));
  NOR2_X1    g14986(.A1(new_n15976_), .A2(new_n15964_), .ZN(new_n15989_));
  NAND3_X1   g14987(.A1(new_n15989_), .A2(new_n15304_), .A3(new_n15336_), .ZN(new_n15990_));
  NAND2_X1   g14988(.A1(new_n15981_), .A2(new_n15303_), .ZN(new_n15991_));
  NAND2_X1   g14989(.A1(new_n15977_), .A2(new_n15979_), .ZN(new_n15992_));
  AOI22_X1   g14990(.A1(new_n15986_), .A2(new_n15291_), .B1(new_n15992_), .B2(new_n15991_), .ZN(new_n15993_));
  INV_X1     g14991(.I(new_n15993_), .ZN(new_n15994_));
  NAND2_X1   g14992(.A1(new_n15994_), .A2(new_n15990_), .ZN(new_n15995_));
  AOI21_X1   g14993(.A1(new_n15988_), .A2(new_n15995_), .B(new_n15975_), .ZN(new_n15996_));
  INV_X1     g14994(.I(new_n15968_), .ZN(new_n15997_));
  NOR2_X1    g14995(.A1(new_n15966_), .A2(new_n15972_), .ZN(new_n15998_));
  NOR2_X1    g14996(.A1(new_n15969_), .A2(new_n15335_), .ZN(new_n15999_));
  NOR2_X1    g14997(.A1(new_n15999_), .A2(new_n15998_), .ZN(new_n16000_));
  AOI21_X1   g14998(.A1(new_n15323_), .A2(new_n15997_), .B(new_n16000_), .ZN(new_n16001_));
  AND4_X2    g14999(.A1(new_n15291_), .A2(new_n15304_), .A3(new_n15336_), .A4(new_n15323_), .Z(new_n16002_));
  NAND2_X1   g15000(.A1(new_n15994_), .A2(new_n16002_), .ZN(new_n16003_));
  NAND2_X1   g15001(.A1(new_n15993_), .A2(new_n15990_), .ZN(new_n16004_));
  AOI21_X1   g15002(.A1(new_n16003_), .A2(new_n16004_), .B(new_n16001_), .ZN(new_n16005_));
  XOR2_X1    g15003(.A1(new_n15305_), .A2(new_n15337_), .Z(new_n16006_));
  NAND2_X1   g15004(.A1(new_n16006_), .A2(new_n15403_), .ZN(new_n16007_));
  NOR3_X1    g15005(.A1(new_n15996_), .A2(new_n16005_), .A3(new_n16007_), .ZN(new_n16008_));
  NAND2_X1   g15006(.A1(new_n15992_), .A2(new_n15991_), .ZN(new_n16009_));
  NAND3_X1   g15007(.A1(new_n16009_), .A2(new_n15304_), .A3(new_n15989_), .ZN(new_n16010_));
  NAND2_X1   g15008(.A1(new_n15987_), .A2(new_n15336_), .ZN(new_n16011_));
  NOR2_X1    g15009(.A1(new_n16010_), .A2(new_n16011_), .ZN(new_n16012_));
  NOR2_X1    g15010(.A1(new_n15993_), .A2(new_n16002_), .ZN(new_n16013_));
  OAI21_X1   g15011(.A1(new_n16012_), .A2(new_n16013_), .B(new_n16001_), .ZN(new_n16014_));
  NOR2_X1    g15012(.A1(new_n15993_), .A2(new_n15990_), .ZN(new_n16015_));
  INV_X1     g15013(.I(new_n16004_), .ZN(new_n16016_));
  OAI21_X1   g15014(.A1(new_n16016_), .A2(new_n16015_), .B(new_n15975_), .ZN(new_n16017_));
  XNOR2_X1   g15015(.A1(new_n15370_), .A2(new_n15402_), .ZN(new_n16018_));
  NOR2_X1    g15016(.A1(new_n15338_), .A2(new_n16018_), .ZN(new_n16019_));
  AOI21_X1   g15017(.A1(new_n16017_), .A2(new_n16014_), .B(new_n16019_), .ZN(new_n16020_));
  OAI21_X1   g15018(.A1(new_n16008_), .A2(new_n16020_), .B(new_n15963_), .ZN(new_n16021_));
  NAND2_X1   g15019(.A1(new_n16017_), .A2(new_n16014_), .ZN(new_n16022_));
  NOR3_X1    g15020(.A1(new_n15996_), .A2(new_n16005_), .A3(new_n16019_), .ZN(new_n16023_));
  AOI21_X1   g15021(.A1(new_n16019_), .A2(new_n16022_), .B(new_n16023_), .ZN(new_n16024_));
  OAI21_X1   g15022(.A1(new_n15963_), .A2(new_n16024_), .B(new_n16021_), .ZN(new_n16025_));
  AOI21_X1   g15023(.A1(new_n15258_), .A2(\A[684] ), .B(new_n15263_), .ZN(new_n16026_));
  XOR2_X1    g15024(.A1(new_n16026_), .A2(new_n15267_), .Z(new_n16027_));
  NOR2_X1    g15025(.A1(new_n16026_), .A2(new_n15267_), .ZN(new_n16028_));
  AOI21_X1   g15026(.A1(new_n16027_), .A2(new_n15269_), .B(new_n16028_), .ZN(new_n16029_));
  INV_X1     g15027(.I(new_n16029_), .ZN(new_n16030_));
  XOR2_X1    g15028(.A1(new_n15265_), .A2(new_n15267_), .Z(new_n16031_));
  NAND2_X1   g15029(.A1(new_n16031_), .A2(new_n15269_), .ZN(new_n16032_));
  INV_X1     g15030(.I(new_n15269_), .ZN(new_n16033_));
  NAND2_X1   g15031(.A1(new_n16027_), .A2(new_n16033_), .ZN(new_n16034_));
  AOI22_X1   g15032(.A1(new_n16030_), .A2(new_n15260_), .B1(new_n16032_), .B2(new_n16034_), .ZN(new_n16035_));
  XOR2_X1    g15033(.A1(new_n15232_), .A2(new_n15236_), .Z(new_n16036_));
  NAND2_X1   g15034(.A1(new_n16036_), .A2(new_n15239_), .ZN(new_n16037_));
  AOI21_X1   g15035(.A1(new_n15225_), .A2(\A[690] ), .B(new_n15230_), .ZN(new_n16038_));
  XOR2_X1    g15036(.A1(new_n16038_), .A2(new_n15236_), .Z(new_n16039_));
  INV_X1     g15037(.I(new_n15226_), .ZN(new_n16040_));
  NAND2_X1   g15038(.A1(new_n16040_), .A2(new_n15217_), .ZN(new_n16041_));
  NAND2_X1   g15039(.A1(new_n16039_), .A2(new_n16041_), .ZN(new_n16042_));
  NAND2_X1   g15040(.A1(new_n16037_), .A2(new_n16042_), .ZN(new_n16043_));
  INV_X1     g15041(.I(new_n15227_), .ZN(new_n16044_));
  XNOR2_X1   g15042(.A1(new_n15250_), .A2(new_n15259_), .ZN(new_n16045_));
  NOR2_X1    g15043(.A1(new_n16044_), .A2(new_n16045_), .ZN(new_n16046_));
  NAND3_X1   g15044(.A1(new_n16046_), .A2(new_n16043_), .A3(new_n15240_), .ZN(new_n16047_));
  NOR2_X1    g15045(.A1(new_n16038_), .A2(new_n15236_), .ZN(new_n16048_));
  INV_X1     g15046(.I(new_n16048_), .ZN(new_n16049_));
  OAI21_X1   g15047(.A1(new_n16036_), .A2(new_n16041_), .B(new_n16049_), .ZN(new_n16050_));
  NAND2_X1   g15048(.A1(new_n16050_), .A2(new_n15227_), .ZN(new_n16051_));
  NAND2_X1   g15049(.A1(new_n16051_), .A2(new_n15270_), .ZN(new_n16052_));
  NOR2_X1    g15050(.A1(new_n16047_), .A2(new_n16052_), .ZN(new_n16053_));
  INV_X1     g15051(.I(new_n15240_), .ZN(new_n16054_));
  INV_X1     g15052(.I(new_n15270_), .ZN(new_n16055_));
  NOR4_X1    g15053(.A1(new_n16055_), .A2(new_n16054_), .A3(new_n16044_), .A4(new_n16045_), .ZN(new_n16056_));
  XOR2_X1    g15054(.A1(new_n16036_), .A2(new_n15239_), .Z(new_n16057_));
  AOI21_X1   g15055(.A1(new_n16039_), .A2(new_n15239_), .B(new_n16048_), .ZN(new_n16058_));
  NOR2_X1    g15056(.A1(new_n16058_), .A2(new_n16044_), .ZN(new_n16059_));
  NOR2_X1    g15057(.A1(new_n16057_), .A2(new_n16059_), .ZN(new_n16060_));
  NOR2_X1    g15058(.A1(new_n16060_), .A2(new_n16056_), .ZN(new_n16061_));
  OAI21_X1   g15059(.A1(new_n16061_), .A2(new_n16053_), .B(new_n16035_), .ZN(new_n16062_));
  NAND2_X1   g15060(.A1(new_n16032_), .A2(new_n16034_), .ZN(new_n16063_));
  OAI21_X1   g15061(.A1(new_n16045_), .A2(new_n16029_), .B(new_n16063_), .ZN(new_n16064_));
  NAND2_X1   g15062(.A1(new_n16051_), .A2(new_n16043_), .ZN(new_n16065_));
  NOR2_X1    g15063(.A1(new_n16065_), .A2(new_n16056_), .ZN(new_n16066_));
  NAND3_X1   g15064(.A1(new_n16046_), .A2(new_n15240_), .A3(new_n15270_), .ZN(new_n16067_));
  NOR2_X1    g15065(.A1(new_n16060_), .A2(new_n16067_), .ZN(new_n16068_));
  OAI21_X1   g15066(.A1(new_n16068_), .A2(new_n16066_), .B(new_n16064_), .ZN(new_n16069_));
  NAND2_X1   g15067(.A1(new_n16062_), .A2(new_n16069_), .ZN(new_n16070_));
  NAND2_X1   g15068(.A1(new_n15209_), .A2(new_n15272_), .ZN(new_n16071_));
  XOR2_X1    g15069(.A1(new_n15193_), .A2(new_n15184_), .Z(new_n16072_));
  AOI21_X1   g15070(.A1(new_n15192_), .A2(\A[696] ), .B(new_n15197_), .ZN(new_n16073_));
  XOR2_X1    g15071(.A1(new_n16073_), .A2(new_n15203_), .Z(new_n16074_));
  NOR2_X1    g15072(.A1(new_n16073_), .A2(new_n15203_), .ZN(new_n16075_));
  AOI21_X1   g15073(.A1(new_n16074_), .A2(new_n15206_), .B(new_n16075_), .ZN(new_n16076_));
  INV_X1     g15074(.I(new_n15193_), .ZN(new_n16077_));
  NAND2_X1   g15075(.A1(new_n16077_), .A2(new_n15184_), .ZN(new_n16078_));
  NOR2_X1    g15076(.A1(new_n16074_), .A2(new_n16078_), .ZN(new_n16079_));
  XOR2_X1    g15077(.A1(new_n15199_), .A2(new_n15203_), .Z(new_n16080_));
  NOR2_X1    g15078(.A1(new_n16080_), .A2(new_n15206_), .ZN(new_n16081_));
  OAI22_X1   g15079(.A1(new_n16072_), .A2(new_n16076_), .B1(new_n16079_), .B2(new_n16081_), .ZN(new_n16082_));
  INV_X1     g15080(.I(new_n16082_), .ZN(new_n16083_));
  XOR2_X1    g15081(.A1(new_n15167_), .A2(new_n15171_), .Z(new_n16084_));
  NAND2_X1   g15082(.A1(new_n16084_), .A2(new_n15174_), .ZN(new_n16085_));
  AOI21_X1   g15083(.A1(new_n15160_), .A2(\A[702] ), .B(new_n15165_), .ZN(new_n16086_));
  XOR2_X1    g15084(.A1(new_n16086_), .A2(new_n15171_), .Z(new_n16087_));
  INV_X1     g15085(.I(new_n15161_), .ZN(new_n16088_));
  NAND2_X1   g15086(.A1(new_n16088_), .A2(new_n15152_), .ZN(new_n16089_));
  NAND2_X1   g15087(.A1(new_n16087_), .A2(new_n16089_), .ZN(new_n16090_));
  NAND2_X1   g15088(.A1(new_n16085_), .A2(new_n16090_), .ZN(new_n16091_));
  XOR2_X1    g15089(.A1(new_n15161_), .A2(new_n15152_), .Z(new_n16092_));
  NOR2_X1    g15090(.A1(new_n16092_), .A2(new_n16072_), .ZN(new_n16093_));
  NAND3_X1   g15091(.A1(new_n16091_), .A2(new_n15175_), .A3(new_n16093_), .ZN(new_n16094_));
  NOR2_X1    g15092(.A1(new_n16086_), .A2(new_n15171_), .ZN(new_n16095_));
  INV_X1     g15093(.I(new_n16095_), .ZN(new_n16096_));
  OAI21_X1   g15094(.A1(new_n16084_), .A2(new_n16089_), .B(new_n16096_), .ZN(new_n16097_));
  NAND2_X1   g15095(.A1(new_n16097_), .A2(new_n15162_), .ZN(new_n16098_));
  NAND2_X1   g15096(.A1(new_n16098_), .A2(new_n15207_), .ZN(new_n16099_));
  NOR2_X1    g15097(.A1(new_n16094_), .A2(new_n16099_), .ZN(new_n16100_));
  AND4_X2    g15098(.A1(new_n15162_), .A2(new_n15175_), .A3(new_n15207_), .A4(new_n15194_), .Z(new_n16101_));
  NOR2_X1    g15099(.A1(new_n16087_), .A2(new_n16089_), .ZN(new_n16102_));
  NOR2_X1    g15100(.A1(new_n16084_), .A2(new_n15174_), .ZN(new_n16103_));
  NOR2_X1    g15101(.A1(new_n16103_), .A2(new_n16102_), .ZN(new_n16104_));
  AOI21_X1   g15102(.A1(new_n16087_), .A2(new_n15174_), .B(new_n16095_), .ZN(new_n16105_));
  NOR2_X1    g15103(.A1(new_n16105_), .A2(new_n16092_), .ZN(new_n16106_));
  NOR2_X1    g15104(.A1(new_n16106_), .A2(new_n16104_), .ZN(new_n16107_));
  NOR2_X1    g15105(.A1(new_n16107_), .A2(new_n16101_), .ZN(new_n16108_));
  OAI21_X1   g15106(.A1(new_n16108_), .A2(new_n16100_), .B(new_n16083_), .ZN(new_n16109_));
  NAND3_X1   g15107(.A1(new_n16093_), .A2(new_n15175_), .A3(new_n15207_), .ZN(new_n16110_));
  NOR2_X1    g15108(.A1(new_n16107_), .A2(new_n16110_), .ZN(new_n16111_));
  NOR3_X1    g15109(.A1(new_n16101_), .A2(new_n16104_), .A3(new_n16106_), .ZN(new_n16112_));
  OAI21_X1   g15110(.A1(new_n16111_), .A2(new_n16112_), .B(new_n16082_), .ZN(new_n16113_));
  AOI21_X1   g15111(.A1(new_n16109_), .A2(new_n16113_), .B(new_n16071_), .ZN(new_n16114_));
  XNOR2_X1   g15112(.A1(new_n15176_), .A2(new_n15208_), .ZN(new_n16115_));
  XNOR2_X1   g15113(.A1(new_n15241_), .A2(new_n15271_), .ZN(new_n16116_));
  NOR2_X1    g15114(.A1(new_n16115_), .A2(new_n16116_), .ZN(new_n16117_));
  NOR3_X1    g15115(.A1(new_n16104_), .A2(new_n16092_), .A3(new_n16072_), .ZN(new_n16118_));
  NAND4_X1   g15116(.A1(new_n16118_), .A2(new_n15175_), .A3(new_n15207_), .A4(new_n16098_), .ZN(new_n16119_));
  NAND2_X1   g15117(.A1(new_n16098_), .A2(new_n16091_), .ZN(new_n16120_));
  NAND2_X1   g15118(.A1(new_n16120_), .A2(new_n16110_), .ZN(new_n16121_));
  AOI21_X1   g15119(.A1(new_n16119_), .A2(new_n16121_), .B(new_n16082_), .ZN(new_n16122_));
  NAND2_X1   g15120(.A1(new_n16120_), .A2(new_n16101_), .ZN(new_n16123_));
  NAND2_X1   g15121(.A1(new_n16107_), .A2(new_n16110_), .ZN(new_n16124_));
  AOI21_X1   g15122(.A1(new_n16124_), .A2(new_n16123_), .B(new_n16083_), .ZN(new_n16125_));
  NOR3_X1    g15123(.A1(new_n16122_), .A2(new_n16125_), .A3(new_n16117_), .ZN(new_n16126_));
  OAI21_X1   g15124(.A1(new_n16126_), .A2(new_n16114_), .B(new_n16070_), .ZN(new_n16127_));
  NOR2_X1    g15125(.A1(new_n16059_), .A2(new_n16055_), .ZN(new_n16128_));
  NAND4_X1   g15126(.A1(new_n16128_), .A2(new_n16043_), .A3(new_n16058_), .A4(new_n16046_), .ZN(new_n16129_));
  NAND2_X1   g15127(.A1(new_n16067_), .A2(new_n16065_), .ZN(new_n16130_));
  AOI21_X1   g15128(.A1(new_n16129_), .A2(new_n16130_), .B(new_n16064_), .ZN(new_n16131_));
  NAND2_X1   g15129(.A1(new_n16060_), .A2(new_n16067_), .ZN(new_n16132_));
  NAND2_X1   g15130(.A1(new_n16065_), .A2(new_n16056_), .ZN(new_n16133_));
  AOI21_X1   g15131(.A1(new_n16132_), .A2(new_n16133_), .B(new_n16035_), .ZN(new_n16134_));
  NOR2_X1    g15132(.A1(new_n16131_), .A2(new_n16134_), .ZN(new_n16135_));
  AOI21_X1   g15133(.A1(new_n16109_), .A2(new_n16113_), .B(new_n16117_), .ZN(new_n16136_));
  NOR3_X1    g15134(.A1(new_n16122_), .A2(new_n16125_), .A3(new_n16071_), .ZN(new_n16137_));
  OAI21_X1   g15135(.A1(new_n16137_), .A2(new_n16136_), .B(new_n16135_), .ZN(new_n16138_));
  XOR2_X1    g15136(.A1(new_n16006_), .A2(new_n15403_), .Z(new_n16139_));
  AND2_X2    g15137(.A1(new_n16139_), .A2(new_n15273_), .Z(new_n16140_));
  NAND3_X1   g15138(.A1(new_n16140_), .A2(new_n16127_), .A3(new_n16138_), .ZN(new_n16141_));
  NAND2_X1   g15139(.A1(new_n16139_), .A2(new_n15273_), .ZN(new_n16142_));
  NAND2_X1   g15140(.A1(new_n16127_), .A2(new_n16138_), .ZN(new_n16143_));
  NAND2_X1   g15141(.A1(new_n16143_), .A2(new_n16142_), .ZN(new_n16144_));
  AOI21_X1   g15142(.A1(new_n16144_), .A2(new_n16141_), .B(new_n16025_), .ZN(new_n16145_));
  NOR2_X1    g15143(.A1(new_n15941_), .A2(new_n15920_), .ZN(new_n16146_));
  NAND3_X1   g15144(.A1(new_n15949_), .A2(new_n15369_), .A3(new_n16146_), .ZN(new_n16147_));
  NAND2_X1   g15145(.A1(new_n15953_), .A2(new_n15401_), .ZN(new_n16148_));
  NOR2_X1    g15146(.A1(new_n16147_), .A2(new_n16148_), .ZN(new_n16149_));
  NOR2_X1    g15147(.A1(new_n15959_), .A2(new_n15947_), .ZN(new_n16150_));
  OAI21_X1   g15148(.A1(new_n16149_), .A2(new_n16150_), .B(new_n15958_), .ZN(new_n16151_));
  NOR2_X1    g15149(.A1(new_n15954_), .A2(new_n15947_), .ZN(new_n16152_));
  NOR2_X1    g15150(.A1(new_n15948_), .A2(new_n15959_), .ZN(new_n16153_));
  OAI21_X1   g15151(.A1(new_n16153_), .A2(new_n16152_), .B(new_n15931_), .ZN(new_n16154_));
  NAND2_X1   g15152(.A1(new_n16154_), .A2(new_n16151_), .ZN(new_n16155_));
  NOR2_X1    g15153(.A1(new_n16008_), .A2(new_n16020_), .ZN(new_n16156_));
  NOR2_X1    g15154(.A1(new_n16156_), .A2(new_n16155_), .ZN(new_n16157_));
  NAND3_X1   g15155(.A1(new_n16017_), .A2(new_n16014_), .A3(new_n16007_), .ZN(new_n16158_));
  OAI21_X1   g15156(.A1(new_n15996_), .A2(new_n16005_), .B(new_n16019_), .ZN(new_n16159_));
  AOI21_X1   g15157(.A1(new_n16158_), .A2(new_n16159_), .B(new_n15963_), .ZN(new_n16160_));
  NOR2_X1    g15158(.A1(new_n16157_), .A2(new_n16160_), .ZN(new_n16161_));
  NAND3_X1   g15159(.A1(new_n16127_), .A2(new_n16138_), .A3(new_n16142_), .ZN(new_n16162_));
  OAI21_X1   g15160(.A1(new_n16122_), .A2(new_n16125_), .B(new_n16117_), .ZN(new_n16163_));
  NAND3_X1   g15161(.A1(new_n16109_), .A2(new_n16113_), .A3(new_n16071_), .ZN(new_n16164_));
  AOI21_X1   g15162(.A1(new_n16163_), .A2(new_n16164_), .B(new_n16135_), .ZN(new_n16165_));
  OAI21_X1   g15163(.A1(new_n16122_), .A2(new_n16125_), .B(new_n16071_), .ZN(new_n16166_));
  NAND3_X1   g15164(.A1(new_n16109_), .A2(new_n16113_), .A3(new_n16117_), .ZN(new_n16167_));
  AOI21_X1   g15165(.A1(new_n16166_), .A2(new_n16167_), .B(new_n16070_), .ZN(new_n16168_));
  OAI21_X1   g15166(.A1(new_n16165_), .A2(new_n16168_), .B(new_n16140_), .ZN(new_n16169_));
  AOI21_X1   g15167(.A1(new_n16162_), .A2(new_n16169_), .B(new_n16161_), .ZN(new_n16170_));
  OR2_X2     g15168(.A1(new_n16145_), .A2(new_n16170_), .Z(new_n16171_));
  XOR2_X1    g15169(.A1(new_n15132_), .A2(new_n15136_), .Z(new_n16172_));
  NAND2_X1   g15170(.A1(new_n16172_), .A2(new_n15139_), .ZN(new_n16173_));
  AOI21_X1   g15171(.A1(new_n15125_), .A2(\A[708] ), .B(new_n15130_), .ZN(new_n16174_));
  XOR2_X1    g15172(.A1(new_n16174_), .A2(new_n15136_), .Z(new_n16175_));
  INV_X1     g15173(.I(new_n15126_), .ZN(new_n16176_));
  NAND2_X1   g15174(.A1(new_n16176_), .A2(new_n15117_), .ZN(new_n16177_));
  NAND2_X1   g15175(.A1(new_n16175_), .A2(new_n16177_), .ZN(new_n16178_));
  NAND2_X1   g15176(.A1(new_n16173_), .A2(new_n16178_), .ZN(new_n16179_));
  NAND2_X1   g15177(.A1(new_n15137_), .A2(new_n15132_), .ZN(new_n16180_));
  OAI21_X1   g15178(.A1(new_n16172_), .A2(new_n16177_), .B(new_n16180_), .ZN(new_n16181_));
  NAND2_X1   g15179(.A1(new_n16181_), .A2(new_n15127_), .ZN(new_n16182_));
  NAND2_X1   g15180(.A1(new_n16182_), .A2(new_n16179_), .ZN(new_n16183_));
  XOR2_X1    g15181(.A1(new_n15100_), .A2(new_n15104_), .Z(new_n16184_));
  XOR2_X1    g15182(.A1(new_n16184_), .A2(new_n15107_), .Z(new_n16185_));
  INV_X1     g15183(.I(new_n15108_), .ZN(new_n16186_));
  NAND2_X1   g15184(.A1(new_n15095_), .A2(new_n15127_), .ZN(new_n16187_));
  NOR3_X1    g15185(.A1(new_n16185_), .A2(new_n16186_), .A3(new_n16187_), .ZN(new_n16188_));
  INV_X1     g15186(.I(new_n15140_), .ZN(new_n16189_));
  INV_X1     g15187(.I(new_n15095_), .ZN(new_n16190_));
  AOI21_X1   g15188(.A1(new_n15093_), .A2(\A[714] ), .B(new_n15098_), .ZN(new_n16191_));
  XOR2_X1    g15189(.A1(new_n16191_), .A2(new_n15104_), .Z(new_n16192_));
  NOR2_X1    g15190(.A1(new_n16191_), .A2(new_n15104_), .ZN(new_n16193_));
  AOI21_X1   g15191(.A1(new_n16192_), .A2(new_n15107_), .B(new_n16193_), .ZN(new_n16194_));
  NOR2_X1    g15192(.A1(new_n16194_), .A2(new_n16190_), .ZN(new_n16195_));
  NOR2_X1    g15193(.A1(new_n16195_), .A2(new_n16189_), .ZN(new_n16196_));
  NAND2_X1   g15194(.A1(new_n16188_), .A2(new_n16196_), .ZN(new_n16197_));
  XOR2_X1    g15195(.A1(new_n15126_), .A2(new_n15117_), .Z(new_n16198_));
  NOR2_X1    g15196(.A1(new_n16190_), .A2(new_n16198_), .ZN(new_n16199_));
  NAND3_X1   g15197(.A1(new_n16199_), .A2(new_n15108_), .A3(new_n15140_), .ZN(new_n16200_));
  NAND2_X1   g15198(.A1(new_n16184_), .A2(new_n15107_), .ZN(new_n16201_));
  INV_X1     g15199(.I(new_n15094_), .ZN(new_n16202_));
  NAND2_X1   g15200(.A1(new_n16202_), .A2(new_n15085_), .ZN(new_n16203_));
  NAND2_X1   g15201(.A1(new_n16192_), .A2(new_n16203_), .ZN(new_n16204_));
  NAND2_X1   g15202(.A1(new_n16201_), .A2(new_n16204_), .ZN(new_n16205_));
  INV_X1     g15203(.I(new_n16193_), .ZN(new_n16206_));
  OAI21_X1   g15204(.A1(new_n16184_), .A2(new_n16203_), .B(new_n16206_), .ZN(new_n16207_));
  NAND2_X1   g15205(.A1(new_n16207_), .A2(new_n15095_), .ZN(new_n16208_));
  NAND2_X1   g15206(.A1(new_n16208_), .A2(new_n16205_), .ZN(new_n16209_));
  NAND2_X1   g15207(.A1(new_n16200_), .A2(new_n16209_), .ZN(new_n16210_));
  AOI21_X1   g15208(.A1(new_n16197_), .A2(new_n16210_), .B(new_n16183_), .ZN(new_n16211_));
  AOI22_X1   g15209(.A1(new_n16181_), .A2(new_n15127_), .B1(new_n16173_), .B2(new_n16178_), .ZN(new_n16212_));
  NOR2_X1    g15210(.A1(new_n16185_), .A2(new_n16195_), .ZN(new_n16213_));
  NAND2_X1   g15211(.A1(new_n16213_), .A2(new_n16200_), .ZN(new_n16214_));
  NOR3_X1    g15212(.A1(new_n16187_), .A2(new_n16186_), .A3(new_n16189_), .ZN(new_n16215_));
  NAND2_X1   g15213(.A1(new_n16209_), .A2(new_n16215_), .ZN(new_n16216_));
  AOI21_X1   g15214(.A1(new_n16214_), .A2(new_n16216_), .B(new_n16212_), .ZN(new_n16217_));
  NOR2_X1    g15215(.A1(new_n16211_), .A2(new_n16217_), .ZN(new_n16218_));
  XNOR2_X1   g15216(.A1(new_n15038_), .A2(new_n15046_), .ZN(new_n16219_));
  XOR2_X1    g15217(.A1(new_n15049_), .A2(new_n15051_), .Z(new_n16220_));
  NOR2_X1    g15218(.A1(new_n15038_), .A2(new_n15046_), .ZN(new_n16221_));
  NOR2_X1    g15219(.A1(new_n15049_), .A2(new_n15051_), .ZN(new_n16222_));
  AOI21_X1   g15220(.A1(new_n16220_), .A2(new_n16221_), .B(new_n16222_), .ZN(new_n16223_));
  INV_X1     g15221(.I(new_n16221_), .ZN(new_n16224_));
  NOR2_X1    g15222(.A1(new_n16220_), .A2(new_n16224_), .ZN(new_n16225_));
  XNOR2_X1   g15223(.A1(new_n15049_), .A2(new_n15051_), .ZN(new_n16226_));
  NOR2_X1    g15224(.A1(new_n16226_), .A2(new_n16221_), .ZN(new_n16227_));
  OAI22_X1   g15225(.A1(new_n16219_), .A2(new_n16223_), .B1(new_n16227_), .B2(new_n16225_), .ZN(new_n16228_));
  XNOR2_X1   g15226(.A1(new_n15072_), .A2(new_n15074_), .ZN(new_n16229_));
  NOR2_X1    g15227(.A1(new_n15061_), .A2(new_n15069_), .ZN(new_n16230_));
  NAND2_X1   g15228(.A1(new_n16229_), .A2(new_n16230_), .ZN(new_n16231_));
  XOR2_X1    g15229(.A1(new_n15072_), .A2(new_n15074_), .Z(new_n16232_));
  INV_X1     g15230(.I(new_n16230_), .ZN(new_n16233_));
  NAND2_X1   g15231(.A1(new_n16232_), .A2(new_n16233_), .ZN(new_n16234_));
  NAND2_X1   g15232(.A1(new_n16231_), .A2(new_n16234_), .ZN(new_n16235_));
  XNOR2_X1   g15233(.A1(new_n15061_), .A2(new_n15069_), .ZN(new_n16236_));
  NOR2_X1    g15234(.A1(new_n16219_), .A2(new_n16236_), .ZN(new_n16237_));
  NOR2_X1    g15235(.A1(new_n15072_), .A2(new_n15074_), .ZN(new_n16238_));
  INV_X1     g15236(.I(new_n16238_), .ZN(new_n16239_));
  OAI21_X1   g15237(.A1(new_n16229_), .A2(new_n16233_), .B(new_n16239_), .ZN(new_n16240_));
  OAI21_X1   g15238(.A1(new_n16235_), .A2(new_n15070_), .B(new_n16240_), .ZN(new_n16241_));
  NAND4_X1   g15239(.A1(new_n16241_), .A2(new_n15052_), .A3(new_n16235_), .A4(new_n16237_), .ZN(new_n16242_));
  AND4_X2    g15240(.A1(new_n15047_), .A2(new_n15070_), .A3(new_n15052_), .A4(new_n15075_), .Z(new_n16243_));
  AOI22_X1   g15241(.A1(new_n16240_), .A2(new_n15070_), .B1(new_n16231_), .B2(new_n16234_), .ZN(new_n16244_));
  NOR2_X1    g15242(.A1(new_n16244_), .A2(new_n16243_), .ZN(new_n16245_));
  INV_X1     g15243(.I(new_n16245_), .ZN(new_n16246_));
  AOI21_X1   g15244(.A1(new_n16242_), .A2(new_n16246_), .B(new_n16228_), .ZN(new_n16247_));
  INV_X1     g15245(.I(new_n16223_), .ZN(new_n16248_));
  NAND2_X1   g15246(.A1(new_n16226_), .A2(new_n16221_), .ZN(new_n16249_));
  NAND2_X1   g15247(.A1(new_n16220_), .A2(new_n16224_), .ZN(new_n16250_));
  AOI22_X1   g15248(.A1(new_n16248_), .A2(new_n15047_), .B1(new_n16249_), .B2(new_n16250_), .ZN(new_n16251_));
  NAND3_X1   g15249(.A1(new_n16237_), .A2(new_n15052_), .A3(new_n15075_), .ZN(new_n16252_));
  NAND2_X1   g15250(.A1(new_n16244_), .A2(new_n16252_), .ZN(new_n16253_));
  NAND2_X1   g15251(.A1(new_n16240_), .A2(new_n15070_), .ZN(new_n16254_));
  NAND2_X1   g15252(.A1(new_n16254_), .A2(new_n16235_), .ZN(new_n16255_));
  NAND2_X1   g15253(.A1(new_n16255_), .A2(new_n16243_), .ZN(new_n16256_));
  AOI21_X1   g15254(.A1(new_n16256_), .A2(new_n16253_), .B(new_n16251_), .ZN(new_n16257_));
  NAND2_X1   g15255(.A1(new_n15142_), .A2(new_n15077_), .ZN(new_n16258_));
  NOR3_X1    g15256(.A1(new_n16247_), .A2(new_n16257_), .A3(new_n16258_), .ZN(new_n16259_));
  NAND3_X1   g15257(.A1(new_n16235_), .A2(new_n15052_), .A3(new_n16237_), .ZN(new_n16260_));
  NAND2_X1   g15258(.A1(new_n16254_), .A2(new_n15075_), .ZN(new_n16261_));
  NOR2_X1    g15259(.A1(new_n16260_), .A2(new_n16261_), .ZN(new_n16262_));
  OAI21_X1   g15260(.A1(new_n16262_), .A2(new_n16245_), .B(new_n16251_), .ZN(new_n16263_));
  NOR2_X1    g15261(.A1(new_n16255_), .A2(new_n16243_), .ZN(new_n16264_));
  NOR2_X1    g15262(.A1(new_n16244_), .A2(new_n16252_), .ZN(new_n16265_));
  OAI21_X1   g15263(.A1(new_n16264_), .A2(new_n16265_), .B(new_n16228_), .ZN(new_n16266_));
  XNOR2_X1   g15264(.A1(new_n15053_), .A2(new_n15076_), .ZN(new_n16267_));
  XNOR2_X1   g15265(.A1(new_n15109_), .A2(new_n15141_), .ZN(new_n16268_));
  NOR2_X1    g15266(.A1(new_n16268_), .A2(new_n16267_), .ZN(new_n16269_));
  AOI21_X1   g15267(.A1(new_n16263_), .A2(new_n16266_), .B(new_n16269_), .ZN(new_n16270_));
  OAI21_X1   g15268(.A1(new_n16259_), .A2(new_n16270_), .B(new_n16218_), .ZN(new_n16271_));
  NAND3_X1   g15269(.A1(new_n16199_), .A2(new_n16205_), .A3(new_n15108_), .ZN(new_n16272_));
  NAND2_X1   g15270(.A1(new_n16208_), .A2(new_n15140_), .ZN(new_n16273_));
  NOR2_X1    g15271(.A1(new_n16272_), .A2(new_n16273_), .ZN(new_n16274_));
  NOR2_X1    g15272(.A1(new_n16213_), .A2(new_n16215_), .ZN(new_n16275_));
  OAI21_X1   g15273(.A1(new_n16275_), .A2(new_n16274_), .B(new_n16212_), .ZN(new_n16276_));
  NOR2_X1    g15274(.A1(new_n16209_), .A2(new_n16215_), .ZN(new_n16277_));
  NOR2_X1    g15275(.A1(new_n16213_), .A2(new_n16200_), .ZN(new_n16278_));
  OAI21_X1   g15276(.A1(new_n16278_), .A2(new_n16277_), .B(new_n16183_), .ZN(new_n16279_));
  NAND2_X1   g15277(.A1(new_n16276_), .A2(new_n16279_), .ZN(new_n16280_));
  NOR3_X1    g15278(.A1(new_n16247_), .A2(new_n16257_), .A3(new_n16269_), .ZN(new_n16281_));
  AOI21_X1   g15279(.A1(new_n16263_), .A2(new_n16266_), .B(new_n16258_), .ZN(new_n16282_));
  OAI21_X1   g15280(.A1(new_n16281_), .A2(new_n16282_), .B(new_n16280_), .ZN(new_n16283_));
  NAND2_X1   g15281(.A1(new_n16283_), .A2(new_n16271_), .ZN(new_n16284_));
  XOR2_X1    g15282(.A1(new_n14995_), .A2(new_n14990_), .Z(new_n16285_));
  INV_X1     g15283(.I(new_n14987_), .ZN(new_n16286_));
  NAND2_X1   g15284(.A1(new_n16286_), .A2(new_n14979_), .ZN(new_n16287_));
  NAND2_X1   g15285(.A1(new_n14974_), .A2(\A[728] ), .ZN(new_n16288_));
  NAND2_X1   g15286(.A1(new_n14977_), .A2(new_n16288_), .ZN(new_n16289_));
  AOI21_X1   g15287(.A1(new_n16289_), .A2(\A[729] ), .B(new_n14993_), .ZN(new_n16290_));
  NOR2_X1    g15288(.A1(new_n14990_), .A2(new_n16290_), .ZN(new_n16291_));
  INV_X1     g15289(.I(new_n16291_), .ZN(new_n16292_));
  OAI21_X1   g15290(.A1(new_n16285_), .A2(new_n16287_), .B(new_n16292_), .ZN(new_n16293_));
  NAND2_X1   g15291(.A1(new_n16285_), .A2(new_n14997_), .ZN(new_n16294_));
  XOR2_X1    g15292(.A1(new_n14990_), .A2(new_n16290_), .Z(new_n16295_));
  NAND2_X1   g15293(.A1(new_n16295_), .A2(new_n16287_), .ZN(new_n16296_));
  AOI22_X1   g15294(.A1(new_n16293_), .A2(new_n14988_), .B1(new_n16294_), .B2(new_n16296_), .ZN(new_n16297_));
  INV_X1     g15295(.I(new_n14998_), .ZN(new_n16298_));
  AOI21_X1   g15296(.A1(new_n15005_), .A2(\A[735] ), .B(new_n15023_), .ZN(new_n16299_));
  XOR2_X1    g15297(.A1(new_n15019_), .A2(new_n16299_), .Z(new_n16300_));
  INV_X1     g15298(.I(new_n15026_), .ZN(new_n16301_));
  NOR2_X1    g15299(.A1(new_n16300_), .A2(new_n16301_), .ZN(new_n16302_));
  XOR2_X1    g15300(.A1(new_n15025_), .A2(new_n15019_), .Z(new_n16303_));
  NOR2_X1    g15301(.A1(new_n16303_), .A2(new_n15026_), .ZN(new_n16304_));
  NOR2_X1    g15302(.A1(new_n16304_), .A2(new_n16302_), .ZN(new_n16305_));
  NAND2_X1   g15303(.A1(new_n14988_), .A2(new_n15017_), .ZN(new_n16306_));
  NOR2_X1    g15304(.A1(new_n15019_), .A2(new_n16299_), .ZN(new_n16307_));
  INV_X1     g15305(.I(new_n16307_), .ZN(new_n16308_));
  OAI21_X1   g15306(.A1(new_n16303_), .A2(new_n16301_), .B(new_n16308_), .ZN(new_n16309_));
  NAND2_X1   g15307(.A1(new_n16309_), .A2(new_n15017_), .ZN(new_n16310_));
  NAND2_X1   g15308(.A1(new_n16310_), .A2(new_n15027_), .ZN(new_n16311_));
  NOR4_X1    g15309(.A1(new_n16311_), .A2(new_n16298_), .A3(new_n16305_), .A4(new_n16306_), .ZN(new_n16312_));
  NAND4_X1   g15310(.A1(new_n14998_), .A2(new_n14988_), .A3(new_n15017_), .A4(new_n15027_), .ZN(new_n16313_));
  INV_X1     g15311(.I(new_n16313_), .ZN(new_n16314_));
  NAND2_X1   g15312(.A1(new_n16303_), .A2(new_n15026_), .ZN(new_n16315_));
  NAND2_X1   g15313(.A1(new_n16300_), .A2(new_n16301_), .ZN(new_n16316_));
  AOI22_X1   g15314(.A1(new_n16309_), .A2(new_n15017_), .B1(new_n16315_), .B2(new_n16316_), .ZN(new_n16317_));
  NOR2_X1    g15315(.A1(new_n16317_), .A2(new_n16314_), .ZN(new_n16318_));
  OAI21_X1   g15316(.A1(new_n16312_), .A2(new_n16318_), .B(new_n16297_), .ZN(new_n16319_));
  INV_X1     g15317(.I(new_n16297_), .ZN(new_n16320_));
  NOR2_X1    g15318(.A1(new_n16317_), .A2(new_n16313_), .ZN(new_n16321_));
  NAND2_X1   g15319(.A1(new_n16315_), .A2(new_n16316_), .ZN(new_n16322_));
  NAND2_X1   g15320(.A1(new_n16310_), .A2(new_n16322_), .ZN(new_n16323_));
  NOR2_X1    g15321(.A1(new_n16323_), .A2(new_n16314_), .ZN(new_n16324_));
  OAI21_X1   g15322(.A1(new_n16324_), .A2(new_n16321_), .B(new_n16320_), .ZN(new_n16325_));
  NAND2_X1   g15323(.A1(new_n16319_), .A2(new_n16325_), .ZN(new_n16326_));
  NAND2_X1   g15324(.A1(new_n14971_), .A2(new_n15029_), .ZN(new_n16327_));
  AOI21_X1   g15325(.A1(new_n14920_), .A2(\A[741] ), .B(new_n14936_), .ZN(new_n16328_));
  XNOR2_X1   g15326(.A1(new_n14933_), .A2(new_n16328_), .ZN(new_n16329_));
  INV_X1     g15327(.I(new_n14939_), .ZN(new_n16330_));
  NOR2_X1    g15328(.A1(new_n14933_), .A2(new_n16328_), .ZN(new_n16331_));
  INV_X1     g15329(.I(new_n16331_), .ZN(new_n16332_));
  OAI21_X1   g15330(.A1(new_n16329_), .A2(new_n16330_), .B(new_n16332_), .ZN(new_n16333_));
  NAND2_X1   g15331(.A1(new_n14934_), .A2(new_n16328_), .ZN(new_n16334_));
  NAND2_X1   g15332(.A1(new_n14938_), .A2(new_n14933_), .ZN(new_n16335_));
  NAND3_X1   g15333(.A1(new_n16334_), .A2(new_n16335_), .A3(new_n14939_), .ZN(new_n16336_));
  NAND2_X1   g15334(.A1(new_n16334_), .A2(new_n16335_), .ZN(new_n16337_));
  NAND2_X1   g15335(.A1(new_n16337_), .A2(new_n16330_), .ZN(new_n16338_));
  AOI22_X1   g15336(.A1(new_n16333_), .A2(new_n14931_), .B1(new_n16338_), .B2(new_n16336_), .ZN(new_n16339_));
  AOI21_X1   g15337(.A1(new_n14955_), .A2(\A[750] ), .B(new_n14960_), .ZN(new_n16340_));
  XOR2_X1    g15338(.A1(new_n14966_), .A2(new_n16340_), .Z(new_n16341_));
  NAND2_X1   g15339(.A1(new_n16341_), .A2(new_n14968_), .ZN(new_n16342_));
  NAND2_X1   g15340(.A1(new_n14966_), .A2(new_n16340_), .ZN(new_n16343_));
  NAND2_X1   g15341(.A1(new_n14944_), .A2(\A[746] ), .ZN(new_n16344_));
  NAND2_X1   g15342(.A1(new_n14947_), .A2(new_n16344_), .ZN(new_n16345_));
  AOI21_X1   g15343(.A1(new_n16345_), .A2(\A[747] ), .B(new_n14964_), .ZN(new_n16346_));
  NAND2_X1   g15344(.A1(new_n14962_), .A2(new_n16346_), .ZN(new_n16347_));
  NAND2_X1   g15345(.A1(new_n16347_), .A2(new_n16343_), .ZN(new_n16348_));
  INV_X1     g15346(.I(new_n14957_), .ZN(new_n16349_));
  NAND2_X1   g15347(.A1(new_n16349_), .A2(new_n14949_), .ZN(new_n16350_));
  NAND2_X1   g15348(.A1(new_n16348_), .A2(new_n16350_), .ZN(new_n16351_));
  NAND2_X1   g15349(.A1(new_n16342_), .A2(new_n16351_), .ZN(new_n16352_));
  XNOR2_X1   g15350(.A1(new_n14922_), .A2(new_n14930_), .ZN(new_n16353_));
  XOR2_X1    g15351(.A1(new_n14949_), .A2(new_n14957_), .Z(new_n16354_));
  NOR2_X1    g15352(.A1(new_n16353_), .A2(new_n16354_), .ZN(new_n16355_));
  NAND3_X1   g15353(.A1(new_n16352_), .A2(new_n14940_), .A3(new_n16355_), .ZN(new_n16356_));
  NOR2_X1    g15354(.A1(new_n16340_), .A2(new_n16346_), .ZN(new_n16357_));
  INV_X1     g15355(.I(new_n16357_), .ZN(new_n16358_));
  OAI21_X1   g15356(.A1(new_n16341_), .A2(new_n16350_), .B(new_n16358_), .ZN(new_n16359_));
  NAND2_X1   g15357(.A1(new_n16359_), .A2(new_n14958_), .ZN(new_n16360_));
  NAND2_X1   g15358(.A1(new_n16360_), .A2(new_n14969_), .ZN(new_n16361_));
  NOR2_X1    g15359(.A1(new_n16356_), .A2(new_n16361_), .ZN(new_n16362_));
  AND4_X2    g15360(.A1(new_n14931_), .A2(new_n14969_), .A3(new_n14940_), .A4(new_n14958_), .Z(new_n16363_));
  AOI22_X1   g15361(.A1(new_n16359_), .A2(new_n14958_), .B1(new_n16342_), .B2(new_n16351_), .ZN(new_n16364_));
  NOR2_X1    g15362(.A1(new_n16363_), .A2(new_n16364_), .ZN(new_n16365_));
  OAI21_X1   g15363(.A1(new_n16362_), .A2(new_n16365_), .B(new_n16339_), .ZN(new_n16366_));
  AOI21_X1   g15364(.A1(new_n16337_), .A2(new_n14939_), .B(new_n16331_), .ZN(new_n16367_));
  INV_X1     g15365(.I(new_n16336_), .ZN(new_n16368_));
  NOR2_X1    g15366(.A1(new_n16329_), .A2(new_n14939_), .ZN(new_n16369_));
  OAI22_X1   g15367(.A1(new_n16367_), .A2(new_n16353_), .B1(new_n16369_), .B2(new_n16368_), .ZN(new_n16370_));
  NAND2_X1   g15368(.A1(new_n16360_), .A2(new_n16352_), .ZN(new_n16371_));
  NOR2_X1    g15369(.A1(new_n16371_), .A2(new_n16363_), .ZN(new_n16372_));
  NAND3_X1   g15370(.A1(new_n16355_), .A2(new_n14940_), .A3(new_n14969_), .ZN(new_n16373_));
  NOR2_X1    g15371(.A1(new_n16364_), .A2(new_n16373_), .ZN(new_n16374_));
  OAI21_X1   g15372(.A1(new_n16372_), .A2(new_n16374_), .B(new_n16370_), .ZN(new_n16375_));
  AOI21_X1   g15373(.A1(new_n16366_), .A2(new_n16375_), .B(new_n16327_), .ZN(new_n16376_));
  XNOR2_X1   g15374(.A1(new_n14970_), .A2(new_n14941_), .ZN(new_n16377_));
  XNOR2_X1   g15375(.A1(new_n14999_), .A2(new_n15028_), .ZN(new_n16378_));
  NOR2_X1    g15376(.A1(new_n16377_), .A2(new_n16378_), .ZN(new_n16379_));
  OAI21_X1   g15377(.A1(new_n16352_), .A2(new_n14958_), .B(new_n16359_), .ZN(new_n16380_));
  NAND4_X1   g15378(.A1(new_n16380_), .A2(new_n14940_), .A3(new_n16352_), .A4(new_n16355_), .ZN(new_n16381_));
  NAND2_X1   g15379(.A1(new_n16371_), .A2(new_n16373_), .ZN(new_n16382_));
  AOI21_X1   g15380(.A1(new_n16381_), .A2(new_n16382_), .B(new_n16370_), .ZN(new_n16383_));
  NAND2_X1   g15381(.A1(new_n16364_), .A2(new_n16373_), .ZN(new_n16384_));
  NAND2_X1   g15382(.A1(new_n16371_), .A2(new_n16363_), .ZN(new_n16385_));
  AOI21_X1   g15383(.A1(new_n16385_), .A2(new_n16384_), .B(new_n16339_), .ZN(new_n16386_));
  NOR3_X1    g15384(.A1(new_n16383_), .A2(new_n16386_), .A3(new_n16379_), .ZN(new_n16387_));
  OAI21_X1   g15385(.A1(new_n16387_), .A2(new_n16376_), .B(new_n16326_), .ZN(new_n16388_));
  NOR2_X1    g15386(.A1(new_n16305_), .A2(new_n16306_), .ZN(new_n16389_));
  NAND4_X1   g15387(.A1(new_n16389_), .A2(new_n14998_), .A3(new_n15027_), .A4(new_n16310_), .ZN(new_n16390_));
  NAND2_X1   g15388(.A1(new_n16323_), .A2(new_n16313_), .ZN(new_n16391_));
  AOI21_X1   g15389(.A1(new_n16390_), .A2(new_n16391_), .B(new_n16320_), .ZN(new_n16392_));
  NAND2_X1   g15390(.A1(new_n16323_), .A2(new_n16314_), .ZN(new_n16393_));
  NAND2_X1   g15391(.A1(new_n16317_), .A2(new_n16313_), .ZN(new_n16394_));
  AOI21_X1   g15392(.A1(new_n16393_), .A2(new_n16394_), .B(new_n16297_), .ZN(new_n16395_));
  NOR2_X1    g15393(.A1(new_n16392_), .A2(new_n16395_), .ZN(new_n16396_));
  AOI21_X1   g15394(.A1(new_n16366_), .A2(new_n16375_), .B(new_n16379_), .ZN(new_n16397_));
  NOR3_X1    g15395(.A1(new_n16383_), .A2(new_n16386_), .A3(new_n16327_), .ZN(new_n16398_));
  OAI21_X1   g15396(.A1(new_n16398_), .A2(new_n16397_), .B(new_n16396_), .ZN(new_n16399_));
  NAND2_X1   g15397(.A1(new_n15143_), .A2(new_n15030_), .ZN(new_n16400_));
  NAND3_X1   g15398(.A1(new_n16399_), .A2(new_n16388_), .A3(new_n16400_), .ZN(new_n16401_));
  INV_X1     g15399(.I(new_n16400_), .ZN(new_n16402_));
  NAND2_X1   g15400(.A1(new_n16399_), .A2(new_n16388_), .ZN(new_n16403_));
  NAND2_X1   g15401(.A1(new_n16403_), .A2(new_n16402_), .ZN(new_n16404_));
  NAND2_X1   g15402(.A1(new_n16404_), .A2(new_n16401_), .ZN(new_n16405_));
  NAND2_X1   g15403(.A1(new_n16405_), .A2(new_n16284_), .ZN(new_n16406_));
  INV_X1     g15404(.I(new_n16284_), .ZN(new_n16407_));
  NAND3_X1   g15405(.A1(new_n16402_), .A2(new_n16388_), .A3(new_n16399_), .ZN(new_n16408_));
  INV_X1     g15406(.I(new_n16408_), .ZN(new_n16409_));
  AOI21_X1   g15407(.A1(new_n16399_), .A2(new_n16388_), .B(new_n16402_), .ZN(new_n16410_));
  OAI21_X1   g15408(.A1(new_n16409_), .A2(new_n16410_), .B(new_n16407_), .ZN(new_n16411_));
  NOR2_X1    g15409(.A1(new_n15144_), .A2(new_n15405_), .ZN(new_n16412_));
  NAND3_X1   g15410(.A1(new_n16406_), .A2(new_n16411_), .A3(new_n16412_), .ZN(new_n16413_));
  AOI21_X1   g15411(.A1(new_n16401_), .A2(new_n16404_), .B(new_n16407_), .ZN(new_n16414_));
  NAND2_X1   g15412(.A1(new_n16403_), .A2(new_n16400_), .ZN(new_n16415_));
  AOI21_X1   g15413(.A1(new_n16415_), .A2(new_n16408_), .B(new_n16284_), .ZN(new_n16416_));
  INV_X1     g15414(.I(new_n16412_), .ZN(new_n16417_));
  OAI21_X1   g15415(.A1(new_n16414_), .A2(new_n16416_), .B(new_n16417_), .ZN(new_n16418_));
  AOI21_X1   g15416(.A1(new_n16418_), .A2(new_n16413_), .B(new_n16171_), .ZN(new_n16419_));
  NOR2_X1    g15417(.A1(new_n16145_), .A2(new_n16170_), .ZN(new_n16420_));
  NAND3_X1   g15418(.A1(new_n16406_), .A2(new_n16411_), .A3(new_n16417_), .ZN(new_n16421_));
  OAI21_X1   g15419(.A1(new_n16414_), .A2(new_n16416_), .B(new_n16412_), .ZN(new_n16422_));
  AOI21_X1   g15420(.A1(new_n16421_), .A2(new_n16422_), .B(new_n16420_), .ZN(new_n16423_));
  NOR2_X1    g15421(.A1(new_n16419_), .A2(new_n16423_), .ZN(new_n16424_));
  NOR3_X1    g15422(.A1(new_n15914_), .A2(new_n15918_), .A3(new_n15408_), .ZN(new_n16425_));
  OAI21_X1   g15423(.A1(new_n16424_), .A2(new_n16425_), .B(new_n15919_), .ZN(new_n16426_));
  NAND2_X1   g15424(.A1(new_n16406_), .A2(new_n16411_), .ZN(new_n16427_));
  AOI22_X1   g15425(.A1(new_n16171_), .A2(new_n16421_), .B1(new_n16427_), .B2(new_n16412_), .ZN(new_n16428_));
  NOR3_X1    g15426(.A1(new_n16140_), .A2(new_n16168_), .A3(new_n16165_), .ZN(new_n16429_));
  OAI21_X1   g15427(.A1(new_n16161_), .A2(new_n16429_), .B(new_n16169_), .ZN(new_n16430_));
  AOI22_X1   g15428(.A1(new_n16155_), .A2(new_n16158_), .B1(new_n16022_), .B2(new_n16019_), .ZN(new_n16431_));
  AOI21_X1   g15429(.A1(new_n15949_), .A2(new_n15356_), .B(new_n15943_), .ZN(new_n16432_));
  XOR2_X1    g15430(.A1(new_n15922_), .A2(new_n15928_), .Z(new_n16433_));
  OAI21_X1   g15431(.A1(new_n16433_), .A2(new_n15920_), .B(new_n15957_), .ZN(new_n16434_));
  NOR2_X1    g15432(.A1(new_n16432_), .A2(new_n16434_), .ZN(new_n16435_));
  OAI21_X1   g15433(.A1(new_n15936_), .A2(new_n15941_), .B(new_n15952_), .ZN(new_n16436_));
  AOI21_X1   g15434(.A1(new_n15930_), .A2(new_n15388_), .B(new_n15924_), .ZN(new_n16437_));
  NOR2_X1    g15435(.A1(new_n16436_), .A2(new_n16437_), .ZN(new_n16438_));
  AOI21_X1   g15436(.A1(new_n15948_), .A2(new_n15954_), .B(new_n15931_), .ZN(new_n16439_));
  OAI22_X1   g15437(.A1(new_n16439_), .A2(new_n16149_), .B1(new_n16435_), .B2(new_n16438_), .ZN(new_n16440_));
  NAND2_X1   g15438(.A1(new_n16436_), .A2(new_n16437_), .ZN(new_n16441_));
  NAND2_X1   g15439(.A1(new_n16432_), .A2(new_n16434_), .ZN(new_n16442_));
  OAI21_X1   g15440(.A1(new_n15959_), .A2(new_n15947_), .B(new_n15958_), .ZN(new_n16443_));
  NAND4_X1   g15441(.A1(new_n16443_), .A2(new_n16442_), .A3(new_n15946_), .A4(new_n16441_), .ZN(new_n16444_));
  NAND2_X1   g15442(.A1(new_n16440_), .A2(new_n16444_), .ZN(new_n16445_));
  OAI21_X1   g15443(.A1(new_n15983_), .A2(new_n15976_), .B(new_n15986_), .ZN(new_n16446_));
  AOI21_X1   g15444(.A1(new_n15974_), .A2(new_n15323_), .B(new_n15968_), .ZN(new_n16447_));
  NAND2_X1   g15445(.A1(new_n16446_), .A2(new_n16447_), .ZN(new_n16448_));
  NAND2_X1   g15446(.A1(new_n15977_), .A2(new_n15303_), .ZN(new_n16449_));
  AOI22_X1   g15447(.A1(new_n16009_), .A2(new_n15291_), .B1(new_n16449_), .B2(new_n15985_), .ZN(new_n16450_));
  OAI21_X1   g15448(.A1(new_n16000_), .A2(new_n15964_), .B(new_n15997_), .ZN(new_n16451_));
  NAND2_X1   g15449(.A1(new_n16450_), .A2(new_n16451_), .ZN(new_n16452_));
  OAI21_X1   g15450(.A1(new_n16002_), .A2(new_n15993_), .B(new_n16001_), .ZN(new_n16453_));
  AOI22_X1   g15451(.A1(new_n16453_), .A2(new_n15988_), .B1(new_n16448_), .B2(new_n16452_), .ZN(new_n16454_));
  NOR2_X1    g15452(.A1(new_n16450_), .A2(new_n16451_), .ZN(new_n16455_));
  NOR2_X1    g15453(.A1(new_n16446_), .A2(new_n16447_), .ZN(new_n16456_));
  NOR2_X1    g15454(.A1(new_n16013_), .A2(new_n15975_), .ZN(new_n16457_));
  NOR4_X1    g15455(.A1(new_n16457_), .A2(new_n16455_), .A3(new_n16456_), .A4(new_n16012_), .ZN(new_n16458_));
  NOR2_X1    g15456(.A1(new_n16454_), .A2(new_n16458_), .ZN(new_n16459_));
  NAND2_X1   g15457(.A1(new_n16445_), .A2(new_n16459_), .ZN(new_n16460_));
  AOI22_X1   g15458(.A1(new_n15946_), .A2(new_n16443_), .B1(new_n16442_), .B2(new_n16441_), .ZN(new_n16461_));
  NOR4_X1    g15459(.A1(new_n16439_), .A2(new_n16435_), .A3(new_n16438_), .A4(new_n16149_), .ZN(new_n16462_));
  NOR2_X1    g15460(.A1(new_n16461_), .A2(new_n16462_), .ZN(new_n16463_));
  OAI22_X1   g15461(.A1(new_n16457_), .A2(new_n16012_), .B1(new_n16455_), .B2(new_n16456_), .ZN(new_n16464_));
  NAND4_X1   g15462(.A1(new_n16453_), .A2(new_n15988_), .A3(new_n16448_), .A4(new_n16452_), .ZN(new_n16465_));
  NAND2_X1   g15463(.A1(new_n16465_), .A2(new_n16464_), .ZN(new_n16466_));
  NAND2_X1   g15464(.A1(new_n16463_), .A2(new_n16466_), .ZN(new_n16467_));
  AOI21_X1   g15465(.A1(new_n16460_), .A2(new_n16467_), .B(new_n16431_), .ZN(new_n16468_));
  OAI21_X1   g15466(.A1(new_n15963_), .A2(new_n16023_), .B(new_n16159_), .ZN(new_n16469_));
  NOR2_X1    g15467(.A1(new_n16463_), .A2(new_n16466_), .ZN(new_n16470_));
  NOR2_X1    g15468(.A1(new_n16445_), .A2(new_n16459_), .ZN(new_n16471_));
  NOR3_X1    g15469(.A1(new_n16471_), .A2(new_n16470_), .A3(new_n16469_), .ZN(new_n16472_));
  NOR2_X1    g15470(.A1(new_n16468_), .A2(new_n16472_), .ZN(new_n16473_));
  OAI21_X1   g15471(.A1(new_n16135_), .A2(new_n16126_), .B(new_n16163_), .ZN(new_n16474_));
  OAI21_X1   g15472(.A1(new_n16057_), .A2(new_n16044_), .B(new_n16050_), .ZN(new_n16475_));
  AOI21_X1   g15473(.A1(new_n16063_), .A2(new_n15260_), .B(new_n16029_), .ZN(new_n16476_));
  NAND2_X1   g15474(.A1(new_n16475_), .A2(new_n16476_), .ZN(new_n16477_));
  AOI21_X1   g15475(.A1(new_n16043_), .A2(new_n15227_), .B(new_n16058_), .ZN(new_n16478_));
  XOR2_X1    g15476(.A1(new_n16027_), .A2(new_n16033_), .Z(new_n16479_));
  OAI21_X1   g15477(.A1(new_n16479_), .A2(new_n16045_), .B(new_n16030_), .ZN(new_n16480_));
  NAND2_X1   g15478(.A1(new_n16480_), .A2(new_n16478_), .ZN(new_n16481_));
  OAI21_X1   g15479(.A1(new_n16060_), .A2(new_n16056_), .B(new_n16035_), .ZN(new_n16482_));
  AOI22_X1   g15480(.A1(new_n16482_), .A2(new_n16129_), .B1(new_n16481_), .B2(new_n16477_), .ZN(new_n16483_));
  NOR2_X1    g15481(.A1(new_n16480_), .A2(new_n16478_), .ZN(new_n16484_));
  NOR2_X1    g15482(.A1(new_n16475_), .A2(new_n16476_), .ZN(new_n16485_));
  AOI21_X1   g15483(.A1(new_n16067_), .A2(new_n16065_), .B(new_n16064_), .ZN(new_n16486_));
  NOR4_X1    g15484(.A1(new_n16486_), .A2(new_n16484_), .A3(new_n16485_), .A4(new_n16053_), .ZN(new_n16487_));
  NOR2_X1    g15485(.A1(new_n16487_), .A2(new_n16483_), .ZN(new_n16488_));
  AOI21_X1   g15486(.A1(new_n16091_), .A2(new_n15162_), .B(new_n16105_), .ZN(new_n16489_));
  INV_X1     g15487(.I(new_n16076_), .ZN(new_n16490_));
  NOR2_X1    g15488(.A1(new_n16081_), .A2(new_n16079_), .ZN(new_n16491_));
  OAI21_X1   g15489(.A1(new_n16491_), .A2(new_n16072_), .B(new_n16490_), .ZN(new_n16492_));
  NOR2_X1    g15490(.A1(new_n16492_), .A2(new_n16489_), .ZN(new_n16493_));
  OAI21_X1   g15491(.A1(new_n16104_), .A2(new_n16092_), .B(new_n16097_), .ZN(new_n16494_));
  NAND2_X1   g15492(.A1(new_n16080_), .A2(new_n15206_), .ZN(new_n16495_));
  NAND2_X1   g15493(.A1(new_n16074_), .A2(new_n16078_), .ZN(new_n16496_));
  NAND2_X1   g15494(.A1(new_n16495_), .A2(new_n16496_), .ZN(new_n16497_));
  AOI21_X1   g15495(.A1(new_n16497_), .A2(new_n15194_), .B(new_n16076_), .ZN(new_n16498_));
  NOR2_X1    g15496(.A1(new_n16494_), .A2(new_n16498_), .ZN(new_n16499_));
  AOI21_X1   g15497(.A1(new_n16120_), .A2(new_n16110_), .B(new_n16082_), .ZN(new_n16500_));
  OAI22_X1   g15498(.A1(new_n16493_), .A2(new_n16499_), .B1(new_n16500_), .B2(new_n16100_), .ZN(new_n16501_));
  NAND2_X1   g15499(.A1(new_n16494_), .A2(new_n16498_), .ZN(new_n16502_));
  NAND2_X1   g15500(.A1(new_n16492_), .A2(new_n16489_), .ZN(new_n16503_));
  OAI21_X1   g15501(.A1(new_n16107_), .A2(new_n16101_), .B(new_n16083_), .ZN(new_n16504_));
  NAND4_X1   g15502(.A1(new_n16504_), .A2(new_n16119_), .A3(new_n16502_), .A4(new_n16503_), .ZN(new_n16505_));
  NAND2_X1   g15503(.A1(new_n16505_), .A2(new_n16501_), .ZN(new_n16506_));
  NOR2_X1    g15504(.A1(new_n16488_), .A2(new_n16506_), .ZN(new_n16507_));
  OAI22_X1   g15505(.A1(new_n16486_), .A2(new_n16053_), .B1(new_n16484_), .B2(new_n16485_), .ZN(new_n16508_));
  NAND4_X1   g15506(.A1(new_n16482_), .A2(new_n16129_), .A3(new_n16481_), .A4(new_n16477_), .ZN(new_n16509_));
  NAND2_X1   g15507(.A1(new_n16508_), .A2(new_n16509_), .ZN(new_n16510_));
  AOI22_X1   g15508(.A1(new_n16504_), .A2(new_n16119_), .B1(new_n16502_), .B2(new_n16503_), .ZN(new_n16511_));
  NOR4_X1    g15509(.A1(new_n16493_), .A2(new_n16499_), .A3(new_n16500_), .A4(new_n16100_), .ZN(new_n16512_));
  NOR2_X1    g15510(.A1(new_n16511_), .A2(new_n16512_), .ZN(new_n16513_));
  NOR2_X1    g15511(.A1(new_n16510_), .A2(new_n16513_), .ZN(new_n16514_));
  OAI21_X1   g15512(.A1(new_n16507_), .A2(new_n16514_), .B(new_n16474_), .ZN(new_n16515_));
  AOI21_X1   g15513(.A1(new_n16070_), .A2(new_n16164_), .B(new_n16114_), .ZN(new_n16516_));
  NAND2_X1   g15514(.A1(new_n16510_), .A2(new_n16513_), .ZN(new_n16517_));
  NAND2_X1   g15515(.A1(new_n16488_), .A2(new_n16506_), .ZN(new_n16518_));
  NAND3_X1   g15516(.A1(new_n16517_), .A2(new_n16518_), .A3(new_n16516_), .ZN(new_n16519_));
  NAND2_X1   g15517(.A1(new_n16515_), .A2(new_n16519_), .ZN(new_n16520_));
  NOR2_X1    g15518(.A1(new_n16473_), .A2(new_n16520_), .ZN(new_n16521_));
  OAI21_X1   g15519(.A1(new_n16471_), .A2(new_n16470_), .B(new_n16469_), .ZN(new_n16522_));
  NAND3_X1   g15520(.A1(new_n16460_), .A2(new_n16467_), .A3(new_n16431_), .ZN(new_n16523_));
  NAND2_X1   g15521(.A1(new_n16522_), .A2(new_n16523_), .ZN(new_n16524_));
  AOI21_X1   g15522(.A1(new_n16517_), .A2(new_n16518_), .B(new_n16516_), .ZN(new_n16525_));
  NOR3_X1    g15523(.A1(new_n16507_), .A2(new_n16514_), .A3(new_n16474_), .ZN(new_n16526_));
  NOR2_X1    g15524(.A1(new_n16526_), .A2(new_n16525_), .ZN(new_n16527_));
  NOR2_X1    g15525(.A1(new_n16527_), .A2(new_n16524_), .ZN(new_n16528_));
  OAI21_X1   g15526(.A1(new_n16528_), .A2(new_n16521_), .B(new_n16430_), .ZN(new_n16529_));
  AOI22_X1   g15527(.A1(new_n16025_), .A2(new_n16162_), .B1(new_n16140_), .B2(new_n16143_), .ZN(new_n16530_));
  NAND2_X1   g15528(.A1(new_n16527_), .A2(new_n16524_), .ZN(new_n16531_));
  NAND2_X1   g15529(.A1(new_n16473_), .A2(new_n16520_), .ZN(new_n16532_));
  NAND3_X1   g15530(.A1(new_n16531_), .A2(new_n16532_), .A3(new_n16530_), .ZN(new_n16533_));
  NAND2_X1   g15531(.A1(new_n16529_), .A2(new_n16533_), .ZN(new_n16534_));
  AOI22_X1   g15532(.A1(new_n16284_), .A2(new_n16401_), .B1(new_n16403_), .B2(new_n16402_), .ZN(new_n16535_));
  NOR2_X1    g15533(.A1(new_n16247_), .A2(new_n16257_), .ZN(new_n16536_));
  OAI22_X1   g15534(.A1(new_n16281_), .A2(new_n16218_), .B1(new_n16536_), .B2(new_n16258_), .ZN(new_n16537_));
  OAI21_X1   g15535(.A1(new_n16185_), .A2(new_n16190_), .B(new_n16207_), .ZN(new_n16538_));
  NAND2_X1   g15536(.A1(new_n16175_), .A2(new_n15139_), .ZN(new_n16539_));
  AOI22_X1   g15537(.A1(new_n16179_), .A2(new_n15127_), .B1(new_n16539_), .B2(new_n16180_), .ZN(new_n16540_));
  NAND2_X1   g15538(.A1(new_n16538_), .A2(new_n16540_), .ZN(new_n16541_));
  AOI21_X1   g15539(.A1(new_n16205_), .A2(new_n15095_), .B(new_n16194_), .ZN(new_n16542_));
  XOR2_X1    g15540(.A1(new_n16175_), .A2(new_n16177_), .Z(new_n16543_));
  OAI21_X1   g15541(.A1(new_n16543_), .A2(new_n16198_), .B(new_n16181_), .ZN(new_n16544_));
  NAND2_X1   g15542(.A1(new_n16544_), .A2(new_n16542_), .ZN(new_n16545_));
  OAI21_X1   g15543(.A1(new_n16213_), .A2(new_n16215_), .B(new_n16212_), .ZN(new_n16546_));
  AOI22_X1   g15544(.A1(new_n16197_), .A2(new_n16546_), .B1(new_n16541_), .B2(new_n16545_), .ZN(new_n16547_));
  NOR2_X1    g15545(.A1(new_n16544_), .A2(new_n16542_), .ZN(new_n16548_));
  NOR2_X1    g15546(.A1(new_n16538_), .A2(new_n16540_), .ZN(new_n16549_));
  AOI21_X1   g15547(.A1(new_n16200_), .A2(new_n16209_), .B(new_n16183_), .ZN(new_n16550_));
  NOR4_X1    g15548(.A1(new_n16549_), .A2(new_n16550_), .A3(new_n16548_), .A4(new_n16274_), .ZN(new_n16551_));
  NOR2_X1    g15549(.A1(new_n16547_), .A2(new_n16551_), .ZN(new_n16552_));
  NAND2_X1   g15550(.A1(new_n16232_), .A2(new_n16230_), .ZN(new_n16553_));
  AOI22_X1   g15551(.A1(new_n16235_), .A2(new_n15070_), .B1(new_n16239_), .B2(new_n16553_), .ZN(new_n16554_));
  NOR2_X1    g15552(.A1(new_n16227_), .A2(new_n16225_), .ZN(new_n16555_));
  OAI21_X1   g15553(.A1(new_n16555_), .A2(new_n16219_), .B(new_n16248_), .ZN(new_n16556_));
  NOR2_X1    g15554(.A1(new_n16554_), .A2(new_n16556_), .ZN(new_n16557_));
  NOR2_X1    g15555(.A1(new_n16232_), .A2(new_n16233_), .ZN(new_n16558_));
  NOR2_X1    g15556(.A1(new_n16229_), .A2(new_n16230_), .ZN(new_n16559_));
  NOR2_X1    g15557(.A1(new_n16559_), .A2(new_n16558_), .ZN(new_n16560_));
  OAI21_X1   g15558(.A1(new_n16560_), .A2(new_n16236_), .B(new_n16240_), .ZN(new_n16561_));
  NAND2_X1   g15559(.A1(new_n16249_), .A2(new_n16250_), .ZN(new_n16562_));
  AOI21_X1   g15560(.A1(new_n16562_), .A2(new_n15047_), .B(new_n16223_), .ZN(new_n16563_));
  NOR2_X1    g15561(.A1(new_n16561_), .A2(new_n16563_), .ZN(new_n16564_));
  AOI21_X1   g15562(.A1(new_n16255_), .A2(new_n16252_), .B(new_n16228_), .ZN(new_n16565_));
  OAI22_X1   g15563(.A1(new_n16557_), .A2(new_n16564_), .B1(new_n16565_), .B2(new_n16262_), .ZN(new_n16566_));
  NAND2_X1   g15564(.A1(new_n16561_), .A2(new_n16563_), .ZN(new_n16567_));
  NAND2_X1   g15565(.A1(new_n16554_), .A2(new_n16556_), .ZN(new_n16568_));
  OAI21_X1   g15566(.A1(new_n16244_), .A2(new_n16243_), .B(new_n16251_), .ZN(new_n16569_));
  NAND4_X1   g15567(.A1(new_n16569_), .A2(new_n16242_), .A3(new_n16568_), .A4(new_n16567_), .ZN(new_n16570_));
  NAND2_X1   g15568(.A1(new_n16570_), .A2(new_n16566_), .ZN(new_n16571_));
  NOR2_X1    g15569(.A1(new_n16552_), .A2(new_n16571_), .ZN(new_n16572_));
  OAI22_X1   g15570(.A1(new_n16548_), .A2(new_n16549_), .B1(new_n16550_), .B2(new_n16274_), .ZN(new_n16573_));
  NAND4_X1   g15571(.A1(new_n16197_), .A2(new_n16541_), .A3(new_n16546_), .A4(new_n16545_), .ZN(new_n16574_));
  NAND2_X1   g15572(.A1(new_n16573_), .A2(new_n16574_), .ZN(new_n16575_));
  AOI22_X1   g15573(.A1(new_n16569_), .A2(new_n16242_), .B1(new_n16568_), .B2(new_n16567_), .ZN(new_n16576_));
  NOR4_X1    g15574(.A1(new_n16565_), .A2(new_n16557_), .A3(new_n16564_), .A4(new_n16262_), .ZN(new_n16577_));
  NOR2_X1    g15575(.A1(new_n16576_), .A2(new_n16577_), .ZN(new_n16578_));
  NOR2_X1    g15576(.A1(new_n16575_), .A2(new_n16578_), .ZN(new_n16579_));
  OAI21_X1   g15577(.A1(new_n16579_), .A2(new_n16572_), .B(new_n16537_), .ZN(new_n16580_));
  NAND3_X1   g15578(.A1(new_n16263_), .A2(new_n16266_), .A3(new_n16258_), .ZN(new_n16581_));
  AOI21_X1   g15579(.A1(new_n16280_), .A2(new_n16581_), .B(new_n16282_), .ZN(new_n16582_));
  NAND2_X1   g15580(.A1(new_n16575_), .A2(new_n16578_), .ZN(new_n16583_));
  NAND2_X1   g15581(.A1(new_n16552_), .A2(new_n16571_), .ZN(new_n16584_));
  NAND3_X1   g15582(.A1(new_n16583_), .A2(new_n16584_), .A3(new_n16582_), .ZN(new_n16585_));
  NAND2_X1   g15583(.A1(new_n16580_), .A2(new_n16585_), .ZN(new_n16586_));
  NAND3_X1   g15584(.A1(new_n16366_), .A2(new_n16375_), .A3(new_n16327_), .ZN(new_n16587_));
  AOI21_X1   g15585(.A1(new_n16326_), .A2(new_n16587_), .B(new_n16376_), .ZN(new_n16588_));
  AOI21_X1   g15586(.A1(new_n16300_), .A2(new_n15026_), .B(new_n16307_), .ZN(new_n16589_));
  AOI21_X1   g15587(.A1(new_n16322_), .A2(new_n15017_), .B(new_n16589_), .ZN(new_n16590_));
  INV_X1     g15588(.I(new_n14988_), .ZN(new_n16591_));
  NOR2_X1    g15589(.A1(new_n16295_), .A2(new_n16287_), .ZN(new_n16592_));
  NOR2_X1    g15590(.A1(new_n16285_), .A2(new_n14997_), .ZN(new_n16593_));
  NOR2_X1    g15591(.A1(new_n16593_), .A2(new_n16592_), .ZN(new_n16594_));
  OAI21_X1   g15592(.A1(new_n16594_), .A2(new_n16591_), .B(new_n16293_), .ZN(new_n16595_));
  NOR2_X1    g15593(.A1(new_n16595_), .A2(new_n16590_), .ZN(new_n16596_));
  INV_X1     g15594(.I(new_n15017_), .ZN(new_n16597_));
  OAI21_X1   g15595(.A1(new_n16305_), .A2(new_n16597_), .B(new_n16309_), .ZN(new_n16598_));
  INV_X1     g15596(.I(new_n16293_), .ZN(new_n16599_));
  NAND2_X1   g15597(.A1(new_n16294_), .A2(new_n16296_), .ZN(new_n16600_));
  AOI21_X1   g15598(.A1(new_n16600_), .A2(new_n14988_), .B(new_n16599_), .ZN(new_n16601_));
  NOR2_X1    g15599(.A1(new_n16601_), .A2(new_n16598_), .ZN(new_n16602_));
  OAI21_X1   g15600(.A1(new_n16317_), .A2(new_n16314_), .B(new_n16297_), .ZN(new_n16603_));
  INV_X1     g15601(.I(new_n16603_), .ZN(new_n16604_));
  OAI22_X1   g15602(.A1(new_n16604_), .A2(new_n16312_), .B1(new_n16596_), .B2(new_n16602_), .ZN(new_n16605_));
  NAND2_X1   g15603(.A1(new_n16601_), .A2(new_n16598_), .ZN(new_n16606_));
  NAND2_X1   g15604(.A1(new_n16595_), .A2(new_n16590_), .ZN(new_n16607_));
  NAND4_X1   g15605(.A1(new_n16390_), .A2(new_n16606_), .A3(new_n16607_), .A4(new_n16603_), .ZN(new_n16608_));
  NAND2_X1   g15606(.A1(new_n16605_), .A2(new_n16608_), .ZN(new_n16609_));
  NOR2_X1    g15607(.A1(new_n16348_), .A2(new_n16350_), .ZN(new_n16610_));
  NOR2_X1    g15608(.A1(new_n16341_), .A2(new_n14968_), .ZN(new_n16611_));
  NOR2_X1    g15609(.A1(new_n16611_), .A2(new_n16610_), .ZN(new_n16612_));
  OAI21_X1   g15610(.A1(new_n16612_), .A2(new_n16354_), .B(new_n16359_), .ZN(new_n16613_));
  NAND2_X1   g15611(.A1(new_n16338_), .A2(new_n16336_), .ZN(new_n16614_));
  AOI21_X1   g15612(.A1(new_n16614_), .A2(new_n14931_), .B(new_n16367_), .ZN(new_n16615_));
  NAND2_X1   g15613(.A1(new_n16613_), .A2(new_n16615_), .ZN(new_n16616_));
  NAND2_X1   g15614(.A1(new_n16348_), .A2(new_n14968_), .ZN(new_n16617_));
  AOI22_X1   g15615(.A1(new_n16352_), .A2(new_n14958_), .B1(new_n16358_), .B2(new_n16617_), .ZN(new_n16618_));
  NOR2_X1    g15616(.A1(new_n16369_), .A2(new_n16368_), .ZN(new_n16619_));
  OAI21_X1   g15617(.A1(new_n16619_), .A2(new_n16353_), .B(new_n16333_), .ZN(new_n16620_));
  NAND2_X1   g15618(.A1(new_n16618_), .A2(new_n16620_), .ZN(new_n16621_));
  OAI21_X1   g15619(.A1(new_n16364_), .A2(new_n16363_), .B(new_n16339_), .ZN(new_n16622_));
  AOI22_X1   g15620(.A1(new_n16616_), .A2(new_n16621_), .B1(new_n16381_), .B2(new_n16622_), .ZN(new_n16623_));
  NOR2_X1    g15621(.A1(new_n16618_), .A2(new_n16620_), .ZN(new_n16624_));
  NOR2_X1    g15622(.A1(new_n16613_), .A2(new_n16615_), .ZN(new_n16625_));
  AOI21_X1   g15623(.A1(new_n16371_), .A2(new_n16373_), .B(new_n16370_), .ZN(new_n16626_));
  NOR4_X1    g15624(.A1(new_n16624_), .A2(new_n16625_), .A3(new_n16626_), .A4(new_n16362_), .ZN(new_n16627_));
  NOR2_X1    g15625(.A1(new_n16623_), .A2(new_n16627_), .ZN(new_n16628_));
  NAND2_X1   g15626(.A1(new_n16609_), .A2(new_n16628_), .ZN(new_n16629_));
  AOI22_X1   g15627(.A1(new_n16606_), .A2(new_n16607_), .B1(new_n16390_), .B2(new_n16603_), .ZN(new_n16630_));
  NOR4_X1    g15628(.A1(new_n16604_), .A2(new_n16596_), .A3(new_n16602_), .A4(new_n16312_), .ZN(new_n16631_));
  NOR2_X1    g15629(.A1(new_n16631_), .A2(new_n16630_), .ZN(new_n16632_));
  OAI22_X1   g15630(.A1(new_n16624_), .A2(new_n16625_), .B1(new_n16626_), .B2(new_n16362_), .ZN(new_n16633_));
  NAND4_X1   g15631(.A1(new_n16621_), .A2(new_n16381_), .A3(new_n16616_), .A4(new_n16622_), .ZN(new_n16634_));
  NAND2_X1   g15632(.A1(new_n16633_), .A2(new_n16634_), .ZN(new_n16635_));
  NAND2_X1   g15633(.A1(new_n16632_), .A2(new_n16635_), .ZN(new_n16636_));
  AOI21_X1   g15634(.A1(new_n16629_), .A2(new_n16636_), .B(new_n16588_), .ZN(new_n16637_));
  NOR2_X1    g15635(.A1(new_n16383_), .A2(new_n16386_), .ZN(new_n16638_));
  OAI22_X1   g15636(.A1(new_n16387_), .A2(new_n16396_), .B1(new_n16638_), .B2(new_n16327_), .ZN(new_n16639_));
  NOR2_X1    g15637(.A1(new_n16632_), .A2(new_n16635_), .ZN(new_n16640_));
  NOR2_X1    g15638(.A1(new_n16609_), .A2(new_n16628_), .ZN(new_n16641_));
  NOR3_X1    g15639(.A1(new_n16639_), .A2(new_n16641_), .A3(new_n16640_), .ZN(new_n16642_));
  NOR2_X1    g15640(.A1(new_n16642_), .A2(new_n16637_), .ZN(new_n16643_));
  NAND2_X1   g15641(.A1(new_n16586_), .A2(new_n16643_), .ZN(new_n16644_));
  AOI21_X1   g15642(.A1(new_n16583_), .A2(new_n16584_), .B(new_n16582_), .ZN(new_n16645_));
  NOR3_X1    g15643(.A1(new_n16537_), .A2(new_n16579_), .A3(new_n16572_), .ZN(new_n16646_));
  NOR2_X1    g15644(.A1(new_n16646_), .A2(new_n16645_), .ZN(new_n16647_));
  OAI21_X1   g15645(.A1(new_n16640_), .A2(new_n16641_), .B(new_n16639_), .ZN(new_n16648_));
  NAND3_X1   g15646(.A1(new_n16629_), .A2(new_n16636_), .A3(new_n16588_), .ZN(new_n16649_));
  NAND2_X1   g15647(.A1(new_n16648_), .A2(new_n16649_), .ZN(new_n16650_));
  NAND2_X1   g15648(.A1(new_n16647_), .A2(new_n16650_), .ZN(new_n16651_));
  AOI21_X1   g15649(.A1(new_n16644_), .A2(new_n16651_), .B(new_n16535_), .ZN(new_n16652_));
  INV_X1     g15650(.I(new_n16535_), .ZN(new_n16653_));
  NOR2_X1    g15651(.A1(new_n16647_), .A2(new_n16650_), .ZN(new_n16654_));
  NOR2_X1    g15652(.A1(new_n16586_), .A2(new_n16643_), .ZN(new_n16655_));
  NOR3_X1    g15653(.A1(new_n16655_), .A2(new_n16654_), .A3(new_n16653_), .ZN(new_n16656_));
  NOR2_X1    g15654(.A1(new_n16652_), .A2(new_n16656_), .ZN(new_n16657_));
  NAND2_X1   g15655(.A1(new_n16534_), .A2(new_n16657_), .ZN(new_n16658_));
  AOI21_X1   g15656(.A1(new_n16531_), .A2(new_n16532_), .B(new_n16530_), .ZN(new_n16659_));
  NOR3_X1    g15657(.A1(new_n16528_), .A2(new_n16521_), .A3(new_n16430_), .ZN(new_n16660_));
  NOR2_X1    g15658(.A1(new_n16659_), .A2(new_n16660_), .ZN(new_n16661_));
  OAI21_X1   g15659(.A1(new_n16655_), .A2(new_n16654_), .B(new_n16653_), .ZN(new_n16662_));
  NAND3_X1   g15660(.A1(new_n16644_), .A2(new_n16651_), .A3(new_n16535_), .ZN(new_n16663_));
  NAND2_X1   g15661(.A1(new_n16662_), .A2(new_n16663_), .ZN(new_n16664_));
  NAND2_X1   g15662(.A1(new_n16661_), .A2(new_n16664_), .ZN(new_n16665_));
  AOI21_X1   g15663(.A1(new_n16658_), .A2(new_n16665_), .B(new_n16428_), .ZN(new_n16666_));
  NOR3_X1    g15664(.A1(new_n16414_), .A2(new_n16416_), .A3(new_n16412_), .ZN(new_n16667_));
  OAI21_X1   g15665(.A1(new_n16420_), .A2(new_n16667_), .B(new_n16422_), .ZN(new_n16668_));
  NOR2_X1    g15666(.A1(new_n16661_), .A2(new_n16664_), .ZN(new_n16669_));
  NOR2_X1    g15667(.A1(new_n16534_), .A2(new_n16657_), .ZN(new_n16670_));
  NOR3_X1    g15668(.A1(new_n16670_), .A2(new_n16669_), .A3(new_n16668_), .ZN(new_n16671_));
  NOR2_X1    g15669(.A1(new_n16666_), .A2(new_n16671_), .ZN(new_n16672_));
  NOR3_X1    g15670(.A1(new_n15902_), .A2(new_n15905_), .A3(new_n15906_), .ZN(new_n16673_));
  OAI21_X1   g15671(.A1(new_n15915_), .A2(new_n16673_), .B(new_n15917_), .ZN(new_n16674_));
  INV_X1     g15672(.I(new_n15629_), .ZN(new_n16675_));
  AOI21_X1   g15673(.A1(new_n15625_), .A2(new_n15616_), .B(new_n15628_), .ZN(new_n16676_));
  OAI21_X1   g15674(.A1(new_n16675_), .A2(new_n16676_), .B(new_n15644_), .ZN(new_n16677_));
  NOR3_X1    g15675(.A1(new_n15633_), .A2(new_n15636_), .A3(new_n15628_), .ZN(new_n16678_));
  AOI21_X1   g15676(.A1(new_n15625_), .A2(new_n15616_), .B(new_n15637_), .ZN(new_n16679_));
  OAI21_X1   g15677(.A1(new_n16678_), .A2(new_n16679_), .B(new_n15574_), .ZN(new_n16680_));
  NAND2_X1   g15678(.A1(new_n16677_), .A2(new_n16680_), .ZN(new_n16681_));
  NAND3_X1   g15679(.A1(new_n16677_), .A2(new_n15527_), .A3(new_n16680_), .ZN(new_n16682_));
  AOI22_X1   g15680(.A1(new_n16682_), .A2(new_n15656_), .B1(new_n16681_), .B2(new_n15528_), .ZN(new_n16683_));
  OAI21_X1   g15681(.A1(new_n15522_), .A2(new_n15653_), .B(new_n15524_), .ZN(new_n16684_));
  OAI21_X1   g15682(.A1(new_n15514_), .A2(new_n15430_), .B(new_n15436_), .ZN(new_n16685_));
  NAND2_X1   g15683(.A1(new_n15412_), .A2(new_n14672_), .ZN(new_n16686_));
  AOI22_X1   g15684(.A1(new_n15416_), .A2(new_n14660_), .B1(new_n16686_), .B2(new_n15417_), .ZN(new_n16687_));
  NAND2_X1   g15685(.A1(new_n16687_), .A2(new_n16685_), .ZN(new_n16688_));
  AOI21_X1   g15686(.A1(new_n15429_), .A2(new_n14628_), .B(new_n15516_), .ZN(new_n16689_));
  NAND2_X1   g15687(.A1(new_n15416_), .A2(new_n14660_), .ZN(new_n16690_));
  NAND2_X1   g15688(.A1(new_n16690_), .A2(new_n15418_), .ZN(new_n16691_));
  NAND2_X1   g15689(.A1(new_n16691_), .A2(new_n16689_), .ZN(new_n16692_));
  NAND2_X1   g15690(.A1(new_n15442_), .A2(new_n15421_), .ZN(new_n16693_));
  AOI22_X1   g15691(.A1(new_n16693_), .A2(new_n15519_), .B1(new_n16692_), .B2(new_n16688_), .ZN(new_n16694_));
  NOR2_X1    g15692(.A1(new_n16691_), .A2(new_n16689_), .ZN(new_n16695_));
  NOR2_X1    g15693(.A1(new_n16687_), .A2(new_n16685_), .ZN(new_n16696_));
  AOI21_X1   g15694(.A1(new_n15440_), .A2(new_n15441_), .B(new_n15420_), .ZN(new_n16697_));
  NOR4_X1    g15695(.A1(new_n16695_), .A2(new_n16697_), .A3(new_n15439_), .A4(new_n16696_), .ZN(new_n16698_));
  NOR2_X1    g15696(.A1(new_n16694_), .A2(new_n16698_), .ZN(new_n16699_));
  NAND2_X1   g15697(.A1(new_n15466_), .A2(new_n14575_), .ZN(new_n16700_));
  AOI22_X1   g15698(.A1(new_n15483_), .A2(new_n14563_), .B1(new_n16700_), .B2(new_n15475_), .ZN(new_n16701_));
  NOR2_X1    g15699(.A1(new_n15462_), .A2(new_n15460_), .ZN(new_n16702_));
  OAI21_X1   g15700(.A1(new_n16702_), .A2(new_n15453_), .B(new_n15487_), .ZN(new_n16703_));
  NOR2_X1    g15701(.A1(new_n16701_), .A2(new_n16703_), .ZN(new_n16704_));
  OAI21_X1   g15702(.A1(new_n15472_), .A2(new_n15464_), .B(new_n15476_), .ZN(new_n16705_));
  NAND2_X1   g15703(.A1(new_n15488_), .A2(new_n15489_), .ZN(new_n16706_));
  AOI21_X1   g15704(.A1(new_n16706_), .A2(new_n14595_), .B(new_n15457_), .ZN(new_n16707_));
  NOR2_X1    g15705(.A1(new_n16705_), .A2(new_n16707_), .ZN(new_n16708_));
  AOI21_X1   g15706(.A1(new_n15484_), .A2(new_n15480_), .B(new_n15463_), .ZN(new_n16709_));
  OAI22_X1   g15707(.A1(new_n16704_), .A2(new_n16708_), .B1(new_n16709_), .B2(new_n15500_), .ZN(new_n16710_));
  NAND2_X1   g15708(.A1(new_n16705_), .A2(new_n16707_), .ZN(new_n16711_));
  NAND2_X1   g15709(.A1(new_n16701_), .A2(new_n16703_), .ZN(new_n16712_));
  OAI21_X1   g15710(.A1(new_n15493_), .A2(new_n15491_), .B(new_n15490_), .ZN(new_n16713_));
  NAND4_X1   g15711(.A1(new_n16713_), .A2(new_n15478_), .A3(new_n16712_), .A4(new_n16711_), .ZN(new_n16714_));
  NAND2_X1   g15712(.A1(new_n16714_), .A2(new_n16710_), .ZN(new_n16715_));
  NOR2_X1    g15713(.A1(new_n16699_), .A2(new_n16715_), .ZN(new_n16716_));
  OAI22_X1   g15714(.A1(new_n16695_), .A2(new_n16696_), .B1(new_n16697_), .B2(new_n15439_), .ZN(new_n16717_));
  NAND4_X1   g15715(.A1(new_n16693_), .A2(new_n16692_), .A3(new_n15519_), .A4(new_n16688_), .ZN(new_n16718_));
  NAND2_X1   g15716(.A1(new_n16718_), .A2(new_n16717_), .ZN(new_n16719_));
  AOI22_X1   g15717(.A1(new_n16713_), .A2(new_n15478_), .B1(new_n16712_), .B2(new_n16711_), .ZN(new_n16720_));
  NOR4_X1    g15718(.A1(new_n16704_), .A2(new_n16708_), .A3(new_n16709_), .A4(new_n15500_), .ZN(new_n16721_));
  NOR2_X1    g15719(.A1(new_n16720_), .A2(new_n16721_), .ZN(new_n16722_));
  NOR2_X1    g15720(.A1(new_n16719_), .A2(new_n16722_), .ZN(new_n16723_));
  OAI21_X1   g15721(.A1(new_n16716_), .A2(new_n16723_), .B(new_n16684_), .ZN(new_n16724_));
  AOI21_X1   g15722(.A1(new_n15452_), .A2(new_n15523_), .B(new_n15654_), .ZN(new_n16725_));
  NAND2_X1   g15723(.A1(new_n16719_), .A2(new_n16722_), .ZN(new_n16726_));
  NAND2_X1   g15724(.A1(new_n16699_), .A2(new_n16715_), .ZN(new_n16727_));
  NAND3_X1   g15725(.A1(new_n16727_), .A2(new_n16726_), .A3(new_n16725_), .ZN(new_n16728_));
  NAND2_X1   g15726(.A1(new_n16724_), .A2(new_n16728_), .ZN(new_n16729_));
  AOI21_X1   g15727(.A1(new_n15574_), .A2(new_n15645_), .B(new_n16679_), .ZN(new_n16730_));
  AOI21_X1   g15728(.A1(new_n15568_), .A2(new_n14514_), .B(new_n15549_), .ZN(new_n16731_));
  OAI21_X1   g15729(.A1(new_n15562_), .A2(new_n15529_), .B(new_n15559_), .ZN(new_n16732_));
  NOR2_X1    g15730(.A1(new_n16732_), .A2(new_n16731_), .ZN(new_n16733_));
  NOR2_X1    g15731(.A1(new_n15550_), .A2(new_n15552_), .ZN(new_n16734_));
  NOR2_X1    g15732(.A1(new_n15551_), .A2(new_n15553_), .ZN(new_n16735_));
  OAI22_X1   g15733(.A1(new_n16735_), .A2(new_n15543_), .B1(new_n15547_), .B2(new_n16734_), .ZN(new_n16736_));
  AOI21_X1   g15734(.A1(new_n15541_), .A2(new_n14532_), .B(new_n15535_), .ZN(new_n16737_));
  NOR2_X1    g15735(.A1(new_n16736_), .A2(new_n16737_), .ZN(new_n16738_));
  AOI21_X1   g15736(.A1(new_n15545_), .A2(new_n15554_), .B(new_n15542_), .ZN(new_n16739_));
  OAI22_X1   g15737(.A1(new_n16739_), .A2(new_n15570_), .B1(new_n16733_), .B2(new_n16738_), .ZN(new_n16740_));
  NAND2_X1   g15738(.A1(new_n16736_), .A2(new_n16737_), .ZN(new_n16741_));
  NAND2_X1   g15739(.A1(new_n16732_), .A2(new_n16731_), .ZN(new_n16742_));
  NAND2_X1   g15740(.A1(new_n15571_), .A2(new_n15563_), .ZN(new_n16743_));
  NAND4_X1   g15741(.A1(new_n16743_), .A2(new_n15642_), .A3(new_n16741_), .A4(new_n16742_), .ZN(new_n16744_));
  NAND2_X1   g15742(.A1(new_n16740_), .A2(new_n16744_), .ZN(new_n16745_));
  XOR2_X1    g15743(.A1(new_n14440_), .A2(new_n15594_), .Z(new_n16746_));
  NOR2_X1    g15744(.A1(new_n16746_), .A2(new_n15595_), .ZN(new_n16747_));
  OAI22_X1   g15745(.A1(new_n15613_), .A2(new_n15604_), .B1(new_n15608_), .B2(new_n16747_), .ZN(new_n16748_));
  NAND2_X1   g15746(.A1(new_n15585_), .A2(new_n15587_), .ZN(new_n16749_));
  AOI21_X1   g15747(.A1(new_n16749_), .A2(new_n14476_), .B(new_n15617_), .ZN(new_n16750_));
  NAND2_X1   g15748(.A1(new_n16748_), .A2(new_n16750_), .ZN(new_n16751_));
  AOI21_X1   g15749(.A1(new_n15603_), .A2(new_n14458_), .B(new_n15609_), .ZN(new_n16752_));
  NOR2_X1    g15750(.A1(new_n15619_), .A2(new_n15618_), .ZN(new_n16753_));
  OAI21_X1   g15751(.A1(new_n16753_), .A2(new_n15605_), .B(new_n15584_), .ZN(new_n16754_));
  NAND2_X1   g15752(.A1(new_n16754_), .A2(new_n16752_), .ZN(new_n16755_));
  OAI21_X1   g15753(.A1(new_n15614_), .A2(new_n15612_), .B(new_n15588_), .ZN(new_n16756_));
  AOI22_X1   g15754(.A1(new_n16751_), .A2(new_n16755_), .B1(new_n16756_), .B2(new_n15631_), .ZN(new_n16757_));
  NOR2_X1    g15755(.A1(new_n16754_), .A2(new_n16752_), .ZN(new_n16758_));
  NOR2_X1    g15756(.A1(new_n16748_), .A2(new_n16750_), .ZN(new_n16759_));
  AOI21_X1   g15757(.A1(new_n15621_), .A2(new_n15623_), .B(new_n15620_), .ZN(new_n16760_));
  NOR4_X1    g15758(.A1(new_n16759_), .A2(new_n16760_), .A3(new_n16758_), .A4(new_n15611_), .ZN(new_n16761_));
  NOR2_X1    g15759(.A1(new_n16761_), .A2(new_n16757_), .ZN(new_n16762_));
  NAND2_X1   g15760(.A1(new_n16745_), .A2(new_n16762_), .ZN(new_n16763_));
  AOI22_X1   g15761(.A1(new_n16743_), .A2(new_n15642_), .B1(new_n16741_), .B2(new_n16742_), .ZN(new_n16764_));
  NOR4_X1    g15762(.A1(new_n16739_), .A2(new_n16733_), .A3(new_n16738_), .A4(new_n15570_), .ZN(new_n16765_));
  NOR2_X1    g15763(.A1(new_n16765_), .A2(new_n16764_), .ZN(new_n16766_));
  OAI22_X1   g15764(.A1(new_n16759_), .A2(new_n16758_), .B1(new_n16760_), .B2(new_n15611_), .ZN(new_n16767_));
  NAND4_X1   g15765(.A1(new_n16751_), .A2(new_n16755_), .A3(new_n16756_), .A4(new_n15631_), .ZN(new_n16768_));
  NAND2_X1   g15766(.A1(new_n16767_), .A2(new_n16768_), .ZN(new_n16769_));
  NAND2_X1   g15767(.A1(new_n16766_), .A2(new_n16769_), .ZN(new_n16770_));
  AOI21_X1   g15768(.A1(new_n16770_), .A2(new_n16763_), .B(new_n16730_), .ZN(new_n16771_));
  OAI21_X1   g15769(.A1(new_n15644_), .A2(new_n16678_), .B(new_n15646_), .ZN(new_n16772_));
  NOR2_X1    g15770(.A1(new_n16766_), .A2(new_n16769_), .ZN(new_n16773_));
  NOR2_X1    g15771(.A1(new_n16745_), .A2(new_n16762_), .ZN(new_n16774_));
  NOR3_X1    g15772(.A1(new_n16773_), .A2(new_n16774_), .A3(new_n16772_), .ZN(new_n16775_));
  NOR2_X1    g15773(.A1(new_n16775_), .A2(new_n16771_), .ZN(new_n16776_));
  NAND2_X1   g15774(.A1(new_n16729_), .A2(new_n16776_), .ZN(new_n16777_));
  AOI21_X1   g15775(.A1(new_n16727_), .A2(new_n16726_), .B(new_n16725_), .ZN(new_n16778_));
  NOR3_X1    g15776(.A1(new_n16716_), .A2(new_n16723_), .A3(new_n16684_), .ZN(new_n16779_));
  NOR2_X1    g15777(.A1(new_n16779_), .A2(new_n16778_), .ZN(new_n16780_));
  OAI21_X1   g15778(.A1(new_n16773_), .A2(new_n16774_), .B(new_n16772_), .ZN(new_n16781_));
  NAND3_X1   g15779(.A1(new_n16770_), .A2(new_n16763_), .A3(new_n16730_), .ZN(new_n16782_));
  NAND2_X1   g15780(.A1(new_n16781_), .A2(new_n16782_), .ZN(new_n16783_));
  NAND2_X1   g15781(.A1(new_n16780_), .A2(new_n16783_), .ZN(new_n16784_));
  AOI21_X1   g15782(.A1(new_n16784_), .A2(new_n16777_), .B(new_n16683_), .ZN(new_n16785_));
  OAI22_X1   g15783(.A1(new_n15526_), .A2(new_n15658_), .B1(new_n15527_), .B2(new_n15648_), .ZN(new_n16786_));
  NOR2_X1    g15784(.A1(new_n16780_), .A2(new_n16783_), .ZN(new_n16787_));
  NOR2_X1    g15785(.A1(new_n16729_), .A2(new_n16776_), .ZN(new_n16788_));
  NOR3_X1    g15786(.A1(new_n16787_), .A2(new_n16788_), .A3(new_n16786_), .ZN(new_n16789_));
  NOR2_X1    g15787(.A1(new_n16785_), .A2(new_n16789_), .ZN(new_n16790_));
  AOI22_X1   g15788(.A1(new_n15780_), .A2(new_n15898_), .B1(new_n15900_), .B2(new_n15899_), .ZN(new_n16791_));
  INV_X1     g15789(.I(new_n16791_), .ZN(new_n16792_));
  NAND3_X1   g15790(.A1(new_n15764_), .A2(new_n15761_), .A3(new_n15755_), .ZN(new_n16793_));
  AOI21_X1   g15791(.A1(new_n15776_), .A2(new_n16793_), .B(new_n15778_), .ZN(new_n16794_));
  NAND2_X1   g15792(.A1(new_n15672_), .A2(new_n14883_), .ZN(new_n16795_));
  AOI22_X1   g15793(.A1(new_n15691_), .A2(new_n14871_), .B1(new_n16795_), .B2(new_n15682_), .ZN(new_n16796_));
  NOR2_X1    g15794(.A1(new_n15669_), .A2(new_n15667_), .ZN(new_n16797_));
  OAI21_X1   g15795(.A1(new_n16797_), .A2(new_n15661_), .B(new_n15695_), .ZN(new_n16798_));
  NOR2_X1    g15796(.A1(new_n16796_), .A2(new_n16798_), .ZN(new_n16799_));
  OAI21_X1   g15797(.A1(new_n15678_), .A2(new_n15686_), .B(new_n15683_), .ZN(new_n16800_));
  NAND2_X1   g15798(.A1(new_n15696_), .A2(new_n15697_), .ZN(new_n16801_));
  AOI21_X1   g15799(.A1(new_n16801_), .A2(new_n14904_), .B(new_n15665_), .ZN(new_n16802_));
  NOR2_X1    g15800(.A1(new_n16800_), .A2(new_n16802_), .ZN(new_n16803_));
  AOI21_X1   g15801(.A1(new_n15688_), .A2(new_n15692_), .B(new_n15670_), .ZN(new_n16804_));
  OAI22_X1   g15802(.A1(new_n15770_), .A2(new_n16804_), .B1(new_n16799_), .B2(new_n16803_), .ZN(new_n16805_));
  NAND2_X1   g15803(.A1(new_n16800_), .A2(new_n16802_), .ZN(new_n16806_));
  NAND2_X1   g15804(.A1(new_n16796_), .A2(new_n16798_), .ZN(new_n16807_));
  OAI21_X1   g15805(.A1(new_n15699_), .A2(new_n15703_), .B(new_n15698_), .ZN(new_n16808_));
  NAND4_X1   g15806(.A1(new_n16808_), .A2(new_n15685_), .A3(new_n16807_), .A4(new_n16806_), .ZN(new_n16809_));
  NAND2_X1   g15807(.A1(new_n16805_), .A2(new_n16809_), .ZN(new_n16810_));
  INV_X1     g15808(.I(new_n15732_), .ZN(new_n16811_));
  NAND2_X1   g15809(.A1(new_n15725_), .A2(new_n14850_), .ZN(new_n16812_));
  NAND2_X1   g15810(.A1(new_n16812_), .A2(new_n16811_), .ZN(new_n16813_));
  OAI21_X1   g15811(.A1(new_n15730_), .A2(new_n15718_), .B(new_n16813_), .ZN(new_n16814_));
  NAND2_X1   g15812(.A1(new_n15748_), .A2(new_n15713_), .ZN(new_n16815_));
  AOI21_X1   g15813(.A1(new_n16815_), .A2(new_n14814_), .B(new_n15710_), .ZN(new_n16816_));
  NAND2_X1   g15814(.A1(new_n16814_), .A2(new_n16816_), .ZN(new_n16817_));
  AOI21_X1   g15815(.A1(new_n15741_), .A2(new_n14840_), .B(new_n15733_), .ZN(new_n16818_));
  NOR2_X1    g15816(.A1(new_n15714_), .A2(new_n15716_), .ZN(new_n16819_));
  OAI21_X1   g15817(.A1(new_n16819_), .A2(new_n15707_), .B(new_n15747_), .ZN(new_n16820_));
  NAND2_X1   g15818(.A1(new_n16820_), .A2(new_n16818_), .ZN(new_n16821_));
  OAI21_X1   g15819(.A1(new_n15750_), .A2(new_n15752_), .B(new_n15749_), .ZN(new_n16822_));
  AOI22_X1   g15820(.A1(new_n15736_), .A2(new_n16822_), .B1(new_n16821_), .B2(new_n16817_), .ZN(new_n16823_));
  NOR2_X1    g15821(.A1(new_n16820_), .A2(new_n16818_), .ZN(new_n16824_));
  NOR2_X1    g15822(.A1(new_n16814_), .A2(new_n16816_), .ZN(new_n16825_));
  AOI21_X1   g15823(.A1(new_n15742_), .A2(new_n15738_), .B(new_n15717_), .ZN(new_n16826_));
  NOR4_X1    g15824(.A1(new_n16826_), .A2(new_n16824_), .A3(new_n16825_), .A4(new_n15759_), .ZN(new_n16827_));
  NOR2_X1    g15825(.A1(new_n16823_), .A2(new_n16827_), .ZN(new_n16828_));
  NAND2_X1   g15826(.A1(new_n16810_), .A2(new_n16828_), .ZN(new_n16829_));
  AOI22_X1   g15827(.A1(new_n16808_), .A2(new_n15685_), .B1(new_n16807_), .B2(new_n16806_), .ZN(new_n16830_));
  NOR4_X1    g15828(.A1(new_n16799_), .A2(new_n16804_), .A3(new_n16803_), .A4(new_n15770_), .ZN(new_n16831_));
  NOR2_X1    g15829(.A1(new_n16830_), .A2(new_n16831_), .ZN(new_n16832_));
  OAI22_X1   g15830(.A1(new_n15759_), .A2(new_n16826_), .B1(new_n16824_), .B2(new_n16825_), .ZN(new_n16833_));
  NAND4_X1   g15831(.A1(new_n15736_), .A2(new_n16821_), .A3(new_n16822_), .A4(new_n16817_), .ZN(new_n16834_));
  NAND2_X1   g15832(.A1(new_n16833_), .A2(new_n16834_), .ZN(new_n16835_));
  NAND2_X1   g15833(.A1(new_n16832_), .A2(new_n16835_), .ZN(new_n16836_));
  AOI21_X1   g15834(.A1(new_n16836_), .A2(new_n16829_), .B(new_n16794_), .ZN(new_n16837_));
  NOR2_X1    g15835(.A1(new_n15744_), .A2(new_n15754_), .ZN(new_n16838_));
  OAI22_X1   g15836(.A1(new_n15777_), .A2(new_n15706_), .B1(new_n16838_), .B2(new_n15755_), .ZN(new_n16839_));
  NOR2_X1    g15837(.A1(new_n16832_), .A2(new_n16835_), .ZN(new_n16840_));
  NOR2_X1    g15838(.A1(new_n16810_), .A2(new_n16828_), .ZN(new_n16841_));
  NOR3_X1    g15839(.A1(new_n16839_), .A2(new_n16840_), .A3(new_n16841_), .ZN(new_n16842_));
  NOR2_X1    g15840(.A1(new_n16842_), .A2(new_n16837_), .ZN(new_n16843_));
  NOR2_X1    g15841(.A1(new_n15880_), .A2(new_n15883_), .ZN(new_n16844_));
  OAI22_X1   g15842(.A1(new_n15893_), .A2(new_n15884_), .B1(new_n16844_), .B2(new_n15822_), .ZN(new_n16845_));
  NOR2_X1    g15843(.A1(new_n15795_), .A2(new_n15796_), .ZN(new_n16846_));
  NOR2_X1    g15844(.A1(new_n15792_), .A2(new_n14793_), .ZN(new_n16847_));
  NOR2_X1    g15845(.A1(new_n16847_), .A2(new_n16846_), .ZN(new_n16848_));
  OAI21_X1   g15846(.A1(new_n16848_), .A2(new_n15800_), .B(new_n15805_), .ZN(new_n16849_));
  NAND2_X1   g15847(.A1(new_n15788_), .A2(new_n15790_), .ZN(new_n16850_));
  AOI21_X1   g15848(.A1(new_n16850_), .A2(new_n14755_), .B(new_n15785_), .ZN(new_n16851_));
  NAND2_X1   g15849(.A1(new_n16849_), .A2(new_n16851_), .ZN(new_n16852_));
  AOI21_X1   g15850(.A1(new_n15795_), .A2(new_n14793_), .B(new_n15803_), .ZN(new_n16853_));
  AOI21_X1   g15851(.A1(new_n15798_), .A2(new_n14784_), .B(new_n16853_), .ZN(new_n16854_));
  NOR2_X1    g15852(.A1(new_n15814_), .A2(new_n15813_), .ZN(new_n16855_));
  OAI21_X1   g15853(.A1(new_n16855_), .A2(new_n15799_), .B(new_n15786_), .ZN(new_n16856_));
  NAND2_X1   g15854(.A1(new_n16856_), .A2(new_n16854_), .ZN(new_n16857_));
  OAI21_X1   g15855(.A1(new_n15810_), .A2(new_n15809_), .B(new_n15791_), .ZN(new_n16858_));
  AOI22_X1   g15856(.A1(new_n16858_), .A2(new_n15887_), .B1(new_n16852_), .B2(new_n16857_), .ZN(new_n16859_));
  NOR2_X1    g15857(.A1(new_n16856_), .A2(new_n16854_), .ZN(new_n16860_));
  NOR2_X1    g15858(.A1(new_n16849_), .A2(new_n16851_), .ZN(new_n16861_));
  AOI21_X1   g15859(.A1(new_n15818_), .A2(new_n15816_), .B(new_n15815_), .ZN(new_n16862_));
  NOR4_X1    g15860(.A1(new_n16860_), .A2(new_n16861_), .A3(new_n16862_), .A4(new_n15808_), .ZN(new_n16863_));
  NOR2_X1    g15861(.A1(new_n16859_), .A2(new_n16863_), .ZN(new_n16864_));
  AOI21_X1   g15862(.A1(new_n15847_), .A2(new_n14724_), .B(new_n15853_), .ZN(new_n16865_));
  NOR2_X1    g15863(.A1(new_n15836_), .A2(new_n15826_), .ZN(new_n16866_));
  NOR2_X1    g15864(.A1(new_n15824_), .A2(new_n14704_), .ZN(new_n16867_));
  NOR2_X1    g15865(.A1(new_n16867_), .A2(new_n16866_), .ZN(new_n16868_));
  OAI21_X1   g15866(.A1(new_n16868_), .A2(new_n15848_), .B(new_n15832_), .ZN(new_n16869_));
  NOR2_X1    g15867(.A1(new_n16869_), .A2(new_n16865_), .ZN(new_n16870_));
  NOR2_X1    g15868(.A1(new_n15867_), .A2(new_n15866_), .ZN(new_n16871_));
  OAI21_X1   g15869(.A1(new_n16871_), .A2(new_n15849_), .B(new_n15859_), .ZN(new_n16872_));
  AOI21_X1   g15870(.A1(new_n15864_), .A2(new_n14694_), .B(new_n15863_), .ZN(new_n16873_));
  NOR2_X1    g15871(.A1(new_n16872_), .A2(new_n16873_), .ZN(new_n16874_));
  NOR2_X1    g15872(.A1(new_n15861_), .A2(new_n15865_), .ZN(new_n16875_));
  OAI22_X1   g15873(.A1(new_n16875_), .A2(new_n15855_), .B1(new_n16870_), .B2(new_n16874_), .ZN(new_n16876_));
  NAND2_X1   g15874(.A1(new_n16872_), .A2(new_n16873_), .ZN(new_n16877_));
  NAND2_X1   g15875(.A1(new_n16869_), .A2(new_n16865_), .ZN(new_n16878_));
  OAI21_X1   g15876(.A1(new_n15856_), .A2(new_n15860_), .B(new_n15838_), .ZN(new_n16879_));
  NAND4_X1   g15877(.A1(new_n15878_), .A2(new_n16878_), .A3(new_n16877_), .A4(new_n16879_), .ZN(new_n16880_));
  NAND2_X1   g15878(.A1(new_n16876_), .A2(new_n16880_), .ZN(new_n16881_));
  NOR2_X1    g15879(.A1(new_n16864_), .A2(new_n16881_), .ZN(new_n16882_));
  OAI22_X1   g15880(.A1(new_n16860_), .A2(new_n16861_), .B1(new_n16862_), .B2(new_n15808_), .ZN(new_n16883_));
  NAND4_X1   g15881(.A1(new_n16858_), .A2(new_n15887_), .A3(new_n16852_), .A4(new_n16857_), .ZN(new_n16884_));
  NAND2_X1   g15882(.A1(new_n16884_), .A2(new_n16883_), .ZN(new_n16885_));
  AOI22_X1   g15883(.A1(new_n15878_), .A2(new_n16879_), .B1(new_n16878_), .B2(new_n16877_), .ZN(new_n16886_));
  NOR4_X1    g15884(.A1(new_n16875_), .A2(new_n16870_), .A3(new_n16874_), .A4(new_n15855_), .ZN(new_n16887_));
  NOR2_X1    g15885(.A1(new_n16887_), .A2(new_n16886_), .ZN(new_n16888_));
  NOR2_X1    g15886(.A1(new_n16885_), .A2(new_n16888_), .ZN(new_n16889_));
  OAI21_X1   g15887(.A1(new_n16889_), .A2(new_n16882_), .B(new_n16845_), .ZN(new_n16890_));
  NAND3_X1   g15888(.A1(new_n15862_), .A2(new_n15872_), .A3(new_n15822_), .ZN(new_n16891_));
  AOI21_X1   g15889(.A1(new_n15821_), .A2(new_n16891_), .B(new_n15873_), .ZN(new_n16892_));
  NAND2_X1   g15890(.A1(new_n16885_), .A2(new_n16888_), .ZN(new_n16893_));
  NAND2_X1   g15891(.A1(new_n16864_), .A2(new_n16881_), .ZN(new_n16894_));
  NAND3_X1   g15892(.A1(new_n16893_), .A2(new_n16894_), .A3(new_n16892_), .ZN(new_n16895_));
  NAND2_X1   g15893(.A1(new_n16890_), .A2(new_n16895_), .ZN(new_n16896_));
  NOR2_X1    g15894(.A1(new_n16843_), .A2(new_n16896_), .ZN(new_n16897_));
  OAI21_X1   g15895(.A1(new_n16840_), .A2(new_n16841_), .B(new_n16839_), .ZN(new_n16898_));
  NAND3_X1   g15896(.A1(new_n16836_), .A2(new_n16829_), .A3(new_n16794_), .ZN(new_n16899_));
  NAND2_X1   g15897(.A1(new_n16898_), .A2(new_n16899_), .ZN(new_n16900_));
  AOI21_X1   g15898(.A1(new_n16893_), .A2(new_n16894_), .B(new_n16892_), .ZN(new_n16901_));
  NOR3_X1    g15899(.A1(new_n16882_), .A2(new_n16889_), .A3(new_n16845_), .ZN(new_n16902_));
  NOR2_X1    g15900(.A1(new_n16902_), .A2(new_n16901_), .ZN(new_n16903_));
  NOR2_X1    g15901(.A1(new_n16900_), .A2(new_n16903_), .ZN(new_n16904_));
  OAI21_X1   g15902(.A1(new_n16904_), .A2(new_n16897_), .B(new_n16792_), .ZN(new_n16905_));
  NAND2_X1   g15903(.A1(new_n16900_), .A2(new_n16903_), .ZN(new_n16906_));
  NAND2_X1   g15904(.A1(new_n16843_), .A2(new_n16896_), .ZN(new_n16907_));
  NAND3_X1   g15905(.A1(new_n16906_), .A2(new_n16907_), .A3(new_n16791_), .ZN(new_n16908_));
  NAND2_X1   g15906(.A1(new_n16905_), .A2(new_n16908_), .ZN(new_n16909_));
  NOR2_X1    g15907(.A1(new_n16790_), .A2(new_n16909_), .ZN(new_n16910_));
  OAI21_X1   g15908(.A1(new_n16787_), .A2(new_n16788_), .B(new_n16786_), .ZN(new_n16911_));
  NAND3_X1   g15909(.A1(new_n16784_), .A2(new_n16777_), .A3(new_n16683_), .ZN(new_n16912_));
  NAND2_X1   g15910(.A1(new_n16911_), .A2(new_n16912_), .ZN(new_n16913_));
  AOI21_X1   g15911(.A1(new_n16906_), .A2(new_n16907_), .B(new_n16791_), .ZN(new_n16914_));
  NOR3_X1    g15912(.A1(new_n16904_), .A2(new_n16897_), .A3(new_n16792_), .ZN(new_n16915_));
  NOR2_X1    g15913(.A1(new_n16914_), .A2(new_n16915_), .ZN(new_n16916_));
  NOR2_X1    g15914(.A1(new_n16913_), .A2(new_n16916_), .ZN(new_n16917_));
  OAI21_X1   g15915(.A1(new_n16917_), .A2(new_n16910_), .B(new_n16674_), .ZN(new_n16918_));
  AOI21_X1   g15916(.A1(new_n15911_), .A2(new_n15910_), .B(new_n15907_), .ZN(new_n16919_));
  AOI21_X1   g15917(.A1(new_n15660_), .A2(new_n15916_), .B(new_n16919_), .ZN(new_n16920_));
  NAND2_X1   g15918(.A1(new_n16913_), .A2(new_n16916_), .ZN(new_n16921_));
  NAND3_X1   g15919(.A1(new_n16909_), .A2(new_n16911_), .A3(new_n16912_), .ZN(new_n16922_));
  NAND3_X1   g15920(.A1(new_n16921_), .A2(new_n16922_), .A3(new_n16920_), .ZN(new_n16923_));
  NAND2_X1   g15921(.A1(new_n16918_), .A2(new_n16923_), .ZN(new_n16924_));
  NOR2_X1    g15922(.A1(new_n16672_), .A2(new_n16924_), .ZN(new_n16925_));
  OAI21_X1   g15923(.A1(new_n16670_), .A2(new_n16669_), .B(new_n16668_), .ZN(new_n16926_));
  NAND3_X1   g15924(.A1(new_n16658_), .A2(new_n16665_), .A3(new_n16428_), .ZN(new_n16927_));
  NAND2_X1   g15925(.A1(new_n16926_), .A2(new_n16927_), .ZN(new_n16928_));
  AOI21_X1   g15926(.A1(new_n16921_), .A2(new_n16922_), .B(new_n16920_), .ZN(new_n16929_));
  NOR3_X1    g15927(.A1(new_n16917_), .A2(new_n16910_), .A3(new_n16674_), .ZN(new_n16930_));
  NOR2_X1    g15928(.A1(new_n16930_), .A2(new_n16929_), .ZN(new_n16931_));
  NOR2_X1    g15929(.A1(new_n16928_), .A2(new_n16931_), .ZN(new_n16932_));
  OAI21_X1   g15930(.A1(new_n16932_), .A2(new_n16925_), .B(new_n16426_), .ZN(new_n16933_));
  OAI21_X1   g15931(.A1(new_n15908_), .A2(new_n15912_), .B(new_n15915_), .ZN(new_n16934_));
  OAI21_X1   g15932(.A1(new_n16919_), .A2(new_n16673_), .B(new_n15660_), .ZN(new_n16935_));
  AOI21_X1   g15933(.A1(new_n16934_), .A2(new_n16935_), .B(new_n15407_), .ZN(new_n16936_));
  INV_X1     g15934(.I(new_n16424_), .ZN(new_n16937_));
  NAND3_X1   g15935(.A1(new_n16934_), .A2(new_n15407_), .A3(new_n16935_), .ZN(new_n16938_));
  AOI21_X1   g15936(.A1(new_n16937_), .A2(new_n16938_), .B(new_n16936_), .ZN(new_n16939_));
  NAND2_X1   g15937(.A1(new_n16928_), .A2(new_n16931_), .ZN(new_n16940_));
  NAND3_X1   g15938(.A1(new_n16924_), .A2(new_n16926_), .A3(new_n16927_), .ZN(new_n16941_));
  NAND3_X1   g15939(.A1(new_n16940_), .A2(new_n16941_), .A3(new_n16939_), .ZN(new_n16942_));
  NAND4_X1   g15940(.A1(new_n14422_), .A2(new_n16933_), .A3(new_n14431_), .A4(new_n16942_), .ZN(new_n16943_));
  XNOR2_X1   g15941(.A1(new_n15406_), .A2(new_n14914_), .ZN(new_n16944_));
  XNOR2_X1   g15942(.A1(new_n12395_), .A2(new_n12912_), .ZN(new_n16945_));
  NOR2_X1    g15943(.A1(new_n16945_), .A2(new_n16944_), .ZN(new_n16946_));
  INV_X1     g15944(.I(new_n16946_), .ZN(new_n16947_));
  NAND3_X1   g15945(.A1(new_n16934_), .A2(new_n15408_), .A3(new_n16935_), .ZN(new_n16948_));
  OAI21_X1   g15946(.A1(new_n15914_), .A2(new_n15918_), .B(new_n15407_), .ZN(new_n16949_));
  AOI21_X1   g15947(.A1(new_n16949_), .A2(new_n16948_), .B(new_n16937_), .ZN(new_n16950_));
  AOI21_X1   g15948(.A1(new_n15919_), .A2(new_n16938_), .B(new_n16424_), .ZN(new_n16951_));
  NOR2_X1    g15949(.A1(new_n16950_), .A2(new_n16951_), .ZN(new_n16952_));
  NAND3_X1   g15950(.A1(new_n14425_), .A2(new_n14424_), .A3(new_n12914_), .ZN(new_n16953_));
  NAND2_X1   g15951(.A1(new_n14426_), .A2(new_n12913_), .ZN(new_n16954_));
  AOI21_X1   g15952(.A1(new_n16954_), .A2(new_n16953_), .B(new_n13933_), .ZN(new_n16955_));
  AOI21_X1   g15953(.A1(new_n14427_), .A2(new_n13422_), .B(new_n13934_), .ZN(new_n16956_));
  NOR2_X1    g15954(.A1(new_n16955_), .A2(new_n16956_), .ZN(new_n16957_));
  NOR3_X1    g15955(.A1(new_n16950_), .A2(new_n16951_), .A3(new_n16946_), .ZN(new_n16958_));
  OAI22_X1   g15956(.A1(new_n16957_), .A2(new_n16958_), .B1(new_n16947_), .B2(new_n16952_), .ZN(new_n16959_));
  INV_X1     g15957(.I(new_n16959_), .ZN(new_n16960_));
  AOI22_X1   g15958(.A1(new_n14422_), .A2(new_n14431_), .B1(new_n16933_), .B2(new_n16942_), .ZN(new_n16961_));
  OAI21_X1   g15959(.A1(new_n16961_), .A2(new_n16960_), .B(new_n16943_), .ZN(new_n16962_));
  NOR2_X1    g15960(.A1(new_n16928_), .A2(new_n16924_), .ZN(new_n16963_));
  AOI21_X1   g15961(.A1(new_n16928_), .A2(new_n16924_), .B(new_n16939_), .ZN(new_n16964_));
  NOR2_X1    g15962(.A1(new_n16964_), .A2(new_n16963_), .ZN(new_n16965_));
  NOR2_X1    g15963(.A1(new_n16913_), .A2(new_n16909_), .ZN(new_n16966_));
  AOI21_X1   g15964(.A1(new_n16913_), .A2(new_n16909_), .B(new_n16920_), .ZN(new_n16967_));
  NAND2_X1   g15965(.A1(new_n16780_), .A2(new_n16776_), .ZN(new_n16968_));
  OAI21_X1   g15966(.A1(new_n16780_), .A2(new_n16776_), .B(new_n16786_), .ZN(new_n16969_));
  NAND2_X1   g15967(.A1(new_n16756_), .A2(new_n15631_), .ZN(new_n16970_));
  NAND3_X1   g15968(.A1(new_n16756_), .A2(new_n15631_), .A3(new_n16748_), .ZN(new_n16971_));
  AOI22_X1   g15969(.A1(new_n16971_), .A2(new_n16750_), .B1(new_n16970_), .B2(new_n16752_), .ZN(new_n16972_));
  OAI21_X1   g15970(.A1(new_n16739_), .A2(new_n15570_), .B(new_n16731_), .ZN(new_n16973_));
  NAND2_X1   g15971(.A1(new_n15642_), .A2(new_n16736_), .ZN(new_n16974_));
  OAI21_X1   g15972(.A1(new_n16974_), .A2(new_n16739_), .B(new_n16737_), .ZN(new_n16975_));
  NAND2_X1   g15973(.A1(new_n16975_), .A2(new_n16973_), .ZN(new_n16976_));
  NOR2_X1    g15974(.A1(new_n16976_), .A2(new_n16972_), .ZN(new_n16977_));
  INV_X1     g15975(.I(new_n16972_), .ZN(new_n16978_));
  NAND2_X1   g15976(.A1(new_n16743_), .A2(new_n15642_), .ZN(new_n16979_));
  NAND3_X1   g15977(.A1(new_n16743_), .A2(new_n15642_), .A3(new_n16736_), .ZN(new_n16980_));
  AOI22_X1   g15978(.A1(new_n16980_), .A2(new_n16737_), .B1(new_n16979_), .B2(new_n16731_), .ZN(new_n16981_));
  NOR2_X1    g15979(.A1(new_n16978_), .A2(new_n16981_), .ZN(new_n16982_));
  NOR2_X1    g15980(.A1(new_n16982_), .A2(new_n16977_), .ZN(new_n16983_));
  NAND2_X1   g15981(.A1(new_n16745_), .A2(new_n16769_), .ZN(new_n16984_));
  NAND2_X1   g15982(.A1(new_n16984_), .A2(new_n16772_), .ZN(new_n16985_));
  INV_X1     g15983(.I(new_n16985_), .ZN(new_n16986_));
  NAND4_X1   g15984(.A1(new_n16740_), .A2(new_n16744_), .A3(new_n16767_), .A4(new_n16768_), .ZN(new_n16987_));
  INV_X1     g15985(.I(new_n16987_), .ZN(new_n16988_));
  AOI21_X1   g15986(.A1(new_n16984_), .A2(new_n16772_), .B(new_n16988_), .ZN(new_n16989_));
  NAND2_X1   g15987(.A1(new_n16978_), .A2(new_n16981_), .ZN(new_n16990_));
  NAND2_X1   g15988(.A1(new_n16976_), .A2(new_n16972_), .ZN(new_n16991_));
  NAND3_X1   g15989(.A1(new_n16990_), .A2(new_n16991_), .A3(new_n16987_), .ZN(new_n16992_));
  OAI22_X1   g15990(.A1(new_n16986_), .A2(new_n16992_), .B1(new_n16989_), .B2(new_n16983_), .ZN(new_n16993_));
  OAI21_X1   g15991(.A1(new_n16709_), .A2(new_n15500_), .B(new_n16701_), .ZN(new_n16994_));
  OAI21_X1   g15992(.A1(new_n15498_), .A2(new_n15499_), .B(new_n16705_), .ZN(new_n16995_));
  OAI21_X1   g15993(.A1(new_n16995_), .A2(new_n16709_), .B(new_n16707_), .ZN(new_n16996_));
  NAND2_X1   g15994(.A1(new_n16996_), .A2(new_n16994_), .ZN(new_n16997_));
  AOI21_X1   g15995(.A1(new_n16693_), .A2(new_n15519_), .B(new_n16685_), .ZN(new_n16998_));
  NOR2_X1    g15996(.A1(new_n15439_), .A2(new_n16689_), .ZN(new_n16999_));
  AOI21_X1   g15997(.A1(new_n16999_), .A2(new_n16693_), .B(new_n16691_), .ZN(new_n17000_));
  NOR2_X1    g15998(.A1(new_n17000_), .A2(new_n16998_), .ZN(new_n17001_));
  NAND2_X1   g15999(.A1(new_n17001_), .A2(new_n16997_), .ZN(new_n17002_));
  INV_X1     g16000(.I(new_n16997_), .ZN(new_n17003_));
  NOR2_X1    g16001(.A1(new_n16697_), .A2(new_n15439_), .ZN(new_n17004_));
  NAND2_X1   g16002(.A1(new_n15519_), .A2(new_n16685_), .ZN(new_n17005_));
  NOR2_X1    g16003(.A1(new_n17005_), .A2(new_n16697_), .ZN(new_n17006_));
  OAI22_X1   g16004(.A1(new_n17006_), .A2(new_n16691_), .B1(new_n16685_), .B2(new_n17004_), .ZN(new_n17007_));
  NAND2_X1   g16005(.A1(new_n17003_), .A2(new_n17007_), .ZN(new_n17008_));
  NAND2_X1   g16006(.A1(new_n17008_), .A2(new_n17002_), .ZN(new_n17009_));
  NAND2_X1   g16007(.A1(new_n16719_), .A2(new_n16715_), .ZN(new_n17010_));
  NAND2_X1   g16008(.A1(new_n17010_), .A2(new_n16684_), .ZN(new_n17011_));
  NOR2_X1    g16009(.A1(new_n16699_), .A2(new_n16722_), .ZN(new_n17012_));
  NAND4_X1   g16010(.A1(new_n16718_), .A2(new_n16717_), .A3(new_n16714_), .A4(new_n16710_), .ZN(new_n17013_));
  OAI21_X1   g16011(.A1(new_n17012_), .A2(new_n16725_), .B(new_n17013_), .ZN(new_n17014_));
  NOR2_X1    g16012(.A1(new_n17003_), .A2(new_n17007_), .ZN(new_n17015_));
  NOR2_X1    g16013(.A1(new_n17001_), .A2(new_n16997_), .ZN(new_n17016_));
  INV_X1     g16014(.I(new_n17013_), .ZN(new_n17017_));
  NOR3_X1    g16015(.A1(new_n17015_), .A2(new_n17017_), .A3(new_n17016_), .ZN(new_n17018_));
  AOI22_X1   g16016(.A1(new_n17018_), .A2(new_n17011_), .B1(new_n17014_), .B2(new_n17009_), .ZN(new_n17019_));
  NAND2_X1   g16017(.A1(new_n16993_), .A2(new_n17019_), .ZN(new_n17020_));
  NAND2_X1   g16018(.A1(new_n16990_), .A2(new_n16991_), .ZN(new_n17021_));
  NOR2_X1    g16019(.A1(new_n16766_), .A2(new_n16762_), .ZN(new_n17022_));
  OAI21_X1   g16020(.A1(new_n17022_), .A2(new_n16730_), .B(new_n16987_), .ZN(new_n17023_));
  NOR3_X1    g16021(.A1(new_n16982_), .A2(new_n16977_), .A3(new_n16988_), .ZN(new_n17024_));
  AOI22_X1   g16022(.A1(new_n17024_), .A2(new_n16985_), .B1(new_n17021_), .B2(new_n17023_), .ZN(new_n17025_));
  NOR2_X1    g16023(.A1(new_n17015_), .A2(new_n17016_), .ZN(new_n17026_));
  NOR2_X1    g16024(.A1(new_n17012_), .A2(new_n16725_), .ZN(new_n17027_));
  AOI21_X1   g16025(.A1(new_n17010_), .A2(new_n16684_), .B(new_n17017_), .ZN(new_n17028_));
  NAND3_X1   g16026(.A1(new_n17008_), .A2(new_n17002_), .A3(new_n17013_), .ZN(new_n17029_));
  OAI22_X1   g16027(.A1(new_n17028_), .A2(new_n17026_), .B1(new_n17029_), .B2(new_n17027_), .ZN(new_n17030_));
  NAND2_X1   g16028(.A1(new_n17030_), .A2(new_n17025_), .ZN(new_n17031_));
  AOI22_X1   g16029(.A1(new_n16969_), .A2(new_n16968_), .B1(new_n17020_), .B2(new_n17031_), .ZN(new_n17032_));
  NOR2_X1    g16030(.A1(new_n16729_), .A2(new_n16783_), .ZN(new_n17033_));
  AOI21_X1   g16031(.A1(new_n16729_), .A2(new_n16783_), .B(new_n16683_), .ZN(new_n17034_));
  NOR2_X1    g16032(.A1(new_n17030_), .A2(new_n17025_), .ZN(new_n17035_));
  NOR2_X1    g16033(.A1(new_n16993_), .A2(new_n17019_), .ZN(new_n17036_));
  NOR4_X1    g16034(.A1(new_n17034_), .A2(new_n17036_), .A3(new_n17035_), .A4(new_n17033_), .ZN(new_n17037_));
  NOR2_X1    g16035(.A1(new_n17032_), .A2(new_n17037_), .ZN(new_n17038_));
  NOR2_X1    g16036(.A1(new_n16900_), .A2(new_n16896_), .ZN(new_n17039_));
  AOI21_X1   g16037(.A1(new_n16900_), .A2(new_n16896_), .B(new_n16791_), .ZN(new_n17040_));
  OAI21_X1   g16038(.A1(new_n16875_), .A2(new_n15855_), .B(new_n16865_), .ZN(new_n17041_));
  OAI21_X1   g16039(.A1(new_n15851_), .A2(new_n15854_), .B(new_n16872_), .ZN(new_n17042_));
  OAI21_X1   g16040(.A1(new_n16875_), .A2(new_n17042_), .B(new_n16873_), .ZN(new_n17043_));
  NAND2_X1   g16041(.A1(new_n17043_), .A2(new_n17041_), .ZN(new_n17044_));
  NAND2_X1   g16042(.A1(new_n16858_), .A2(new_n15887_), .ZN(new_n17045_));
  NAND3_X1   g16043(.A1(new_n16858_), .A2(new_n15887_), .A3(new_n16849_), .ZN(new_n17046_));
  AOI22_X1   g16044(.A1(new_n17046_), .A2(new_n16851_), .B1(new_n17045_), .B2(new_n16854_), .ZN(new_n17047_));
  NAND2_X1   g16045(.A1(new_n17047_), .A2(new_n17044_), .ZN(new_n17048_));
  INV_X1     g16046(.I(new_n17044_), .ZN(new_n17049_));
  OAI21_X1   g16047(.A1(new_n16862_), .A2(new_n15808_), .B(new_n16854_), .ZN(new_n17050_));
  NAND2_X1   g16048(.A1(new_n17046_), .A2(new_n16851_), .ZN(new_n17051_));
  NAND2_X1   g16049(.A1(new_n17051_), .A2(new_n17050_), .ZN(new_n17052_));
  NAND2_X1   g16050(.A1(new_n17052_), .A2(new_n17049_), .ZN(new_n17053_));
  NAND2_X1   g16051(.A1(new_n17053_), .A2(new_n17048_), .ZN(new_n17054_));
  NAND2_X1   g16052(.A1(new_n16885_), .A2(new_n16881_), .ZN(new_n17055_));
  NAND2_X1   g16053(.A1(new_n17055_), .A2(new_n16845_), .ZN(new_n17056_));
  NOR2_X1    g16054(.A1(new_n16864_), .A2(new_n16888_), .ZN(new_n17057_));
  NAND4_X1   g16055(.A1(new_n16884_), .A2(new_n16876_), .A3(new_n16883_), .A4(new_n16880_), .ZN(new_n17058_));
  OAI21_X1   g16056(.A1(new_n17057_), .A2(new_n16892_), .B(new_n17058_), .ZN(new_n17059_));
  NOR2_X1    g16057(.A1(new_n17052_), .A2(new_n17049_), .ZN(new_n17060_));
  NOR2_X1    g16058(.A1(new_n17047_), .A2(new_n17044_), .ZN(new_n17061_));
  INV_X1     g16059(.I(new_n17058_), .ZN(new_n17062_));
  NOR3_X1    g16060(.A1(new_n17060_), .A2(new_n17061_), .A3(new_n17062_), .ZN(new_n17063_));
  AOI22_X1   g16061(.A1(new_n17063_), .A2(new_n17056_), .B1(new_n17054_), .B2(new_n17059_), .ZN(new_n17064_));
  OAI21_X1   g16062(.A1(new_n16826_), .A2(new_n15759_), .B(new_n16818_), .ZN(new_n17065_));
  OAI21_X1   g16063(.A1(new_n15757_), .A2(new_n15758_), .B(new_n16814_), .ZN(new_n17066_));
  OAI21_X1   g16064(.A1(new_n17066_), .A2(new_n16826_), .B(new_n16816_), .ZN(new_n17067_));
  NAND2_X1   g16065(.A1(new_n17067_), .A2(new_n17065_), .ZN(new_n17068_));
  OAI21_X1   g16066(.A1(new_n16804_), .A2(new_n15770_), .B(new_n16796_), .ZN(new_n17069_));
  OAI21_X1   g16067(.A1(new_n15768_), .A2(new_n15769_), .B(new_n16800_), .ZN(new_n17070_));
  OAI21_X1   g16068(.A1(new_n17070_), .A2(new_n16804_), .B(new_n16802_), .ZN(new_n17071_));
  NAND3_X1   g16069(.A1(new_n17068_), .A2(new_n17069_), .A3(new_n17071_), .ZN(new_n17072_));
  NAND2_X1   g16070(.A1(new_n17071_), .A2(new_n17069_), .ZN(new_n17073_));
  NAND3_X1   g16071(.A1(new_n17073_), .A2(new_n17065_), .A3(new_n17067_), .ZN(new_n17074_));
  NAND2_X1   g16072(.A1(new_n17072_), .A2(new_n17074_), .ZN(new_n17075_));
  INV_X1     g16073(.I(new_n17075_), .ZN(new_n17076_));
  NOR2_X1    g16074(.A1(new_n16832_), .A2(new_n16828_), .ZN(new_n17077_));
  NOR2_X1    g16075(.A1(new_n17077_), .A2(new_n16794_), .ZN(new_n17078_));
  NAND2_X1   g16076(.A1(new_n16810_), .A2(new_n16835_), .ZN(new_n17079_));
  NAND4_X1   g16077(.A1(new_n16805_), .A2(new_n16809_), .A3(new_n16833_), .A4(new_n16834_), .ZN(new_n17080_));
  INV_X1     g16078(.I(new_n17080_), .ZN(new_n17081_));
  AOI21_X1   g16079(.A1(new_n16839_), .A2(new_n17079_), .B(new_n17081_), .ZN(new_n17082_));
  NAND3_X1   g16080(.A1(new_n17072_), .A2(new_n17074_), .A3(new_n17080_), .ZN(new_n17083_));
  OAI22_X1   g16081(.A1(new_n17082_), .A2(new_n17076_), .B1(new_n17078_), .B2(new_n17083_), .ZN(new_n17084_));
  NOR2_X1    g16082(.A1(new_n17064_), .A2(new_n17084_), .ZN(new_n17085_));
  NOR2_X1    g16083(.A1(new_n17060_), .A2(new_n17061_), .ZN(new_n17086_));
  INV_X1     g16084(.I(new_n17056_), .ZN(new_n17087_));
  AOI21_X1   g16085(.A1(new_n16845_), .A2(new_n17055_), .B(new_n17062_), .ZN(new_n17088_));
  NAND3_X1   g16086(.A1(new_n17053_), .A2(new_n17048_), .A3(new_n17058_), .ZN(new_n17089_));
  OAI22_X1   g16087(.A1(new_n17087_), .A2(new_n17089_), .B1(new_n17086_), .B2(new_n17088_), .ZN(new_n17090_));
  NAND2_X1   g16088(.A1(new_n16839_), .A2(new_n17079_), .ZN(new_n17091_));
  OAI21_X1   g16089(.A1(new_n17077_), .A2(new_n16794_), .B(new_n17080_), .ZN(new_n17092_));
  INV_X1     g16090(.I(new_n17083_), .ZN(new_n17093_));
  AOI22_X1   g16091(.A1(new_n17093_), .A2(new_n17091_), .B1(new_n17075_), .B2(new_n17092_), .ZN(new_n17094_));
  NOR2_X1    g16092(.A1(new_n17090_), .A2(new_n17094_), .ZN(new_n17095_));
  OAI22_X1   g16093(.A1(new_n17085_), .A2(new_n17095_), .B1(new_n17039_), .B2(new_n17040_), .ZN(new_n17096_));
  NOR2_X1    g16094(.A1(new_n17040_), .A2(new_n17039_), .ZN(new_n17097_));
  NAND2_X1   g16095(.A1(new_n17090_), .A2(new_n17094_), .ZN(new_n17098_));
  NAND2_X1   g16096(.A1(new_n17064_), .A2(new_n17084_), .ZN(new_n17099_));
  NAND3_X1   g16097(.A1(new_n17097_), .A2(new_n17098_), .A3(new_n17099_), .ZN(new_n17100_));
  NAND2_X1   g16098(.A1(new_n17100_), .A2(new_n17096_), .ZN(new_n17101_));
  NOR2_X1    g16099(.A1(new_n17101_), .A2(new_n17038_), .ZN(new_n17102_));
  OAI22_X1   g16100(.A1(new_n17033_), .A2(new_n17034_), .B1(new_n17036_), .B2(new_n17035_), .ZN(new_n17103_));
  NAND4_X1   g16101(.A1(new_n16969_), .A2(new_n17020_), .A3(new_n17031_), .A4(new_n16968_), .ZN(new_n17104_));
  NAND2_X1   g16102(.A1(new_n17103_), .A2(new_n17104_), .ZN(new_n17105_));
  NAND2_X1   g16103(.A1(new_n16843_), .A2(new_n16903_), .ZN(new_n17106_));
  INV_X1     g16104(.I(new_n17040_), .ZN(new_n17107_));
  AOI22_X1   g16105(.A1(new_n17107_), .A2(new_n17106_), .B1(new_n17098_), .B2(new_n17099_), .ZN(new_n17108_));
  NOR2_X1    g16106(.A1(new_n16843_), .A2(new_n16903_), .ZN(new_n17109_));
  OAI21_X1   g16107(.A1(new_n16791_), .A2(new_n17109_), .B(new_n17106_), .ZN(new_n17110_));
  NOR3_X1    g16108(.A1(new_n17110_), .A2(new_n17085_), .A3(new_n17095_), .ZN(new_n17111_));
  NOR2_X1    g16109(.A1(new_n17108_), .A2(new_n17111_), .ZN(new_n17112_));
  NOR2_X1    g16110(.A1(new_n17112_), .A2(new_n17105_), .ZN(new_n17113_));
  OAI22_X1   g16111(.A1(new_n17113_), .A2(new_n17102_), .B1(new_n16967_), .B2(new_n16966_), .ZN(new_n17114_));
  NAND2_X1   g16112(.A1(new_n16790_), .A2(new_n16916_), .ZN(new_n17115_));
  OAI21_X1   g16113(.A1(new_n16790_), .A2(new_n16916_), .B(new_n16674_), .ZN(new_n17116_));
  NAND2_X1   g16114(.A1(new_n17112_), .A2(new_n17105_), .ZN(new_n17117_));
  NAND2_X1   g16115(.A1(new_n17101_), .A2(new_n17038_), .ZN(new_n17118_));
  NAND4_X1   g16116(.A1(new_n17117_), .A2(new_n17118_), .A3(new_n17116_), .A4(new_n17115_), .ZN(new_n17119_));
  NAND2_X1   g16117(.A1(new_n17114_), .A2(new_n17119_), .ZN(new_n17120_));
  NAND2_X1   g16118(.A1(new_n16661_), .A2(new_n16657_), .ZN(new_n17121_));
  OAI21_X1   g16119(.A1(new_n16661_), .A2(new_n16657_), .B(new_n16668_), .ZN(new_n17122_));
  NOR2_X1    g16120(.A1(new_n16586_), .A2(new_n16650_), .ZN(new_n17123_));
  AOI21_X1   g16121(.A1(new_n16586_), .A2(new_n16650_), .B(new_n16535_), .ZN(new_n17124_));
  NAND2_X1   g16122(.A1(new_n16381_), .A2(new_n16622_), .ZN(new_n17125_));
  NAND2_X1   g16123(.A1(new_n17125_), .A2(new_n16618_), .ZN(new_n17126_));
  NAND3_X1   g16124(.A1(new_n16381_), .A2(new_n16613_), .A3(new_n16622_), .ZN(new_n17127_));
  NAND2_X1   g16125(.A1(new_n17127_), .A2(new_n16615_), .ZN(new_n17128_));
  NAND2_X1   g16126(.A1(new_n17128_), .A2(new_n17126_), .ZN(new_n17129_));
  NAND2_X1   g16127(.A1(new_n16390_), .A2(new_n16603_), .ZN(new_n17130_));
  NAND3_X1   g16128(.A1(new_n16390_), .A2(new_n16603_), .A3(new_n16598_), .ZN(new_n17131_));
  AOI22_X1   g16129(.A1(new_n17131_), .A2(new_n16601_), .B1(new_n17130_), .B2(new_n16590_), .ZN(new_n17132_));
  NAND2_X1   g16130(.A1(new_n17129_), .A2(new_n17132_), .ZN(new_n17133_));
  AOI22_X1   g16131(.A1(new_n17127_), .A2(new_n16615_), .B1(new_n17125_), .B2(new_n16618_), .ZN(new_n17134_));
  INV_X1     g16132(.I(new_n17132_), .ZN(new_n17135_));
  NAND2_X1   g16133(.A1(new_n17135_), .A2(new_n17134_), .ZN(new_n17136_));
  NAND2_X1   g16134(.A1(new_n17136_), .A2(new_n17133_), .ZN(new_n17137_));
  NOR2_X1    g16135(.A1(new_n16632_), .A2(new_n16628_), .ZN(new_n17138_));
  NOR2_X1    g16136(.A1(new_n17138_), .A2(new_n16588_), .ZN(new_n17139_));
  INV_X1     g16137(.I(new_n17139_), .ZN(new_n17140_));
  NAND4_X1   g16138(.A1(new_n16605_), .A2(new_n16608_), .A3(new_n16633_), .A4(new_n16634_), .ZN(new_n17141_));
  OAI21_X1   g16139(.A1(new_n17138_), .A2(new_n16588_), .B(new_n17141_), .ZN(new_n17142_));
  NOR2_X1    g16140(.A1(new_n17135_), .A2(new_n17134_), .ZN(new_n17143_));
  NOR2_X1    g16141(.A1(new_n17129_), .A2(new_n17132_), .ZN(new_n17144_));
  INV_X1     g16142(.I(new_n17141_), .ZN(new_n17145_));
  NOR3_X1    g16143(.A1(new_n17143_), .A2(new_n17144_), .A3(new_n17145_), .ZN(new_n17146_));
  AOI22_X1   g16144(.A1(new_n17140_), .A2(new_n17146_), .B1(new_n17137_), .B2(new_n17142_), .ZN(new_n17147_));
  NOR2_X1    g16145(.A1(new_n16565_), .A2(new_n16262_), .ZN(new_n17148_));
  NOR3_X1    g16146(.A1(new_n16565_), .A2(new_n16262_), .A3(new_n16554_), .ZN(new_n17149_));
  OAI22_X1   g16147(.A1(new_n17149_), .A2(new_n16556_), .B1(new_n17148_), .B2(new_n16561_), .ZN(new_n17150_));
  INV_X1     g16148(.I(new_n17150_), .ZN(new_n17151_));
  NAND2_X1   g16149(.A1(new_n16546_), .A2(new_n16197_), .ZN(new_n17152_));
  NAND2_X1   g16150(.A1(new_n17152_), .A2(new_n16542_), .ZN(new_n17153_));
  NAND3_X1   g16151(.A1(new_n16546_), .A2(new_n16197_), .A3(new_n16538_), .ZN(new_n17154_));
  NAND2_X1   g16152(.A1(new_n17154_), .A2(new_n16540_), .ZN(new_n17155_));
  NAND2_X1   g16153(.A1(new_n17155_), .A2(new_n17153_), .ZN(new_n17156_));
  NOR2_X1    g16154(.A1(new_n17151_), .A2(new_n17156_), .ZN(new_n17157_));
  AOI22_X1   g16155(.A1(new_n17154_), .A2(new_n16540_), .B1(new_n17152_), .B2(new_n16542_), .ZN(new_n17158_));
  NOR2_X1    g16156(.A1(new_n17158_), .A2(new_n17150_), .ZN(new_n17159_));
  NOR2_X1    g16157(.A1(new_n17157_), .A2(new_n17159_), .ZN(new_n17160_));
  NAND2_X1   g16158(.A1(new_n16575_), .A2(new_n16571_), .ZN(new_n17161_));
  NAND2_X1   g16159(.A1(new_n16537_), .A2(new_n17161_), .ZN(new_n17162_));
  INV_X1     g16160(.I(new_n17162_), .ZN(new_n17163_));
  NAND4_X1   g16161(.A1(new_n16573_), .A2(new_n16574_), .A3(new_n16570_), .A4(new_n16566_), .ZN(new_n17164_));
  INV_X1     g16162(.I(new_n17164_), .ZN(new_n17165_));
  AOI21_X1   g16163(.A1(new_n17161_), .A2(new_n16537_), .B(new_n17165_), .ZN(new_n17166_));
  NAND2_X1   g16164(.A1(new_n17158_), .A2(new_n17150_), .ZN(new_n17167_));
  INV_X1     g16165(.I(new_n17159_), .ZN(new_n17168_));
  NAND3_X1   g16166(.A1(new_n17168_), .A2(new_n17167_), .A3(new_n17164_), .ZN(new_n17169_));
  OAI22_X1   g16167(.A1(new_n17163_), .A2(new_n17169_), .B1(new_n17166_), .B2(new_n17160_), .ZN(new_n17170_));
  NOR2_X1    g16168(.A1(new_n17170_), .A2(new_n17147_), .ZN(new_n17171_));
  NOR2_X1    g16169(.A1(new_n17143_), .A2(new_n17144_), .ZN(new_n17172_));
  NAND2_X1   g16170(.A1(new_n16609_), .A2(new_n16635_), .ZN(new_n17173_));
  AOI21_X1   g16171(.A1(new_n17173_), .A2(new_n16639_), .B(new_n17145_), .ZN(new_n17174_));
  NAND3_X1   g16172(.A1(new_n17136_), .A2(new_n17133_), .A3(new_n17141_), .ZN(new_n17175_));
  OAI22_X1   g16173(.A1(new_n17139_), .A2(new_n17175_), .B1(new_n17174_), .B2(new_n17172_), .ZN(new_n17176_));
  NAND2_X1   g16174(.A1(new_n17168_), .A2(new_n17167_), .ZN(new_n17177_));
  NOR2_X1    g16175(.A1(new_n16552_), .A2(new_n16578_), .ZN(new_n17178_));
  OAI21_X1   g16176(.A1(new_n17178_), .A2(new_n16582_), .B(new_n17164_), .ZN(new_n17179_));
  NOR3_X1    g16177(.A1(new_n17157_), .A2(new_n17159_), .A3(new_n17165_), .ZN(new_n17180_));
  AOI22_X1   g16178(.A1(new_n17180_), .A2(new_n17162_), .B1(new_n17177_), .B2(new_n17179_), .ZN(new_n17181_));
  NOR2_X1    g16179(.A1(new_n17181_), .A2(new_n17176_), .ZN(new_n17182_));
  OAI22_X1   g16180(.A1(new_n17171_), .A2(new_n17182_), .B1(new_n17123_), .B2(new_n17124_), .ZN(new_n17183_));
  NOR2_X1    g16181(.A1(new_n17124_), .A2(new_n17123_), .ZN(new_n17184_));
  NAND2_X1   g16182(.A1(new_n17181_), .A2(new_n17176_), .ZN(new_n17185_));
  NAND2_X1   g16183(.A1(new_n17170_), .A2(new_n17147_), .ZN(new_n17186_));
  NAND3_X1   g16184(.A1(new_n17184_), .A2(new_n17185_), .A3(new_n17186_), .ZN(new_n17187_));
  NAND2_X1   g16185(.A1(new_n17187_), .A2(new_n17183_), .ZN(new_n17188_));
  NAND2_X1   g16186(.A1(new_n16473_), .A2(new_n16527_), .ZN(new_n17189_));
  OAI21_X1   g16187(.A1(new_n16473_), .A2(new_n16527_), .B(new_n16430_), .ZN(new_n17190_));
  NOR2_X1    g16188(.A1(new_n16500_), .A2(new_n16100_), .ZN(new_n17191_));
  NOR3_X1    g16189(.A1(new_n16500_), .A2(new_n16100_), .A3(new_n16489_), .ZN(new_n17192_));
  OAI22_X1   g16190(.A1(new_n17192_), .A2(new_n16492_), .B1(new_n17191_), .B2(new_n16494_), .ZN(new_n17193_));
  INV_X1     g16191(.I(new_n17193_), .ZN(new_n17194_));
  NAND2_X1   g16192(.A1(new_n16482_), .A2(new_n16129_), .ZN(new_n17195_));
  NAND2_X1   g16193(.A1(new_n17195_), .A2(new_n16478_), .ZN(new_n17196_));
  NAND3_X1   g16194(.A1(new_n16482_), .A2(new_n16129_), .A3(new_n16475_), .ZN(new_n17197_));
  NAND2_X1   g16195(.A1(new_n17197_), .A2(new_n16476_), .ZN(new_n17198_));
  NAND2_X1   g16196(.A1(new_n17198_), .A2(new_n17196_), .ZN(new_n17199_));
  NOR2_X1    g16197(.A1(new_n17199_), .A2(new_n17194_), .ZN(new_n17200_));
  AOI22_X1   g16198(.A1(new_n17197_), .A2(new_n16476_), .B1(new_n17195_), .B2(new_n16478_), .ZN(new_n17201_));
  NOR2_X1    g16199(.A1(new_n17201_), .A2(new_n17193_), .ZN(new_n17202_));
  NOR2_X1    g16200(.A1(new_n17200_), .A2(new_n17202_), .ZN(new_n17203_));
  NOR2_X1    g16201(.A1(new_n16488_), .A2(new_n16513_), .ZN(new_n17204_));
  NOR2_X1    g16202(.A1(new_n17204_), .A2(new_n16516_), .ZN(new_n17205_));
  NAND2_X1   g16203(.A1(new_n16510_), .A2(new_n16506_), .ZN(new_n17206_));
  NOR4_X1    g16204(.A1(new_n16487_), .A2(new_n16483_), .A3(new_n16511_), .A4(new_n16512_), .ZN(new_n17207_));
  AOI21_X1   g16205(.A1(new_n16474_), .A2(new_n17206_), .B(new_n17207_), .ZN(new_n17208_));
  NAND2_X1   g16206(.A1(new_n17201_), .A2(new_n17193_), .ZN(new_n17209_));
  NAND2_X1   g16207(.A1(new_n17199_), .A2(new_n17194_), .ZN(new_n17210_));
  NAND4_X1   g16208(.A1(new_n16508_), .A2(new_n16509_), .A3(new_n16505_), .A4(new_n16501_), .ZN(new_n17211_));
  NAND3_X1   g16209(.A1(new_n17210_), .A2(new_n17209_), .A3(new_n17211_), .ZN(new_n17212_));
  OAI22_X1   g16210(.A1(new_n17212_), .A2(new_n17205_), .B1(new_n17203_), .B2(new_n17208_), .ZN(new_n17213_));
  OAI21_X1   g16211(.A1(new_n16457_), .A2(new_n16012_), .B(new_n16450_), .ZN(new_n17214_));
  OAI21_X1   g16212(.A1(new_n16010_), .A2(new_n16011_), .B(new_n16446_), .ZN(new_n17215_));
  OAI21_X1   g16213(.A1(new_n16457_), .A2(new_n17215_), .B(new_n16447_), .ZN(new_n17216_));
  NAND2_X1   g16214(.A1(new_n17216_), .A2(new_n17214_), .ZN(new_n17217_));
  NAND2_X1   g16215(.A1(new_n16443_), .A2(new_n15946_), .ZN(new_n17218_));
  NAND3_X1   g16216(.A1(new_n16443_), .A2(new_n15946_), .A3(new_n16436_), .ZN(new_n17219_));
  AOI22_X1   g16217(.A1(new_n17219_), .A2(new_n16437_), .B1(new_n17218_), .B2(new_n16432_), .ZN(new_n17220_));
  NAND2_X1   g16218(.A1(new_n17220_), .A2(new_n17217_), .ZN(new_n17221_));
  AND2_X2    g16219(.A1(new_n17216_), .A2(new_n17214_), .Z(new_n17222_));
  OAI21_X1   g16220(.A1(new_n16439_), .A2(new_n16149_), .B(new_n16432_), .ZN(new_n17223_));
  NAND2_X1   g16221(.A1(new_n15946_), .A2(new_n16436_), .ZN(new_n17224_));
  OAI21_X1   g16222(.A1(new_n17224_), .A2(new_n16439_), .B(new_n16437_), .ZN(new_n17225_));
  NAND2_X1   g16223(.A1(new_n17225_), .A2(new_n17223_), .ZN(new_n17226_));
  NAND2_X1   g16224(.A1(new_n17222_), .A2(new_n17226_), .ZN(new_n17227_));
  NAND2_X1   g16225(.A1(new_n17227_), .A2(new_n17221_), .ZN(new_n17228_));
  OAI22_X1   g16226(.A1(new_n16461_), .A2(new_n16462_), .B1(new_n16454_), .B2(new_n16458_), .ZN(new_n17229_));
  NAND2_X1   g16227(.A1(new_n16469_), .A2(new_n17229_), .ZN(new_n17230_));
  NOR2_X1    g16228(.A1(new_n16463_), .A2(new_n16459_), .ZN(new_n17231_));
  NAND4_X1   g16229(.A1(new_n16440_), .A2(new_n16444_), .A3(new_n16465_), .A4(new_n16464_), .ZN(new_n17232_));
  OAI21_X1   g16230(.A1(new_n17231_), .A2(new_n16431_), .B(new_n17232_), .ZN(new_n17233_));
  NOR2_X1    g16231(.A1(new_n17222_), .A2(new_n17226_), .ZN(new_n17234_));
  NOR2_X1    g16232(.A1(new_n17220_), .A2(new_n17217_), .ZN(new_n17235_));
  NOR4_X1    g16233(.A1(new_n16461_), .A2(new_n16454_), .A3(new_n16462_), .A4(new_n16458_), .ZN(new_n17236_));
  NOR3_X1    g16234(.A1(new_n17234_), .A2(new_n17235_), .A3(new_n17236_), .ZN(new_n17237_));
  AOI22_X1   g16235(.A1(new_n17237_), .A2(new_n17230_), .B1(new_n17228_), .B2(new_n17233_), .ZN(new_n17238_));
  NAND2_X1   g16236(.A1(new_n17213_), .A2(new_n17238_), .ZN(new_n17239_));
  NAND2_X1   g16237(.A1(new_n17210_), .A2(new_n17209_), .ZN(new_n17240_));
  NAND2_X1   g16238(.A1(new_n16474_), .A2(new_n17206_), .ZN(new_n17241_));
  OAI21_X1   g16239(.A1(new_n17204_), .A2(new_n16516_), .B(new_n17211_), .ZN(new_n17242_));
  NOR3_X1    g16240(.A1(new_n17200_), .A2(new_n17202_), .A3(new_n17207_), .ZN(new_n17243_));
  AOI22_X1   g16241(.A1(new_n17243_), .A2(new_n17241_), .B1(new_n17240_), .B2(new_n17242_), .ZN(new_n17244_));
  NOR2_X1    g16242(.A1(new_n17234_), .A2(new_n17235_), .ZN(new_n17245_));
  NOR2_X1    g16243(.A1(new_n17231_), .A2(new_n16431_), .ZN(new_n17246_));
  AOI21_X1   g16244(.A1(new_n16469_), .A2(new_n17229_), .B(new_n17236_), .ZN(new_n17247_));
  NAND3_X1   g16245(.A1(new_n17227_), .A2(new_n17221_), .A3(new_n17232_), .ZN(new_n17248_));
  OAI22_X1   g16246(.A1(new_n17248_), .A2(new_n17246_), .B1(new_n17245_), .B2(new_n17247_), .ZN(new_n17249_));
  NAND2_X1   g16247(.A1(new_n17244_), .A2(new_n17249_), .ZN(new_n17250_));
  AOI22_X1   g16248(.A1(new_n17189_), .A2(new_n17190_), .B1(new_n17239_), .B2(new_n17250_), .ZN(new_n17251_));
  NOR2_X1    g16249(.A1(new_n16524_), .A2(new_n16520_), .ZN(new_n17252_));
  AOI21_X1   g16250(.A1(new_n16524_), .A2(new_n16520_), .B(new_n16530_), .ZN(new_n17253_));
  NOR2_X1    g16251(.A1(new_n17244_), .A2(new_n17249_), .ZN(new_n17254_));
  NOR2_X1    g16252(.A1(new_n17213_), .A2(new_n17238_), .ZN(new_n17255_));
  NOR4_X1    g16253(.A1(new_n17253_), .A2(new_n17255_), .A3(new_n17254_), .A4(new_n17252_), .ZN(new_n17256_));
  NOR2_X1    g16254(.A1(new_n17251_), .A2(new_n17256_), .ZN(new_n17257_));
  NAND2_X1   g16255(.A1(new_n17257_), .A2(new_n17188_), .ZN(new_n17258_));
  NAND2_X1   g16256(.A1(new_n16647_), .A2(new_n16643_), .ZN(new_n17259_));
  INV_X1     g16257(.I(new_n17124_), .ZN(new_n17260_));
  AOI22_X1   g16258(.A1(new_n17260_), .A2(new_n17259_), .B1(new_n17186_), .B2(new_n17185_), .ZN(new_n17261_));
  NOR4_X1    g16259(.A1(new_n17171_), .A2(new_n17182_), .A3(new_n17123_), .A4(new_n17124_), .ZN(new_n17262_));
  NOR2_X1    g16260(.A1(new_n17261_), .A2(new_n17262_), .ZN(new_n17263_));
  OAI22_X1   g16261(.A1(new_n17254_), .A2(new_n17255_), .B1(new_n17253_), .B2(new_n17252_), .ZN(new_n17264_));
  NAND4_X1   g16262(.A1(new_n17190_), .A2(new_n17239_), .A3(new_n17250_), .A4(new_n17189_), .ZN(new_n17265_));
  NAND2_X1   g16263(.A1(new_n17264_), .A2(new_n17265_), .ZN(new_n17266_));
  NAND2_X1   g16264(.A1(new_n17263_), .A2(new_n17266_), .ZN(new_n17267_));
  AOI22_X1   g16265(.A1(new_n17258_), .A2(new_n17267_), .B1(new_n17121_), .B2(new_n17122_), .ZN(new_n17268_));
  NOR2_X1    g16266(.A1(new_n16534_), .A2(new_n16664_), .ZN(new_n17269_));
  AOI21_X1   g16267(.A1(new_n16534_), .A2(new_n16664_), .B(new_n16428_), .ZN(new_n17270_));
  NOR2_X1    g16268(.A1(new_n17263_), .A2(new_n17266_), .ZN(new_n17271_));
  NOR2_X1    g16269(.A1(new_n17257_), .A2(new_n17188_), .ZN(new_n17272_));
  NOR4_X1    g16270(.A1(new_n17272_), .A2(new_n17271_), .A3(new_n17269_), .A4(new_n17270_), .ZN(new_n17273_));
  NOR2_X1    g16271(.A1(new_n17268_), .A2(new_n17273_), .ZN(new_n17274_));
  NAND2_X1   g16272(.A1(new_n17274_), .A2(new_n17120_), .ZN(new_n17275_));
  AOI22_X1   g16273(.A1(new_n17117_), .A2(new_n17118_), .B1(new_n17116_), .B2(new_n17115_), .ZN(new_n17276_));
  NAND2_X1   g16274(.A1(new_n17116_), .A2(new_n17115_), .ZN(new_n17277_));
  NOR3_X1    g16275(.A1(new_n17277_), .A2(new_n17102_), .A3(new_n17113_), .ZN(new_n17278_));
  NOR2_X1    g16276(.A1(new_n17278_), .A2(new_n17276_), .ZN(new_n17279_));
  OAI22_X1   g16277(.A1(new_n17272_), .A2(new_n17271_), .B1(new_n17270_), .B2(new_n17269_), .ZN(new_n17280_));
  NAND4_X1   g16278(.A1(new_n17258_), .A2(new_n17267_), .A3(new_n17121_), .A4(new_n17122_), .ZN(new_n17281_));
  NAND2_X1   g16279(.A1(new_n17280_), .A2(new_n17281_), .ZN(new_n17282_));
  NAND2_X1   g16280(.A1(new_n17279_), .A2(new_n17282_), .ZN(new_n17283_));
  AOI21_X1   g16281(.A1(new_n17283_), .A2(new_n17275_), .B(new_n16965_), .ZN(new_n17284_));
  NAND2_X1   g16282(.A1(new_n16672_), .A2(new_n16931_), .ZN(new_n17285_));
  OAI21_X1   g16283(.A1(new_n16672_), .A2(new_n16931_), .B(new_n16426_), .ZN(new_n17286_));
  NAND2_X1   g16284(.A1(new_n17286_), .A2(new_n17285_), .ZN(new_n17287_));
  NOR2_X1    g16285(.A1(new_n17279_), .A2(new_n17282_), .ZN(new_n17288_));
  NOR2_X1    g16286(.A1(new_n17274_), .A2(new_n17120_), .ZN(new_n17289_));
  NOR3_X1    g16287(.A1(new_n17287_), .A2(new_n17288_), .A3(new_n17289_), .ZN(new_n17290_));
  NOR2_X1    g16288(.A1(new_n17290_), .A2(new_n17284_), .ZN(new_n17291_));
  NOR2_X1    g16289(.A1(new_n14417_), .A2(new_n14413_), .ZN(new_n17292_));
  AOI21_X1   g16290(.A1(new_n14417_), .A2(new_n14413_), .B(new_n14428_), .ZN(new_n17293_));
  NAND2_X1   g16291(.A1(new_n14286_), .A2(new_n14405_), .ZN(new_n17294_));
  OAI21_X1   g16292(.A1(new_n14286_), .A2(new_n14405_), .B(new_n14173_), .ZN(new_n17295_));
  NOR2_X1    g16293(.A1(new_n14388_), .A2(new_n14384_), .ZN(new_n17296_));
  AOI21_X1   g16294(.A1(new_n14388_), .A2(new_n14384_), .B(new_n14394_), .ZN(new_n17297_));
  AOI21_X1   g16295(.A1(new_n13372_), .A2(new_n14368_), .B(new_n14360_), .ZN(new_n17298_));
  NOR2_X1    g16296(.A1(new_n13353_), .A2(new_n14356_), .ZN(new_n17299_));
  AOI21_X1   g16297(.A1(new_n17299_), .A2(new_n14368_), .B(new_n14358_), .ZN(new_n17300_));
  NOR2_X1    g16298(.A1(new_n17300_), .A2(new_n17298_), .ZN(new_n17301_));
  INV_X1     g16299(.I(new_n17301_), .ZN(new_n17302_));
  NAND2_X1   g16300(.A1(new_n14349_), .A2(new_n13385_), .ZN(new_n17303_));
  NAND3_X1   g16301(.A1(new_n14349_), .A2(new_n13385_), .A3(new_n14338_), .ZN(new_n17304_));
  AOI22_X1   g16302(.A1(new_n17304_), .A2(new_n14341_), .B1(new_n17303_), .B2(new_n14343_), .ZN(new_n17305_));
  NAND2_X1   g16303(.A1(new_n17302_), .A2(new_n17305_), .ZN(new_n17306_));
  OAI21_X1   g16304(.A1(new_n14353_), .A2(new_n13301_), .B(new_n14343_), .ZN(new_n17307_));
  NAND2_X1   g16305(.A1(new_n17304_), .A2(new_n14341_), .ZN(new_n17308_));
  NAND2_X1   g16306(.A1(new_n17308_), .A2(new_n17307_), .ZN(new_n17309_));
  NAND2_X1   g16307(.A1(new_n17309_), .A2(new_n17301_), .ZN(new_n17310_));
  NAND2_X1   g16308(.A1(new_n17310_), .A2(new_n17306_), .ZN(new_n17311_));
  NAND2_X1   g16309(.A1(new_n14374_), .A2(new_n14370_), .ZN(new_n17312_));
  NAND2_X1   g16310(.A1(new_n17312_), .A2(new_n14337_), .ZN(new_n17313_));
  NOR2_X1    g16311(.A1(new_n14355_), .A2(new_n14377_), .ZN(new_n17314_));
  NAND4_X1   g16312(.A1(new_n14372_), .A2(new_n14373_), .A3(new_n14369_), .A4(new_n14365_), .ZN(new_n17315_));
  OAI21_X1   g16313(.A1(new_n17314_), .A2(new_n14380_), .B(new_n17315_), .ZN(new_n17316_));
  NOR2_X1    g16314(.A1(new_n17309_), .A2(new_n17301_), .ZN(new_n17317_));
  NOR2_X1    g16315(.A1(new_n17302_), .A2(new_n17305_), .ZN(new_n17318_));
  NOR4_X1    g16316(.A1(new_n14354_), .A2(new_n14350_), .A3(new_n14375_), .A4(new_n14376_), .ZN(new_n17319_));
  NOR3_X1    g16317(.A1(new_n17317_), .A2(new_n17318_), .A3(new_n17319_), .ZN(new_n17320_));
  AOI22_X1   g16318(.A1(new_n17320_), .A2(new_n17313_), .B1(new_n17311_), .B2(new_n17316_), .ZN(new_n17321_));
  OAI21_X1   g16319(.A1(new_n14319_), .A2(new_n13244_), .B(new_n14311_), .ZN(new_n17322_));
  OAI21_X1   g16320(.A1(new_n13242_), .A2(new_n13243_), .B(new_n14306_), .ZN(new_n17323_));
  OAI21_X1   g16321(.A1(new_n17323_), .A2(new_n14319_), .B(new_n14308_), .ZN(new_n17324_));
  NAND2_X1   g16322(.A1(new_n17324_), .A2(new_n17322_), .ZN(new_n17325_));
  INV_X1     g16323(.I(new_n17325_), .ZN(new_n17326_));
  OAI21_X1   g16324(.A1(new_n14299_), .A2(new_n13261_), .B(new_n14291_), .ZN(new_n17327_));
  AOI21_X1   g16325(.A1(new_n13182_), .A2(new_n13188_), .B(new_n14291_), .ZN(new_n17328_));
  INV_X1     g16326(.I(new_n17328_), .ZN(new_n17329_));
  OAI21_X1   g16327(.A1(new_n17329_), .A2(new_n14299_), .B(new_n14297_), .ZN(new_n17330_));
  NAND2_X1   g16328(.A1(new_n17330_), .A2(new_n17327_), .ZN(new_n17331_));
  NOR2_X1    g16329(.A1(new_n17326_), .A2(new_n17331_), .ZN(new_n17332_));
  NAND2_X1   g16330(.A1(new_n14303_), .A2(new_n13189_), .ZN(new_n17333_));
  NAND2_X1   g16331(.A1(new_n17328_), .A2(new_n14303_), .ZN(new_n17334_));
  AOI22_X1   g16332(.A1(new_n17334_), .A2(new_n14297_), .B1(new_n17333_), .B2(new_n14291_), .ZN(new_n17335_));
  NOR2_X1    g16333(.A1(new_n17335_), .A2(new_n17325_), .ZN(new_n17336_));
  NOR2_X1    g16334(.A1(new_n17332_), .A2(new_n17336_), .ZN(new_n17337_));
  NOR2_X1    g16335(.A1(new_n14325_), .A2(new_n14321_), .ZN(new_n17338_));
  NOR2_X1    g16336(.A1(new_n17338_), .A2(new_n14290_), .ZN(new_n17339_));
  NAND2_X1   g16337(.A1(new_n14305_), .A2(new_n14328_), .ZN(new_n17340_));
  NAND4_X1   g16338(.A1(new_n14300_), .A2(new_n14326_), .A3(new_n14327_), .A4(new_n14304_), .ZN(new_n17341_));
  INV_X1     g16339(.I(new_n17341_), .ZN(new_n17342_));
  AOI21_X1   g16340(.A1(new_n14332_), .A2(new_n17340_), .B(new_n17342_), .ZN(new_n17343_));
  NAND2_X1   g16341(.A1(new_n17335_), .A2(new_n17325_), .ZN(new_n17344_));
  NAND2_X1   g16342(.A1(new_n17326_), .A2(new_n17331_), .ZN(new_n17345_));
  NAND3_X1   g16343(.A1(new_n17345_), .A2(new_n17344_), .A3(new_n17341_), .ZN(new_n17346_));
  OAI22_X1   g16344(.A1(new_n17337_), .A2(new_n17343_), .B1(new_n17346_), .B2(new_n17339_), .ZN(new_n17347_));
  NOR2_X1    g16345(.A1(new_n17347_), .A2(new_n17321_), .ZN(new_n17348_));
  NOR2_X1    g16346(.A1(new_n17317_), .A2(new_n17318_), .ZN(new_n17349_));
  NOR2_X1    g16347(.A1(new_n17314_), .A2(new_n14380_), .ZN(new_n17350_));
  AOI21_X1   g16348(.A1(new_n17312_), .A2(new_n14337_), .B(new_n17319_), .ZN(new_n17351_));
  NAND3_X1   g16349(.A1(new_n17310_), .A2(new_n17306_), .A3(new_n17315_), .ZN(new_n17352_));
  OAI22_X1   g16350(.A1(new_n17350_), .A2(new_n17352_), .B1(new_n17349_), .B2(new_n17351_), .ZN(new_n17353_));
  NAND2_X1   g16351(.A1(new_n17345_), .A2(new_n17344_), .ZN(new_n17354_));
  NAND2_X1   g16352(.A1(new_n14332_), .A2(new_n17340_), .ZN(new_n17355_));
  OAI21_X1   g16353(.A1(new_n17338_), .A2(new_n14290_), .B(new_n17341_), .ZN(new_n17356_));
  NOR3_X1    g16354(.A1(new_n17332_), .A2(new_n17342_), .A3(new_n17336_), .ZN(new_n17357_));
  AOI22_X1   g16355(.A1(new_n17357_), .A2(new_n17355_), .B1(new_n17354_), .B2(new_n17356_), .ZN(new_n17358_));
  NOR2_X1    g16356(.A1(new_n17358_), .A2(new_n17353_), .ZN(new_n17359_));
  OAI22_X1   g16357(.A1(new_n17348_), .A2(new_n17359_), .B1(new_n17297_), .B2(new_n17296_), .ZN(new_n17360_));
  NAND2_X1   g16358(.A1(new_n14336_), .A2(new_n14391_), .ZN(new_n17361_));
  OAI21_X1   g16359(.A1(new_n14336_), .A2(new_n14391_), .B(new_n14288_), .ZN(new_n17362_));
  NAND2_X1   g16360(.A1(new_n17358_), .A2(new_n17353_), .ZN(new_n17363_));
  NAND2_X1   g16361(.A1(new_n17347_), .A2(new_n17321_), .ZN(new_n17364_));
  NAND4_X1   g16362(.A1(new_n17362_), .A2(new_n17363_), .A3(new_n17364_), .A4(new_n17361_), .ZN(new_n17365_));
  NAND2_X1   g16363(.A1(new_n17365_), .A2(new_n17360_), .ZN(new_n17366_));
  NAND2_X1   g16364(.A1(new_n14275_), .A2(new_n14271_), .ZN(new_n17367_));
  OAI21_X1   g16365(.A1(new_n14275_), .A2(new_n14271_), .B(new_n14282_), .ZN(new_n17368_));
  NAND2_X1   g16366(.A1(new_n14251_), .A2(new_n13116_), .ZN(new_n17369_));
  NAND3_X1   g16367(.A1(new_n14251_), .A2(new_n13116_), .A3(new_n14240_), .ZN(new_n17370_));
  AOI22_X1   g16368(.A1(new_n17370_), .A2(new_n14244_), .B1(new_n17369_), .B2(new_n14246_), .ZN(new_n17371_));
  AOI21_X1   g16369(.A1(new_n13125_), .A2(new_n14232_), .B(new_n14227_), .ZN(new_n17372_));
  NAND3_X1   g16370(.A1(new_n13125_), .A2(new_n14232_), .A3(new_n14227_), .ZN(new_n17373_));
  AOI21_X1   g16371(.A1(new_n17373_), .A2(new_n14230_), .B(new_n17372_), .ZN(new_n17374_));
  INV_X1     g16372(.I(new_n17374_), .ZN(new_n17375_));
  NOR2_X1    g16373(.A1(new_n17375_), .A2(new_n17371_), .ZN(new_n17376_));
  OAI21_X1   g16374(.A1(new_n13098_), .A2(new_n14255_), .B(new_n14246_), .ZN(new_n17377_));
  NAND2_X1   g16375(.A1(new_n13116_), .A2(new_n14240_), .ZN(new_n17378_));
  OAI21_X1   g16376(.A1(new_n17378_), .A2(new_n14255_), .B(new_n14244_), .ZN(new_n17379_));
  NAND2_X1   g16377(.A1(new_n17379_), .A2(new_n17377_), .ZN(new_n17380_));
  NOR2_X1    g16378(.A1(new_n17380_), .A2(new_n17374_), .ZN(new_n17381_));
  NOR2_X1    g16379(.A1(new_n17376_), .A2(new_n17381_), .ZN(new_n17382_));
  NOR2_X1    g16380(.A1(new_n14261_), .A2(new_n14257_), .ZN(new_n17383_));
  NOR2_X1    g16381(.A1(new_n17383_), .A2(new_n14219_), .ZN(new_n17384_));
  NAND2_X1   g16382(.A1(new_n14238_), .A2(new_n14264_), .ZN(new_n17385_));
  NOR4_X1    g16383(.A1(new_n14260_), .A2(new_n14259_), .A3(new_n14252_), .A4(new_n14256_), .ZN(new_n17386_));
  AOI21_X1   g16384(.A1(new_n17385_), .A2(new_n14267_), .B(new_n17386_), .ZN(new_n17387_));
  NAND2_X1   g16385(.A1(new_n17380_), .A2(new_n17374_), .ZN(new_n17388_));
  NAND2_X1   g16386(.A1(new_n17375_), .A2(new_n17371_), .ZN(new_n17389_));
  NAND4_X1   g16387(.A1(new_n14234_), .A2(new_n14262_), .A3(new_n14263_), .A4(new_n14237_), .ZN(new_n17390_));
  NAND3_X1   g16388(.A1(new_n17389_), .A2(new_n17388_), .A3(new_n17390_), .ZN(new_n17391_));
  OAI22_X1   g16389(.A1(new_n17384_), .A2(new_n17391_), .B1(new_n17382_), .B2(new_n17387_), .ZN(new_n17392_));
  NOR2_X1    g16390(.A1(new_n14198_), .A2(new_n12979_), .ZN(new_n17393_));
  NOR3_X1    g16391(.A1(new_n14198_), .A2(new_n12979_), .A3(new_n14190_), .ZN(new_n17394_));
  OAI22_X1   g16392(.A1(new_n17394_), .A2(new_n14192_), .B1(new_n17393_), .B2(new_n14194_), .ZN(new_n17395_));
  NAND2_X1   g16393(.A1(new_n14182_), .A2(new_n12939_), .ZN(new_n17396_));
  AOI21_X1   g16394(.A1(new_n12932_), .A2(new_n12938_), .B(new_n14179_), .ZN(new_n17397_));
  NAND2_X1   g16395(.A1(new_n17397_), .A2(new_n14182_), .ZN(new_n17398_));
  AOI22_X1   g16396(.A1(new_n17398_), .A2(new_n14177_), .B1(new_n17396_), .B2(new_n14179_), .ZN(new_n17399_));
  NAND2_X1   g16397(.A1(new_n17399_), .A2(new_n17395_), .ZN(new_n17400_));
  INV_X1     g16398(.I(new_n17395_), .ZN(new_n17401_));
  OAI21_X1   g16399(.A1(new_n14186_), .A2(new_n13006_), .B(new_n14179_), .ZN(new_n17402_));
  NAND2_X1   g16400(.A1(new_n12939_), .A2(new_n14176_), .ZN(new_n17403_));
  OAI21_X1   g16401(.A1(new_n17403_), .A2(new_n14186_), .B(new_n14177_), .ZN(new_n17404_));
  NAND2_X1   g16402(.A1(new_n17404_), .A2(new_n17402_), .ZN(new_n17405_));
  NAND2_X1   g16403(.A1(new_n17401_), .A2(new_n17405_), .ZN(new_n17406_));
  NAND2_X1   g16404(.A1(new_n17406_), .A2(new_n17400_), .ZN(new_n17407_));
  OAI22_X1   g16405(.A1(new_n14183_), .A2(new_n14187_), .B1(new_n14209_), .B2(new_n14210_), .ZN(new_n17408_));
  NAND2_X1   g16406(.A1(new_n14175_), .A2(new_n17408_), .ZN(new_n17409_));
  AOI22_X1   g16407(.A1(new_n14206_), .A2(new_n14207_), .B1(new_n14199_), .B2(new_n14203_), .ZN(new_n17410_));
  NAND4_X1   g16408(.A1(new_n14206_), .A2(new_n14207_), .A3(new_n14199_), .A4(new_n14203_), .ZN(new_n17411_));
  OAI21_X1   g16409(.A1(new_n14214_), .A2(new_n17410_), .B(new_n17411_), .ZN(new_n17412_));
  NOR2_X1    g16410(.A1(new_n17401_), .A2(new_n17405_), .ZN(new_n17413_));
  NOR2_X1    g16411(.A1(new_n17399_), .A2(new_n17395_), .ZN(new_n17414_));
  NOR4_X1    g16412(.A1(new_n14183_), .A2(new_n14187_), .A3(new_n14209_), .A4(new_n14210_), .ZN(new_n17415_));
  NOR3_X1    g16413(.A1(new_n17413_), .A2(new_n17414_), .A3(new_n17415_), .ZN(new_n17416_));
  AOI22_X1   g16414(.A1(new_n17416_), .A2(new_n17409_), .B1(new_n17407_), .B2(new_n17412_), .ZN(new_n17417_));
  NAND2_X1   g16415(.A1(new_n17392_), .A2(new_n17417_), .ZN(new_n17418_));
  NAND2_X1   g16416(.A1(new_n17389_), .A2(new_n17388_), .ZN(new_n17419_));
  NAND2_X1   g16417(.A1(new_n17385_), .A2(new_n14267_), .ZN(new_n17420_));
  OAI21_X1   g16418(.A1(new_n17383_), .A2(new_n14219_), .B(new_n17390_), .ZN(new_n17421_));
  NOR3_X1    g16419(.A1(new_n17376_), .A2(new_n17381_), .A3(new_n17386_), .ZN(new_n17422_));
  AOI22_X1   g16420(.A1(new_n17422_), .A2(new_n17420_), .B1(new_n17419_), .B2(new_n17421_), .ZN(new_n17423_));
  NOR2_X1    g16421(.A1(new_n17413_), .A2(new_n17414_), .ZN(new_n17424_));
  NOR2_X1    g16422(.A1(new_n14214_), .A2(new_n17410_), .ZN(new_n17425_));
  AOI21_X1   g16423(.A1(new_n14175_), .A2(new_n17408_), .B(new_n17415_), .ZN(new_n17426_));
  NAND3_X1   g16424(.A1(new_n17406_), .A2(new_n17400_), .A3(new_n17411_), .ZN(new_n17427_));
  OAI22_X1   g16425(.A1(new_n17427_), .A2(new_n17425_), .B1(new_n17424_), .B2(new_n17426_), .ZN(new_n17428_));
  NAND2_X1   g16426(.A1(new_n17428_), .A2(new_n17423_), .ZN(new_n17429_));
  AOI22_X1   g16427(.A1(new_n17418_), .A2(new_n17429_), .B1(new_n17368_), .B2(new_n17367_), .ZN(new_n17430_));
  NOR2_X1    g16428(.A1(new_n14218_), .A2(new_n14278_), .ZN(new_n17431_));
  AOI21_X1   g16429(.A1(new_n14218_), .A2(new_n14278_), .B(new_n14174_), .ZN(new_n17432_));
  NOR2_X1    g16430(.A1(new_n17428_), .A2(new_n17423_), .ZN(new_n17433_));
  NOR2_X1    g16431(.A1(new_n17392_), .A2(new_n17417_), .ZN(new_n17434_));
  NOR4_X1    g16432(.A1(new_n17433_), .A2(new_n17434_), .A3(new_n17432_), .A4(new_n17431_), .ZN(new_n17435_));
  NOR2_X1    g16433(.A1(new_n17435_), .A2(new_n17430_), .ZN(new_n17436_));
  NAND2_X1   g16434(.A1(new_n17366_), .A2(new_n17436_), .ZN(new_n17437_));
  AOI22_X1   g16435(.A1(new_n17362_), .A2(new_n17361_), .B1(new_n17363_), .B2(new_n17364_), .ZN(new_n17438_));
  NOR4_X1    g16436(.A1(new_n17297_), .A2(new_n17348_), .A3(new_n17359_), .A4(new_n17296_), .ZN(new_n17439_));
  NOR2_X1    g16437(.A1(new_n17438_), .A2(new_n17439_), .ZN(new_n17440_));
  OAI22_X1   g16438(.A1(new_n17433_), .A2(new_n17434_), .B1(new_n17432_), .B2(new_n17431_), .ZN(new_n17441_));
  NAND4_X1   g16439(.A1(new_n17418_), .A2(new_n17429_), .A3(new_n17368_), .A4(new_n17367_), .ZN(new_n17442_));
  NAND2_X1   g16440(.A1(new_n17441_), .A2(new_n17442_), .ZN(new_n17443_));
  NAND2_X1   g16441(.A1(new_n17440_), .A2(new_n17443_), .ZN(new_n17444_));
  AOI22_X1   g16442(.A1(new_n17437_), .A2(new_n17444_), .B1(new_n17294_), .B2(new_n17295_), .ZN(new_n17445_));
  NOR2_X1    g16443(.A1(new_n14402_), .A2(new_n14398_), .ZN(new_n17446_));
  AOI21_X1   g16444(.A1(new_n14402_), .A2(new_n14398_), .B(new_n14409_), .ZN(new_n17447_));
  NOR2_X1    g16445(.A1(new_n17440_), .A2(new_n17443_), .ZN(new_n17448_));
  NOR2_X1    g16446(.A1(new_n17366_), .A2(new_n17436_), .ZN(new_n17449_));
  NOR4_X1    g16447(.A1(new_n17449_), .A2(new_n17448_), .A3(new_n17446_), .A4(new_n17447_), .ZN(new_n17450_));
  NOR2_X1    g16448(.A1(new_n17445_), .A2(new_n17450_), .ZN(new_n17451_));
  NOR2_X1    g16449(.A1(new_n14047_), .A2(new_n14164_), .ZN(new_n17452_));
  AOI21_X1   g16450(.A1(new_n14047_), .A2(new_n14164_), .B(new_n13938_), .ZN(new_n17453_));
  NAND2_X1   g16451(.A1(new_n14146_), .A2(new_n14142_), .ZN(new_n17454_));
  OAI21_X1   g16452(.A1(new_n14146_), .A2(new_n14142_), .B(new_n14153_), .ZN(new_n17455_));
  NAND2_X1   g16453(.A1(new_n14122_), .A2(new_n13871_), .ZN(new_n17456_));
  NAND3_X1   g16454(.A1(new_n14122_), .A2(new_n13871_), .A3(new_n14111_), .ZN(new_n17457_));
  AOI22_X1   g16455(.A1(new_n17457_), .A2(new_n14115_), .B1(new_n17456_), .B2(new_n14117_), .ZN(new_n17458_));
  AOI21_X1   g16456(.A1(new_n14107_), .A2(new_n13880_), .B(new_n14098_), .ZN(new_n17459_));
  INV_X1     g16457(.I(new_n17459_), .ZN(new_n17460_));
  NAND3_X1   g16458(.A1(new_n14107_), .A2(new_n13880_), .A3(new_n14098_), .ZN(new_n17461_));
  NAND2_X1   g16459(.A1(new_n17461_), .A2(new_n14101_), .ZN(new_n17462_));
  NAND2_X1   g16460(.A1(new_n17462_), .A2(new_n17460_), .ZN(new_n17463_));
  NOR2_X1    g16461(.A1(new_n17463_), .A2(new_n17458_), .ZN(new_n17464_));
  OAI21_X1   g16462(.A1(new_n13851_), .A2(new_n14126_), .B(new_n14117_), .ZN(new_n17465_));
  NAND2_X1   g16463(.A1(new_n13871_), .A2(new_n14111_), .ZN(new_n17466_));
  OAI21_X1   g16464(.A1(new_n17466_), .A2(new_n14126_), .B(new_n14115_), .ZN(new_n17467_));
  NAND2_X1   g16465(.A1(new_n17467_), .A2(new_n17465_), .ZN(new_n17468_));
  AOI21_X1   g16466(.A1(new_n17461_), .A2(new_n14101_), .B(new_n17459_), .ZN(new_n17469_));
  NOR2_X1    g16467(.A1(new_n17468_), .A2(new_n17469_), .ZN(new_n17470_));
  NOR2_X1    g16468(.A1(new_n17464_), .A2(new_n17470_), .ZN(new_n17471_));
  NAND2_X1   g16469(.A1(new_n14109_), .A2(new_n14135_), .ZN(new_n17472_));
  NAND2_X1   g16470(.A1(new_n17472_), .A2(new_n14138_), .ZN(new_n17473_));
  INV_X1     g16471(.I(new_n17473_), .ZN(new_n17474_));
  NOR4_X1    g16472(.A1(new_n14131_), .A2(new_n14130_), .A3(new_n14123_), .A4(new_n14127_), .ZN(new_n17475_));
  AOI21_X1   g16473(.A1(new_n17472_), .A2(new_n14138_), .B(new_n17475_), .ZN(new_n17476_));
  NAND2_X1   g16474(.A1(new_n17468_), .A2(new_n17469_), .ZN(new_n17477_));
  NAND2_X1   g16475(.A1(new_n17463_), .A2(new_n17458_), .ZN(new_n17478_));
  NAND4_X1   g16476(.A1(new_n14104_), .A2(new_n14133_), .A3(new_n14108_), .A4(new_n14134_), .ZN(new_n17479_));
  NAND3_X1   g16477(.A1(new_n17478_), .A2(new_n17477_), .A3(new_n17479_), .ZN(new_n17480_));
  OAI22_X1   g16478(.A1(new_n17474_), .A2(new_n17480_), .B1(new_n17471_), .B2(new_n17476_), .ZN(new_n17481_));
  OAI21_X1   g16479(.A1(new_n14071_), .A2(new_n13761_), .B(new_n14065_), .ZN(new_n17482_));
  OAI21_X1   g16480(.A1(new_n13759_), .A2(new_n13760_), .B(new_n14068_), .ZN(new_n17483_));
  OAI21_X1   g16481(.A1(new_n14071_), .A2(new_n17483_), .B(new_n14069_), .ZN(new_n17484_));
  NAND2_X1   g16482(.A1(new_n17484_), .A2(new_n17482_), .ZN(new_n17485_));
  NAND2_X1   g16483(.A1(new_n14057_), .A2(new_n13698_), .ZN(new_n17486_));
  NAND3_X1   g16484(.A1(new_n14057_), .A2(new_n13698_), .A3(new_n14051_), .ZN(new_n17487_));
  AOI22_X1   g16485(.A1(new_n17487_), .A2(new_n14052_), .B1(new_n17486_), .B2(new_n14054_), .ZN(new_n17488_));
  NAND2_X1   g16486(.A1(new_n17488_), .A2(new_n17485_), .ZN(new_n17489_));
  AND2_X2    g16487(.A1(new_n17484_), .A2(new_n17482_), .Z(new_n17490_));
  NOR2_X1    g16488(.A1(new_n14061_), .A2(new_n13909_), .ZN(new_n17491_));
  NOR3_X1    g16489(.A1(new_n14061_), .A2(new_n13909_), .A3(new_n14054_), .ZN(new_n17492_));
  OAI22_X1   g16490(.A1(new_n17492_), .A2(new_n14055_), .B1(new_n17491_), .B2(new_n14051_), .ZN(new_n17493_));
  NAND2_X1   g16491(.A1(new_n17490_), .A2(new_n17493_), .ZN(new_n17494_));
  NAND2_X1   g16492(.A1(new_n17494_), .A2(new_n17489_), .ZN(new_n17495_));
  NAND2_X1   g16493(.A1(new_n14081_), .A2(new_n14077_), .ZN(new_n17496_));
  NAND2_X1   g16494(.A1(new_n17496_), .A2(new_n14050_), .ZN(new_n17497_));
  AOI22_X1   g16495(.A1(new_n14079_), .A2(new_n14080_), .B1(new_n14076_), .B2(new_n14072_), .ZN(new_n17498_));
  NAND4_X1   g16496(.A1(new_n14079_), .A2(new_n14076_), .A3(new_n14080_), .A4(new_n14072_), .ZN(new_n17499_));
  OAI21_X1   g16497(.A1(new_n14088_), .A2(new_n17498_), .B(new_n17499_), .ZN(new_n17500_));
  NOR2_X1    g16498(.A1(new_n17490_), .A2(new_n17493_), .ZN(new_n17501_));
  NOR2_X1    g16499(.A1(new_n17488_), .A2(new_n17485_), .ZN(new_n17502_));
  NOR4_X1    g16500(.A1(new_n14082_), .A2(new_n14058_), .A3(new_n14062_), .A4(new_n14083_), .ZN(new_n17503_));
  NOR3_X1    g16501(.A1(new_n17501_), .A2(new_n17502_), .A3(new_n17503_), .ZN(new_n17504_));
  AOI22_X1   g16502(.A1(new_n17504_), .A2(new_n17497_), .B1(new_n17495_), .B2(new_n17500_), .ZN(new_n17505_));
  NAND2_X1   g16503(.A1(new_n17481_), .A2(new_n17505_), .ZN(new_n17506_));
  NAND2_X1   g16504(.A1(new_n17478_), .A2(new_n17477_), .ZN(new_n17507_));
  NOR2_X1    g16505(.A1(new_n14132_), .A2(new_n14128_), .ZN(new_n17508_));
  OAI21_X1   g16506(.A1(new_n17508_), .A2(new_n14093_), .B(new_n17479_), .ZN(new_n17509_));
  NOR3_X1    g16507(.A1(new_n17464_), .A2(new_n17470_), .A3(new_n17475_), .ZN(new_n17510_));
  AOI22_X1   g16508(.A1(new_n17510_), .A2(new_n17473_), .B1(new_n17507_), .B2(new_n17509_), .ZN(new_n17511_));
  NOR2_X1    g16509(.A1(new_n17501_), .A2(new_n17502_), .ZN(new_n17512_));
  INV_X1     g16510(.I(new_n17497_), .ZN(new_n17513_));
  AOI21_X1   g16511(.A1(new_n17496_), .A2(new_n14050_), .B(new_n17503_), .ZN(new_n17514_));
  NAND3_X1   g16512(.A1(new_n17494_), .A2(new_n17489_), .A3(new_n17499_), .ZN(new_n17515_));
  OAI22_X1   g16513(.A1(new_n17513_), .A2(new_n17515_), .B1(new_n17514_), .B2(new_n17512_), .ZN(new_n17516_));
  NAND2_X1   g16514(.A1(new_n17516_), .A2(new_n17511_), .ZN(new_n17517_));
  AOI22_X1   g16515(.A1(new_n17517_), .A2(new_n17506_), .B1(new_n17455_), .B2(new_n17454_), .ZN(new_n17518_));
  NOR2_X1    g16516(.A1(new_n14092_), .A2(new_n14149_), .ZN(new_n17519_));
  AOI21_X1   g16517(.A1(new_n14092_), .A2(new_n14149_), .B(new_n14048_), .ZN(new_n17520_));
  NOR2_X1    g16518(.A1(new_n17516_), .A2(new_n17511_), .ZN(new_n17521_));
  NOR2_X1    g16519(.A1(new_n17481_), .A2(new_n17505_), .ZN(new_n17522_));
  NOR4_X1    g16520(.A1(new_n17521_), .A2(new_n17520_), .A3(new_n17522_), .A4(new_n17519_), .ZN(new_n17523_));
  NOR2_X1    g16521(.A1(new_n17523_), .A2(new_n17518_), .ZN(new_n17524_));
  NOR2_X1    g16522(.A1(new_n14036_), .A2(new_n14032_), .ZN(new_n17525_));
  AOI22_X1   g16523(.A1(new_n14034_), .A2(new_n14035_), .B1(new_n14027_), .B2(new_n14031_), .ZN(new_n17526_));
  NOR2_X1    g16524(.A1(new_n17526_), .A2(new_n14043_), .ZN(new_n17527_));
  OAI21_X1   g16525(.A1(new_n13611_), .A2(new_n14012_), .B(new_n14000_), .ZN(new_n17528_));
  NAND2_X1   g16526(.A1(new_n13631_), .A2(new_n14006_), .ZN(new_n17529_));
  OAI21_X1   g16527(.A1(new_n17529_), .A2(new_n14012_), .B(new_n14010_), .ZN(new_n17530_));
  NAND2_X1   g16528(.A1(new_n17530_), .A2(new_n17528_), .ZN(new_n17531_));
  NAND2_X1   g16529(.A1(new_n13993_), .A2(new_n13641_), .ZN(new_n17532_));
  NAND3_X1   g16530(.A1(new_n13993_), .A2(new_n13641_), .A3(new_n13987_), .ZN(new_n17533_));
  AOI22_X1   g16531(.A1(new_n17533_), .A2(new_n13988_), .B1(new_n17532_), .B2(new_n13990_), .ZN(new_n17534_));
  NAND2_X1   g16532(.A1(new_n17534_), .A2(new_n17531_), .ZN(new_n17535_));
  NAND2_X1   g16533(.A1(new_n14016_), .A2(new_n13631_), .ZN(new_n17536_));
  NAND3_X1   g16534(.A1(new_n14016_), .A2(new_n13631_), .A3(new_n14006_), .ZN(new_n17537_));
  AOI22_X1   g16535(.A1(new_n17537_), .A2(new_n14010_), .B1(new_n17536_), .B2(new_n14000_), .ZN(new_n17538_));
  NOR2_X1    g16536(.A1(new_n13997_), .A2(new_n13560_), .ZN(new_n17539_));
  OAI21_X1   g16537(.A1(new_n13552_), .A2(new_n13559_), .B(new_n13987_), .ZN(new_n17540_));
  NOR2_X1    g16538(.A1(new_n17540_), .A2(new_n13997_), .ZN(new_n17541_));
  OAI22_X1   g16539(.A1(new_n17541_), .A2(new_n13991_), .B1(new_n17539_), .B2(new_n13987_), .ZN(new_n17542_));
  NAND2_X1   g16540(.A1(new_n17542_), .A2(new_n17538_), .ZN(new_n17543_));
  NAND2_X1   g16541(.A1(new_n17535_), .A2(new_n17543_), .ZN(new_n17544_));
  AOI22_X1   g16542(.A1(new_n14020_), .A2(new_n14021_), .B1(new_n14013_), .B2(new_n14017_), .ZN(new_n17545_));
  NOR2_X1    g16543(.A1(new_n14028_), .A2(new_n17545_), .ZN(new_n17546_));
  INV_X1     g16544(.I(new_n17546_), .ZN(new_n17547_));
  NAND4_X1   g16545(.A1(new_n14020_), .A2(new_n14021_), .A3(new_n14013_), .A4(new_n14017_), .ZN(new_n17548_));
  OAI21_X1   g16546(.A1(new_n14028_), .A2(new_n17545_), .B(new_n17548_), .ZN(new_n17549_));
  NOR2_X1    g16547(.A1(new_n17542_), .A2(new_n17538_), .ZN(new_n17550_));
  NOR2_X1    g16548(.A1(new_n17534_), .A2(new_n17531_), .ZN(new_n17551_));
  NOR4_X1    g16549(.A1(new_n13994_), .A2(new_n13998_), .A3(new_n14023_), .A4(new_n14024_), .ZN(new_n17552_));
  NOR3_X1    g16550(.A1(new_n17551_), .A2(new_n17550_), .A3(new_n17552_), .ZN(new_n17553_));
  AOI22_X1   g16551(.A1(new_n17547_), .A2(new_n17553_), .B1(new_n17544_), .B2(new_n17549_), .ZN(new_n17554_));
  NAND2_X1   g16552(.A1(new_n13494_), .A2(new_n13965_), .ZN(new_n17555_));
  NAND3_X1   g16553(.A1(new_n13494_), .A2(new_n13965_), .A3(new_n13955_), .ZN(new_n17556_));
  AOI22_X1   g16554(.A1(new_n17556_), .A2(new_n13958_), .B1(new_n17555_), .B2(new_n13961_), .ZN(new_n17557_));
  OAI21_X1   g16555(.A1(new_n13948_), .A2(new_n13521_), .B(new_n13942_), .ZN(new_n17558_));
  OAI21_X1   g16556(.A1(new_n13519_), .A2(new_n13520_), .B(new_n13945_), .ZN(new_n17559_));
  OAI21_X1   g16557(.A1(new_n17559_), .A2(new_n13948_), .B(new_n13946_), .ZN(new_n17560_));
  NAND2_X1   g16558(.A1(new_n17560_), .A2(new_n17558_), .ZN(new_n17561_));
  NOR2_X1    g16559(.A1(new_n17557_), .A2(new_n17561_), .ZN(new_n17562_));
  OAI21_X1   g16560(.A1(new_n13969_), .A2(new_n13531_), .B(new_n13961_), .ZN(new_n17563_));
  OAI21_X1   g16561(.A1(new_n13529_), .A2(new_n13530_), .B(new_n13955_), .ZN(new_n17564_));
  OAI21_X1   g16562(.A1(new_n13969_), .A2(new_n17564_), .B(new_n13958_), .ZN(new_n17565_));
  NAND2_X1   g16563(.A1(new_n17565_), .A2(new_n17563_), .ZN(new_n17566_));
  NAND2_X1   g16564(.A1(new_n13952_), .A2(new_n13448_), .ZN(new_n17567_));
  NAND3_X1   g16565(.A1(new_n13952_), .A2(new_n13448_), .A3(new_n13945_), .ZN(new_n17568_));
  AOI22_X1   g16566(.A1(new_n17568_), .A2(new_n13946_), .B1(new_n17567_), .B2(new_n13942_), .ZN(new_n17569_));
  NOR2_X1    g16567(.A1(new_n17569_), .A2(new_n17566_), .ZN(new_n17570_));
  NOR2_X1    g16568(.A1(new_n17570_), .A2(new_n17562_), .ZN(new_n17571_));
  AOI22_X1   g16569(.A1(new_n13949_), .A2(new_n13953_), .B1(new_n13976_), .B2(new_n13977_), .ZN(new_n17572_));
  NOR2_X1    g16570(.A1(new_n13941_), .A2(new_n17572_), .ZN(new_n17573_));
  OAI22_X1   g16571(.A1(new_n13973_), .A2(new_n13974_), .B1(new_n13970_), .B2(new_n13966_), .ZN(new_n17574_));
  NOR4_X1    g16572(.A1(new_n13973_), .A2(new_n13974_), .A3(new_n13970_), .A4(new_n13966_), .ZN(new_n17575_));
  AOI21_X1   g16573(.A1(new_n13981_), .A2(new_n17574_), .B(new_n17575_), .ZN(new_n17576_));
  NAND2_X1   g16574(.A1(new_n17569_), .A2(new_n17566_), .ZN(new_n17577_));
  NAND2_X1   g16575(.A1(new_n17557_), .A2(new_n17561_), .ZN(new_n17578_));
  NAND4_X1   g16576(.A1(new_n13949_), .A2(new_n13953_), .A3(new_n13976_), .A4(new_n13977_), .ZN(new_n17579_));
  NAND3_X1   g16577(.A1(new_n17577_), .A2(new_n17578_), .A3(new_n17579_), .ZN(new_n17580_));
  OAI22_X1   g16578(.A1(new_n17571_), .A2(new_n17576_), .B1(new_n17580_), .B2(new_n17573_), .ZN(new_n17581_));
  NOR2_X1    g16579(.A1(new_n17554_), .A2(new_n17581_), .ZN(new_n17582_));
  NOR2_X1    g16580(.A1(new_n17551_), .A2(new_n17550_), .ZN(new_n17583_));
  NAND2_X1   g16581(.A1(new_n14022_), .A2(new_n14018_), .ZN(new_n17584_));
  AOI21_X1   g16582(.A1(new_n17584_), .A2(new_n13986_), .B(new_n17552_), .ZN(new_n17585_));
  NAND3_X1   g16583(.A1(new_n17535_), .A2(new_n17543_), .A3(new_n17548_), .ZN(new_n17586_));
  OAI22_X1   g16584(.A1(new_n17546_), .A2(new_n17586_), .B1(new_n17583_), .B2(new_n17585_), .ZN(new_n17587_));
  NAND2_X1   g16585(.A1(new_n17577_), .A2(new_n17578_), .ZN(new_n17588_));
  NAND2_X1   g16586(.A1(new_n13981_), .A2(new_n17574_), .ZN(new_n17589_));
  OAI21_X1   g16587(.A1(new_n13941_), .A2(new_n17572_), .B(new_n17579_), .ZN(new_n17590_));
  NOR3_X1    g16588(.A1(new_n17570_), .A2(new_n17562_), .A3(new_n17575_), .ZN(new_n17591_));
  AOI22_X1   g16589(.A1(new_n17591_), .A2(new_n17589_), .B1(new_n17588_), .B2(new_n17590_), .ZN(new_n17592_));
  NOR2_X1    g16590(.A1(new_n17587_), .A2(new_n17592_), .ZN(new_n17593_));
  OAI22_X1   g16591(.A1(new_n17525_), .A2(new_n17527_), .B1(new_n17582_), .B2(new_n17593_), .ZN(new_n17594_));
  NAND2_X1   g16592(.A1(new_n13985_), .A2(new_n14039_), .ZN(new_n17595_));
  OAI21_X1   g16593(.A1(new_n13985_), .A2(new_n14039_), .B(new_n13940_), .ZN(new_n17596_));
  NAND2_X1   g16594(.A1(new_n17587_), .A2(new_n17592_), .ZN(new_n17597_));
  NAND2_X1   g16595(.A1(new_n17554_), .A2(new_n17581_), .ZN(new_n17598_));
  NAND4_X1   g16596(.A1(new_n17596_), .A2(new_n17598_), .A3(new_n17597_), .A4(new_n17595_), .ZN(new_n17599_));
  NAND2_X1   g16597(.A1(new_n17594_), .A2(new_n17599_), .ZN(new_n17600_));
  NOR2_X1    g16598(.A1(new_n17524_), .A2(new_n17600_), .ZN(new_n17601_));
  OAI22_X1   g16599(.A1(new_n17521_), .A2(new_n17522_), .B1(new_n17520_), .B2(new_n17519_), .ZN(new_n17602_));
  NAND4_X1   g16600(.A1(new_n17517_), .A2(new_n17455_), .A3(new_n17506_), .A4(new_n17454_), .ZN(new_n17603_));
  NAND2_X1   g16601(.A1(new_n17602_), .A2(new_n17603_), .ZN(new_n17604_));
  AOI22_X1   g16602(.A1(new_n17597_), .A2(new_n17598_), .B1(new_n17596_), .B2(new_n17595_), .ZN(new_n17605_));
  NOR4_X1    g16603(.A1(new_n17527_), .A2(new_n17582_), .A3(new_n17593_), .A4(new_n17525_), .ZN(new_n17606_));
  NOR2_X1    g16604(.A1(new_n17605_), .A2(new_n17606_), .ZN(new_n17607_));
  NOR2_X1    g16605(.A1(new_n17604_), .A2(new_n17607_), .ZN(new_n17608_));
  OAI22_X1   g16606(.A1(new_n17608_), .A2(new_n17601_), .B1(new_n17453_), .B2(new_n17452_), .ZN(new_n17609_));
  NAND2_X1   g16607(.A1(new_n14161_), .A2(new_n14157_), .ZN(new_n17610_));
  OAI21_X1   g16608(.A1(new_n14161_), .A2(new_n14157_), .B(new_n14167_), .ZN(new_n17611_));
  NAND2_X1   g16609(.A1(new_n17604_), .A2(new_n17607_), .ZN(new_n17612_));
  NAND2_X1   g16610(.A1(new_n17524_), .A2(new_n17600_), .ZN(new_n17613_));
  NAND4_X1   g16611(.A1(new_n17612_), .A2(new_n17613_), .A3(new_n17610_), .A4(new_n17611_), .ZN(new_n17614_));
  NAND2_X1   g16612(.A1(new_n17609_), .A2(new_n17614_), .ZN(new_n17615_));
  NOR2_X1    g16613(.A1(new_n17451_), .A2(new_n17615_), .ZN(new_n17616_));
  OAI22_X1   g16614(.A1(new_n17449_), .A2(new_n17448_), .B1(new_n17446_), .B2(new_n17447_), .ZN(new_n17617_));
  NAND4_X1   g16615(.A1(new_n17437_), .A2(new_n17444_), .A3(new_n17294_), .A4(new_n17295_), .ZN(new_n17618_));
  NAND2_X1   g16616(.A1(new_n17617_), .A2(new_n17618_), .ZN(new_n17619_));
  AOI22_X1   g16617(.A1(new_n17612_), .A2(new_n17613_), .B1(new_n17610_), .B2(new_n17611_), .ZN(new_n17620_));
  NOR4_X1    g16618(.A1(new_n17608_), .A2(new_n17601_), .A3(new_n17453_), .A4(new_n17452_), .ZN(new_n17621_));
  NOR2_X1    g16619(.A1(new_n17620_), .A2(new_n17621_), .ZN(new_n17622_));
  NOR2_X1    g16620(.A1(new_n17622_), .A2(new_n17619_), .ZN(new_n17623_));
  OAI22_X1   g16621(.A1(new_n17623_), .A2(new_n17616_), .B1(new_n17292_), .B2(new_n17293_), .ZN(new_n17624_));
  NOR2_X1    g16622(.A1(new_n17293_), .A2(new_n17292_), .ZN(new_n17625_));
  NAND2_X1   g16623(.A1(new_n17622_), .A2(new_n17619_), .ZN(new_n17626_));
  NAND2_X1   g16624(.A1(new_n17451_), .A2(new_n17615_), .ZN(new_n17627_));
  NAND3_X1   g16625(.A1(new_n17625_), .A2(new_n17626_), .A3(new_n17627_), .ZN(new_n17628_));
  NAND2_X1   g16626(.A1(new_n17624_), .A2(new_n17628_), .ZN(new_n17629_));
  NOR2_X1    g16627(.A1(new_n17291_), .A2(new_n17629_), .ZN(new_n17630_));
  OAI21_X1   g16628(.A1(new_n17288_), .A2(new_n17289_), .B(new_n17287_), .ZN(new_n17631_));
  NAND3_X1   g16629(.A1(new_n17275_), .A2(new_n17283_), .A3(new_n16965_), .ZN(new_n17632_));
  NAND2_X1   g16630(.A1(new_n17631_), .A2(new_n17632_), .ZN(new_n17633_));
  AOI21_X1   g16631(.A1(new_n17626_), .A2(new_n17627_), .B(new_n17625_), .ZN(new_n17634_));
  NOR4_X1    g16632(.A1(new_n17623_), .A2(new_n17616_), .A3(new_n17292_), .A4(new_n17293_), .ZN(new_n17635_));
  NOR2_X1    g16633(.A1(new_n17634_), .A2(new_n17635_), .ZN(new_n17636_));
  NOR2_X1    g16634(.A1(new_n17636_), .A2(new_n17633_), .ZN(new_n17637_));
  OAI21_X1   g16635(.A1(new_n17637_), .A2(new_n17630_), .B(new_n16962_), .ZN(new_n17638_));
  NAND2_X1   g16636(.A1(new_n14422_), .A2(new_n14431_), .ZN(new_n17639_));
  NAND2_X1   g16637(.A1(new_n16933_), .A2(new_n16942_), .ZN(new_n17640_));
  NOR2_X1    g16638(.A1(new_n17639_), .A2(new_n17640_), .ZN(new_n17641_));
  NAND2_X1   g16639(.A1(new_n17639_), .A2(new_n17640_), .ZN(new_n17642_));
  AOI21_X1   g16640(.A1(new_n16959_), .A2(new_n17642_), .B(new_n17641_), .ZN(new_n17643_));
  NAND2_X1   g16641(.A1(new_n17636_), .A2(new_n17633_), .ZN(new_n17644_));
  NAND2_X1   g16642(.A1(new_n17291_), .A2(new_n17629_), .ZN(new_n17645_));
  NAND3_X1   g16643(.A1(new_n17643_), .A2(new_n17644_), .A3(new_n17645_), .ZN(new_n17646_));
  NAND2_X1   g16644(.A1(new_n17646_), .A2(new_n17638_), .ZN(new_n17647_));
  NOR3_X1    g16645(.A1(new_n11873_), .A2(new_n11879_), .A3(new_n17647_), .ZN(new_n17648_));
  NAND3_X1   g16646(.A1(new_n10670_), .A2(new_n10676_), .A3(new_n10696_), .ZN(new_n17649_));
  OAI21_X1   g16647(.A1(new_n10698_), .A2(new_n10697_), .B(new_n4171_), .ZN(new_n17650_));
  AOI21_X1   g16648(.A1(new_n17650_), .A2(new_n17649_), .B(new_n11874_), .ZN(new_n17651_));
  NAND3_X1   g16649(.A1(new_n17650_), .A2(new_n17649_), .A3(new_n11874_), .ZN(new_n17652_));
  AOI21_X1   g16650(.A1(new_n16940_), .A2(new_n16941_), .B(new_n16939_), .ZN(new_n17653_));
  NOR3_X1    g16651(.A1(new_n16932_), .A2(new_n16925_), .A3(new_n16426_), .ZN(new_n17654_));
  NOR2_X1    g16652(.A1(new_n17654_), .A2(new_n17653_), .ZN(new_n17655_));
  NAND2_X1   g16653(.A1(new_n17639_), .A2(new_n17655_), .ZN(new_n17656_));
  NAND3_X1   g16654(.A1(new_n17640_), .A2(new_n14422_), .A3(new_n14431_), .ZN(new_n17657_));
  AOI21_X1   g16655(.A1(new_n17656_), .A2(new_n17657_), .B(new_n16960_), .ZN(new_n17658_));
  AOI21_X1   g16656(.A1(new_n14429_), .A2(new_n14430_), .B(new_n14428_), .ZN(new_n17659_));
  NOR3_X1    g16657(.A1(new_n14421_), .A2(new_n14414_), .A3(new_n13936_), .ZN(new_n17660_));
  NOR2_X1    g16658(.A1(new_n17659_), .A2(new_n17660_), .ZN(new_n17661_));
  NOR2_X1    g16659(.A1(new_n17661_), .A2(new_n17640_), .ZN(new_n17662_));
  NOR2_X1    g16660(.A1(new_n17639_), .A2(new_n17655_), .ZN(new_n17663_));
  NOR3_X1    g16661(.A1(new_n17663_), .A2(new_n17662_), .A3(new_n16959_), .ZN(new_n17664_));
  NOR2_X1    g16662(.A1(new_n17664_), .A2(new_n17658_), .ZN(new_n17665_));
  NAND2_X1   g16663(.A1(new_n17652_), .A2(new_n17665_), .ZN(new_n17666_));
  XNOR2_X1   g16664(.A1(new_n16945_), .A2(new_n16944_), .ZN(new_n17667_));
  INV_X1     g16665(.I(new_n10681_), .ZN(new_n17668_));
  NOR2_X1    g16666(.A1(new_n10678_), .A2(new_n17668_), .ZN(new_n17669_));
  NAND2_X1   g16667(.A1(new_n10678_), .A2(new_n17668_), .ZN(new_n17670_));
  INV_X1     g16668(.I(new_n17670_), .ZN(new_n17671_));
  NOR2_X1    g16669(.A1(new_n17671_), .A2(new_n17669_), .ZN(new_n17672_));
  NOR2_X1    g16670(.A1(new_n17672_), .A2(new_n17667_), .ZN(new_n17673_));
  INV_X1     g16671(.I(new_n17673_), .ZN(new_n17674_));
  INV_X1     g16672(.I(new_n10682_), .ZN(new_n17675_));
  NOR3_X1    g16673(.A1(new_n10685_), .A2(new_n10686_), .A3(new_n17675_), .ZN(new_n17676_));
  OAI21_X1   g16674(.A1(new_n10685_), .A2(new_n10686_), .B(new_n17675_), .ZN(new_n17677_));
  INV_X1     g16675(.I(new_n17677_), .ZN(new_n17678_));
  OAI21_X1   g16676(.A1(new_n17678_), .A2(new_n17676_), .B(new_n10693_), .ZN(new_n17679_));
  INV_X1     g16677(.I(new_n10685_), .ZN(new_n17680_));
  OAI21_X1   g16678(.A1(new_n9668_), .A2(new_n10671_), .B(new_n10672_), .ZN(new_n17681_));
  AOI21_X1   g16679(.A1(new_n17680_), .A2(new_n17681_), .B(new_n17675_), .ZN(new_n17682_));
  OAI21_X1   g16680(.A1(new_n17682_), .A2(new_n10694_), .B(new_n10692_), .ZN(new_n17683_));
  AOI21_X1   g16681(.A1(new_n17679_), .A2(new_n17683_), .B(new_n17674_), .ZN(new_n17684_));
  NOR2_X1    g16682(.A1(new_n16952_), .A2(new_n16946_), .ZN(new_n17685_));
  NOR3_X1    g16683(.A1(new_n16950_), .A2(new_n16951_), .A3(new_n16947_), .ZN(new_n17686_));
  OAI21_X1   g16684(.A1(new_n17685_), .A2(new_n17686_), .B(new_n16957_), .ZN(new_n17687_));
  NOR2_X1    g16685(.A1(new_n16952_), .A2(new_n16947_), .ZN(new_n17688_));
  OAI22_X1   g16686(.A1(new_n17688_), .A2(new_n16958_), .B1(new_n16955_), .B2(new_n16956_), .ZN(new_n17689_));
  NAND2_X1   g16687(.A1(new_n17689_), .A2(new_n17687_), .ZN(new_n17690_));
  NAND3_X1   g16688(.A1(new_n17679_), .A2(new_n17683_), .A3(new_n17674_), .ZN(new_n17691_));
  AOI21_X1   g16689(.A1(new_n17690_), .A2(new_n17691_), .B(new_n17684_), .ZN(new_n17692_));
  NOR3_X1    g16690(.A1(new_n10698_), .A2(new_n10697_), .A3(new_n4171_), .ZN(new_n17693_));
  AOI21_X1   g16691(.A1(new_n10670_), .A2(new_n10676_), .B(new_n10696_), .ZN(new_n17694_));
  OAI21_X1   g16692(.A1(new_n17693_), .A2(new_n17694_), .B(new_n10695_), .ZN(new_n17695_));
  AOI21_X1   g16693(.A1(new_n17695_), .A2(new_n17652_), .B(new_n17665_), .ZN(new_n17696_));
  OAI22_X1   g16694(.A1(new_n17696_), .A2(new_n17692_), .B1(new_n17666_), .B2(new_n17651_), .ZN(new_n17697_));
  OAI21_X1   g16695(.A1(new_n11873_), .A2(new_n11879_), .B(new_n17647_), .ZN(new_n17698_));
  AOI21_X1   g16696(.A1(new_n17697_), .A2(new_n17698_), .B(new_n17648_), .ZN(new_n17699_));
  OAI22_X1   g16697(.A1(new_n17634_), .A2(new_n17635_), .B1(new_n17290_), .B2(new_n17284_), .ZN(new_n17700_));
  NOR4_X1    g16698(.A1(new_n17290_), .A2(new_n17634_), .A3(new_n17284_), .A4(new_n17635_), .ZN(new_n17701_));
  AOI21_X1   g16699(.A1(new_n16962_), .A2(new_n17700_), .B(new_n17701_), .ZN(new_n17702_));
  NOR2_X1    g16700(.A1(new_n17619_), .A2(new_n17615_), .ZN(new_n17703_));
  NAND2_X1   g16701(.A1(new_n14171_), .A2(new_n14420_), .ZN(new_n17704_));
  OAI21_X1   g16702(.A1(new_n14171_), .A2(new_n14420_), .B(new_n13936_), .ZN(new_n17705_));
  AOI22_X1   g16703(.A1(new_n17705_), .A2(new_n17704_), .B1(new_n17619_), .B2(new_n17615_), .ZN(new_n17706_));
  NOR2_X1    g16704(.A1(new_n17604_), .A2(new_n17600_), .ZN(new_n17707_));
  AOI22_X1   g16705(.A1(new_n17611_), .A2(new_n17610_), .B1(new_n17604_), .B2(new_n17600_), .ZN(new_n17708_));
  NOR2_X1    g16706(.A1(new_n17554_), .A2(new_n17592_), .ZN(new_n17709_));
  AOI21_X1   g16707(.A1(new_n17595_), .A2(new_n17596_), .B(new_n17709_), .ZN(new_n17710_));
  NAND2_X1   g16708(.A1(new_n17596_), .A2(new_n17595_), .ZN(new_n17711_));
  NOR2_X1    g16709(.A1(new_n17583_), .A2(new_n17585_), .ZN(new_n17712_));
  NOR2_X1    g16710(.A1(new_n17586_), .A2(new_n17546_), .ZN(new_n17713_));
  NOR2_X1    g16711(.A1(new_n17576_), .A2(new_n17571_), .ZN(new_n17714_));
  NOR2_X1    g16712(.A1(new_n17580_), .A2(new_n17573_), .ZN(new_n17715_));
  NOR4_X1    g16713(.A1(new_n17712_), .A2(new_n17713_), .A3(new_n17714_), .A4(new_n17715_), .ZN(new_n17716_));
  INV_X1     g16714(.I(new_n17709_), .ZN(new_n17717_));
  AOI21_X1   g16715(.A1(new_n17711_), .A2(new_n17717_), .B(new_n17716_), .ZN(new_n17718_));
  NAND2_X1   g16716(.A1(new_n17534_), .A2(new_n17538_), .ZN(new_n17719_));
  NOR2_X1    g16717(.A1(new_n17534_), .A2(new_n17538_), .ZN(new_n17720_));
  AOI21_X1   g16718(.A1(new_n17549_), .A2(new_n17719_), .B(new_n17720_), .ZN(new_n17721_));
  INV_X1     g16719(.I(new_n17721_), .ZN(new_n17722_));
  NAND2_X1   g16720(.A1(new_n17569_), .A2(new_n17557_), .ZN(new_n17723_));
  NOR2_X1    g16721(.A1(new_n17569_), .A2(new_n17557_), .ZN(new_n17724_));
  AOI21_X1   g16722(.A1(new_n17590_), .A2(new_n17723_), .B(new_n17724_), .ZN(new_n17725_));
  NAND2_X1   g16723(.A1(new_n17722_), .A2(new_n17725_), .ZN(new_n17726_));
  INV_X1     g16724(.I(new_n17725_), .ZN(new_n17727_));
  NAND2_X1   g16725(.A1(new_n17727_), .A2(new_n17721_), .ZN(new_n17728_));
  NAND2_X1   g16726(.A1(new_n17726_), .A2(new_n17728_), .ZN(new_n17729_));
  INV_X1     g16727(.I(new_n17729_), .ZN(new_n17730_));
  OR4_X2     g16728(.A1(new_n17712_), .A2(new_n17714_), .A3(new_n17713_), .A4(new_n17715_), .Z(new_n17731_));
  NAND3_X1   g16729(.A1(new_n17731_), .A2(new_n17728_), .A3(new_n17726_), .ZN(new_n17732_));
  OAI22_X1   g16730(.A1(new_n17718_), .A2(new_n17730_), .B1(new_n17732_), .B2(new_n17710_), .ZN(new_n17733_));
  NAND2_X1   g16731(.A1(new_n17455_), .A2(new_n17454_), .ZN(new_n17734_));
  NOR2_X1    g16732(.A1(new_n17511_), .A2(new_n17505_), .ZN(new_n17735_));
  INV_X1     g16733(.I(new_n17735_), .ZN(new_n17736_));
  NAND2_X1   g16734(.A1(new_n17734_), .A2(new_n17736_), .ZN(new_n17737_));
  NOR2_X1    g16735(.A1(new_n17520_), .A2(new_n17519_), .ZN(new_n17738_));
  NAND2_X1   g16736(.A1(new_n17507_), .A2(new_n17509_), .ZN(new_n17739_));
  NAND2_X1   g16737(.A1(new_n17510_), .A2(new_n17473_), .ZN(new_n17740_));
  NAND2_X1   g16738(.A1(new_n17495_), .A2(new_n17500_), .ZN(new_n17741_));
  NAND2_X1   g16739(.A1(new_n17504_), .A2(new_n17497_), .ZN(new_n17742_));
  NAND4_X1   g16740(.A1(new_n17740_), .A2(new_n17742_), .A3(new_n17739_), .A4(new_n17741_), .ZN(new_n17743_));
  OAI21_X1   g16741(.A1(new_n17738_), .A2(new_n17735_), .B(new_n17743_), .ZN(new_n17744_));
  NAND2_X1   g16742(.A1(new_n17458_), .A2(new_n17469_), .ZN(new_n17745_));
  NOR2_X1    g16743(.A1(new_n17458_), .A2(new_n17469_), .ZN(new_n17746_));
  AOI21_X1   g16744(.A1(new_n17509_), .A2(new_n17745_), .B(new_n17746_), .ZN(new_n17747_));
  NAND2_X1   g16745(.A1(new_n17490_), .A2(new_n17488_), .ZN(new_n17748_));
  NOR2_X1    g16746(.A1(new_n17490_), .A2(new_n17488_), .ZN(new_n17749_));
  AOI21_X1   g16747(.A1(new_n17500_), .A2(new_n17748_), .B(new_n17749_), .ZN(new_n17750_));
  INV_X1     g16748(.I(new_n17750_), .ZN(new_n17751_));
  NOR2_X1    g16749(.A1(new_n17751_), .A2(new_n17747_), .ZN(new_n17752_));
  INV_X1     g16750(.I(new_n17747_), .ZN(new_n17753_));
  NOR2_X1    g16751(.A1(new_n17753_), .A2(new_n17750_), .ZN(new_n17754_));
  NOR2_X1    g16752(.A1(new_n17754_), .A2(new_n17752_), .ZN(new_n17755_));
  INV_X1     g16753(.I(new_n17755_), .ZN(new_n17756_));
  INV_X1     g16754(.I(new_n17743_), .ZN(new_n17757_));
  NOR3_X1    g16755(.A1(new_n17757_), .A2(new_n17752_), .A3(new_n17754_), .ZN(new_n17758_));
  AOI22_X1   g16756(.A1(new_n17744_), .A2(new_n17756_), .B1(new_n17737_), .B2(new_n17758_), .ZN(new_n17759_));
  NOR2_X1    g16757(.A1(new_n17759_), .A2(new_n17733_), .ZN(new_n17760_));
  NAND2_X1   g16758(.A1(new_n17711_), .A2(new_n17717_), .ZN(new_n17761_));
  NOR2_X1    g16759(.A1(new_n17527_), .A2(new_n17525_), .ZN(new_n17762_));
  OAI21_X1   g16760(.A1(new_n17762_), .A2(new_n17709_), .B(new_n17731_), .ZN(new_n17763_));
  INV_X1     g16761(.I(new_n17726_), .ZN(new_n17764_));
  NOR2_X1    g16762(.A1(new_n17722_), .A2(new_n17725_), .ZN(new_n17765_));
  NOR3_X1    g16763(.A1(new_n17764_), .A2(new_n17716_), .A3(new_n17765_), .ZN(new_n17766_));
  AOI22_X1   g16764(.A1(new_n17763_), .A2(new_n17729_), .B1(new_n17761_), .B2(new_n17766_), .ZN(new_n17767_));
  NOR2_X1    g16765(.A1(new_n17738_), .A2(new_n17735_), .ZN(new_n17768_));
  AOI21_X1   g16766(.A1(new_n17734_), .A2(new_n17736_), .B(new_n17757_), .ZN(new_n17769_));
  INV_X1     g16767(.I(new_n17752_), .ZN(new_n17770_));
  INV_X1     g16768(.I(new_n17754_), .ZN(new_n17771_));
  NAND3_X1   g16769(.A1(new_n17771_), .A2(new_n17770_), .A3(new_n17743_), .ZN(new_n17772_));
  OAI22_X1   g16770(.A1(new_n17769_), .A2(new_n17755_), .B1(new_n17768_), .B2(new_n17772_), .ZN(new_n17773_));
  NOR2_X1    g16771(.A1(new_n17773_), .A2(new_n17767_), .ZN(new_n17774_));
  OAI22_X1   g16772(.A1(new_n17708_), .A2(new_n17707_), .B1(new_n17774_), .B2(new_n17760_), .ZN(new_n17775_));
  INV_X1     g16773(.I(new_n17707_), .ZN(new_n17776_));
  OAI22_X1   g16774(.A1(new_n17518_), .A2(new_n17523_), .B1(new_n17605_), .B2(new_n17606_), .ZN(new_n17777_));
  OAI21_X1   g16775(.A1(new_n17453_), .A2(new_n17452_), .B(new_n17777_), .ZN(new_n17778_));
  NAND2_X1   g16776(.A1(new_n17773_), .A2(new_n17767_), .ZN(new_n17779_));
  NAND2_X1   g16777(.A1(new_n17759_), .A2(new_n17733_), .ZN(new_n17780_));
  NAND4_X1   g16778(.A1(new_n17778_), .A2(new_n17779_), .A3(new_n17780_), .A4(new_n17776_), .ZN(new_n17781_));
  NAND2_X1   g16779(.A1(new_n17775_), .A2(new_n17781_), .ZN(new_n17782_));
  NAND2_X1   g16780(.A1(new_n17440_), .A2(new_n17436_), .ZN(new_n17783_));
  OAI22_X1   g16781(.A1(new_n17447_), .A2(new_n17446_), .B1(new_n17440_), .B2(new_n17436_), .ZN(new_n17784_));
  NAND2_X1   g16782(.A1(new_n17368_), .A2(new_n17367_), .ZN(new_n17785_));
  NAND2_X1   g16783(.A1(new_n17428_), .A2(new_n17392_), .ZN(new_n17786_));
  NAND2_X1   g16784(.A1(new_n17785_), .A2(new_n17786_), .ZN(new_n17787_));
  NOR2_X1    g16785(.A1(new_n17432_), .A2(new_n17431_), .ZN(new_n17788_));
  NOR2_X1    g16786(.A1(new_n17382_), .A2(new_n17387_), .ZN(new_n17789_));
  NOR2_X1    g16787(.A1(new_n17391_), .A2(new_n17384_), .ZN(new_n17790_));
  NOR2_X1    g16788(.A1(new_n17424_), .A2(new_n17426_), .ZN(new_n17791_));
  NOR2_X1    g16789(.A1(new_n17427_), .A2(new_n17425_), .ZN(new_n17792_));
  OR4_X2     g16790(.A1(new_n17789_), .A2(new_n17792_), .A3(new_n17790_), .A4(new_n17791_), .Z(new_n17793_));
  NOR2_X1    g16791(.A1(new_n17417_), .A2(new_n17423_), .ZN(new_n17794_));
  OAI21_X1   g16792(.A1(new_n17788_), .A2(new_n17794_), .B(new_n17793_), .ZN(new_n17795_));
  NAND2_X1   g16793(.A1(new_n17371_), .A2(new_n17374_), .ZN(new_n17796_));
  NOR2_X1    g16794(.A1(new_n17371_), .A2(new_n17374_), .ZN(new_n17797_));
  AOI21_X1   g16795(.A1(new_n17421_), .A2(new_n17796_), .B(new_n17797_), .ZN(new_n17798_));
  INV_X1     g16796(.I(new_n17798_), .ZN(new_n17799_));
  AOI22_X1   g16797(.A1(new_n17409_), .A2(new_n17411_), .B1(new_n17401_), .B2(new_n17399_), .ZN(new_n17800_));
  NOR2_X1    g16798(.A1(new_n17401_), .A2(new_n17399_), .ZN(new_n17801_));
  NOR2_X1    g16799(.A1(new_n17800_), .A2(new_n17801_), .ZN(new_n17802_));
  NAND2_X1   g16800(.A1(new_n17802_), .A2(new_n17799_), .ZN(new_n17803_));
  OAI21_X1   g16801(.A1(new_n17395_), .A2(new_n17405_), .B(new_n17412_), .ZN(new_n17804_));
  INV_X1     g16802(.I(new_n17801_), .ZN(new_n17805_));
  NAND2_X1   g16803(.A1(new_n17804_), .A2(new_n17805_), .ZN(new_n17806_));
  NAND2_X1   g16804(.A1(new_n17806_), .A2(new_n17798_), .ZN(new_n17807_));
  NAND2_X1   g16805(.A1(new_n17803_), .A2(new_n17807_), .ZN(new_n17808_));
  NOR4_X1    g16806(.A1(new_n17790_), .A2(new_n17792_), .A3(new_n17791_), .A4(new_n17789_), .ZN(new_n17809_));
  NOR2_X1    g16807(.A1(new_n17806_), .A2(new_n17798_), .ZN(new_n17810_));
  NOR2_X1    g16808(.A1(new_n17802_), .A2(new_n17799_), .ZN(new_n17811_));
  NOR3_X1    g16809(.A1(new_n17811_), .A2(new_n17810_), .A3(new_n17809_), .ZN(new_n17812_));
  AOI22_X1   g16810(.A1(new_n17795_), .A2(new_n17808_), .B1(new_n17787_), .B2(new_n17812_), .ZN(new_n17813_));
  NOR2_X1    g16811(.A1(new_n17297_), .A2(new_n17296_), .ZN(new_n17814_));
  NOR2_X1    g16812(.A1(new_n17358_), .A2(new_n17321_), .ZN(new_n17815_));
  NOR2_X1    g16813(.A1(new_n17814_), .A2(new_n17815_), .ZN(new_n17816_));
  NOR2_X1    g16814(.A1(new_n14336_), .A2(new_n14391_), .ZN(new_n17817_));
  OAI21_X1   g16815(.A1(new_n14394_), .A2(new_n17817_), .B(new_n17361_), .ZN(new_n17818_));
  NAND2_X1   g16816(.A1(new_n17311_), .A2(new_n17316_), .ZN(new_n17819_));
  NAND2_X1   g16817(.A1(new_n17320_), .A2(new_n17313_), .ZN(new_n17820_));
  NAND2_X1   g16818(.A1(new_n17354_), .A2(new_n17356_), .ZN(new_n17821_));
  NAND2_X1   g16819(.A1(new_n17357_), .A2(new_n17355_), .ZN(new_n17822_));
  NAND4_X1   g16820(.A1(new_n17822_), .A2(new_n17820_), .A3(new_n17821_), .A4(new_n17819_), .ZN(new_n17823_));
  INV_X1     g16821(.I(new_n17823_), .ZN(new_n17824_));
  INV_X1     g16822(.I(new_n17815_), .ZN(new_n17825_));
  AOI21_X1   g16823(.A1(new_n17818_), .A2(new_n17825_), .B(new_n17824_), .ZN(new_n17826_));
  NAND2_X1   g16824(.A1(new_n17305_), .A2(new_n17301_), .ZN(new_n17827_));
  NOR2_X1    g16825(.A1(new_n17305_), .A2(new_n17301_), .ZN(new_n17828_));
  AOI21_X1   g16826(.A1(new_n17316_), .A2(new_n17827_), .B(new_n17828_), .ZN(new_n17829_));
  NOR2_X1    g16827(.A1(new_n17331_), .A2(new_n17325_), .ZN(new_n17830_));
  NOR2_X1    g16828(.A1(new_n17326_), .A2(new_n17335_), .ZN(new_n17831_));
  INV_X1     g16829(.I(new_n17831_), .ZN(new_n17832_));
  OAI21_X1   g16830(.A1(new_n17343_), .A2(new_n17830_), .B(new_n17832_), .ZN(new_n17833_));
  NOR2_X1    g16831(.A1(new_n17833_), .A2(new_n17829_), .ZN(new_n17834_));
  NAND2_X1   g16832(.A1(new_n17833_), .A2(new_n17829_), .ZN(new_n17835_));
  INV_X1     g16833(.I(new_n17835_), .ZN(new_n17836_));
  NOR2_X1    g16834(.A1(new_n17836_), .A2(new_n17834_), .ZN(new_n17837_));
  INV_X1     g16835(.I(new_n17834_), .ZN(new_n17838_));
  NAND3_X1   g16836(.A1(new_n17838_), .A2(new_n17835_), .A3(new_n17823_), .ZN(new_n17839_));
  OAI22_X1   g16837(.A1(new_n17826_), .A2(new_n17837_), .B1(new_n17816_), .B2(new_n17839_), .ZN(new_n17840_));
  NAND2_X1   g16838(.A1(new_n17840_), .A2(new_n17813_), .ZN(new_n17841_));
  NOR2_X1    g16839(.A1(new_n17788_), .A2(new_n17794_), .ZN(new_n17842_));
  AOI21_X1   g16840(.A1(new_n17785_), .A2(new_n17786_), .B(new_n17809_), .ZN(new_n17843_));
  INV_X1     g16841(.I(new_n17808_), .ZN(new_n17844_));
  NAND3_X1   g16842(.A1(new_n17793_), .A2(new_n17803_), .A3(new_n17807_), .ZN(new_n17845_));
  OAI22_X1   g16843(.A1(new_n17844_), .A2(new_n17843_), .B1(new_n17842_), .B2(new_n17845_), .ZN(new_n17846_));
  NAND2_X1   g16844(.A1(new_n17818_), .A2(new_n17825_), .ZN(new_n17847_));
  OAI21_X1   g16845(.A1(new_n17814_), .A2(new_n17815_), .B(new_n17823_), .ZN(new_n17848_));
  INV_X1     g16846(.I(new_n17837_), .ZN(new_n17849_));
  NOR3_X1    g16847(.A1(new_n17824_), .A2(new_n17836_), .A3(new_n17834_), .ZN(new_n17850_));
  AOI22_X1   g16848(.A1(new_n17848_), .A2(new_n17849_), .B1(new_n17847_), .B2(new_n17850_), .ZN(new_n17851_));
  NAND2_X1   g16849(.A1(new_n17851_), .A2(new_n17846_), .ZN(new_n17852_));
  AOI22_X1   g16850(.A1(new_n17783_), .A2(new_n17784_), .B1(new_n17852_), .B2(new_n17841_), .ZN(new_n17853_));
  NOR2_X1    g16851(.A1(new_n17366_), .A2(new_n17443_), .ZN(new_n17854_));
  AOI22_X1   g16852(.A1(new_n17295_), .A2(new_n17294_), .B1(new_n17366_), .B2(new_n17443_), .ZN(new_n17855_));
  NOR2_X1    g16853(.A1(new_n17851_), .A2(new_n17846_), .ZN(new_n17856_));
  NOR2_X1    g16854(.A1(new_n17840_), .A2(new_n17813_), .ZN(new_n17857_));
  NOR4_X1    g16855(.A1(new_n17856_), .A2(new_n17857_), .A3(new_n17855_), .A4(new_n17854_), .ZN(new_n17858_));
  NOR2_X1    g16856(.A1(new_n17853_), .A2(new_n17858_), .ZN(new_n17859_));
  NOR2_X1    g16857(.A1(new_n17859_), .A2(new_n17782_), .ZN(new_n17860_));
  AOI22_X1   g16858(.A1(new_n17778_), .A2(new_n17776_), .B1(new_n17779_), .B2(new_n17780_), .ZN(new_n17861_));
  NOR4_X1    g16859(.A1(new_n17708_), .A2(new_n17774_), .A3(new_n17760_), .A4(new_n17707_), .ZN(new_n17862_));
  NOR2_X1    g16860(.A1(new_n17861_), .A2(new_n17862_), .ZN(new_n17863_));
  OAI22_X1   g16861(.A1(new_n17856_), .A2(new_n17857_), .B1(new_n17855_), .B2(new_n17854_), .ZN(new_n17864_));
  NAND4_X1   g16862(.A1(new_n17784_), .A2(new_n17852_), .A3(new_n17841_), .A4(new_n17783_), .ZN(new_n17865_));
  NAND2_X1   g16863(.A1(new_n17864_), .A2(new_n17865_), .ZN(new_n17866_));
  NOR2_X1    g16864(.A1(new_n17863_), .A2(new_n17866_), .ZN(new_n17867_));
  OAI22_X1   g16865(.A1(new_n17860_), .A2(new_n17867_), .B1(new_n17703_), .B2(new_n17706_), .ZN(new_n17868_));
  NOR2_X1    g16866(.A1(new_n17706_), .A2(new_n17703_), .ZN(new_n17869_));
  NAND2_X1   g16867(.A1(new_n17863_), .A2(new_n17866_), .ZN(new_n17870_));
  NAND2_X1   g16868(.A1(new_n17859_), .A2(new_n17782_), .ZN(new_n17871_));
  NAND3_X1   g16869(.A1(new_n17869_), .A2(new_n17870_), .A3(new_n17871_), .ZN(new_n17872_));
  NAND2_X1   g16870(.A1(new_n17872_), .A2(new_n17868_), .ZN(new_n17873_));
  OAI22_X1   g16871(.A1(new_n17279_), .A2(new_n17274_), .B1(new_n16964_), .B2(new_n16963_), .ZN(new_n17874_));
  NAND2_X1   g16872(.A1(new_n17279_), .A2(new_n17274_), .ZN(new_n17875_));
  NOR2_X1    g16873(.A1(new_n17188_), .A2(new_n17266_), .ZN(new_n17876_));
  AOI22_X1   g16874(.A1(new_n17122_), .A2(new_n17121_), .B1(new_n17188_), .B2(new_n17266_), .ZN(new_n17877_));
  NOR2_X1    g16875(.A1(new_n17253_), .A2(new_n17252_), .ZN(new_n17878_));
  NOR2_X1    g16876(.A1(new_n17244_), .A2(new_n17238_), .ZN(new_n17879_));
  NOR2_X1    g16877(.A1(new_n17878_), .A2(new_n17879_), .ZN(new_n17880_));
  NAND2_X1   g16878(.A1(new_n17190_), .A2(new_n17189_), .ZN(new_n17881_));
  NOR2_X1    g16879(.A1(new_n17203_), .A2(new_n17208_), .ZN(new_n17882_));
  NOR2_X1    g16880(.A1(new_n17212_), .A2(new_n17205_), .ZN(new_n17883_));
  NOR2_X1    g16881(.A1(new_n17245_), .A2(new_n17247_), .ZN(new_n17884_));
  NOR2_X1    g16882(.A1(new_n17248_), .A2(new_n17246_), .ZN(new_n17885_));
  NOR4_X1    g16883(.A1(new_n17883_), .A2(new_n17882_), .A3(new_n17885_), .A4(new_n17884_), .ZN(new_n17886_));
  INV_X1     g16884(.I(new_n17879_), .ZN(new_n17887_));
  AOI21_X1   g16885(.A1(new_n17881_), .A2(new_n17887_), .B(new_n17886_), .ZN(new_n17888_));
  NAND2_X1   g16886(.A1(new_n17194_), .A2(new_n17201_), .ZN(new_n17889_));
  NOR2_X1    g16887(.A1(new_n17194_), .A2(new_n17201_), .ZN(new_n17890_));
  AOI21_X1   g16888(.A1(new_n17242_), .A2(new_n17889_), .B(new_n17890_), .ZN(new_n17891_));
  NOR2_X1    g16889(.A1(new_n17226_), .A2(new_n17217_), .ZN(new_n17892_));
  NOR2_X1    g16890(.A1(new_n17247_), .A2(new_n17892_), .ZN(new_n17893_));
  INV_X1     g16891(.I(new_n17893_), .ZN(new_n17894_));
  NAND2_X1   g16892(.A1(new_n17226_), .A2(new_n17217_), .ZN(new_n17895_));
  NAND2_X1   g16893(.A1(new_n17894_), .A2(new_n17895_), .ZN(new_n17896_));
  NOR2_X1    g16894(.A1(new_n17896_), .A2(new_n17891_), .ZN(new_n17897_));
  INV_X1     g16895(.I(new_n17891_), .ZN(new_n17898_));
  AOI21_X1   g16896(.A1(new_n17217_), .A2(new_n17226_), .B(new_n17893_), .ZN(new_n17899_));
  NOR2_X1    g16897(.A1(new_n17899_), .A2(new_n17898_), .ZN(new_n17900_));
  NOR2_X1    g16898(.A1(new_n17897_), .A2(new_n17900_), .ZN(new_n17901_));
  INV_X1     g16899(.I(new_n17886_), .ZN(new_n17902_));
  NAND2_X1   g16900(.A1(new_n17899_), .A2(new_n17898_), .ZN(new_n17903_));
  NAND2_X1   g16901(.A1(new_n17896_), .A2(new_n17891_), .ZN(new_n17904_));
  NAND3_X1   g16902(.A1(new_n17902_), .A2(new_n17904_), .A3(new_n17903_), .ZN(new_n17905_));
  OAI22_X1   g16903(.A1(new_n17888_), .A2(new_n17901_), .B1(new_n17880_), .B2(new_n17905_), .ZN(new_n17906_));
  NAND2_X1   g16904(.A1(new_n17134_), .A2(new_n17132_), .ZN(new_n17907_));
  NOR2_X1    g16905(.A1(new_n17134_), .A2(new_n17132_), .ZN(new_n17908_));
  AOI21_X1   g16906(.A1(new_n17142_), .A2(new_n17907_), .B(new_n17908_), .ZN(new_n17909_));
  NAND2_X1   g16907(.A1(new_n17151_), .A2(new_n17158_), .ZN(new_n17910_));
  NOR2_X1    g16908(.A1(new_n17151_), .A2(new_n17158_), .ZN(new_n17911_));
  AOI21_X1   g16909(.A1(new_n17179_), .A2(new_n17910_), .B(new_n17911_), .ZN(new_n17912_));
  INV_X1     g16910(.I(new_n17912_), .ZN(new_n17913_));
  NOR2_X1    g16911(.A1(new_n17913_), .A2(new_n17909_), .ZN(new_n17914_));
  INV_X1     g16912(.I(new_n17909_), .ZN(new_n17915_));
  NOR2_X1    g16913(.A1(new_n17915_), .A2(new_n17912_), .ZN(new_n17916_));
  NOR2_X1    g16914(.A1(new_n17914_), .A2(new_n17916_), .ZN(new_n17917_));
  INV_X1     g16915(.I(new_n17917_), .ZN(new_n17918_));
  NOR2_X1    g16916(.A1(new_n16647_), .A2(new_n16643_), .ZN(new_n17919_));
  OAI21_X1   g16917(.A1(new_n16535_), .A2(new_n17919_), .B(new_n17259_), .ZN(new_n17920_));
  NAND2_X1   g16918(.A1(new_n17170_), .A2(new_n17176_), .ZN(new_n17921_));
  NAND2_X1   g16919(.A1(new_n17920_), .A2(new_n17921_), .ZN(new_n17922_));
  NOR2_X1    g16920(.A1(new_n17181_), .A2(new_n17147_), .ZN(new_n17923_));
  NAND2_X1   g16921(.A1(new_n17137_), .A2(new_n17142_), .ZN(new_n17924_));
  NAND2_X1   g16922(.A1(new_n17140_), .A2(new_n17146_), .ZN(new_n17925_));
  NAND2_X1   g16923(.A1(new_n17177_), .A2(new_n17179_), .ZN(new_n17926_));
  NAND2_X1   g16924(.A1(new_n17180_), .A2(new_n17162_), .ZN(new_n17927_));
  NAND4_X1   g16925(.A1(new_n17925_), .A2(new_n17927_), .A3(new_n17926_), .A4(new_n17924_), .ZN(new_n17928_));
  OAI21_X1   g16926(.A1(new_n17184_), .A2(new_n17923_), .B(new_n17928_), .ZN(new_n17929_));
  INV_X1     g16927(.I(new_n17928_), .ZN(new_n17930_));
  NOR3_X1    g16928(.A1(new_n17930_), .A2(new_n17916_), .A3(new_n17914_), .ZN(new_n17931_));
  AOI22_X1   g16929(.A1(new_n17922_), .A2(new_n17931_), .B1(new_n17929_), .B2(new_n17918_), .ZN(new_n17932_));
  NOR2_X1    g16930(.A1(new_n17906_), .A2(new_n17932_), .ZN(new_n17933_));
  NAND2_X1   g16931(.A1(new_n17881_), .A2(new_n17887_), .ZN(new_n17934_));
  OAI21_X1   g16932(.A1(new_n17878_), .A2(new_n17879_), .B(new_n17902_), .ZN(new_n17935_));
  NAND2_X1   g16933(.A1(new_n17904_), .A2(new_n17903_), .ZN(new_n17936_));
  NOR3_X1    g16934(.A1(new_n17897_), .A2(new_n17900_), .A3(new_n17886_), .ZN(new_n17937_));
  AOI22_X1   g16935(.A1(new_n17935_), .A2(new_n17936_), .B1(new_n17934_), .B2(new_n17937_), .ZN(new_n17938_));
  NOR2_X1    g16936(.A1(new_n17184_), .A2(new_n17923_), .ZN(new_n17939_));
  AOI21_X1   g16937(.A1(new_n17920_), .A2(new_n17921_), .B(new_n17930_), .ZN(new_n17940_));
  INV_X1     g16938(.I(new_n17914_), .ZN(new_n17941_));
  NAND2_X1   g16939(.A1(new_n17913_), .A2(new_n17909_), .ZN(new_n17942_));
  NAND3_X1   g16940(.A1(new_n17941_), .A2(new_n17942_), .A3(new_n17928_), .ZN(new_n17943_));
  OAI22_X1   g16941(.A1(new_n17940_), .A2(new_n17917_), .B1(new_n17939_), .B2(new_n17943_), .ZN(new_n17944_));
  NOR2_X1    g16942(.A1(new_n17938_), .A2(new_n17944_), .ZN(new_n17945_));
  OAI22_X1   g16943(.A1(new_n17945_), .A2(new_n17933_), .B1(new_n17877_), .B2(new_n17876_), .ZN(new_n17946_));
  NAND2_X1   g16944(.A1(new_n17263_), .A2(new_n17257_), .ZN(new_n17947_));
  OAI22_X1   g16945(.A1(new_n17270_), .A2(new_n17269_), .B1(new_n17263_), .B2(new_n17257_), .ZN(new_n17948_));
  NAND2_X1   g16946(.A1(new_n17938_), .A2(new_n17944_), .ZN(new_n17949_));
  NAND2_X1   g16947(.A1(new_n17906_), .A2(new_n17932_), .ZN(new_n17950_));
  NAND4_X1   g16948(.A1(new_n17948_), .A2(new_n17949_), .A3(new_n17950_), .A4(new_n17947_), .ZN(new_n17951_));
  NAND2_X1   g16949(.A1(new_n17951_), .A2(new_n17946_), .ZN(new_n17952_));
  OAI22_X1   g16950(.A1(new_n17108_), .A2(new_n17111_), .B1(new_n17032_), .B2(new_n17037_), .ZN(new_n17953_));
  OAI21_X1   g16951(.A1(new_n16967_), .A2(new_n16966_), .B(new_n17953_), .ZN(new_n17954_));
  NAND2_X1   g16952(.A1(new_n17112_), .A2(new_n17038_), .ZN(new_n17955_));
  NAND2_X1   g16953(.A1(new_n17003_), .A2(new_n17001_), .ZN(new_n17956_));
  NOR2_X1    g16954(.A1(new_n17003_), .A2(new_n17001_), .ZN(new_n17957_));
  AOI21_X1   g16955(.A1(new_n17014_), .A2(new_n17956_), .B(new_n17957_), .ZN(new_n17958_));
  NAND2_X1   g16956(.A1(new_n16981_), .A2(new_n16972_), .ZN(new_n17959_));
  NOR2_X1    g16957(.A1(new_n16981_), .A2(new_n16972_), .ZN(new_n17960_));
  AOI21_X1   g16958(.A1(new_n17023_), .A2(new_n17959_), .B(new_n17960_), .ZN(new_n17961_));
  INV_X1     g16959(.I(new_n17961_), .ZN(new_n17962_));
  NOR2_X1    g16960(.A1(new_n17962_), .A2(new_n17958_), .ZN(new_n17963_));
  INV_X1     g16961(.I(new_n17958_), .ZN(new_n17964_));
  NOR2_X1    g16962(.A1(new_n17964_), .A2(new_n17961_), .ZN(new_n17965_));
  NOR2_X1    g16963(.A1(new_n17965_), .A2(new_n17963_), .ZN(new_n17966_));
  NOR2_X1    g16964(.A1(new_n17019_), .A2(new_n17025_), .ZN(new_n17967_));
  AOI21_X1   g16965(.A1(new_n16969_), .A2(new_n16968_), .B(new_n17967_), .ZN(new_n17968_));
  NOR2_X1    g16966(.A1(new_n16780_), .A2(new_n16776_), .ZN(new_n17969_));
  OAI21_X1   g16967(.A1(new_n16683_), .A2(new_n17969_), .B(new_n16968_), .ZN(new_n17970_));
  INV_X1     g16968(.I(new_n17967_), .ZN(new_n17971_));
  NAND2_X1   g16969(.A1(new_n17021_), .A2(new_n17023_), .ZN(new_n17972_));
  NAND2_X1   g16970(.A1(new_n17024_), .A2(new_n16985_), .ZN(new_n17973_));
  NAND2_X1   g16971(.A1(new_n17014_), .A2(new_n17009_), .ZN(new_n17974_));
  NAND2_X1   g16972(.A1(new_n17018_), .A2(new_n17011_), .ZN(new_n17975_));
  NAND4_X1   g16973(.A1(new_n17973_), .A2(new_n17975_), .A3(new_n17974_), .A4(new_n17972_), .ZN(new_n17976_));
  INV_X1     g16974(.I(new_n17976_), .ZN(new_n17977_));
  AOI21_X1   g16975(.A1(new_n17970_), .A2(new_n17971_), .B(new_n17977_), .ZN(new_n17978_));
  NAND2_X1   g16976(.A1(new_n17964_), .A2(new_n17961_), .ZN(new_n17979_));
  NAND2_X1   g16977(.A1(new_n17962_), .A2(new_n17958_), .ZN(new_n17980_));
  NAND3_X1   g16978(.A1(new_n17979_), .A2(new_n17980_), .A3(new_n17976_), .ZN(new_n17981_));
  OAI22_X1   g16979(.A1(new_n17978_), .A2(new_n17966_), .B1(new_n17968_), .B2(new_n17981_), .ZN(new_n17982_));
  NAND2_X1   g16980(.A1(new_n17049_), .A2(new_n17047_), .ZN(new_n17983_));
  NOR2_X1    g16981(.A1(new_n17049_), .A2(new_n17047_), .ZN(new_n17984_));
  AOI21_X1   g16982(.A1(new_n17059_), .A2(new_n17983_), .B(new_n17984_), .ZN(new_n17985_));
  NAND4_X1   g16983(.A1(new_n17071_), .A2(new_n17067_), .A3(new_n17069_), .A4(new_n17065_), .ZN(new_n17986_));
  AOI22_X1   g16984(.A1(new_n17065_), .A2(new_n17067_), .B1(new_n17071_), .B2(new_n17069_), .ZN(new_n17987_));
  AOI21_X1   g16985(.A1(new_n17092_), .A2(new_n17986_), .B(new_n17987_), .ZN(new_n17988_));
  INV_X1     g16986(.I(new_n17988_), .ZN(new_n17989_));
  NOR2_X1    g16987(.A1(new_n17989_), .A2(new_n17985_), .ZN(new_n17990_));
  INV_X1     g16988(.I(new_n17985_), .ZN(new_n17991_));
  NOR2_X1    g16989(.A1(new_n17991_), .A2(new_n17988_), .ZN(new_n17992_));
  NOR2_X1    g16990(.A1(new_n17990_), .A2(new_n17992_), .ZN(new_n17993_));
  INV_X1     g16991(.I(new_n17993_), .ZN(new_n17994_));
  NAND2_X1   g16992(.A1(new_n17090_), .A2(new_n17084_), .ZN(new_n17995_));
  NAND2_X1   g16993(.A1(new_n17110_), .A2(new_n17995_), .ZN(new_n17996_));
  NOR2_X1    g16994(.A1(new_n17064_), .A2(new_n17094_), .ZN(new_n17997_));
  NAND2_X1   g16995(.A1(new_n17054_), .A2(new_n17059_), .ZN(new_n17998_));
  NAND2_X1   g16996(.A1(new_n17063_), .A2(new_n17056_), .ZN(new_n17999_));
  NAND2_X1   g16997(.A1(new_n17092_), .A2(new_n17075_), .ZN(new_n18000_));
  NAND2_X1   g16998(.A1(new_n17093_), .A2(new_n17091_), .ZN(new_n18001_));
  NAND4_X1   g16999(.A1(new_n17999_), .A2(new_n18001_), .A3(new_n17998_), .A4(new_n18000_), .ZN(new_n18002_));
  OAI21_X1   g17000(.A1(new_n17097_), .A2(new_n17997_), .B(new_n18002_), .ZN(new_n18003_));
  INV_X1     g17001(.I(new_n18002_), .ZN(new_n18004_));
  NOR3_X1    g17002(.A1(new_n18004_), .A2(new_n17992_), .A3(new_n17990_), .ZN(new_n18005_));
  AOI22_X1   g17003(.A1(new_n17994_), .A2(new_n18003_), .B1(new_n18005_), .B2(new_n17996_), .ZN(new_n18006_));
  NAND2_X1   g17004(.A1(new_n18006_), .A2(new_n17982_), .ZN(new_n18007_));
  INV_X1     g17005(.I(new_n17966_), .ZN(new_n18008_));
  NAND2_X1   g17006(.A1(new_n17970_), .A2(new_n17971_), .ZN(new_n18009_));
  NOR2_X1    g17007(.A1(new_n17034_), .A2(new_n17033_), .ZN(new_n18010_));
  OAI21_X1   g17008(.A1(new_n18010_), .A2(new_n17967_), .B(new_n17976_), .ZN(new_n18011_));
  NOR3_X1    g17009(.A1(new_n17977_), .A2(new_n17963_), .A3(new_n17965_), .ZN(new_n18012_));
  AOI22_X1   g17010(.A1(new_n18011_), .A2(new_n18008_), .B1(new_n18009_), .B2(new_n18012_), .ZN(new_n18013_));
  NOR2_X1    g17011(.A1(new_n17097_), .A2(new_n17997_), .ZN(new_n18014_));
  AOI21_X1   g17012(.A1(new_n17110_), .A2(new_n17995_), .B(new_n18004_), .ZN(new_n18015_));
  NAND2_X1   g17013(.A1(new_n17991_), .A2(new_n17988_), .ZN(new_n18016_));
  NAND2_X1   g17014(.A1(new_n17989_), .A2(new_n17985_), .ZN(new_n18017_));
  NAND3_X1   g17015(.A1(new_n18002_), .A2(new_n18017_), .A3(new_n18016_), .ZN(new_n18018_));
  OAI22_X1   g17016(.A1(new_n18015_), .A2(new_n17993_), .B1(new_n18014_), .B2(new_n18018_), .ZN(new_n18019_));
  NAND2_X1   g17017(.A1(new_n18013_), .A2(new_n18019_), .ZN(new_n18020_));
  AOI22_X1   g17018(.A1(new_n17954_), .A2(new_n17955_), .B1(new_n18020_), .B2(new_n18007_), .ZN(new_n18021_));
  AOI22_X1   g17019(.A1(new_n17116_), .A2(new_n17115_), .B1(new_n17105_), .B2(new_n17101_), .ZN(new_n18022_));
  NOR2_X1    g17020(.A1(new_n17101_), .A2(new_n17105_), .ZN(new_n18023_));
  NOR2_X1    g17021(.A1(new_n18013_), .A2(new_n18019_), .ZN(new_n18024_));
  NOR2_X1    g17022(.A1(new_n18006_), .A2(new_n17982_), .ZN(new_n18025_));
  NOR4_X1    g17023(.A1(new_n18022_), .A2(new_n18024_), .A3(new_n18025_), .A4(new_n18023_), .ZN(new_n18026_));
  NOR2_X1    g17024(.A1(new_n18021_), .A2(new_n18026_), .ZN(new_n18027_));
  NAND2_X1   g17025(.A1(new_n17952_), .A2(new_n18027_), .ZN(new_n18028_));
  AOI22_X1   g17026(.A1(new_n17948_), .A2(new_n17947_), .B1(new_n17949_), .B2(new_n17950_), .ZN(new_n18029_));
  NOR4_X1    g17027(.A1(new_n17945_), .A2(new_n17933_), .A3(new_n17877_), .A4(new_n17876_), .ZN(new_n18030_));
  NOR2_X1    g17028(.A1(new_n18029_), .A2(new_n18030_), .ZN(new_n18031_));
  OAI22_X1   g17029(.A1(new_n18022_), .A2(new_n18023_), .B1(new_n18024_), .B2(new_n18025_), .ZN(new_n18032_));
  NAND4_X1   g17030(.A1(new_n17954_), .A2(new_n18020_), .A3(new_n18007_), .A4(new_n17955_), .ZN(new_n18033_));
  NAND2_X1   g17031(.A1(new_n18032_), .A2(new_n18033_), .ZN(new_n18034_));
  NAND2_X1   g17032(.A1(new_n18031_), .A2(new_n18034_), .ZN(new_n18035_));
  AOI22_X1   g17033(.A1(new_n18028_), .A2(new_n18035_), .B1(new_n17874_), .B2(new_n17875_), .ZN(new_n18036_));
  AOI22_X1   g17034(.A1(new_n17286_), .A2(new_n17285_), .B1(new_n17282_), .B2(new_n17120_), .ZN(new_n18037_));
  NOR2_X1    g17035(.A1(new_n17282_), .A2(new_n17120_), .ZN(new_n18038_));
  NOR2_X1    g17036(.A1(new_n18031_), .A2(new_n18034_), .ZN(new_n18039_));
  NOR2_X1    g17037(.A1(new_n17952_), .A2(new_n18027_), .ZN(new_n18040_));
  NOR4_X1    g17038(.A1(new_n18040_), .A2(new_n18039_), .A3(new_n18037_), .A4(new_n18038_), .ZN(new_n18041_));
  NOR2_X1    g17039(.A1(new_n18036_), .A2(new_n18041_), .ZN(new_n18042_));
  NAND2_X1   g17040(.A1(new_n17873_), .A2(new_n18042_), .ZN(new_n18043_));
  NAND2_X1   g17041(.A1(new_n17451_), .A2(new_n17622_), .ZN(new_n18044_));
  OAI22_X1   g17042(.A1(new_n17293_), .A2(new_n17292_), .B1(new_n17451_), .B2(new_n17622_), .ZN(new_n18045_));
  AOI22_X1   g17043(.A1(new_n17871_), .A2(new_n17870_), .B1(new_n18044_), .B2(new_n18045_), .ZN(new_n18046_));
  NOR4_X1    g17044(.A1(new_n17860_), .A2(new_n17867_), .A3(new_n17703_), .A4(new_n17706_), .ZN(new_n18047_));
  NOR2_X1    g17045(.A1(new_n18046_), .A2(new_n18047_), .ZN(new_n18048_));
  OAI22_X1   g17046(.A1(new_n18040_), .A2(new_n18039_), .B1(new_n18037_), .B2(new_n18038_), .ZN(new_n18049_));
  NAND4_X1   g17047(.A1(new_n18028_), .A2(new_n18035_), .A3(new_n17874_), .A4(new_n17875_), .ZN(new_n18050_));
  NAND2_X1   g17048(.A1(new_n18049_), .A2(new_n18050_), .ZN(new_n18051_));
  NAND2_X1   g17049(.A1(new_n18048_), .A2(new_n18051_), .ZN(new_n18052_));
  AOI21_X1   g17050(.A1(new_n18043_), .A2(new_n18052_), .B(new_n17702_), .ZN(new_n18053_));
  AOI22_X1   g17051(.A1(new_n17631_), .A2(new_n17632_), .B1(new_n17624_), .B2(new_n17628_), .ZN(new_n18054_));
  NAND4_X1   g17052(.A1(new_n17631_), .A2(new_n17632_), .A3(new_n17624_), .A4(new_n17628_), .ZN(new_n18055_));
  OAI21_X1   g17053(.A1(new_n17643_), .A2(new_n18054_), .B(new_n18055_), .ZN(new_n18056_));
  NOR2_X1    g17054(.A1(new_n18048_), .A2(new_n18051_), .ZN(new_n18057_));
  NOR2_X1    g17055(.A1(new_n17873_), .A2(new_n18042_), .ZN(new_n18058_));
  NOR3_X1    g17056(.A1(new_n18056_), .A2(new_n18058_), .A3(new_n18057_), .ZN(new_n18059_));
  NOR2_X1    g17057(.A1(new_n18059_), .A2(new_n18053_), .ZN(new_n18060_));
  AOI21_X1   g17058(.A1(new_n11856_), .A2(new_n11855_), .B(new_n11616_), .ZN(new_n18061_));
  NAND3_X1   g17059(.A1(new_n11856_), .A2(new_n11855_), .A3(new_n11616_), .ZN(new_n18062_));
  OAI21_X1   g17060(.A1(new_n11461_), .A2(new_n18061_), .B(new_n18062_), .ZN(new_n18063_));
  NAND2_X1   g17061(.A1(new_n11628_), .A2(new_n11630_), .ZN(new_n18064_));
  NOR2_X1    g17062(.A1(new_n11628_), .A2(new_n11630_), .ZN(new_n18065_));
  AOI21_X1   g17063(.A1(new_n11636_), .A2(new_n18064_), .B(new_n18065_), .ZN(new_n18066_));
  NOR2_X1    g17064(.A1(new_n11645_), .A2(new_n11650_), .ZN(new_n18067_));
  NAND2_X1   g17065(.A1(new_n11645_), .A2(new_n11650_), .ZN(new_n18068_));
  OAI21_X1   g17066(.A1(new_n11660_), .A2(new_n18067_), .B(new_n18068_), .ZN(new_n18069_));
  NOR2_X1    g17067(.A1(new_n18066_), .A2(new_n18069_), .ZN(new_n18070_));
  NAND2_X1   g17068(.A1(new_n18066_), .A2(new_n18069_), .ZN(new_n18071_));
  INV_X1     g17069(.I(new_n18071_), .ZN(new_n18072_));
  NOR2_X1    g17070(.A1(new_n18072_), .A2(new_n18070_), .ZN(new_n18073_));
  NOR2_X1    g17071(.A1(new_n11672_), .A2(new_n11641_), .ZN(new_n18074_));
  NOR2_X1    g17072(.A1(new_n11677_), .A2(new_n18074_), .ZN(new_n18075_));
  AOI22_X1   g17073(.A1(new_n11634_), .A2(new_n11635_), .B1(new_n11629_), .B2(new_n11631_), .ZN(new_n18076_));
  INV_X1     g17074(.I(new_n11667_), .ZN(new_n18077_));
  NOR2_X1    g17075(.A1(new_n11654_), .A2(new_n11660_), .ZN(new_n18078_));
  NOR2_X1    g17076(.A1(new_n11663_), .A2(new_n11657_), .ZN(new_n18079_));
  NOR4_X1    g17077(.A1(new_n18079_), .A2(new_n18077_), .A3(new_n18078_), .A4(new_n18076_), .ZN(new_n18080_));
  NOR2_X1    g17078(.A1(new_n18075_), .A2(new_n18080_), .ZN(new_n18081_));
  INV_X1     g17079(.I(new_n18070_), .ZN(new_n18082_));
  INV_X1     g17080(.I(new_n18080_), .ZN(new_n18083_));
  NAND3_X1   g17081(.A1(new_n18083_), .A2(new_n18082_), .A3(new_n18071_), .ZN(new_n18084_));
  OAI22_X1   g17082(.A1(new_n18081_), .A2(new_n18073_), .B1(new_n18075_), .B2(new_n18084_), .ZN(new_n18085_));
  NOR2_X1    g17083(.A1(new_n11815_), .A2(new_n11813_), .ZN(new_n18086_));
  NOR2_X1    g17084(.A1(new_n3784_), .A2(new_n3776_), .ZN(new_n18087_));
  OAI21_X1   g17085(.A1(new_n18087_), .A2(new_n3869_), .B(new_n3881_), .ZN(new_n18088_));
  AOI22_X1   g17086(.A1(new_n18088_), .A2(new_n11830_), .B1(new_n11815_), .B2(new_n11813_), .ZN(new_n18089_));
  NAND2_X1   g17087(.A1(new_n11759_), .A2(new_n11806_), .ZN(new_n18090_));
  AOI21_X1   g17088(.A1(new_n11799_), .A2(new_n11792_), .B(new_n11771_), .ZN(new_n18091_));
  OAI21_X1   g17089(.A1(new_n11810_), .A2(new_n18091_), .B(new_n11800_), .ZN(new_n18092_));
  AOI22_X1   g17090(.A1(new_n11797_), .A2(new_n11798_), .B1(new_n11774_), .B2(new_n11786_), .ZN(new_n18093_));
  NOR2_X1    g17091(.A1(new_n11774_), .A2(new_n11786_), .ZN(new_n18094_));
  NOR3_X1    g17092(.A1(new_n18093_), .A2(new_n11765_), .A3(new_n18094_), .ZN(new_n18095_));
  OAI22_X1   g17093(.A1(new_n11790_), .A2(new_n11791_), .B1(new_n11783_), .B2(new_n11778_), .ZN(new_n18096_));
  INV_X1     g17094(.I(new_n18094_), .ZN(new_n18097_));
  AOI21_X1   g17095(.A1(new_n18096_), .A2(new_n18097_), .B(new_n11801_), .ZN(new_n18098_));
  NOR2_X1    g17096(.A1(new_n18095_), .A2(new_n18098_), .ZN(new_n18099_));
  OAI21_X1   g17097(.A1(new_n18098_), .A2(new_n18095_), .B(new_n11800_), .ZN(new_n18100_));
  INV_X1     g17098(.I(new_n18100_), .ZN(new_n18101_));
  AOI22_X1   g17099(.A1(new_n18101_), .A2(new_n18090_), .B1(new_n18092_), .B2(new_n18099_), .ZN(new_n18102_));
  NAND3_X1   g17100(.A1(new_n11693_), .A2(new_n11686_), .A3(new_n11688_), .ZN(new_n18103_));
  NAND2_X1   g17101(.A1(new_n11705_), .A2(new_n18103_), .ZN(new_n18104_));
  NAND2_X1   g17102(.A1(new_n11689_), .A2(new_n11698_), .ZN(new_n18105_));
  NAND2_X1   g17103(.A1(new_n18104_), .A2(new_n18105_), .ZN(new_n18106_));
  OAI21_X1   g17104(.A1(new_n11723_), .A2(new_n11719_), .B(new_n11748_), .ZN(new_n18107_));
  NAND2_X1   g17105(.A1(new_n11719_), .A2(new_n11723_), .ZN(new_n18108_));
  NAND3_X1   g17106(.A1(new_n18106_), .A2(new_n18107_), .A3(new_n18108_), .ZN(new_n18109_));
  NOR2_X1    g17107(.A1(new_n11719_), .A2(new_n11723_), .ZN(new_n18110_));
  OAI21_X1   g17108(.A1(new_n11734_), .A2(new_n18110_), .B(new_n18108_), .ZN(new_n18111_));
  NAND3_X1   g17109(.A1(new_n18111_), .A2(new_n18104_), .A3(new_n18105_), .ZN(new_n18112_));
  NAND2_X1   g17110(.A1(new_n18109_), .A2(new_n18112_), .ZN(new_n18113_));
  INV_X1     g17111(.I(new_n18113_), .ZN(new_n18114_));
  AOI22_X1   g17112(.A1(new_n11753_), .A2(new_n11682_), .B1(new_n11745_), .B2(new_n11739_), .ZN(new_n18115_));
  NAND2_X1   g17113(.A1(new_n11739_), .A2(new_n11745_), .ZN(new_n18116_));
  NAND2_X1   g17114(.A1(new_n11700_), .A2(new_n11705_), .ZN(new_n18117_));
  INV_X1     g17115(.I(new_n18117_), .ZN(new_n18118_));
  NOR2_X1    g17116(.A1(new_n11744_), .A2(new_n11742_), .ZN(new_n18119_));
  NOR2_X1    g17117(.A1(new_n11729_), .A2(new_n11734_), .ZN(new_n18120_));
  NOR2_X1    g17118(.A1(new_n11738_), .A2(new_n11731_), .ZN(new_n18121_));
  NOR4_X1    g17119(.A1(new_n18118_), .A2(new_n18120_), .A3(new_n18121_), .A4(new_n18119_), .ZN(new_n18122_));
  AOI21_X1   g17120(.A1(new_n11826_), .A2(new_n18116_), .B(new_n18122_), .ZN(new_n18123_));
  NAND2_X1   g17121(.A1(new_n11709_), .A2(new_n11703_), .ZN(new_n18124_));
  NAND2_X1   g17122(.A1(new_n11746_), .A2(new_n11748_), .ZN(new_n18125_));
  NAND2_X1   g17123(.A1(new_n11749_), .A2(new_n11747_), .ZN(new_n18126_));
  NAND4_X1   g17124(.A1(new_n18126_), .A2(new_n18125_), .A3(new_n18124_), .A4(new_n18117_), .ZN(new_n18127_));
  NAND3_X1   g17125(.A1(new_n18109_), .A2(new_n18127_), .A3(new_n18112_), .ZN(new_n18128_));
  OAI22_X1   g17126(.A1(new_n18114_), .A2(new_n18123_), .B1(new_n18115_), .B2(new_n18128_), .ZN(new_n18129_));
  NOR2_X1    g17127(.A1(new_n18129_), .A2(new_n18102_), .ZN(new_n18130_));
  NOR2_X1    g17128(.A1(new_n11810_), .A2(new_n18091_), .ZN(new_n18131_));
  INV_X1     g17129(.I(new_n11800_), .ZN(new_n18132_));
  AOI21_X1   g17130(.A1(new_n11759_), .A2(new_n11806_), .B(new_n18132_), .ZN(new_n18133_));
  INV_X1     g17131(.I(new_n18099_), .ZN(new_n18134_));
  OAI22_X1   g17132(.A1(new_n18133_), .A2(new_n18134_), .B1(new_n18131_), .B2(new_n18100_), .ZN(new_n18135_));
  OAI21_X1   g17133(.A1(new_n18115_), .A2(new_n18122_), .B(new_n18113_), .ZN(new_n18136_));
  NOR2_X1    g17134(.A1(new_n18115_), .A2(new_n18128_), .ZN(new_n18137_));
  INV_X1     g17135(.I(new_n18137_), .ZN(new_n18138_));
  AOI21_X1   g17136(.A1(new_n18138_), .A2(new_n18136_), .B(new_n18135_), .ZN(new_n18139_));
  OAI22_X1   g17137(.A1(new_n18089_), .A2(new_n18086_), .B1(new_n18139_), .B2(new_n18130_), .ZN(new_n18140_));
  NAND2_X1   g17138(.A1(new_n11828_), .A2(new_n11818_), .ZN(new_n18141_));
  NAND2_X1   g17139(.A1(new_n3871_), .A2(new_n3872_), .ZN(new_n18142_));
  AOI21_X1   g17140(.A1(new_n18142_), .A2(new_n3875_), .B(new_n3675_), .ZN(new_n18143_));
  OAI22_X1   g17141(.A1(new_n18143_), .A2(new_n11820_), .B1(new_n11828_), .B2(new_n11818_), .ZN(new_n18144_));
  NAND3_X1   g17142(.A1(new_n18138_), .A2(new_n18135_), .A3(new_n18136_), .ZN(new_n18145_));
  NAND2_X1   g17143(.A1(new_n18129_), .A2(new_n18102_), .ZN(new_n18146_));
  NAND4_X1   g17144(.A1(new_n18144_), .A2(new_n18145_), .A3(new_n18146_), .A4(new_n18141_), .ZN(new_n18147_));
  AOI21_X1   g17145(.A1(new_n18140_), .A2(new_n18147_), .B(new_n18085_), .ZN(new_n18148_));
  INV_X1     g17146(.I(new_n18073_), .ZN(new_n18149_));
  NAND2_X1   g17147(.A1(new_n11668_), .A2(new_n11664_), .ZN(new_n18150_));
  NAND2_X1   g17148(.A1(new_n11619_), .A2(new_n18150_), .ZN(new_n18151_));
  NAND2_X1   g17149(.A1(new_n18151_), .A2(new_n18083_), .ZN(new_n18152_));
  NOR3_X1    g17150(.A1(new_n18072_), .A2(new_n18080_), .A3(new_n18070_), .ZN(new_n18153_));
  AOI22_X1   g17151(.A1(new_n18152_), .A2(new_n18149_), .B1(new_n18151_), .B2(new_n18153_), .ZN(new_n18154_));
  AOI22_X1   g17152(.A1(new_n18144_), .A2(new_n18141_), .B1(new_n18145_), .B2(new_n18146_), .ZN(new_n18155_));
  NOR4_X1    g17153(.A1(new_n18089_), .A2(new_n18086_), .A3(new_n18139_), .A4(new_n18130_), .ZN(new_n18156_));
  NOR3_X1    g17154(.A1(new_n18156_), .A2(new_n18155_), .A3(new_n18154_), .ZN(new_n18157_));
  AOI21_X1   g17155(.A1(new_n11833_), .A2(new_n11823_), .B(new_n11837_), .ZN(new_n18158_));
  NAND3_X1   g17156(.A1(new_n11833_), .A2(new_n11823_), .A3(new_n11837_), .ZN(new_n18159_));
  OAI21_X1   g17157(.A1(new_n11849_), .A2(new_n18158_), .B(new_n18159_), .ZN(new_n18160_));
  NOR3_X1    g17158(.A1(new_n18160_), .A2(new_n18148_), .A3(new_n18157_), .ZN(new_n18161_));
  OAI21_X1   g17159(.A1(new_n18156_), .A2(new_n18155_), .B(new_n18154_), .ZN(new_n18162_));
  NAND3_X1   g17160(.A1(new_n18140_), .A2(new_n18147_), .A3(new_n18085_), .ZN(new_n18163_));
  OAI21_X1   g17161(.A1(new_n11839_), .A2(new_n11838_), .B(new_n11681_), .ZN(new_n18164_));
  NAND2_X1   g17162(.A1(new_n18164_), .A2(new_n11843_), .ZN(new_n18165_));
  AOI22_X1   g17163(.A1(new_n18165_), .A2(new_n18159_), .B1(new_n18162_), .B2(new_n18163_), .ZN(new_n18166_));
  NOR2_X1    g17164(.A1(new_n11529_), .A2(new_n11607_), .ZN(new_n18167_));
  NAND2_X1   g17165(.A1(new_n11529_), .A2(new_n11607_), .ZN(new_n18168_));
  AOI21_X1   g17166(.A1(new_n11612_), .A2(new_n18168_), .B(new_n18167_), .ZN(new_n18169_));
  OAI22_X1   g17167(.A1(new_n11543_), .A2(new_n11546_), .B1(new_n11536_), .B2(new_n11551_), .ZN(new_n18170_));
  NAND2_X1   g17168(.A1(new_n11551_), .A2(new_n11536_), .ZN(new_n18171_));
  NAND2_X1   g17169(.A1(new_n18170_), .A2(new_n18171_), .ZN(new_n18172_));
  NOR2_X1    g17170(.A1(new_n11558_), .A2(new_n11569_), .ZN(new_n18173_));
  NOR2_X1    g17171(.A1(new_n11590_), .A2(new_n18173_), .ZN(new_n18174_));
  AOI21_X1   g17172(.A1(new_n11558_), .A2(new_n11569_), .B(new_n18174_), .ZN(new_n18175_));
  NAND2_X1   g17173(.A1(new_n18175_), .A2(new_n18172_), .ZN(new_n18176_));
  AND2_X2    g17174(.A1(new_n18170_), .A2(new_n18171_), .Z(new_n18177_));
  INV_X1     g17175(.I(new_n18174_), .ZN(new_n18178_));
  NAND2_X1   g17176(.A1(new_n11558_), .A2(new_n11569_), .ZN(new_n18179_));
  NAND2_X1   g17177(.A1(new_n18178_), .A2(new_n18179_), .ZN(new_n18180_));
  NAND2_X1   g17178(.A1(new_n18177_), .A2(new_n18180_), .ZN(new_n18181_));
  NAND2_X1   g17179(.A1(new_n18181_), .A2(new_n18176_), .ZN(new_n18182_));
  NOR2_X1    g17180(.A1(new_n11596_), .A2(new_n11595_), .ZN(new_n18183_));
  NOR2_X1    g17181(.A1(new_n11587_), .A2(new_n11581_), .ZN(new_n18184_));
  NAND2_X1   g17182(.A1(new_n11585_), .A2(new_n11583_), .ZN(new_n18185_));
  NAND2_X1   g17183(.A1(new_n11586_), .A2(new_n11584_), .ZN(new_n18186_));
  NAND2_X1   g17184(.A1(new_n11571_), .A2(new_n11576_), .ZN(new_n18187_));
  NAND2_X1   g17185(.A1(new_n11580_), .A2(new_n11573_), .ZN(new_n18188_));
  NAND4_X1   g17186(.A1(new_n18185_), .A2(new_n18186_), .A3(new_n18187_), .A4(new_n18188_), .ZN(new_n18189_));
  OAI21_X1   g17187(.A1(new_n18183_), .A2(new_n18184_), .B(new_n18189_), .ZN(new_n18190_));
  NAND2_X1   g17188(.A1(new_n18190_), .A2(new_n18182_), .ZN(new_n18191_));
  OAI22_X1   g17189(.A1(new_n11596_), .A2(new_n11595_), .B1(new_n11587_), .B2(new_n11581_), .ZN(new_n18192_));
  NOR2_X1    g17190(.A1(new_n18177_), .A2(new_n18180_), .ZN(new_n18193_));
  NOR2_X1    g17191(.A1(new_n18175_), .A2(new_n18172_), .ZN(new_n18194_));
  INV_X1     g17192(.I(new_n18189_), .ZN(new_n18195_));
  NOR3_X1    g17193(.A1(new_n18193_), .A2(new_n18194_), .A3(new_n18195_), .ZN(new_n18196_));
  NAND2_X1   g17194(.A1(new_n18196_), .A2(new_n18192_), .ZN(new_n18197_));
  NAND2_X1   g17195(.A1(new_n18197_), .A2(new_n18191_), .ZN(new_n18198_));
  INV_X1     g17196(.I(new_n11474_), .ZN(new_n18199_));
  NOR2_X1    g17197(.A1(new_n18199_), .A2(new_n11470_), .ZN(new_n18200_));
  NAND2_X1   g17198(.A1(new_n18199_), .A2(new_n11470_), .ZN(new_n18201_));
  OAI21_X1   g17199(.A1(new_n11517_), .A2(new_n18200_), .B(new_n18201_), .ZN(new_n18202_));
  AOI21_X1   g17200(.A1(new_n4021_), .A2(new_n11506_), .B(new_n11510_), .ZN(new_n18203_));
  NOR2_X1    g17201(.A1(new_n11491_), .A2(new_n11499_), .ZN(new_n18204_));
  NAND2_X1   g17202(.A1(new_n11491_), .A2(new_n11499_), .ZN(new_n18205_));
  OAI21_X1   g17203(.A1(new_n18203_), .A2(new_n18204_), .B(new_n18205_), .ZN(new_n18206_));
  INV_X1     g17204(.I(new_n18206_), .ZN(new_n18207_));
  NAND2_X1   g17205(.A1(new_n18207_), .A2(new_n18202_), .ZN(new_n18208_));
  INV_X1     g17206(.I(new_n18202_), .ZN(new_n18209_));
  NAND2_X1   g17207(.A1(new_n18209_), .A2(new_n18206_), .ZN(new_n18210_));
  NAND2_X1   g17208(.A1(new_n18210_), .A2(new_n18208_), .ZN(new_n18211_));
  NAND2_X1   g17209(.A1(new_n11525_), .A2(new_n11523_), .ZN(new_n18212_));
  NOR2_X1    g17210(.A1(new_n11486_), .A2(new_n11520_), .ZN(new_n18213_));
  INV_X1     g17211(.I(new_n18213_), .ZN(new_n18214_));
  NAND2_X1   g17212(.A1(new_n18212_), .A2(new_n18214_), .ZN(new_n18215_));
  NOR2_X1    g17213(.A1(new_n11466_), .A2(new_n11465_), .ZN(new_n18216_));
  NOR2_X1    g17214(.A1(new_n11517_), .A2(new_n11515_), .ZN(new_n18217_));
  NOR2_X1    g17215(.A1(new_n11518_), .A2(new_n11516_), .ZN(new_n18218_));
  AOI22_X1   g17216(.A1(new_n11507_), .A2(new_n11503_), .B1(new_n11494_), .B2(new_n11500_), .ZN(new_n18219_));
  NOR2_X1    g17217(.A1(new_n11502_), .A2(new_n4064_), .ZN(new_n18220_));
  NOR3_X1    g17218(.A1(new_n11501_), .A2(new_n18220_), .A3(new_n11510_), .ZN(new_n18221_));
  NOR4_X1    g17219(.A1(new_n18217_), .A2(new_n18218_), .A3(new_n18221_), .A4(new_n18219_), .ZN(new_n18222_));
  INV_X1     g17220(.I(new_n18222_), .ZN(new_n18223_));
  OAI21_X1   g17221(.A1(new_n18216_), .A2(new_n18213_), .B(new_n18223_), .ZN(new_n18224_));
  NOR2_X1    g17222(.A1(new_n18211_), .A2(new_n18222_), .ZN(new_n18225_));
  AOI22_X1   g17223(.A1(new_n18225_), .A2(new_n18215_), .B1(new_n18224_), .B2(new_n18211_), .ZN(new_n18226_));
  NAND2_X1   g17224(.A1(new_n18198_), .A2(new_n18226_), .ZN(new_n18227_));
  AOI22_X1   g17225(.A1(new_n18196_), .A2(new_n18192_), .B1(new_n18190_), .B2(new_n18182_), .ZN(new_n18228_));
  INV_X1     g17226(.I(new_n18211_), .ZN(new_n18229_));
  NOR2_X1    g17227(.A1(new_n18216_), .A2(new_n18213_), .ZN(new_n18230_));
  AOI21_X1   g17228(.A1(new_n18212_), .A2(new_n18214_), .B(new_n18222_), .ZN(new_n18231_));
  NAND3_X1   g17229(.A1(new_n18223_), .A2(new_n18210_), .A3(new_n18208_), .ZN(new_n18232_));
  OAI22_X1   g17230(.A1(new_n18229_), .A2(new_n18231_), .B1(new_n18230_), .B2(new_n18232_), .ZN(new_n18233_));
  NAND2_X1   g17231(.A1(new_n18233_), .A2(new_n18228_), .ZN(new_n18234_));
  AOI21_X1   g17232(.A1(new_n18227_), .A2(new_n18234_), .B(new_n18169_), .ZN(new_n18235_));
  NAND2_X1   g17233(.A1(new_n11604_), .A2(new_n11600_), .ZN(new_n18236_));
  NOR2_X1    g17234(.A1(new_n11604_), .A2(new_n11600_), .ZN(new_n18237_));
  OAI21_X1   g17235(.A1(new_n11464_), .A2(new_n18237_), .B(new_n18236_), .ZN(new_n18238_));
  NOR2_X1    g17236(.A1(new_n18233_), .A2(new_n18228_), .ZN(new_n18239_));
  NOR2_X1    g17237(.A1(new_n18198_), .A2(new_n18226_), .ZN(new_n18240_));
  NOR3_X1    g17238(.A1(new_n18238_), .A2(new_n18240_), .A3(new_n18239_), .ZN(new_n18241_));
  NOR2_X1    g17239(.A1(new_n18235_), .A2(new_n18241_), .ZN(new_n18242_));
  NOR3_X1    g17240(.A1(new_n18166_), .A2(new_n18161_), .A3(new_n18242_), .ZN(new_n18243_));
  NOR2_X1    g17241(.A1(new_n11838_), .A2(new_n11681_), .ZN(new_n18244_));
  AOI22_X1   g17242(.A1(new_n18164_), .A2(new_n11843_), .B1(new_n18244_), .B2(new_n11833_), .ZN(new_n18245_));
  NAND3_X1   g17243(.A1(new_n18245_), .A2(new_n18162_), .A3(new_n18163_), .ZN(new_n18246_));
  OAI21_X1   g17244(.A1(new_n18148_), .A2(new_n18157_), .B(new_n18160_), .ZN(new_n18247_));
  OAI21_X1   g17245(.A1(new_n18239_), .A2(new_n18240_), .B(new_n18238_), .ZN(new_n18248_));
  NAND3_X1   g17246(.A1(new_n18169_), .A2(new_n18227_), .A3(new_n18234_), .ZN(new_n18249_));
  NAND2_X1   g17247(.A1(new_n18248_), .A2(new_n18249_), .ZN(new_n18250_));
  AOI21_X1   g17248(.A1(new_n18247_), .A2(new_n18246_), .B(new_n18250_), .ZN(new_n18251_));
  OAI21_X1   g17249(.A1(new_n18243_), .A2(new_n18251_), .B(new_n18063_), .ZN(new_n18252_));
  OAI21_X1   g17250(.A1(new_n11850_), .A2(new_n11844_), .B(new_n11854_), .ZN(new_n18253_));
  NOR2_X1    g17251(.A1(new_n11844_), .A2(new_n11854_), .ZN(new_n18254_));
  AOI22_X1   g17252(.A1(new_n11861_), .A2(new_n18253_), .B1(new_n11856_), .B2(new_n18254_), .ZN(new_n18255_));
  NAND3_X1   g17253(.A1(new_n18247_), .A2(new_n18246_), .A3(new_n18250_), .ZN(new_n18256_));
  OAI21_X1   g17254(.A1(new_n18166_), .A2(new_n18161_), .B(new_n18242_), .ZN(new_n18257_));
  NAND3_X1   g17255(.A1(new_n18255_), .A2(new_n18256_), .A3(new_n18257_), .ZN(new_n18258_));
  NAND2_X1   g17256(.A1(new_n18252_), .A2(new_n18258_), .ZN(new_n18259_));
  NOR4_X1    g17257(.A1(new_n11436_), .A2(new_n11445_), .A3(new_n11442_), .A4(new_n11446_), .ZN(new_n18260_));
  OAI21_X1   g17258(.A1(new_n10170_), .A2(new_n10668_), .B(new_n9669_), .ZN(new_n18261_));
  AOI22_X1   g17259(.A1(new_n18261_), .A2(new_n11453_), .B1(new_n11070_), .B2(new_n11450_), .ZN(new_n18262_));
  NAND2_X1   g17260(.A1(new_n11429_), .A2(new_n11425_), .ZN(new_n18263_));
  AOI21_X1   g17261(.A1(new_n9914_), .A2(new_n10163_), .B(new_n9671_), .ZN(new_n18264_));
  OAI22_X1   g17262(.A1(new_n18264_), .A2(new_n11071_), .B1(new_n11429_), .B2(new_n11425_), .ZN(new_n18265_));
  NOR2_X1    g17263(.A1(new_n11329_), .A2(new_n11417_), .ZN(new_n18266_));
  AOI22_X1   g17264(.A1(new_n11253_), .A2(new_n11252_), .B1(new_n11329_), .B2(new_n11417_), .ZN(new_n18267_));
  NAND2_X1   g17265(.A1(new_n11347_), .A2(new_n11335_), .ZN(new_n18268_));
  NOR2_X1    g17266(.A1(new_n11347_), .A2(new_n11335_), .ZN(new_n18269_));
  AOI21_X1   g17267(.A1(new_n11391_), .A2(new_n18268_), .B(new_n18269_), .ZN(new_n18270_));
  INV_X1     g17268(.I(new_n18270_), .ZN(new_n18271_));
  NAND2_X1   g17269(.A1(new_n11371_), .A2(new_n11367_), .ZN(new_n18272_));
  NOR2_X1    g17270(.A1(new_n11371_), .A2(new_n11367_), .ZN(new_n18273_));
  AOI21_X1   g17271(.A1(new_n11382_), .A2(new_n18272_), .B(new_n18273_), .ZN(new_n18274_));
  NAND2_X1   g17272(.A1(new_n18271_), .A2(new_n18274_), .ZN(new_n18275_));
  INV_X1     g17273(.I(new_n18274_), .ZN(new_n18276_));
  NAND2_X1   g17274(.A1(new_n18276_), .A2(new_n18270_), .ZN(new_n18277_));
  NAND2_X1   g17275(.A1(new_n18277_), .A2(new_n18275_), .ZN(new_n18278_));
  NAND2_X1   g17276(.A1(new_n11359_), .A2(new_n11398_), .ZN(new_n18279_));
  NAND2_X1   g17277(.A1(new_n11402_), .A2(new_n18279_), .ZN(new_n18280_));
  NAND2_X1   g17278(.A1(new_n11389_), .A2(new_n11391_), .ZN(new_n18281_));
  NAND2_X1   g17279(.A1(new_n11392_), .A2(new_n11390_), .ZN(new_n18282_));
  NAND2_X1   g17280(.A1(new_n11382_), .A2(new_n11377_), .ZN(new_n18283_));
  NAND2_X1   g17281(.A1(new_n11386_), .A2(new_n11379_), .ZN(new_n18284_));
  NAND4_X1   g17282(.A1(new_n18282_), .A2(new_n18281_), .A3(new_n18284_), .A4(new_n18283_), .ZN(new_n18285_));
  NAND2_X1   g17283(.A1(new_n18280_), .A2(new_n18285_), .ZN(new_n18286_));
  NAND3_X1   g17284(.A1(new_n18275_), .A2(new_n18277_), .A3(new_n18285_), .ZN(new_n18287_));
  INV_X1     g17285(.I(new_n18287_), .ZN(new_n18288_));
  AOI22_X1   g17286(.A1(new_n18286_), .A2(new_n18278_), .B1(new_n18288_), .B2(new_n18280_), .ZN(new_n18289_));
  NAND2_X1   g17287(.A1(new_n11267_), .A2(new_n11263_), .ZN(new_n18290_));
  NOR2_X1    g17288(.A1(new_n11267_), .A2(new_n11263_), .ZN(new_n18291_));
  AOI21_X1   g17289(.A1(new_n11277_), .A2(new_n18290_), .B(new_n18291_), .ZN(new_n18292_));
  NAND2_X1   g17290(.A1(new_n11286_), .A2(new_n11299_), .ZN(new_n18293_));
  NOR2_X1    g17291(.A1(new_n11286_), .A2(new_n11299_), .ZN(new_n18294_));
  AOI21_X1   g17292(.A1(new_n11320_), .A2(new_n18293_), .B(new_n18294_), .ZN(new_n18295_));
  INV_X1     g17293(.I(new_n18295_), .ZN(new_n18296_));
  NOR2_X1    g17294(.A1(new_n18296_), .A2(new_n18292_), .ZN(new_n18297_));
  INV_X1     g17295(.I(new_n18292_), .ZN(new_n18298_));
  NOR2_X1    g17296(.A1(new_n18298_), .A2(new_n18295_), .ZN(new_n18299_));
  NOR2_X1    g17297(.A1(new_n18297_), .A2(new_n18299_), .ZN(new_n18300_));
  NOR2_X1    g17298(.A1(new_n11282_), .A2(new_n11322_), .ZN(new_n18301_));
  AOI21_X1   g17299(.A1(new_n11254_), .A2(new_n11325_), .B(new_n18301_), .ZN(new_n18302_));
  INV_X1     g17300(.I(new_n18301_), .ZN(new_n18303_));
  NAND2_X1   g17301(.A1(new_n11272_), .A2(new_n11277_), .ZN(new_n18304_));
  NAND2_X1   g17302(.A1(new_n11281_), .A2(new_n11274_), .ZN(new_n18305_));
  NAND2_X1   g17303(.A1(new_n11320_), .A2(new_n11318_), .ZN(new_n18306_));
  NAND2_X1   g17304(.A1(new_n11321_), .A2(new_n11319_), .ZN(new_n18307_));
  NAND4_X1   g17305(.A1(new_n18305_), .A2(new_n18304_), .A3(new_n18307_), .A4(new_n18306_), .ZN(new_n18308_));
  INV_X1     g17306(.I(new_n18308_), .ZN(new_n18309_));
  AOI21_X1   g17307(.A1(new_n11410_), .A2(new_n18303_), .B(new_n18309_), .ZN(new_n18310_));
  NAND2_X1   g17308(.A1(new_n18298_), .A2(new_n18295_), .ZN(new_n18311_));
  NAND2_X1   g17309(.A1(new_n18296_), .A2(new_n18292_), .ZN(new_n18312_));
  NAND3_X1   g17310(.A1(new_n18311_), .A2(new_n18312_), .A3(new_n18308_), .ZN(new_n18313_));
  OAI22_X1   g17311(.A1(new_n18310_), .A2(new_n18300_), .B1(new_n18302_), .B2(new_n18313_), .ZN(new_n18314_));
  NOR2_X1    g17312(.A1(new_n18289_), .A2(new_n18314_), .ZN(new_n18315_));
  INV_X1     g17313(.I(new_n18278_), .ZN(new_n18316_));
  AOI22_X1   g17314(.A1(new_n11331_), .A2(new_n11330_), .B1(new_n11359_), .B2(new_n11398_), .ZN(new_n18317_));
  INV_X1     g17315(.I(new_n18285_), .ZN(new_n18318_));
  AOI21_X1   g17316(.A1(new_n11402_), .A2(new_n18279_), .B(new_n18318_), .ZN(new_n18319_));
  OAI22_X1   g17317(.A1(new_n18319_), .A2(new_n18316_), .B1(new_n18317_), .B2(new_n18287_), .ZN(new_n18320_));
  INV_X1     g17318(.I(new_n18300_), .ZN(new_n18321_));
  NAND2_X1   g17319(.A1(new_n18303_), .A2(new_n11410_), .ZN(new_n18322_));
  NOR2_X1    g17320(.A1(new_n11256_), .A2(new_n11255_), .ZN(new_n18323_));
  OAI21_X1   g17321(.A1(new_n18323_), .A2(new_n18301_), .B(new_n18308_), .ZN(new_n18324_));
  NOR3_X1    g17322(.A1(new_n18309_), .A2(new_n18297_), .A3(new_n18299_), .ZN(new_n18325_));
  AOI22_X1   g17323(.A1(new_n18324_), .A2(new_n18321_), .B1(new_n18325_), .B2(new_n18322_), .ZN(new_n18326_));
  NOR2_X1    g17324(.A1(new_n18326_), .A2(new_n18320_), .ZN(new_n18327_));
  OAI22_X1   g17325(.A1(new_n18266_), .A2(new_n18267_), .B1(new_n18315_), .B2(new_n18327_), .ZN(new_n18328_));
  INV_X1     g17326(.I(new_n18266_), .ZN(new_n18329_));
  OAI22_X1   g17327(.A1(new_n11431_), .A2(new_n11430_), .B1(new_n11412_), .B2(new_n11406_), .ZN(new_n18330_));
  NAND2_X1   g17328(.A1(new_n18326_), .A2(new_n18320_), .ZN(new_n18331_));
  NAND2_X1   g17329(.A1(new_n18286_), .A2(new_n18278_), .ZN(new_n18332_));
  NAND2_X1   g17330(.A1(new_n18288_), .A2(new_n18280_), .ZN(new_n18333_));
  NAND3_X1   g17331(.A1(new_n18314_), .A2(new_n18332_), .A3(new_n18333_), .ZN(new_n18334_));
  NAND4_X1   g17332(.A1(new_n18330_), .A2(new_n18331_), .A3(new_n18334_), .A4(new_n18329_), .ZN(new_n18335_));
  NAND2_X1   g17333(.A1(new_n18328_), .A2(new_n18335_), .ZN(new_n18336_));
  NOR2_X1    g17334(.A1(new_n11241_), .A2(new_n11235_), .ZN(new_n18337_));
  INV_X1     g17335(.I(new_n18337_), .ZN(new_n18338_));
  NOR2_X1    g17336(.A1(new_n10028_), .A2(new_n10148_), .ZN(new_n18339_));
  AOI21_X1   g17337(.A1(new_n10028_), .A2(new_n10148_), .B(new_n9915_), .ZN(new_n18340_));
  OAI22_X1   g17338(.A1(new_n11150_), .A2(new_n11155_), .B1(new_n11242_), .B2(new_n11243_), .ZN(new_n18341_));
  OAI21_X1   g17339(.A1(new_n18340_), .A2(new_n18339_), .B(new_n18341_), .ZN(new_n18342_));
  NAND2_X1   g17340(.A1(new_n11171_), .A2(new_n11166_), .ZN(new_n18343_));
  NOR2_X1    g17341(.A1(new_n11171_), .A2(new_n11166_), .ZN(new_n18344_));
  AOI21_X1   g17342(.A1(new_n11182_), .A2(new_n18343_), .B(new_n18344_), .ZN(new_n18345_));
  NAND2_X1   g17343(.A1(new_n11191_), .A2(new_n11204_), .ZN(new_n18346_));
  NOR2_X1    g17344(.A1(new_n11191_), .A2(new_n11204_), .ZN(new_n18347_));
  AOI21_X1   g17345(.A1(new_n11225_), .A2(new_n18346_), .B(new_n18347_), .ZN(new_n18348_));
  XOR2_X1    g17346(.A1(new_n18348_), .A2(new_n18345_), .Z(new_n18349_));
  INV_X1     g17347(.I(new_n18349_), .ZN(new_n18350_));
  NOR2_X1    g17348(.A1(new_n11227_), .A2(new_n11187_), .ZN(new_n18351_));
  AOI21_X1   g17349(.A1(new_n11230_), .A2(new_n11231_), .B(new_n18351_), .ZN(new_n18352_));
  AOI22_X1   g17350(.A1(new_n10016_), .A2(new_n10017_), .B1(new_n10009_), .B2(new_n10013_), .ZN(new_n18353_));
  OAI21_X1   g17351(.A1(new_n10024_), .A2(new_n18353_), .B(new_n11230_), .ZN(new_n18354_));
  NAND2_X1   g17352(.A1(new_n11216_), .A2(new_n11222_), .ZN(new_n18355_));
  NOR2_X1    g17353(.A1(new_n11218_), .A2(new_n11220_), .ZN(new_n18356_));
  NOR2_X1    g17354(.A1(new_n11221_), .A2(new_n11219_), .ZN(new_n18357_));
  NOR2_X1    g17355(.A1(new_n11206_), .A2(new_n11211_), .ZN(new_n18358_));
  NOR2_X1    g17356(.A1(new_n11215_), .A2(new_n11208_), .ZN(new_n18359_));
  NOR4_X1    g17357(.A1(new_n18359_), .A2(new_n18358_), .A3(new_n18356_), .A4(new_n18357_), .ZN(new_n18360_));
  AOI21_X1   g17358(.A1(new_n18354_), .A2(new_n18355_), .B(new_n18360_), .ZN(new_n18361_));
  INV_X1     g17359(.I(new_n18345_), .ZN(new_n18362_));
  NAND2_X1   g17360(.A1(new_n18362_), .A2(new_n18348_), .ZN(new_n18363_));
  INV_X1     g17361(.I(new_n18348_), .ZN(new_n18364_));
  NAND2_X1   g17362(.A1(new_n18364_), .A2(new_n18345_), .ZN(new_n18365_));
  NAND2_X1   g17363(.A1(new_n11177_), .A2(new_n11182_), .ZN(new_n18366_));
  NAND2_X1   g17364(.A1(new_n11186_), .A2(new_n11179_), .ZN(new_n18367_));
  NAND2_X1   g17365(.A1(new_n11223_), .A2(new_n11225_), .ZN(new_n18368_));
  NAND2_X1   g17366(.A1(new_n11226_), .A2(new_n11224_), .ZN(new_n18369_));
  NAND4_X1   g17367(.A1(new_n18369_), .A2(new_n18367_), .A3(new_n18368_), .A4(new_n18366_), .ZN(new_n18370_));
  NAND3_X1   g17368(.A1(new_n18365_), .A2(new_n18363_), .A3(new_n18370_), .ZN(new_n18371_));
  OAI22_X1   g17369(.A1(new_n18361_), .A2(new_n18350_), .B1(new_n18352_), .B2(new_n18371_), .ZN(new_n18372_));
  NAND2_X1   g17370(.A1(new_n11109_), .A2(new_n11148_), .ZN(new_n18373_));
  NAND2_X1   g17371(.A1(new_n11152_), .A2(new_n18373_), .ZN(new_n18374_));
  AOI21_X1   g17372(.A1(new_n10137_), .A2(new_n11078_), .B(new_n11237_), .ZN(new_n18375_));
  NOR2_X1    g17373(.A1(new_n11143_), .A2(new_n11137_), .ZN(new_n18376_));
  NAND2_X1   g17374(.A1(new_n11141_), .A2(new_n11139_), .ZN(new_n18377_));
  NAND2_X1   g17375(.A1(new_n11142_), .A2(new_n11140_), .ZN(new_n18378_));
  NAND2_X1   g17376(.A1(new_n11132_), .A2(new_n11127_), .ZN(new_n18379_));
  NAND2_X1   g17377(.A1(new_n11136_), .A2(new_n11129_), .ZN(new_n18380_));
  NAND4_X1   g17378(.A1(new_n18378_), .A2(new_n18377_), .A3(new_n18380_), .A4(new_n18379_), .ZN(new_n18381_));
  OAI21_X1   g17379(.A1(new_n18375_), .A2(new_n18376_), .B(new_n18381_), .ZN(new_n18382_));
  NAND2_X1   g17380(.A1(new_n11121_), .A2(new_n11117_), .ZN(new_n18383_));
  NOR2_X1    g17381(.A1(new_n11121_), .A2(new_n11117_), .ZN(new_n18384_));
  AOI21_X1   g17382(.A1(new_n11132_), .A2(new_n18383_), .B(new_n18384_), .ZN(new_n18385_));
  NOR2_X1    g17383(.A1(new_n11086_), .A2(new_n11091_), .ZN(new_n18386_));
  NOR2_X1    g17384(.A1(new_n11082_), .A2(new_n11095_), .ZN(new_n18387_));
  INV_X1     g17385(.I(new_n18387_), .ZN(new_n18388_));
  OAI21_X1   g17386(.A1(new_n11104_), .A2(new_n18386_), .B(new_n18388_), .ZN(new_n18389_));
  NOR2_X1    g17387(.A1(new_n18389_), .A2(new_n18385_), .ZN(new_n18390_));
  INV_X1     g17388(.I(new_n18390_), .ZN(new_n18391_));
  NAND2_X1   g17389(.A1(new_n18389_), .A2(new_n18385_), .ZN(new_n18392_));
  NAND2_X1   g17390(.A1(new_n18391_), .A2(new_n18392_), .ZN(new_n18393_));
  NOR2_X1    g17391(.A1(new_n11104_), .A2(new_n11097_), .ZN(new_n18394_));
  NOR2_X1    g17392(.A1(new_n11108_), .A2(new_n11099_), .ZN(new_n18395_));
  NOR2_X1    g17393(.A1(new_n11146_), .A2(new_n11144_), .ZN(new_n18396_));
  NOR2_X1    g17394(.A1(new_n11147_), .A2(new_n11145_), .ZN(new_n18397_));
  NOR4_X1    g17395(.A1(new_n18394_), .A2(new_n18395_), .A3(new_n18396_), .A4(new_n18397_), .ZN(new_n18398_));
  INV_X1     g17396(.I(new_n18392_), .ZN(new_n18399_));
  NOR3_X1    g17397(.A1(new_n18399_), .A2(new_n18398_), .A3(new_n18390_), .ZN(new_n18400_));
  AOI22_X1   g17398(.A1(new_n18382_), .A2(new_n18393_), .B1(new_n18400_), .B2(new_n18374_), .ZN(new_n18401_));
  NAND2_X1   g17399(.A1(new_n18401_), .A2(new_n18372_), .ZN(new_n18402_));
  NAND2_X1   g17400(.A1(new_n18354_), .A2(new_n18355_), .ZN(new_n18403_));
  NOR2_X1    g17401(.A1(new_n11158_), .A2(new_n11157_), .ZN(new_n18404_));
  OAI21_X1   g17402(.A1(new_n18404_), .A2(new_n18351_), .B(new_n18370_), .ZN(new_n18405_));
  NOR2_X1    g17403(.A1(new_n18349_), .A2(new_n18360_), .ZN(new_n18406_));
  AOI22_X1   g17404(.A1(new_n18405_), .A2(new_n18349_), .B1(new_n18406_), .B2(new_n18403_), .ZN(new_n18407_));
  NOR2_X1    g17405(.A1(new_n18375_), .A2(new_n18376_), .ZN(new_n18408_));
  AOI21_X1   g17406(.A1(new_n11152_), .A2(new_n18373_), .B(new_n18398_), .ZN(new_n18409_));
  NOR2_X1    g17407(.A1(new_n18399_), .A2(new_n18390_), .ZN(new_n18410_));
  NAND3_X1   g17408(.A1(new_n18391_), .A2(new_n18381_), .A3(new_n18392_), .ZN(new_n18411_));
  OAI22_X1   g17409(.A1(new_n18409_), .A2(new_n18410_), .B1(new_n18408_), .B2(new_n18411_), .ZN(new_n18412_));
  NAND2_X1   g17410(.A1(new_n18407_), .A2(new_n18412_), .ZN(new_n18413_));
  AOI22_X1   g17411(.A1(new_n18342_), .A2(new_n18338_), .B1(new_n18413_), .B2(new_n18402_), .ZN(new_n18414_));
  AOI22_X1   g17412(.A1(new_n11239_), .A2(new_n11240_), .B1(new_n11229_), .B2(new_n11234_), .ZN(new_n18415_));
  AOI21_X1   g17413(.A1(new_n11247_), .A2(new_n11074_), .B(new_n18415_), .ZN(new_n18416_));
  NOR2_X1    g17414(.A1(new_n18407_), .A2(new_n18412_), .ZN(new_n18417_));
  NOR2_X1    g17415(.A1(new_n18401_), .A2(new_n18372_), .ZN(new_n18418_));
  NOR4_X1    g17416(.A1(new_n18416_), .A2(new_n18417_), .A3(new_n18337_), .A4(new_n18418_), .ZN(new_n18419_));
  NOR2_X1    g17417(.A1(new_n18414_), .A2(new_n18419_), .ZN(new_n18420_));
  NAND2_X1   g17418(.A1(new_n18336_), .A2(new_n18420_), .ZN(new_n18421_));
  OAI22_X1   g17419(.A1(new_n18416_), .A2(new_n18337_), .B1(new_n18417_), .B2(new_n18418_), .ZN(new_n18422_));
  NAND4_X1   g17420(.A1(new_n18342_), .A2(new_n18338_), .A3(new_n18413_), .A4(new_n18402_), .ZN(new_n18423_));
  NAND2_X1   g17421(.A1(new_n18422_), .A2(new_n18423_), .ZN(new_n18424_));
  NAND3_X1   g17422(.A1(new_n18424_), .A2(new_n18328_), .A3(new_n18335_), .ZN(new_n18425_));
  AOI22_X1   g17423(.A1(new_n18263_), .A2(new_n18265_), .B1(new_n18421_), .B2(new_n18425_), .ZN(new_n18426_));
  AOI22_X1   g17424(.A1(new_n11246_), .A2(new_n11250_), .B1(new_n11432_), .B2(new_n11433_), .ZN(new_n18427_));
  OAI21_X1   g17425(.A1(new_n11073_), .A2(new_n18427_), .B(new_n18263_), .ZN(new_n18428_));
  NAND2_X1   g17426(.A1(new_n11329_), .A2(new_n11417_), .ZN(new_n18429_));
  AOI21_X1   g17427(.A1(new_n11421_), .A2(new_n18429_), .B(new_n18266_), .ZN(new_n18430_));
  AOI21_X1   g17428(.A1(new_n18331_), .A2(new_n18334_), .B(new_n18430_), .ZN(new_n18431_));
  NOR4_X1    g17429(.A1(new_n18267_), .A2(new_n18315_), .A3(new_n18327_), .A4(new_n18266_), .ZN(new_n18432_));
  NOR2_X1    g17430(.A1(new_n18431_), .A2(new_n18432_), .ZN(new_n18433_));
  NOR2_X1    g17431(.A1(new_n18433_), .A2(new_n18424_), .ZN(new_n18434_));
  NOR2_X1    g17432(.A1(new_n18336_), .A2(new_n18420_), .ZN(new_n18435_));
  NOR3_X1    g17433(.A1(new_n18428_), .A2(new_n18434_), .A3(new_n18435_), .ZN(new_n18436_));
  NOR2_X1    g17434(.A1(new_n18436_), .A2(new_n18426_), .ZN(new_n18437_));
  NOR2_X1    g17435(.A1(new_n11056_), .A2(new_n11052_), .ZN(new_n18438_));
  NAND2_X1   g17436(.A1(new_n11065_), .A2(new_n10172_), .ZN(new_n18439_));
  AOI22_X1   g17437(.A1(new_n11054_), .A2(new_n11055_), .B1(new_n11046_), .B2(new_n11051_), .ZN(new_n18440_));
  AOI21_X1   g17438(.A1(new_n18439_), .A2(new_n10704_), .B(new_n18440_), .ZN(new_n18441_));
  NOR2_X1    g17439(.A1(new_n11035_), .A2(new_n11041_), .ZN(new_n18442_));
  INV_X1     g17440(.I(new_n18442_), .ZN(new_n18443_));
  OAI22_X1   g17441(.A1(new_n10880_), .A2(new_n10879_), .B1(new_n10956_), .B2(new_n11044_), .ZN(new_n18444_));
  NAND2_X1   g17442(.A1(new_n10967_), .A2(new_n10971_), .ZN(new_n18445_));
  NOR2_X1    g17443(.A1(new_n10967_), .A2(new_n10971_), .ZN(new_n18446_));
  AOI21_X1   g17444(.A1(new_n10982_), .A2(new_n18445_), .B(new_n18446_), .ZN(new_n18447_));
  INV_X1     g17445(.I(new_n18447_), .ZN(new_n18448_));
  NAND2_X1   g17446(.A1(new_n11004_), .A2(new_n10991_), .ZN(new_n18449_));
  NOR2_X1    g17447(.A1(new_n11004_), .A2(new_n10991_), .ZN(new_n18450_));
  AOI21_X1   g17448(.A1(new_n11025_), .A2(new_n18449_), .B(new_n18450_), .ZN(new_n18451_));
  NAND2_X1   g17449(.A1(new_n18448_), .A2(new_n18451_), .ZN(new_n18452_));
  INV_X1     g17450(.I(new_n18451_), .ZN(new_n18453_));
  NAND2_X1   g17451(.A1(new_n18453_), .A2(new_n18447_), .ZN(new_n18454_));
  NAND2_X1   g17452(.A1(new_n18454_), .A2(new_n18452_), .ZN(new_n18455_));
  INV_X1     g17453(.I(new_n18455_), .ZN(new_n18456_));
  NOR2_X1    g17454(.A1(new_n10987_), .A2(new_n11027_), .ZN(new_n18457_));
  AOI21_X1   g17455(.A1(new_n11030_), .A2(new_n11031_), .B(new_n18457_), .ZN(new_n18458_));
  OAI21_X1   g17456(.A1(new_n10278_), .A2(new_n10958_), .B(new_n11030_), .ZN(new_n18459_));
  INV_X1     g17457(.I(new_n18457_), .ZN(new_n18460_));
  NAND2_X1   g17458(.A1(new_n10977_), .A2(new_n10982_), .ZN(new_n18461_));
  NAND2_X1   g17459(.A1(new_n10986_), .A2(new_n10979_), .ZN(new_n18462_));
  NAND2_X1   g17460(.A1(new_n11025_), .A2(new_n11023_), .ZN(new_n18463_));
  NAND2_X1   g17461(.A1(new_n11026_), .A2(new_n11024_), .ZN(new_n18464_));
  AND4_X2    g17462(.A1(new_n18461_), .A2(new_n18462_), .A3(new_n18463_), .A4(new_n18464_), .Z(new_n18465_));
  AOI21_X1   g17463(.A1(new_n18460_), .A2(new_n18459_), .B(new_n18465_), .ZN(new_n18466_));
  NAND4_X1   g17464(.A1(new_n18461_), .A2(new_n18462_), .A3(new_n18464_), .A4(new_n18463_), .ZN(new_n18467_));
  NAND3_X1   g17465(.A1(new_n18454_), .A2(new_n18452_), .A3(new_n18467_), .ZN(new_n18468_));
  OAI22_X1   g17466(.A1(new_n18466_), .A2(new_n18456_), .B1(new_n18458_), .B2(new_n18468_), .ZN(new_n18469_));
  NAND2_X1   g17467(.A1(new_n10909_), .A2(new_n10948_), .ZN(new_n18470_));
  NAND2_X1   g17468(.A1(new_n10952_), .A2(new_n18470_), .ZN(new_n18471_));
  NOR2_X1    g17469(.A1(new_n11038_), .A2(new_n11037_), .ZN(new_n18472_));
  NOR2_X1    g17470(.A1(new_n10943_), .A2(new_n10937_), .ZN(new_n18473_));
  NAND2_X1   g17471(.A1(new_n10941_), .A2(new_n10939_), .ZN(new_n18474_));
  NAND2_X1   g17472(.A1(new_n10942_), .A2(new_n10940_), .ZN(new_n18475_));
  NAND2_X1   g17473(.A1(new_n10927_), .A2(new_n10932_), .ZN(new_n18476_));
  NAND2_X1   g17474(.A1(new_n10936_), .A2(new_n10929_), .ZN(new_n18477_));
  NAND4_X1   g17475(.A1(new_n18475_), .A2(new_n18474_), .A3(new_n18477_), .A4(new_n18476_), .ZN(new_n18478_));
  OAI21_X1   g17476(.A1(new_n18472_), .A2(new_n18473_), .B(new_n18478_), .ZN(new_n18479_));
  NAND2_X1   g17477(.A1(new_n10921_), .A2(new_n10917_), .ZN(new_n18480_));
  NOR2_X1    g17478(.A1(new_n10921_), .A2(new_n10917_), .ZN(new_n18481_));
  AOI21_X1   g17479(.A1(new_n10932_), .A2(new_n18480_), .B(new_n18481_), .ZN(new_n18482_));
  INV_X1     g17480(.I(new_n18482_), .ZN(new_n18483_));
  NAND2_X1   g17481(.A1(new_n10885_), .A2(new_n10897_), .ZN(new_n18484_));
  NOR2_X1    g17482(.A1(new_n10885_), .A2(new_n10897_), .ZN(new_n18485_));
  AOI21_X1   g17483(.A1(new_n10941_), .A2(new_n18484_), .B(new_n18485_), .ZN(new_n18486_));
  NAND2_X1   g17484(.A1(new_n18483_), .A2(new_n18486_), .ZN(new_n18487_));
  INV_X1     g17485(.I(new_n18486_), .ZN(new_n18488_));
  NAND2_X1   g17486(.A1(new_n18488_), .A2(new_n18482_), .ZN(new_n18489_));
  NAND2_X1   g17487(.A1(new_n18489_), .A2(new_n18487_), .ZN(new_n18490_));
  AND4_X2    g17488(.A1(new_n18474_), .A2(new_n18475_), .A3(new_n18476_), .A4(new_n18477_), .Z(new_n18491_));
  INV_X1     g17489(.I(new_n18487_), .ZN(new_n18492_));
  NOR2_X1    g17490(.A1(new_n18483_), .A2(new_n18486_), .ZN(new_n18493_));
  NOR3_X1    g17491(.A1(new_n18492_), .A2(new_n18491_), .A3(new_n18493_), .ZN(new_n18494_));
  AOI22_X1   g17492(.A1(new_n18479_), .A2(new_n18490_), .B1(new_n18494_), .B2(new_n18471_), .ZN(new_n18495_));
  NAND2_X1   g17493(.A1(new_n18495_), .A2(new_n18469_), .ZN(new_n18496_));
  OAI21_X1   g17494(.A1(new_n18458_), .A2(new_n18465_), .B(new_n18455_), .ZN(new_n18497_));
  NAND2_X1   g17495(.A1(new_n18460_), .A2(new_n18459_), .ZN(new_n18498_));
  AND3_X2    g17496(.A1(new_n18454_), .A2(new_n18452_), .A3(new_n18467_), .Z(new_n18499_));
  NAND2_X1   g17497(.A1(new_n18499_), .A2(new_n18498_), .ZN(new_n18500_));
  AOI21_X1   g17498(.A1(new_n10881_), .A2(new_n10882_), .B(new_n18473_), .ZN(new_n18501_));
  AOI21_X1   g17499(.A1(new_n10952_), .A2(new_n18470_), .B(new_n18491_), .ZN(new_n18502_));
  NOR2_X1    g17500(.A1(new_n18492_), .A2(new_n18493_), .ZN(new_n18503_));
  NAND3_X1   g17501(.A1(new_n18489_), .A2(new_n18478_), .A3(new_n18487_), .ZN(new_n18504_));
  OAI22_X1   g17502(.A1(new_n18502_), .A2(new_n18503_), .B1(new_n18501_), .B2(new_n18504_), .ZN(new_n18505_));
  NAND3_X1   g17503(.A1(new_n18505_), .A2(new_n18497_), .A3(new_n18500_), .ZN(new_n18506_));
  AOI22_X1   g17504(.A1(new_n18444_), .A2(new_n18443_), .B1(new_n18496_), .B2(new_n18506_), .ZN(new_n18507_));
  AOI22_X1   g17505(.A1(new_n11048_), .A2(new_n11047_), .B1(new_n11041_), .B2(new_n11035_), .ZN(new_n18508_));
  NOR2_X1    g17506(.A1(new_n10959_), .A2(new_n10957_), .ZN(new_n18509_));
  OAI21_X1   g17507(.A1(new_n18509_), .A2(new_n18457_), .B(new_n18467_), .ZN(new_n18510_));
  AOI22_X1   g17508(.A1(new_n18510_), .A2(new_n18455_), .B1(new_n18498_), .B2(new_n18499_), .ZN(new_n18511_));
  NOR2_X1    g17509(.A1(new_n18511_), .A2(new_n18505_), .ZN(new_n18512_));
  NOR2_X1    g17510(.A1(new_n18495_), .A2(new_n18469_), .ZN(new_n18513_));
  NOR4_X1    g17511(.A1(new_n18508_), .A2(new_n18512_), .A3(new_n18513_), .A4(new_n18442_), .ZN(new_n18514_));
  NOR2_X1    g17512(.A1(new_n18514_), .A2(new_n18507_), .ZN(new_n18515_));
  NOR2_X1    g17513(.A1(new_n10784_), .A2(new_n10870_), .ZN(new_n18516_));
  AOI22_X1   g17514(.A1(new_n10708_), .A2(new_n10707_), .B1(new_n10784_), .B2(new_n10870_), .ZN(new_n18517_));
  NAND2_X1   g17515(.A1(new_n10789_), .A2(new_n10802_), .ZN(new_n18518_));
  NOR2_X1    g17516(.A1(new_n10789_), .A2(new_n10802_), .ZN(new_n18519_));
  AOI21_X1   g17517(.A1(new_n10846_), .A2(new_n18518_), .B(new_n18519_), .ZN(new_n18520_));
  NAND2_X1   g17518(.A1(new_n10826_), .A2(new_n10822_), .ZN(new_n18521_));
  NOR2_X1    g17519(.A1(new_n10826_), .A2(new_n10822_), .ZN(new_n18522_));
  AOI21_X1   g17520(.A1(new_n10837_), .A2(new_n18521_), .B(new_n18522_), .ZN(new_n18523_));
  INV_X1     g17521(.I(new_n18523_), .ZN(new_n18524_));
  NOR2_X1    g17522(.A1(new_n18524_), .A2(new_n18520_), .ZN(new_n18525_));
  INV_X1     g17523(.I(new_n18520_), .ZN(new_n18526_));
  NOR2_X1    g17524(.A1(new_n18526_), .A2(new_n18523_), .ZN(new_n18527_));
  NOR2_X1    g17525(.A1(new_n18525_), .A2(new_n18527_), .ZN(new_n18528_));
  INV_X1     g17526(.I(new_n18528_), .ZN(new_n18529_));
  AOI22_X1   g17527(.A1(new_n10454_), .A2(new_n10458_), .B1(new_n10511_), .B2(new_n10512_), .ZN(new_n18530_));
  OAI21_X1   g17528(.A1(new_n10411_), .A2(new_n18530_), .B(new_n10785_), .ZN(new_n18531_));
  NAND2_X1   g17529(.A1(new_n10853_), .A2(new_n10814_), .ZN(new_n18532_));
  NAND2_X1   g17530(.A1(new_n18531_), .A2(new_n18532_), .ZN(new_n18533_));
  NOR2_X1    g17531(.A1(new_n10857_), .A2(new_n10856_), .ZN(new_n18534_));
  NOR2_X1    g17532(.A1(new_n10842_), .A2(new_n10848_), .ZN(new_n18535_));
  NAND2_X1   g17533(.A1(new_n10844_), .A2(new_n10846_), .ZN(new_n18536_));
  NAND2_X1   g17534(.A1(new_n10847_), .A2(new_n10845_), .ZN(new_n18537_));
  NAND2_X1   g17535(.A1(new_n10837_), .A2(new_n10832_), .ZN(new_n18538_));
  NAND2_X1   g17536(.A1(new_n10841_), .A2(new_n10834_), .ZN(new_n18539_));
  NAND4_X1   g17537(.A1(new_n18538_), .A2(new_n18539_), .A3(new_n18537_), .A4(new_n18536_), .ZN(new_n18540_));
  OAI21_X1   g17538(.A1(new_n18534_), .A2(new_n18535_), .B(new_n18540_), .ZN(new_n18541_));
  AND4_X2    g17539(.A1(new_n18536_), .A2(new_n18539_), .A3(new_n18538_), .A4(new_n18537_), .Z(new_n18542_));
  NOR3_X1    g17540(.A1(new_n18542_), .A2(new_n18525_), .A3(new_n18527_), .ZN(new_n18543_));
  AOI22_X1   g17541(.A1(new_n18541_), .A2(new_n18529_), .B1(new_n18533_), .B2(new_n18543_), .ZN(new_n18544_));
  NOR2_X1    g17542(.A1(new_n10737_), .A2(new_n10777_), .ZN(new_n18545_));
  AOI21_X1   g17543(.A1(new_n10780_), .A2(new_n10709_), .B(new_n18545_), .ZN(new_n18546_));
  NAND2_X1   g17544(.A1(new_n10772_), .A2(new_n10766_), .ZN(new_n18547_));
  NOR2_X1    g17545(.A1(new_n10770_), .A2(new_n10768_), .ZN(new_n18548_));
  NOR2_X1    g17546(.A1(new_n10771_), .A2(new_n10769_), .ZN(new_n18549_));
  NOR2_X1    g17547(.A1(new_n10761_), .A2(new_n10756_), .ZN(new_n18550_));
  NOR2_X1    g17548(.A1(new_n10765_), .A2(new_n10758_), .ZN(new_n18551_));
  NOR4_X1    g17549(.A1(new_n18548_), .A2(new_n18549_), .A3(new_n18550_), .A4(new_n18551_), .ZN(new_n18552_));
  AOI21_X1   g17550(.A1(new_n10865_), .A2(new_n18547_), .B(new_n18552_), .ZN(new_n18553_));
  NAND2_X1   g17551(.A1(new_n10741_), .A2(new_n10754_), .ZN(new_n18554_));
  NOR2_X1    g17552(.A1(new_n10741_), .A2(new_n10754_), .ZN(new_n18555_));
  AOI21_X1   g17553(.A1(new_n10775_), .A2(new_n18554_), .B(new_n18555_), .ZN(new_n18556_));
  NOR2_X1    g17554(.A1(new_n10725_), .A2(new_n10715_), .ZN(new_n18557_));
  NOR2_X1    g17555(.A1(new_n10721_), .A2(new_n10719_), .ZN(new_n18558_));
  INV_X1     g17556(.I(new_n18558_), .ZN(new_n18559_));
  OAI21_X1   g17557(.A1(new_n10770_), .A2(new_n18557_), .B(new_n18559_), .ZN(new_n18560_));
  NOR2_X1    g17558(.A1(new_n18560_), .A2(new_n18556_), .ZN(new_n18561_));
  NAND2_X1   g17559(.A1(new_n18560_), .A2(new_n18556_), .ZN(new_n18562_));
  INV_X1     g17560(.I(new_n18562_), .ZN(new_n18563_));
  NOR2_X1    g17561(.A1(new_n18563_), .A2(new_n18561_), .ZN(new_n18564_));
  NAND2_X1   g17562(.A1(new_n10727_), .A2(new_n10732_), .ZN(new_n18565_));
  NAND2_X1   g17563(.A1(new_n10736_), .A2(new_n10730_), .ZN(new_n18566_));
  NAND2_X1   g17564(.A1(new_n10773_), .A2(new_n10775_), .ZN(new_n18567_));
  NAND2_X1   g17565(.A1(new_n10776_), .A2(new_n10774_), .ZN(new_n18568_));
  NAND4_X1   g17566(.A1(new_n18566_), .A2(new_n18565_), .A3(new_n18568_), .A4(new_n18567_), .ZN(new_n18569_));
  INV_X1     g17567(.I(new_n18556_), .ZN(new_n18570_));
  INV_X1     g17568(.I(new_n18557_), .ZN(new_n18571_));
  AOI21_X1   g17569(.A1(new_n10732_), .A2(new_n18571_), .B(new_n18558_), .ZN(new_n18572_));
  NAND2_X1   g17570(.A1(new_n18570_), .A2(new_n18572_), .ZN(new_n18573_));
  NAND3_X1   g17571(.A1(new_n18573_), .A2(new_n18569_), .A3(new_n18562_), .ZN(new_n18574_));
  OAI22_X1   g17572(.A1(new_n18553_), .A2(new_n18564_), .B1(new_n18546_), .B2(new_n18574_), .ZN(new_n18575_));
  NOR2_X1    g17573(.A1(new_n18544_), .A2(new_n18575_), .ZN(new_n18576_));
  AOI21_X1   g17574(.A1(new_n10786_), .A2(new_n10785_), .B(new_n18535_), .ZN(new_n18577_));
  AOI21_X1   g17575(.A1(new_n18531_), .A2(new_n18532_), .B(new_n18542_), .ZN(new_n18578_));
  NAND2_X1   g17576(.A1(new_n18526_), .A2(new_n18523_), .ZN(new_n18579_));
  NAND2_X1   g17577(.A1(new_n18524_), .A2(new_n18520_), .ZN(new_n18580_));
  NAND3_X1   g17578(.A1(new_n18580_), .A2(new_n18579_), .A3(new_n18540_), .ZN(new_n18581_));
  OAI22_X1   g17579(.A1(new_n18578_), .A2(new_n18528_), .B1(new_n18577_), .B2(new_n18581_), .ZN(new_n18582_));
  NAND2_X1   g17580(.A1(new_n10865_), .A2(new_n18547_), .ZN(new_n18583_));
  NOR2_X1    g17581(.A1(new_n10711_), .A2(new_n10710_), .ZN(new_n18584_));
  OAI21_X1   g17582(.A1(new_n18584_), .A2(new_n18545_), .B(new_n18569_), .ZN(new_n18585_));
  NAND2_X1   g17583(.A1(new_n18573_), .A2(new_n18562_), .ZN(new_n18586_));
  NOR3_X1    g17584(.A1(new_n18563_), .A2(new_n18552_), .A3(new_n18561_), .ZN(new_n18587_));
  AOI22_X1   g17585(.A1(new_n18585_), .A2(new_n18586_), .B1(new_n18583_), .B2(new_n18587_), .ZN(new_n18588_));
  NOR2_X1    g17586(.A1(new_n18588_), .A2(new_n18582_), .ZN(new_n18589_));
  OAI22_X1   g17587(.A1(new_n18517_), .A2(new_n18516_), .B1(new_n18589_), .B2(new_n18576_), .ZN(new_n18590_));
  INV_X1     g17588(.I(new_n18516_), .ZN(new_n18591_));
  INV_X1     g17589(.I(new_n10707_), .ZN(new_n18592_));
  AOI21_X1   g17590(.A1(new_n10636_), .A2(new_n10632_), .B(new_n10642_), .ZN(new_n18593_));
  OAI22_X1   g17591(.A1(new_n10863_), .A2(new_n10866_), .B1(new_n10855_), .B2(new_n10860_), .ZN(new_n18594_));
  OAI21_X1   g17592(.A1(new_n18592_), .A2(new_n18593_), .B(new_n18594_), .ZN(new_n18595_));
  NAND2_X1   g17593(.A1(new_n18588_), .A2(new_n18582_), .ZN(new_n18596_));
  NAND2_X1   g17594(.A1(new_n18541_), .A2(new_n18529_), .ZN(new_n18597_));
  NAND2_X1   g17595(.A1(new_n18543_), .A2(new_n18533_), .ZN(new_n18598_));
  NAND3_X1   g17596(.A1(new_n18575_), .A2(new_n18597_), .A3(new_n18598_), .ZN(new_n18599_));
  NAND4_X1   g17597(.A1(new_n18595_), .A2(new_n18591_), .A3(new_n18596_), .A4(new_n18599_), .ZN(new_n18600_));
  NAND2_X1   g17598(.A1(new_n18590_), .A2(new_n18600_), .ZN(new_n18601_));
  NOR2_X1    g17599(.A1(new_n18515_), .A2(new_n18601_), .ZN(new_n18602_));
  OAI22_X1   g17600(.A1(new_n18508_), .A2(new_n18442_), .B1(new_n18512_), .B2(new_n18513_), .ZN(new_n18603_));
  NAND4_X1   g17601(.A1(new_n18444_), .A2(new_n18496_), .A3(new_n18443_), .A4(new_n18506_), .ZN(new_n18604_));
  NAND2_X1   g17602(.A1(new_n18603_), .A2(new_n18604_), .ZN(new_n18605_));
  AOI22_X1   g17603(.A1(new_n18595_), .A2(new_n18591_), .B1(new_n18596_), .B2(new_n18599_), .ZN(new_n18606_));
  NOR4_X1    g17604(.A1(new_n18517_), .A2(new_n18576_), .A3(new_n18589_), .A4(new_n18516_), .ZN(new_n18607_));
  NOR2_X1    g17605(.A1(new_n18607_), .A2(new_n18606_), .ZN(new_n18608_));
  NOR2_X1    g17606(.A1(new_n18605_), .A2(new_n18608_), .ZN(new_n18609_));
  OAI22_X1   g17607(.A1(new_n18602_), .A2(new_n18609_), .B1(new_n18441_), .B2(new_n18438_), .ZN(new_n18610_));
  NAND2_X1   g17608(.A1(new_n11061_), .A2(new_n10878_), .ZN(new_n18611_));
  AOI21_X1   g17609(.A1(new_n10650_), .A2(new_n10646_), .B(new_n10657_), .ZN(new_n18612_));
  OAI22_X1   g17610(.A1(new_n18612_), .A2(new_n11064_), .B1(new_n10878_), .B2(new_n11061_), .ZN(new_n18613_));
  NAND2_X1   g17611(.A1(new_n18605_), .A2(new_n18608_), .ZN(new_n18614_));
  NAND2_X1   g17612(.A1(new_n18515_), .A2(new_n18601_), .ZN(new_n18615_));
  NAND4_X1   g17613(.A1(new_n18614_), .A2(new_n18615_), .A3(new_n18613_), .A4(new_n18611_), .ZN(new_n18616_));
  NAND2_X1   g17614(.A1(new_n18610_), .A2(new_n18616_), .ZN(new_n18617_));
  NOR2_X1    g17615(.A1(new_n18437_), .A2(new_n18617_), .ZN(new_n18618_));
  NOR2_X1    g17616(.A1(new_n11251_), .A2(new_n11434_), .ZN(new_n18619_));
  OAI21_X1   g17617(.A1(new_n10156_), .A2(new_n10160_), .B(new_n10166_), .ZN(new_n18620_));
  AOI21_X1   g17618(.A1(new_n18620_), .A2(new_n11437_), .B(new_n18427_), .ZN(new_n18621_));
  OAI22_X1   g17619(.A1(new_n18434_), .A2(new_n18435_), .B1(new_n18621_), .B2(new_n18619_), .ZN(new_n18622_));
  NAND4_X1   g17620(.A1(new_n18265_), .A2(new_n18421_), .A3(new_n18425_), .A4(new_n18263_), .ZN(new_n18623_));
  NAND2_X1   g17621(.A1(new_n18622_), .A2(new_n18623_), .ZN(new_n18624_));
  AOI22_X1   g17622(.A1(new_n18614_), .A2(new_n18615_), .B1(new_n18613_), .B2(new_n18611_), .ZN(new_n18625_));
  NOR4_X1    g17623(.A1(new_n18602_), .A2(new_n18609_), .A3(new_n18441_), .A4(new_n18438_), .ZN(new_n18626_));
  NOR2_X1    g17624(.A1(new_n18626_), .A2(new_n18625_), .ZN(new_n18627_));
  NOR2_X1    g17625(.A1(new_n18627_), .A2(new_n18624_), .ZN(new_n18628_));
  OAI22_X1   g17626(.A1(new_n18618_), .A2(new_n18628_), .B1(new_n18262_), .B2(new_n18260_), .ZN(new_n18629_));
  OAI22_X1   g17627(.A1(new_n11436_), .A2(new_n11442_), .B1(new_n11445_), .B2(new_n11446_), .ZN(new_n18630_));
  AOI21_X1   g17628(.A1(new_n11455_), .A2(new_n18630_), .B(new_n18260_), .ZN(new_n18631_));
  NAND2_X1   g17629(.A1(new_n18627_), .A2(new_n18624_), .ZN(new_n18632_));
  NAND3_X1   g17630(.A1(new_n18617_), .A2(new_n18622_), .A3(new_n18623_), .ZN(new_n18633_));
  NAND3_X1   g17631(.A1(new_n18631_), .A2(new_n18632_), .A3(new_n18633_), .ZN(new_n18634_));
  AOI21_X1   g17632(.A1(new_n18629_), .A2(new_n18634_), .B(new_n18259_), .ZN(new_n18635_));
  AOI21_X1   g17633(.A1(new_n18256_), .A2(new_n18257_), .B(new_n18255_), .ZN(new_n18636_));
  NOR3_X1    g17634(.A1(new_n18063_), .A2(new_n18251_), .A3(new_n18243_), .ZN(new_n18637_));
  NOR2_X1    g17635(.A1(new_n18636_), .A2(new_n18637_), .ZN(new_n18638_));
  AOI21_X1   g17636(.A1(new_n18632_), .A2(new_n18633_), .B(new_n18631_), .ZN(new_n18639_));
  NAND4_X1   g17637(.A1(new_n11063_), .A2(new_n11448_), .A3(new_n11449_), .A4(new_n11069_), .ZN(new_n18640_));
  AOI22_X1   g17638(.A1(new_n11448_), .A2(new_n11449_), .B1(new_n11063_), .B2(new_n11069_), .ZN(new_n18641_));
  OAI21_X1   g17639(.A1(new_n10703_), .A2(new_n18641_), .B(new_n18640_), .ZN(new_n18642_));
  NOR3_X1    g17640(.A1(new_n18642_), .A2(new_n18618_), .A3(new_n18628_), .ZN(new_n18643_));
  NOR3_X1    g17641(.A1(new_n18639_), .A2(new_n18643_), .A3(new_n18638_), .ZN(new_n18644_));
  NOR3_X1    g17642(.A1(new_n11452_), .A2(new_n11458_), .A3(new_n11871_), .ZN(new_n18645_));
  NOR3_X1    g17643(.A1(new_n10698_), .A2(new_n10697_), .A3(new_n10696_), .ZN(new_n18646_));
  AOI21_X1   g17644(.A1(new_n10695_), .A2(new_n10699_), .B(new_n18646_), .ZN(new_n18647_));
  AOI21_X1   g17645(.A1(new_n11868_), .A2(new_n11867_), .B(new_n11865_), .ZN(new_n18648_));
  NOR2_X1    g17646(.A1(new_n18647_), .A2(new_n18648_), .ZN(new_n18649_));
  OAI22_X1   g17647(.A1(new_n18649_), .A2(new_n18645_), .B1(new_n18644_), .B2(new_n18635_), .ZN(new_n18650_));
  OAI21_X1   g17648(.A1(new_n18639_), .A2(new_n18643_), .B(new_n18638_), .ZN(new_n18651_));
  NAND3_X1   g17649(.A1(new_n18629_), .A2(new_n18634_), .A3(new_n18259_), .ZN(new_n18652_));
  OAI21_X1   g17650(.A1(new_n11452_), .A2(new_n11458_), .B(new_n11871_), .ZN(new_n18653_));
  AOI21_X1   g17651(.A1(new_n11876_), .A2(new_n18653_), .B(new_n18645_), .ZN(new_n18654_));
  NAND3_X1   g17652(.A1(new_n18654_), .A2(new_n18651_), .A3(new_n18652_), .ZN(new_n18655_));
  AOI21_X1   g17653(.A1(new_n18650_), .A2(new_n18655_), .B(new_n18060_), .ZN(new_n18656_));
  NAND3_X1   g17654(.A1(new_n18650_), .A2(new_n18655_), .A3(new_n18060_), .ZN(new_n18657_));
  OAI21_X1   g17655(.A1(new_n17699_), .A2(new_n18656_), .B(new_n18657_), .ZN(new_n18658_));
  NAND4_X1   g17656(.A1(new_n17872_), .A2(new_n17868_), .A3(new_n18049_), .A4(new_n18050_), .ZN(new_n18659_));
  AOI22_X1   g17657(.A1(new_n17872_), .A2(new_n17868_), .B1(new_n18049_), .B2(new_n18050_), .ZN(new_n18660_));
  OAI21_X1   g17658(.A1(new_n17702_), .A2(new_n18660_), .B(new_n18659_), .ZN(new_n18661_));
  NOR2_X1    g17659(.A1(new_n17952_), .A2(new_n18034_), .ZN(new_n18662_));
  INV_X1     g17660(.I(new_n18662_), .ZN(new_n18663_));
  OAI22_X1   g17661(.A1(new_n18037_), .A2(new_n18038_), .B1(new_n18031_), .B2(new_n18027_), .ZN(new_n18664_));
  NAND2_X1   g17662(.A1(new_n17059_), .A2(new_n17983_), .ZN(new_n18665_));
  NAND2_X1   g17663(.A1(new_n17092_), .A2(new_n17986_), .ZN(new_n18666_));
  NOR2_X1    g17664(.A1(new_n17984_), .A2(new_n17987_), .ZN(new_n18667_));
  NAND3_X1   g17665(.A1(new_n18665_), .A2(new_n18666_), .A3(new_n18667_), .ZN(new_n18668_));
  NOR2_X1    g17666(.A1(new_n17988_), .A2(new_n17985_), .ZN(new_n18669_));
  AOI21_X1   g17667(.A1(new_n18003_), .A2(new_n18668_), .B(new_n18669_), .ZN(new_n18670_));
  INV_X1     g17668(.I(new_n18670_), .ZN(new_n18671_));
  NOR2_X1    g17669(.A1(new_n17958_), .A2(new_n17961_), .ZN(new_n18672_));
  NAND2_X1   g17670(.A1(new_n17014_), .A2(new_n17956_), .ZN(new_n18673_));
  NAND2_X1   g17671(.A1(new_n17023_), .A2(new_n17959_), .ZN(new_n18674_));
  NOR2_X1    g17672(.A1(new_n17957_), .A2(new_n17960_), .ZN(new_n18675_));
  NAND3_X1   g17673(.A1(new_n18674_), .A2(new_n18673_), .A3(new_n18675_), .ZN(new_n18676_));
  AOI21_X1   g17674(.A1(new_n18011_), .A2(new_n18676_), .B(new_n18672_), .ZN(new_n18677_));
  NAND2_X1   g17675(.A1(new_n18671_), .A2(new_n18677_), .ZN(new_n18678_));
  INV_X1     g17676(.I(new_n18678_), .ZN(new_n18679_));
  NOR2_X1    g17677(.A1(new_n18671_), .A2(new_n18677_), .ZN(new_n18680_));
  NOR2_X1    g17678(.A1(new_n18679_), .A2(new_n18680_), .ZN(new_n18681_));
  NOR2_X1    g17679(.A1(new_n18022_), .A2(new_n18023_), .ZN(new_n18682_));
  NOR2_X1    g17680(.A1(new_n18013_), .A2(new_n18006_), .ZN(new_n18683_));
  NOR2_X1    g17681(.A1(new_n18682_), .A2(new_n18683_), .ZN(new_n18684_));
  NAND2_X1   g17682(.A1(new_n17954_), .A2(new_n17955_), .ZN(new_n18685_));
  INV_X1     g17683(.I(new_n18683_), .ZN(new_n18686_));
  NOR2_X1    g17684(.A1(new_n17978_), .A2(new_n17966_), .ZN(new_n18687_));
  NOR2_X1    g17685(.A1(new_n17968_), .A2(new_n17981_), .ZN(new_n18688_));
  NOR2_X1    g17686(.A1(new_n18015_), .A2(new_n17993_), .ZN(new_n18689_));
  NOR2_X1    g17687(.A1(new_n18014_), .A2(new_n18018_), .ZN(new_n18690_));
  NOR4_X1    g17688(.A1(new_n18689_), .A2(new_n18687_), .A3(new_n18688_), .A4(new_n18690_), .ZN(new_n18691_));
  AOI21_X1   g17689(.A1(new_n18685_), .A2(new_n18686_), .B(new_n18691_), .ZN(new_n18692_));
  INV_X1     g17690(.I(new_n18680_), .ZN(new_n18693_));
  INV_X1     g17691(.I(new_n18691_), .ZN(new_n18694_));
  NAND3_X1   g17692(.A1(new_n18693_), .A2(new_n18694_), .A3(new_n18678_), .ZN(new_n18695_));
  OAI22_X1   g17693(.A1(new_n18692_), .A2(new_n18681_), .B1(new_n18684_), .B2(new_n18695_), .ZN(new_n18696_));
  NAND2_X1   g17694(.A1(new_n17142_), .A2(new_n17907_), .ZN(new_n18697_));
  NAND2_X1   g17695(.A1(new_n17179_), .A2(new_n17910_), .ZN(new_n18698_));
  NOR2_X1    g17696(.A1(new_n17911_), .A2(new_n17908_), .ZN(new_n18699_));
  NAND3_X1   g17697(.A1(new_n18697_), .A2(new_n18698_), .A3(new_n18699_), .ZN(new_n18700_));
  NOR2_X1    g17698(.A1(new_n17912_), .A2(new_n17909_), .ZN(new_n18701_));
  AOI21_X1   g17699(.A1(new_n17929_), .A2(new_n18700_), .B(new_n18701_), .ZN(new_n18702_));
  INV_X1     g17700(.I(new_n18702_), .ZN(new_n18703_));
  NAND2_X1   g17701(.A1(new_n17242_), .A2(new_n17889_), .ZN(new_n18704_));
  INV_X1     g17702(.I(new_n17890_), .ZN(new_n18705_));
  NAND4_X1   g17703(.A1(new_n17894_), .A2(new_n18704_), .A3(new_n18705_), .A4(new_n17895_), .ZN(new_n18706_));
  AOI22_X1   g17704(.A1(new_n17935_), .A2(new_n18706_), .B1(new_n17898_), .B2(new_n17896_), .ZN(new_n18707_));
  NAND2_X1   g17705(.A1(new_n18703_), .A2(new_n18707_), .ZN(new_n18708_));
  INV_X1     g17706(.I(new_n18707_), .ZN(new_n18709_));
  NAND2_X1   g17707(.A1(new_n18709_), .A2(new_n18702_), .ZN(new_n18710_));
  NAND2_X1   g17708(.A1(new_n18710_), .A2(new_n18708_), .ZN(new_n18711_));
  NAND2_X1   g17709(.A1(new_n17948_), .A2(new_n17947_), .ZN(new_n18712_));
  NOR2_X1    g17710(.A1(new_n17938_), .A2(new_n17932_), .ZN(new_n18713_));
  INV_X1     g17711(.I(new_n18713_), .ZN(new_n18714_));
  NAND2_X1   g17712(.A1(new_n18712_), .A2(new_n18714_), .ZN(new_n18715_));
  NOR2_X1    g17713(.A1(new_n17877_), .A2(new_n17876_), .ZN(new_n18716_));
  NOR2_X1    g17714(.A1(new_n17888_), .A2(new_n17901_), .ZN(new_n18717_));
  NOR2_X1    g17715(.A1(new_n17880_), .A2(new_n17905_), .ZN(new_n18718_));
  NOR2_X1    g17716(.A1(new_n17940_), .A2(new_n17917_), .ZN(new_n18719_));
  NOR2_X1    g17717(.A1(new_n17943_), .A2(new_n17939_), .ZN(new_n18720_));
  NOR4_X1    g17718(.A1(new_n18717_), .A2(new_n18719_), .A3(new_n18718_), .A4(new_n18720_), .ZN(new_n18721_));
  INV_X1     g17719(.I(new_n18721_), .ZN(new_n18722_));
  OAI21_X1   g17720(.A1(new_n18716_), .A2(new_n18713_), .B(new_n18722_), .ZN(new_n18723_));
  INV_X1     g17721(.I(new_n18708_), .ZN(new_n18724_));
  NOR2_X1    g17722(.A1(new_n18703_), .A2(new_n18707_), .ZN(new_n18725_));
  NOR3_X1    g17723(.A1(new_n18724_), .A2(new_n18725_), .A3(new_n18721_), .ZN(new_n18726_));
  AOI22_X1   g17724(.A1(new_n18711_), .A2(new_n18723_), .B1(new_n18715_), .B2(new_n18726_), .ZN(new_n18727_));
  NAND2_X1   g17725(.A1(new_n18727_), .A2(new_n18696_), .ZN(new_n18728_));
  NAND2_X1   g17726(.A1(new_n18693_), .A2(new_n18678_), .ZN(new_n18729_));
  NAND2_X1   g17727(.A1(new_n18685_), .A2(new_n18686_), .ZN(new_n18730_));
  OAI21_X1   g17728(.A1(new_n18682_), .A2(new_n18683_), .B(new_n18694_), .ZN(new_n18731_));
  NOR3_X1    g17729(.A1(new_n18679_), .A2(new_n18691_), .A3(new_n18680_), .ZN(new_n18732_));
  AOI22_X1   g17730(.A1(new_n18731_), .A2(new_n18729_), .B1(new_n18730_), .B2(new_n18732_), .ZN(new_n18733_));
  NOR2_X1    g17731(.A1(new_n18724_), .A2(new_n18725_), .ZN(new_n18734_));
  NOR2_X1    g17732(.A1(new_n18716_), .A2(new_n18713_), .ZN(new_n18735_));
  AOI21_X1   g17733(.A1(new_n18712_), .A2(new_n18714_), .B(new_n18721_), .ZN(new_n18736_));
  NAND3_X1   g17734(.A1(new_n18722_), .A2(new_n18710_), .A3(new_n18708_), .ZN(new_n18737_));
  OAI22_X1   g17735(.A1(new_n18736_), .A2(new_n18734_), .B1(new_n18735_), .B2(new_n18737_), .ZN(new_n18738_));
  NAND2_X1   g17736(.A1(new_n18733_), .A2(new_n18738_), .ZN(new_n18739_));
  AOI22_X1   g17737(.A1(new_n18728_), .A2(new_n18739_), .B1(new_n18664_), .B2(new_n18663_), .ZN(new_n18740_));
  AOI22_X1   g17738(.A1(new_n17874_), .A2(new_n17875_), .B1(new_n17952_), .B2(new_n18034_), .ZN(new_n18741_));
  NOR2_X1    g17739(.A1(new_n18733_), .A2(new_n18738_), .ZN(new_n18742_));
  NOR2_X1    g17740(.A1(new_n18727_), .A2(new_n18696_), .ZN(new_n18743_));
  NOR4_X1    g17741(.A1(new_n18742_), .A2(new_n18743_), .A3(new_n18741_), .A4(new_n18662_), .ZN(new_n18744_));
  NOR2_X1    g17742(.A1(new_n18740_), .A2(new_n18744_), .ZN(new_n18745_));
  NAND2_X1   g17743(.A1(new_n17859_), .A2(new_n17863_), .ZN(new_n18746_));
  INV_X1     g17744(.I(new_n18746_), .ZN(new_n18747_));
  AOI22_X1   g17745(.A1(new_n17775_), .A2(new_n17781_), .B1(new_n17864_), .B2(new_n17865_), .ZN(new_n18748_));
  AOI21_X1   g17746(.A1(new_n18045_), .A2(new_n18044_), .B(new_n18748_), .ZN(new_n18749_));
  INV_X1     g17747(.I(new_n17829_), .ZN(new_n18750_));
  AOI21_X1   g17748(.A1(new_n17301_), .A2(new_n17305_), .B(new_n17351_), .ZN(new_n18751_));
  NOR2_X1    g17749(.A1(new_n17343_), .A2(new_n17830_), .ZN(new_n18752_));
  OR4_X2     g17750(.A1(new_n18751_), .A2(new_n18752_), .A3(new_n17828_), .A4(new_n17831_), .Z(new_n18753_));
  AOI22_X1   g17751(.A1(new_n17848_), .A2(new_n18753_), .B1(new_n18750_), .B2(new_n17833_), .ZN(new_n18754_));
  INV_X1     g17752(.I(new_n18754_), .ZN(new_n18755_));
  NOR2_X1    g17753(.A1(new_n17802_), .A2(new_n17798_), .ZN(new_n18756_));
  NAND2_X1   g17754(.A1(new_n17421_), .A2(new_n17796_), .ZN(new_n18757_));
  INV_X1     g17755(.I(new_n17797_), .ZN(new_n18758_));
  NAND4_X1   g17756(.A1(new_n17804_), .A2(new_n18757_), .A3(new_n18758_), .A4(new_n17805_), .ZN(new_n18759_));
  AOI21_X1   g17757(.A1(new_n17795_), .A2(new_n18759_), .B(new_n18756_), .ZN(new_n18760_));
  NAND2_X1   g17758(.A1(new_n18755_), .A2(new_n18760_), .ZN(new_n18761_));
  INV_X1     g17759(.I(new_n18760_), .ZN(new_n18762_));
  NAND2_X1   g17760(.A1(new_n18762_), .A2(new_n18754_), .ZN(new_n18763_));
  NAND2_X1   g17761(.A1(new_n18761_), .A2(new_n18763_), .ZN(new_n18764_));
  NAND2_X1   g17762(.A1(new_n17784_), .A2(new_n17783_), .ZN(new_n18765_));
  NOR2_X1    g17763(.A1(new_n17851_), .A2(new_n17813_), .ZN(new_n18766_));
  INV_X1     g17764(.I(new_n18766_), .ZN(new_n18767_));
  NAND2_X1   g17765(.A1(new_n18765_), .A2(new_n18767_), .ZN(new_n18768_));
  NOR2_X1    g17766(.A1(new_n17855_), .A2(new_n17854_), .ZN(new_n18769_));
  NOR2_X1    g17767(.A1(new_n17844_), .A2(new_n17843_), .ZN(new_n18770_));
  NOR2_X1    g17768(.A1(new_n17842_), .A2(new_n17845_), .ZN(new_n18771_));
  NOR2_X1    g17769(.A1(new_n17826_), .A2(new_n17837_), .ZN(new_n18772_));
  NOR2_X1    g17770(.A1(new_n17816_), .A2(new_n17839_), .ZN(new_n18773_));
  NOR4_X1    g17771(.A1(new_n18770_), .A2(new_n18772_), .A3(new_n18773_), .A4(new_n18771_), .ZN(new_n18774_));
  INV_X1     g17772(.I(new_n18774_), .ZN(new_n18775_));
  OAI21_X1   g17773(.A1(new_n18769_), .A2(new_n18766_), .B(new_n18775_), .ZN(new_n18776_));
  NOR2_X1    g17774(.A1(new_n18762_), .A2(new_n18754_), .ZN(new_n18777_));
  NOR2_X1    g17775(.A1(new_n18755_), .A2(new_n18760_), .ZN(new_n18778_));
  NOR3_X1    g17776(.A1(new_n18778_), .A2(new_n18777_), .A3(new_n18774_), .ZN(new_n18779_));
  AOI22_X1   g17777(.A1(new_n18776_), .A2(new_n18764_), .B1(new_n18768_), .B2(new_n18779_), .ZN(new_n18780_));
  NOR2_X1    g17778(.A1(new_n17747_), .A2(new_n17750_), .ZN(new_n18781_));
  NAND2_X1   g17779(.A1(new_n17509_), .A2(new_n17745_), .ZN(new_n18782_));
  NAND2_X1   g17780(.A1(new_n17500_), .A2(new_n17748_), .ZN(new_n18783_));
  NOR2_X1    g17781(.A1(new_n17749_), .A2(new_n17746_), .ZN(new_n18784_));
  NAND3_X1   g17782(.A1(new_n18783_), .A2(new_n18782_), .A3(new_n18784_), .ZN(new_n18785_));
  AOI21_X1   g17783(.A1(new_n17744_), .A2(new_n18785_), .B(new_n18781_), .ZN(new_n18786_));
  NOR2_X1    g17784(.A1(new_n17721_), .A2(new_n17725_), .ZN(new_n18787_));
  NAND2_X1   g17785(.A1(new_n17549_), .A2(new_n17719_), .ZN(new_n18788_));
  NAND2_X1   g17786(.A1(new_n17590_), .A2(new_n17723_), .ZN(new_n18789_));
  NOR2_X1    g17787(.A1(new_n17724_), .A2(new_n17720_), .ZN(new_n18790_));
  NAND3_X1   g17788(.A1(new_n18789_), .A2(new_n18788_), .A3(new_n18790_), .ZN(new_n18791_));
  AOI21_X1   g17789(.A1(new_n17763_), .A2(new_n18791_), .B(new_n18787_), .ZN(new_n18792_));
  INV_X1     g17790(.I(new_n18792_), .ZN(new_n18793_));
  NOR2_X1    g17791(.A1(new_n18793_), .A2(new_n18786_), .ZN(new_n18794_));
  INV_X1     g17792(.I(new_n18786_), .ZN(new_n18795_));
  NOR2_X1    g17793(.A1(new_n18795_), .A2(new_n18792_), .ZN(new_n18796_));
  NOR2_X1    g17794(.A1(new_n18796_), .A2(new_n18794_), .ZN(new_n18797_));
  AOI22_X1   g17795(.A1(new_n17778_), .A2(new_n17776_), .B1(new_n17733_), .B2(new_n17773_), .ZN(new_n18798_));
  NOR2_X1    g17796(.A1(new_n17718_), .A2(new_n17730_), .ZN(new_n18799_));
  NOR2_X1    g17797(.A1(new_n17732_), .A2(new_n17710_), .ZN(new_n18800_));
  NOR2_X1    g17798(.A1(new_n17769_), .A2(new_n17755_), .ZN(new_n18801_));
  NOR2_X1    g17799(.A1(new_n17768_), .A2(new_n17772_), .ZN(new_n18802_));
  NOR4_X1    g17800(.A1(new_n18801_), .A2(new_n18802_), .A3(new_n18799_), .A4(new_n18800_), .ZN(new_n18803_));
  NOR2_X1    g17801(.A1(new_n18798_), .A2(new_n18803_), .ZN(new_n18804_));
  NAND2_X1   g17802(.A1(new_n18795_), .A2(new_n18792_), .ZN(new_n18805_));
  NAND2_X1   g17803(.A1(new_n18793_), .A2(new_n18786_), .ZN(new_n18806_));
  INV_X1     g17804(.I(new_n18803_), .ZN(new_n18807_));
  NAND3_X1   g17805(.A1(new_n18807_), .A2(new_n18806_), .A3(new_n18805_), .ZN(new_n18808_));
  OAI22_X1   g17806(.A1(new_n18804_), .A2(new_n18797_), .B1(new_n18798_), .B2(new_n18808_), .ZN(new_n18809_));
  NOR2_X1    g17807(.A1(new_n18809_), .A2(new_n18780_), .ZN(new_n18810_));
  NOR2_X1    g17808(.A1(new_n18778_), .A2(new_n18777_), .ZN(new_n18811_));
  NOR2_X1    g17809(.A1(new_n18769_), .A2(new_n18766_), .ZN(new_n18812_));
  AOI21_X1   g17810(.A1(new_n18765_), .A2(new_n18767_), .B(new_n18774_), .ZN(new_n18813_));
  NAND3_X1   g17811(.A1(new_n18775_), .A2(new_n18761_), .A3(new_n18763_), .ZN(new_n18814_));
  OAI22_X1   g17812(.A1(new_n18813_), .A2(new_n18811_), .B1(new_n18812_), .B2(new_n18814_), .ZN(new_n18815_));
  INV_X1     g17813(.I(new_n18797_), .ZN(new_n18816_));
  OAI22_X1   g17814(.A1(new_n17708_), .A2(new_n17707_), .B1(new_n17767_), .B2(new_n17759_), .ZN(new_n18817_));
  NAND2_X1   g17815(.A1(new_n18817_), .A2(new_n18807_), .ZN(new_n18818_));
  NOR3_X1    g17816(.A1(new_n18796_), .A2(new_n18794_), .A3(new_n18803_), .ZN(new_n18819_));
  AOI22_X1   g17817(.A1(new_n18818_), .A2(new_n18816_), .B1(new_n18817_), .B2(new_n18819_), .ZN(new_n18820_));
  NOR2_X1    g17818(.A1(new_n18820_), .A2(new_n18815_), .ZN(new_n18821_));
  OAI22_X1   g17819(.A1(new_n18810_), .A2(new_n18821_), .B1(new_n18749_), .B2(new_n18747_), .ZN(new_n18822_));
  OAI22_X1   g17820(.A1(new_n17706_), .A2(new_n17703_), .B1(new_n17863_), .B2(new_n17859_), .ZN(new_n18823_));
  NAND2_X1   g17821(.A1(new_n18820_), .A2(new_n18815_), .ZN(new_n18824_));
  NAND2_X1   g17822(.A1(new_n18809_), .A2(new_n18780_), .ZN(new_n18825_));
  NAND4_X1   g17823(.A1(new_n18823_), .A2(new_n18825_), .A3(new_n18824_), .A4(new_n18746_), .ZN(new_n18826_));
  NAND2_X1   g17824(.A1(new_n18822_), .A2(new_n18826_), .ZN(new_n18827_));
  NOR2_X1    g17825(.A1(new_n18745_), .A2(new_n18827_), .ZN(new_n18828_));
  OAI22_X1   g17826(.A1(new_n18742_), .A2(new_n18743_), .B1(new_n18741_), .B2(new_n18662_), .ZN(new_n18829_));
  NAND4_X1   g17827(.A1(new_n18728_), .A2(new_n18739_), .A3(new_n18664_), .A4(new_n18663_), .ZN(new_n18830_));
  NAND2_X1   g17828(.A1(new_n18829_), .A2(new_n18830_), .ZN(new_n18831_));
  AOI22_X1   g17829(.A1(new_n18824_), .A2(new_n18825_), .B1(new_n18823_), .B2(new_n18746_), .ZN(new_n18832_));
  NOR4_X1    g17830(.A1(new_n18810_), .A2(new_n18821_), .A3(new_n18749_), .A4(new_n18747_), .ZN(new_n18833_));
  NOR2_X1    g17831(.A1(new_n18832_), .A2(new_n18833_), .ZN(new_n18834_));
  NOR2_X1    g17832(.A1(new_n18831_), .A2(new_n18834_), .ZN(new_n18835_));
  OAI21_X1   g17833(.A1(new_n18835_), .A2(new_n18828_), .B(new_n18661_), .ZN(new_n18836_));
  NOR2_X1    g17834(.A1(new_n17873_), .A2(new_n18051_), .ZN(new_n18837_));
  NAND2_X1   g17835(.A1(new_n17873_), .A2(new_n18051_), .ZN(new_n18838_));
  AOI21_X1   g17836(.A1(new_n18056_), .A2(new_n18838_), .B(new_n18837_), .ZN(new_n18839_));
  NAND2_X1   g17837(.A1(new_n18831_), .A2(new_n18834_), .ZN(new_n18840_));
  NAND2_X1   g17838(.A1(new_n18745_), .A2(new_n18827_), .ZN(new_n18841_));
  NAND3_X1   g17839(.A1(new_n18839_), .A2(new_n18840_), .A3(new_n18841_), .ZN(new_n18842_));
  NAND2_X1   g17840(.A1(new_n18842_), .A2(new_n18836_), .ZN(new_n18843_));
  NAND4_X1   g17841(.A1(new_n18622_), .A2(new_n18610_), .A3(new_n18623_), .A4(new_n18616_), .ZN(new_n18844_));
  OAI22_X1   g17842(.A1(new_n18426_), .A2(new_n18436_), .B1(new_n18626_), .B2(new_n18625_), .ZN(new_n18845_));
  OAI21_X1   g17843(.A1(new_n18262_), .A2(new_n18260_), .B(new_n18845_), .ZN(new_n18846_));
  NAND2_X1   g17844(.A1(new_n18515_), .A2(new_n18608_), .ZN(new_n18847_));
  INV_X1     g17845(.I(new_n18847_), .ZN(new_n18848_));
  AOI22_X1   g17846(.A1(new_n18603_), .A2(new_n18604_), .B1(new_n18590_), .B2(new_n18600_), .ZN(new_n18849_));
  AOI21_X1   g17847(.A1(new_n18613_), .A2(new_n18611_), .B(new_n18849_), .ZN(new_n18850_));
  NAND2_X1   g17848(.A1(new_n10775_), .A2(new_n18554_), .ZN(new_n18851_));
  INV_X1     g17849(.I(new_n18555_), .ZN(new_n18852_));
  NAND2_X1   g17850(.A1(new_n10732_), .A2(new_n18571_), .ZN(new_n18853_));
  NAND4_X1   g17851(.A1(new_n18853_), .A2(new_n18851_), .A3(new_n18852_), .A4(new_n18559_), .ZN(new_n18854_));
  INV_X1     g17852(.I(new_n18854_), .ZN(new_n18855_));
  NAND2_X1   g17853(.A1(new_n18570_), .A2(new_n18560_), .ZN(new_n18856_));
  OAI21_X1   g17854(.A1(new_n18553_), .A2(new_n18855_), .B(new_n18856_), .ZN(new_n18857_));
  NAND2_X1   g17855(.A1(new_n18524_), .A2(new_n18526_), .ZN(new_n18858_));
  NAND2_X1   g17856(.A1(new_n10846_), .A2(new_n18518_), .ZN(new_n18859_));
  INV_X1     g17857(.I(new_n18519_), .ZN(new_n18860_));
  NAND2_X1   g17858(.A1(new_n10837_), .A2(new_n18521_), .ZN(new_n18861_));
  INV_X1     g17859(.I(new_n18522_), .ZN(new_n18862_));
  NAND4_X1   g17860(.A1(new_n18861_), .A2(new_n18859_), .A3(new_n18860_), .A4(new_n18862_), .ZN(new_n18863_));
  NAND2_X1   g17861(.A1(new_n18541_), .A2(new_n18863_), .ZN(new_n18864_));
  NAND3_X1   g17862(.A1(new_n18864_), .A2(new_n18857_), .A3(new_n18858_), .ZN(new_n18865_));
  NAND2_X1   g17863(.A1(new_n18585_), .A2(new_n18854_), .ZN(new_n18866_));
  INV_X1     g17864(.I(new_n18863_), .ZN(new_n18867_));
  OAI21_X1   g17865(.A1(new_n18578_), .A2(new_n18867_), .B(new_n18858_), .ZN(new_n18868_));
  NAND3_X1   g17866(.A1(new_n18866_), .A2(new_n18868_), .A3(new_n18856_), .ZN(new_n18869_));
  NAND2_X1   g17867(.A1(new_n18869_), .A2(new_n18865_), .ZN(new_n18870_));
  AOI21_X1   g17868(.A1(new_n10874_), .A2(new_n18594_), .B(new_n18516_), .ZN(new_n18871_));
  NOR2_X1    g17869(.A1(new_n18588_), .A2(new_n18544_), .ZN(new_n18872_));
  NAND2_X1   g17870(.A1(new_n18585_), .A2(new_n18586_), .ZN(new_n18873_));
  AOI22_X1   g17871(.A1(new_n18543_), .A2(new_n18533_), .B1(new_n18583_), .B2(new_n18587_), .ZN(new_n18874_));
  NAND3_X1   g17872(.A1(new_n18874_), .A2(new_n18597_), .A3(new_n18873_), .ZN(new_n18875_));
  OAI21_X1   g17873(.A1(new_n18871_), .A2(new_n18872_), .B(new_n18875_), .ZN(new_n18876_));
  NAND2_X1   g17874(.A1(new_n18876_), .A2(new_n18870_), .ZN(new_n18877_));
  XNOR2_X1   g17875(.A1(new_n18868_), .A2(new_n18857_), .ZN(new_n18878_));
  NAND2_X1   g17876(.A1(new_n18582_), .A2(new_n18575_), .ZN(new_n18879_));
  OAI21_X1   g17877(.A1(new_n18517_), .A2(new_n18516_), .B(new_n18879_), .ZN(new_n18880_));
  NAND3_X1   g17878(.A1(new_n18880_), .A2(new_n18878_), .A3(new_n18875_), .ZN(new_n18881_));
  NAND2_X1   g17879(.A1(new_n18877_), .A2(new_n18881_), .ZN(new_n18882_));
  NAND2_X1   g17880(.A1(new_n10932_), .A2(new_n18480_), .ZN(new_n18883_));
  INV_X1     g17881(.I(new_n18481_), .ZN(new_n18884_));
  NAND2_X1   g17882(.A1(new_n10941_), .A2(new_n18484_), .ZN(new_n18885_));
  INV_X1     g17883(.I(new_n18485_), .ZN(new_n18886_));
  NAND4_X1   g17884(.A1(new_n18885_), .A2(new_n18883_), .A3(new_n18884_), .A4(new_n18886_), .ZN(new_n18887_));
  INV_X1     g17885(.I(new_n18887_), .ZN(new_n18888_));
  NOR2_X1    g17886(.A1(new_n18486_), .A2(new_n18482_), .ZN(new_n18889_));
  INV_X1     g17887(.I(new_n18889_), .ZN(new_n18890_));
  OAI21_X1   g17888(.A1(new_n18502_), .A2(new_n18888_), .B(new_n18890_), .ZN(new_n18891_));
  NOR2_X1    g17889(.A1(new_n18451_), .A2(new_n18447_), .ZN(new_n18892_));
  NAND2_X1   g17890(.A1(new_n10982_), .A2(new_n18445_), .ZN(new_n18893_));
  INV_X1     g17891(.I(new_n18446_), .ZN(new_n18894_));
  NAND2_X1   g17892(.A1(new_n11025_), .A2(new_n18449_), .ZN(new_n18895_));
  INV_X1     g17893(.I(new_n18450_), .ZN(new_n18896_));
  NAND4_X1   g17894(.A1(new_n18895_), .A2(new_n18893_), .A3(new_n18894_), .A4(new_n18896_), .ZN(new_n18897_));
  AOI21_X1   g17895(.A1(new_n18510_), .A2(new_n18897_), .B(new_n18892_), .ZN(new_n18898_));
  NAND2_X1   g17896(.A1(new_n18898_), .A2(new_n18891_), .ZN(new_n18899_));
  AOI21_X1   g17897(.A1(new_n18479_), .A2(new_n18887_), .B(new_n18889_), .ZN(new_n18900_));
  INV_X1     g17898(.I(new_n18892_), .ZN(new_n18901_));
  INV_X1     g17899(.I(new_n18897_), .ZN(new_n18902_));
  OAI21_X1   g17900(.A1(new_n18466_), .A2(new_n18902_), .B(new_n18901_), .ZN(new_n18903_));
  NAND2_X1   g17901(.A1(new_n18900_), .A2(new_n18903_), .ZN(new_n18904_));
  NAND2_X1   g17902(.A1(new_n18899_), .A2(new_n18904_), .ZN(new_n18905_));
  NAND2_X1   g17903(.A1(new_n18469_), .A2(new_n18505_), .ZN(new_n18906_));
  OAI21_X1   g17904(.A1(new_n18508_), .A2(new_n18442_), .B(new_n18906_), .ZN(new_n18907_));
  NAND2_X1   g17905(.A1(new_n11035_), .A2(new_n11041_), .ZN(new_n18908_));
  AOI21_X1   g17906(.A1(new_n11059_), .A2(new_n18908_), .B(new_n18442_), .ZN(new_n18909_));
  NOR2_X1    g17907(.A1(new_n18511_), .A2(new_n18495_), .ZN(new_n18910_));
  NAND2_X1   g17908(.A1(new_n18479_), .A2(new_n18490_), .ZN(new_n18911_));
  NOR2_X1    g17909(.A1(new_n18458_), .A2(new_n18468_), .ZN(new_n18912_));
  NOR2_X1    g17910(.A1(new_n18501_), .A2(new_n18504_), .ZN(new_n18913_));
  NOR2_X1    g17911(.A1(new_n18912_), .A2(new_n18913_), .ZN(new_n18914_));
  NAND3_X1   g17912(.A1(new_n18914_), .A2(new_n18497_), .A3(new_n18911_), .ZN(new_n18915_));
  OAI21_X1   g17913(.A1(new_n18909_), .A2(new_n18910_), .B(new_n18915_), .ZN(new_n18916_));
  NOR2_X1    g17914(.A1(new_n18900_), .A2(new_n18903_), .ZN(new_n18917_));
  NOR2_X1    g17915(.A1(new_n18898_), .A2(new_n18891_), .ZN(new_n18918_));
  INV_X1     g17916(.I(new_n18497_), .ZN(new_n18919_));
  NOR2_X1    g17917(.A1(new_n18502_), .A2(new_n18503_), .ZN(new_n18920_));
  NOR4_X1    g17918(.A1(new_n18919_), .A2(new_n18920_), .A3(new_n18912_), .A4(new_n18913_), .ZN(new_n18921_));
  NOR3_X1    g17919(.A1(new_n18921_), .A2(new_n18918_), .A3(new_n18917_), .ZN(new_n18922_));
  AOI22_X1   g17920(.A1(new_n18916_), .A2(new_n18905_), .B1(new_n18907_), .B2(new_n18922_), .ZN(new_n18923_));
  NAND2_X1   g17921(.A1(new_n18882_), .A2(new_n18923_), .ZN(new_n18924_));
  INV_X1     g17922(.I(new_n18924_), .ZN(new_n18925_));
  NOR2_X1    g17923(.A1(new_n18882_), .A2(new_n18923_), .ZN(new_n18926_));
  OAI22_X1   g17924(.A1(new_n18925_), .A2(new_n18926_), .B1(new_n18850_), .B2(new_n18848_), .ZN(new_n18927_));
  OAI22_X1   g17925(.A1(new_n18441_), .A2(new_n18438_), .B1(new_n18515_), .B2(new_n18608_), .ZN(new_n18928_));
  AOI21_X1   g17926(.A1(new_n18880_), .A2(new_n18875_), .B(new_n18878_), .ZN(new_n18929_));
  NOR2_X1    g17927(.A1(new_n18871_), .A2(new_n18872_), .ZN(new_n18930_));
  INV_X1     g17928(.I(new_n18875_), .ZN(new_n18931_));
  NOR3_X1    g17929(.A1(new_n18930_), .A2(new_n18870_), .A3(new_n18931_), .ZN(new_n18932_));
  NOR2_X1    g17930(.A1(new_n18932_), .A2(new_n18929_), .ZN(new_n18933_));
  NAND2_X1   g17931(.A1(new_n18916_), .A2(new_n18905_), .ZN(new_n18934_));
  NAND2_X1   g17932(.A1(new_n18907_), .A2(new_n18922_), .ZN(new_n18935_));
  NAND2_X1   g17933(.A1(new_n18934_), .A2(new_n18935_), .ZN(new_n18936_));
  NAND2_X1   g17934(.A1(new_n18933_), .A2(new_n18936_), .ZN(new_n18937_));
  NAND4_X1   g17935(.A1(new_n18928_), .A2(new_n18847_), .A3(new_n18937_), .A4(new_n18924_), .ZN(new_n18938_));
  NAND2_X1   g17936(.A1(new_n18927_), .A2(new_n18938_), .ZN(new_n18939_));
  NAND2_X1   g17937(.A1(new_n18433_), .A2(new_n18420_), .ZN(new_n18940_));
  NAND2_X1   g17938(.A1(new_n18336_), .A2(new_n18424_), .ZN(new_n18941_));
  OAI21_X1   g17939(.A1(new_n18619_), .A2(new_n18621_), .B(new_n18941_), .ZN(new_n18942_));
  NAND2_X1   g17940(.A1(new_n11132_), .A2(new_n18383_), .ZN(new_n18943_));
  INV_X1     g17941(.I(new_n18384_), .ZN(new_n18944_));
  INV_X1     g17942(.I(new_n18386_), .ZN(new_n18945_));
  NAND2_X1   g17943(.A1(new_n11141_), .A2(new_n18945_), .ZN(new_n18946_));
  NAND4_X1   g17944(.A1(new_n18946_), .A2(new_n18943_), .A3(new_n18944_), .A4(new_n18388_), .ZN(new_n18947_));
  AOI21_X1   g17945(.A1(new_n11141_), .A2(new_n18945_), .B(new_n18387_), .ZN(new_n18948_));
  NOR2_X1    g17946(.A1(new_n18948_), .A2(new_n18385_), .ZN(new_n18949_));
  AOI21_X1   g17947(.A1(new_n18382_), .A2(new_n18947_), .B(new_n18949_), .ZN(new_n18950_));
  NOR2_X1    g17948(.A1(new_n18348_), .A2(new_n18345_), .ZN(new_n18951_));
  INV_X1     g17949(.I(new_n18951_), .ZN(new_n18952_));
  NAND2_X1   g17950(.A1(new_n11182_), .A2(new_n18343_), .ZN(new_n18953_));
  INV_X1     g17951(.I(new_n18344_), .ZN(new_n18954_));
  NAND2_X1   g17952(.A1(new_n11225_), .A2(new_n18346_), .ZN(new_n18955_));
  INV_X1     g17953(.I(new_n18347_), .ZN(new_n18956_));
  NAND4_X1   g17954(.A1(new_n18955_), .A2(new_n18953_), .A3(new_n18954_), .A4(new_n18956_), .ZN(new_n18957_));
  INV_X1     g17955(.I(new_n18957_), .ZN(new_n18958_));
  OAI21_X1   g17956(.A1(new_n18361_), .A2(new_n18958_), .B(new_n18952_), .ZN(new_n18959_));
  NOR2_X1    g17957(.A1(new_n18950_), .A2(new_n18959_), .ZN(new_n18960_));
  NAND2_X1   g17958(.A1(new_n18950_), .A2(new_n18959_), .ZN(new_n18961_));
  INV_X1     g17959(.I(new_n18961_), .ZN(new_n18962_));
  NOR2_X1    g17960(.A1(new_n18962_), .A2(new_n18960_), .ZN(new_n18963_));
  AOI22_X1   g17961(.A1(new_n18342_), .A2(new_n18338_), .B1(new_n18372_), .B2(new_n18412_), .ZN(new_n18964_));
  NAND2_X1   g17962(.A1(new_n18342_), .A2(new_n18338_), .ZN(new_n18965_));
  NAND2_X1   g17963(.A1(new_n18412_), .A2(new_n18372_), .ZN(new_n18966_));
  NOR2_X1    g17964(.A1(new_n18361_), .A2(new_n18350_), .ZN(new_n18967_));
  NOR2_X1    g17965(.A1(new_n18352_), .A2(new_n18371_), .ZN(new_n18968_));
  NOR2_X1    g17966(.A1(new_n18409_), .A2(new_n18410_), .ZN(new_n18969_));
  NOR2_X1    g17967(.A1(new_n18408_), .A2(new_n18411_), .ZN(new_n18970_));
  NOR4_X1    g17968(.A1(new_n18967_), .A2(new_n18969_), .A3(new_n18970_), .A4(new_n18968_), .ZN(new_n18971_));
  AOI21_X1   g17969(.A1(new_n18965_), .A2(new_n18966_), .B(new_n18971_), .ZN(new_n18972_));
  INV_X1     g17970(.I(new_n18960_), .ZN(new_n18973_));
  INV_X1     g17971(.I(new_n18971_), .ZN(new_n18974_));
  NAND3_X1   g17972(.A1(new_n18974_), .A2(new_n18973_), .A3(new_n18961_), .ZN(new_n18975_));
  OAI22_X1   g17973(.A1(new_n18972_), .A2(new_n18963_), .B1(new_n18964_), .B2(new_n18975_), .ZN(new_n18976_));
  NAND2_X1   g17974(.A1(new_n11277_), .A2(new_n18290_), .ZN(new_n18977_));
  INV_X1     g17975(.I(new_n18291_), .ZN(new_n18978_));
  NAND2_X1   g17976(.A1(new_n11320_), .A2(new_n18293_), .ZN(new_n18979_));
  INV_X1     g17977(.I(new_n18294_), .ZN(new_n18980_));
  NAND4_X1   g17978(.A1(new_n18979_), .A2(new_n18977_), .A3(new_n18978_), .A4(new_n18980_), .ZN(new_n18981_));
  INV_X1     g17979(.I(new_n18981_), .ZN(new_n18982_));
  NAND2_X1   g17980(.A1(new_n18296_), .A2(new_n18298_), .ZN(new_n18983_));
  OAI21_X1   g17981(.A1(new_n18310_), .A2(new_n18982_), .B(new_n18983_), .ZN(new_n18984_));
  NAND2_X1   g17982(.A1(new_n11391_), .A2(new_n18268_), .ZN(new_n18985_));
  INV_X1     g17983(.I(new_n18269_), .ZN(new_n18986_));
  NAND2_X1   g17984(.A1(new_n11382_), .A2(new_n18272_), .ZN(new_n18987_));
  INV_X1     g17985(.I(new_n18273_), .ZN(new_n18988_));
  NAND4_X1   g17986(.A1(new_n18987_), .A2(new_n18985_), .A3(new_n18986_), .A4(new_n18988_), .ZN(new_n18989_));
  INV_X1     g17987(.I(new_n18989_), .ZN(new_n18990_));
  NOR2_X1    g17988(.A1(new_n18274_), .A2(new_n18270_), .ZN(new_n18991_));
  INV_X1     g17989(.I(new_n18991_), .ZN(new_n18992_));
  OAI21_X1   g17990(.A1(new_n18319_), .A2(new_n18990_), .B(new_n18992_), .ZN(new_n18993_));
  XOR2_X1    g17991(.A1(new_n18993_), .A2(new_n18984_), .Z(new_n18994_));
  NAND2_X1   g17992(.A1(new_n18314_), .A2(new_n18320_), .ZN(new_n18995_));
  OAI21_X1   g17993(.A1(new_n18267_), .A2(new_n18266_), .B(new_n18995_), .ZN(new_n18996_));
  NOR2_X1    g17994(.A1(new_n18289_), .A2(new_n18326_), .ZN(new_n18997_));
  NAND2_X1   g17995(.A1(new_n18324_), .A2(new_n18321_), .ZN(new_n18998_));
  NAND2_X1   g17996(.A1(new_n18325_), .A2(new_n18322_), .ZN(new_n18999_));
  NAND4_X1   g17997(.A1(new_n18332_), .A2(new_n18998_), .A3(new_n18333_), .A4(new_n18999_), .ZN(new_n19000_));
  OAI21_X1   g17998(.A1(new_n18430_), .A2(new_n18997_), .B(new_n19000_), .ZN(new_n19001_));
  AOI22_X1   g17999(.A1(new_n18324_), .A2(new_n18981_), .B1(new_n18298_), .B2(new_n18296_), .ZN(new_n19002_));
  NOR2_X1    g18000(.A1(new_n19002_), .A2(new_n18993_), .ZN(new_n19003_));
  INV_X1     g18001(.I(new_n18993_), .ZN(new_n19004_));
  NOR2_X1    g18002(.A1(new_n19004_), .A2(new_n18984_), .ZN(new_n19005_));
  AND4_X2    g18003(.A1(new_n18332_), .A2(new_n18998_), .A3(new_n18333_), .A4(new_n18999_), .Z(new_n19006_));
  NOR3_X1    g18004(.A1(new_n19006_), .A2(new_n19005_), .A3(new_n19003_), .ZN(new_n19007_));
  AOI22_X1   g18005(.A1(new_n19007_), .A2(new_n18996_), .B1(new_n19001_), .B2(new_n18994_), .ZN(new_n19008_));
  NAND2_X1   g18006(.A1(new_n18976_), .A2(new_n19008_), .ZN(new_n19009_));
  INV_X1     g18007(.I(new_n18963_), .ZN(new_n19010_));
  OAI21_X1   g18008(.A1(new_n18416_), .A2(new_n18337_), .B(new_n18966_), .ZN(new_n19011_));
  NAND2_X1   g18009(.A1(new_n19011_), .A2(new_n18974_), .ZN(new_n19012_));
  NOR3_X1    g18010(.A1(new_n18962_), .A2(new_n18971_), .A3(new_n18960_), .ZN(new_n19013_));
  AOI22_X1   g18011(.A1(new_n19012_), .A2(new_n19010_), .B1(new_n19011_), .B2(new_n19013_), .ZN(new_n19014_));
  NAND2_X1   g18012(.A1(new_n19001_), .A2(new_n18994_), .ZN(new_n19015_));
  NOR2_X1    g18013(.A1(new_n19005_), .A2(new_n19003_), .ZN(new_n19016_));
  NAND3_X1   g18014(.A1(new_n18996_), .A2(new_n19016_), .A3(new_n19000_), .ZN(new_n19017_));
  NAND2_X1   g18015(.A1(new_n19015_), .A2(new_n19017_), .ZN(new_n19018_));
  NAND2_X1   g18016(.A1(new_n19018_), .A2(new_n19014_), .ZN(new_n19019_));
  AOI22_X1   g18017(.A1(new_n18942_), .A2(new_n18940_), .B1(new_n19009_), .B2(new_n19019_), .ZN(new_n19020_));
  NOR2_X1    g18018(.A1(new_n18336_), .A2(new_n18424_), .ZN(new_n19021_));
  AOI22_X1   g18019(.A1(new_n18328_), .A2(new_n18335_), .B1(new_n18422_), .B2(new_n18423_), .ZN(new_n19022_));
  AOI21_X1   g18020(.A1(new_n18265_), .A2(new_n18263_), .B(new_n19022_), .ZN(new_n19023_));
  NOR2_X1    g18021(.A1(new_n19018_), .A2(new_n19014_), .ZN(new_n19024_));
  NOR2_X1    g18022(.A1(new_n18976_), .A2(new_n19008_), .ZN(new_n19025_));
  NOR4_X1    g18023(.A1(new_n19023_), .A2(new_n19024_), .A3(new_n19025_), .A4(new_n19021_), .ZN(new_n19026_));
  NOR2_X1    g18024(.A1(new_n19020_), .A2(new_n19026_), .ZN(new_n19027_));
  NAND2_X1   g18025(.A1(new_n18939_), .A2(new_n19027_), .ZN(new_n19028_));
  AOI22_X1   g18026(.A1(new_n18928_), .A2(new_n18847_), .B1(new_n18937_), .B2(new_n18924_), .ZN(new_n19029_));
  NAND2_X1   g18027(.A1(new_n11056_), .A2(new_n11052_), .ZN(new_n19030_));
  AOI21_X1   g18028(.A1(new_n10706_), .A2(new_n19030_), .B(new_n18438_), .ZN(new_n19031_));
  OAI21_X1   g18029(.A1(new_n19031_), .A2(new_n18849_), .B(new_n18847_), .ZN(new_n19032_));
  NOR3_X1    g18030(.A1(new_n19032_), .A2(new_n18925_), .A3(new_n18926_), .ZN(new_n19033_));
  NOR2_X1    g18031(.A1(new_n19033_), .A2(new_n19029_), .ZN(new_n19034_));
  OAI22_X1   g18032(.A1(new_n19023_), .A2(new_n19021_), .B1(new_n19024_), .B2(new_n19025_), .ZN(new_n19035_));
  NAND4_X1   g18033(.A1(new_n18942_), .A2(new_n18940_), .A3(new_n19019_), .A4(new_n19009_), .ZN(new_n19036_));
  NAND2_X1   g18034(.A1(new_n19036_), .A2(new_n19035_), .ZN(new_n19037_));
  NAND2_X1   g18035(.A1(new_n19034_), .A2(new_n19037_), .ZN(new_n19038_));
  AOI22_X1   g18036(.A1(new_n19028_), .A2(new_n19038_), .B1(new_n18846_), .B2(new_n18844_), .ZN(new_n19039_));
  AOI22_X1   g18037(.A1(new_n18622_), .A2(new_n18623_), .B1(new_n18610_), .B2(new_n18616_), .ZN(new_n19040_));
  OAI21_X1   g18038(.A1(new_n18631_), .A2(new_n19040_), .B(new_n18844_), .ZN(new_n19041_));
  NOR2_X1    g18039(.A1(new_n19034_), .A2(new_n19037_), .ZN(new_n19042_));
  NOR2_X1    g18040(.A1(new_n18939_), .A2(new_n19027_), .ZN(new_n19043_));
  NOR3_X1    g18041(.A1(new_n19041_), .A2(new_n19043_), .A3(new_n19042_), .ZN(new_n19044_));
  INV_X1     g18042(.I(new_n18191_), .ZN(new_n19045_));
  INV_X1     g18043(.I(new_n18197_), .ZN(new_n19046_));
  NOR2_X1    g18044(.A1(new_n18229_), .A2(new_n18231_), .ZN(new_n19047_));
  NOR2_X1    g18045(.A1(new_n18230_), .A2(new_n18232_), .ZN(new_n19048_));
  NOR4_X1    g18046(.A1(new_n19046_), .A2(new_n19045_), .A3(new_n19047_), .A4(new_n19048_), .ZN(new_n19049_));
  INV_X1     g18047(.I(new_n19049_), .ZN(new_n19050_));
  NAND2_X1   g18048(.A1(new_n18198_), .A2(new_n18233_), .ZN(new_n19051_));
  NAND2_X1   g18049(.A1(new_n18238_), .A2(new_n19051_), .ZN(new_n19052_));
  NAND2_X1   g18050(.A1(new_n19052_), .A2(new_n19050_), .ZN(new_n19053_));
  NOR2_X1    g18051(.A1(new_n11517_), .A2(new_n18200_), .ZN(new_n19054_));
  NAND2_X1   g18052(.A1(new_n18205_), .A2(new_n18201_), .ZN(new_n19055_));
  NOR2_X1    g18053(.A1(new_n19054_), .A2(new_n19055_), .ZN(new_n19056_));
  OAI21_X1   g18054(.A1(new_n18203_), .A2(new_n18204_), .B(new_n19056_), .ZN(new_n19057_));
  AOI22_X1   g18055(.A1(new_n18224_), .A2(new_n19057_), .B1(new_n18202_), .B2(new_n18206_), .ZN(new_n19058_));
  NAND4_X1   g18056(.A1(new_n18178_), .A2(new_n18170_), .A3(new_n18171_), .A4(new_n18179_), .ZN(new_n19059_));
  NOR2_X1    g18057(.A1(new_n18177_), .A2(new_n18175_), .ZN(new_n19060_));
  AOI21_X1   g18058(.A1(new_n18190_), .A2(new_n19059_), .B(new_n19060_), .ZN(new_n19061_));
  INV_X1     g18059(.I(new_n19061_), .ZN(new_n19062_));
  NOR2_X1    g18060(.A1(new_n19062_), .A2(new_n19058_), .ZN(new_n19063_));
  INV_X1     g18061(.I(new_n19063_), .ZN(new_n19064_));
  NAND2_X1   g18062(.A1(new_n19062_), .A2(new_n19058_), .ZN(new_n19065_));
  NAND2_X1   g18063(.A1(new_n19064_), .A2(new_n19065_), .ZN(new_n19066_));
  NAND2_X1   g18064(.A1(new_n19053_), .A2(new_n19066_), .ZN(new_n19067_));
  INV_X1     g18065(.I(new_n19065_), .ZN(new_n19068_));
  NOR3_X1    g18066(.A1(new_n19068_), .A2(new_n19049_), .A3(new_n19063_), .ZN(new_n19069_));
  NAND2_X1   g18067(.A1(new_n19069_), .A2(new_n19052_), .ZN(new_n19070_));
  NAND2_X1   g18068(.A1(new_n19067_), .A2(new_n19070_), .ZN(new_n19071_));
  NAND3_X1   g18069(.A1(new_n18140_), .A2(new_n18147_), .A3(new_n18154_), .ZN(new_n19072_));
  AOI21_X1   g18070(.A1(new_n18140_), .A2(new_n18147_), .B(new_n18154_), .ZN(new_n19073_));
  OAI21_X1   g18071(.A1(new_n18245_), .A2(new_n19073_), .B(new_n19072_), .ZN(new_n19074_));
  NAND4_X1   g18072(.A1(new_n18107_), .A2(new_n18104_), .A3(new_n18105_), .A4(new_n18108_), .ZN(new_n19075_));
  OAI21_X1   g18073(.A1(new_n18115_), .A2(new_n18122_), .B(new_n19075_), .ZN(new_n19076_));
  NAND2_X1   g18074(.A1(new_n18106_), .A2(new_n18111_), .ZN(new_n19077_));
  INV_X1     g18075(.I(new_n18098_), .ZN(new_n19078_));
  OAI21_X1   g18076(.A1(new_n18133_), .A2(new_n18095_), .B(new_n19078_), .ZN(new_n19079_));
  AOI21_X1   g18077(.A1(new_n19076_), .A2(new_n19077_), .B(new_n19079_), .ZN(new_n19080_));
  NAND3_X1   g18078(.A1(new_n19079_), .A2(new_n19076_), .A3(new_n19077_), .ZN(new_n19081_));
  INV_X1     g18079(.I(new_n19081_), .ZN(new_n19082_));
  NOR2_X1    g18080(.A1(new_n19082_), .A2(new_n19080_), .ZN(new_n19083_));
  NOR2_X1    g18081(.A1(new_n11828_), .A2(new_n11818_), .ZN(new_n19084_));
  OAI21_X1   g18082(.A1(new_n11822_), .A2(new_n19084_), .B(new_n18141_), .ZN(new_n19085_));
  NAND2_X1   g18083(.A1(new_n18129_), .A2(new_n18135_), .ZN(new_n19086_));
  NOR2_X1    g18084(.A1(new_n18133_), .A2(new_n18134_), .ZN(new_n19087_));
  NOR2_X1    g18085(.A1(new_n18131_), .A2(new_n18100_), .ZN(new_n19088_));
  NOR2_X1    g18086(.A1(new_n18114_), .A2(new_n18123_), .ZN(new_n19089_));
  NOR4_X1    g18087(.A1(new_n19089_), .A2(new_n18137_), .A3(new_n19087_), .A4(new_n19088_), .ZN(new_n19090_));
  AOI21_X1   g18088(.A1(new_n19085_), .A2(new_n19086_), .B(new_n19090_), .ZN(new_n19091_));
  NOR2_X1    g18089(.A1(new_n19091_), .A2(new_n19083_), .ZN(new_n19092_));
  NAND2_X1   g18090(.A1(new_n19076_), .A2(new_n19077_), .ZN(new_n19093_));
  INV_X1     g18091(.I(new_n19079_), .ZN(new_n19094_));
  NAND2_X1   g18092(.A1(new_n19093_), .A2(new_n19094_), .ZN(new_n19095_));
  NAND2_X1   g18093(.A1(new_n19095_), .A2(new_n19081_), .ZN(new_n19096_));
  NAND2_X1   g18094(.A1(new_n19085_), .A2(new_n19086_), .ZN(new_n19097_));
  NAND2_X1   g18095(.A1(new_n11815_), .A2(new_n11813_), .ZN(new_n19098_));
  AOI21_X1   g18096(.A1(new_n11832_), .A2(new_n19098_), .B(new_n18086_), .ZN(new_n19099_));
  AOI21_X1   g18097(.A1(new_n18138_), .A2(new_n18136_), .B(new_n18102_), .ZN(new_n19100_));
  NOR3_X1    g18098(.A1(new_n19087_), .A2(new_n18137_), .A3(new_n19088_), .ZN(new_n19101_));
  NAND2_X1   g18099(.A1(new_n19101_), .A2(new_n18136_), .ZN(new_n19102_));
  OAI21_X1   g18100(.A1(new_n19099_), .A2(new_n19100_), .B(new_n19102_), .ZN(new_n19103_));
  NOR3_X1    g18101(.A1(new_n19082_), .A2(new_n19090_), .A3(new_n19080_), .ZN(new_n19104_));
  AOI22_X1   g18102(.A1(new_n19103_), .A2(new_n19096_), .B1(new_n19097_), .B2(new_n19104_), .ZN(new_n19105_));
  INV_X1     g18103(.I(new_n18066_), .ZN(new_n19106_));
  NAND2_X1   g18104(.A1(new_n11636_), .A2(new_n18064_), .ZN(new_n19107_));
  INV_X1     g18105(.I(new_n18065_), .ZN(new_n19108_));
  NOR2_X1    g18106(.A1(new_n11660_), .A2(new_n18067_), .ZN(new_n19109_));
  INV_X1     g18107(.I(new_n19109_), .ZN(new_n19110_));
  NAND4_X1   g18108(.A1(new_n19110_), .A2(new_n19107_), .A3(new_n19108_), .A4(new_n18068_), .ZN(new_n19111_));
  AOI22_X1   g18109(.A1(new_n18152_), .A2(new_n19111_), .B1(new_n19106_), .B2(new_n18069_), .ZN(new_n19112_));
  NOR2_X1    g18110(.A1(new_n19099_), .A2(new_n19100_), .ZN(new_n19113_));
  NAND3_X1   g18111(.A1(new_n19102_), .A2(new_n19095_), .A3(new_n19081_), .ZN(new_n19114_));
  OAI21_X1   g18112(.A1(new_n19113_), .A2(new_n19114_), .B(new_n19112_), .ZN(new_n19115_));
  OAI22_X1   g18113(.A1(new_n19105_), .A2(new_n19112_), .B1(new_n19092_), .B2(new_n19115_), .ZN(new_n19116_));
  NAND2_X1   g18114(.A1(new_n19116_), .A2(new_n19074_), .ZN(new_n19117_));
  OAI21_X1   g18115(.A1(new_n18156_), .A2(new_n18155_), .B(new_n18085_), .ZN(new_n19118_));
  NAND2_X1   g18116(.A1(new_n18160_), .A2(new_n19118_), .ZN(new_n19119_));
  NOR2_X1    g18117(.A1(new_n19113_), .A2(new_n19114_), .ZN(new_n19120_));
  INV_X1     g18118(.I(new_n19112_), .ZN(new_n19121_));
  OAI21_X1   g18119(.A1(new_n19092_), .A2(new_n19120_), .B(new_n19121_), .ZN(new_n19122_));
  NAND2_X1   g18120(.A1(new_n19103_), .A2(new_n19096_), .ZN(new_n19123_));
  NAND2_X1   g18121(.A1(new_n19097_), .A2(new_n19104_), .ZN(new_n19124_));
  NAND3_X1   g18122(.A1(new_n19123_), .A2(new_n19124_), .A3(new_n19112_), .ZN(new_n19125_));
  NAND4_X1   g18123(.A1(new_n19119_), .A2(new_n19122_), .A3(new_n19125_), .A4(new_n19072_), .ZN(new_n19126_));
  AOI21_X1   g18124(.A1(new_n19117_), .A2(new_n19126_), .B(new_n19071_), .ZN(new_n19127_));
  AOI22_X1   g18125(.A1(new_n19053_), .A2(new_n19066_), .B1(new_n19069_), .B2(new_n19052_), .ZN(new_n19128_));
  NOR3_X1    g18126(.A1(new_n18156_), .A2(new_n18155_), .A3(new_n18085_), .ZN(new_n19129_));
  AOI21_X1   g18127(.A1(new_n18160_), .A2(new_n19118_), .B(new_n19129_), .ZN(new_n19130_));
  AOI21_X1   g18128(.A1(new_n19122_), .A2(new_n19125_), .B(new_n19130_), .ZN(new_n19131_));
  AOI21_X1   g18129(.A1(new_n18165_), .A2(new_n18159_), .B(new_n19073_), .ZN(new_n19132_));
  NOR2_X1    g18130(.A1(new_n19105_), .A2(new_n19112_), .ZN(new_n19133_));
  NOR2_X1    g18131(.A1(new_n19092_), .A2(new_n19115_), .ZN(new_n19134_));
  NOR4_X1    g18132(.A1(new_n19133_), .A2(new_n19132_), .A3(new_n19129_), .A4(new_n19134_), .ZN(new_n19135_));
  NOR3_X1    g18133(.A1(new_n19131_), .A2(new_n19135_), .A3(new_n19128_), .ZN(new_n19136_));
  AOI21_X1   g18134(.A1(new_n18247_), .A2(new_n18246_), .B(new_n18242_), .ZN(new_n19137_));
  NAND3_X1   g18135(.A1(new_n18247_), .A2(new_n18246_), .A3(new_n18242_), .ZN(new_n19138_));
  OAI21_X1   g18136(.A1(new_n18255_), .A2(new_n19137_), .B(new_n19138_), .ZN(new_n19139_));
  NOR3_X1    g18137(.A1(new_n19139_), .A2(new_n19127_), .A3(new_n19136_), .ZN(new_n19140_));
  OAI21_X1   g18138(.A1(new_n19131_), .A2(new_n19135_), .B(new_n19128_), .ZN(new_n19141_));
  NAND3_X1   g18139(.A1(new_n19071_), .A2(new_n19117_), .A3(new_n19126_), .ZN(new_n19142_));
  OAI21_X1   g18140(.A1(new_n18166_), .A2(new_n18161_), .B(new_n18250_), .ZN(new_n19143_));
  NOR3_X1    g18141(.A1(new_n18166_), .A2(new_n18161_), .A3(new_n18250_), .ZN(new_n19144_));
  AOI21_X1   g18142(.A1(new_n18063_), .A2(new_n19143_), .B(new_n19144_), .ZN(new_n19145_));
  AOI21_X1   g18143(.A1(new_n19141_), .A2(new_n19142_), .B(new_n19145_), .ZN(new_n19146_));
  NOR2_X1    g18144(.A1(new_n19146_), .A2(new_n19140_), .ZN(new_n19147_));
  OAI21_X1   g18145(.A1(new_n19039_), .A2(new_n19044_), .B(new_n19147_), .ZN(new_n19148_));
  OAI21_X1   g18146(.A1(new_n19042_), .A2(new_n19043_), .B(new_n19041_), .ZN(new_n19149_));
  NOR2_X1    g18147(.A1(new_n18624_), .A2(new_n18617_), .ZN(new_n19150_));
  AOI21_X1   g18148(.A1(new_n18642_), .A2(new_n18845_), .B(new_n19150_), .ZN(new_n19151_));
  NAND3_X1   g18149(.A1(new_n19151_), .A2(new_n19028_), .A3(new_n19038_), .ZN(new_n19152_));
  NAND3_X1   g18150(.A1(new_n19145_), .A2(new_n19141_), .A3(new_n19142_), .ZN(new_n19153_));
  OAI21_X1   g18151(.A1(new_n19127_), .A2(new_n19136_), .B(new_n19139_), .ZN(new_n19154_));
  NAND2_X1   g18152(.A1(new_n19154_), .A2(new_n19153_), .ZN(new_n19155_));
  NAND3_X1   g18153(.A1(new_n19149_), .A2(new_n19152_), .A3(new_n19155_), .ZN(new_n19156_));
  NAND3_X1   g18154(.A1(new_n18629_), .A2(new_n18634_), .A3(new_n18638_), .ZN(new_n19157_));
  NAND3_X1   g18155(.A1(new_n11868_), .A2(new_n11867_), .A3(new_n11865_), .ZN(new_n19158_));
  OAI21_X1   g18156(.A1(new_n18647_), .A2(new_n18648_), .B(new_n19158_), .ZN(new_n19159_));
  OAI21_X1   g18157(.A1(new_n18639_), .A2(new_n18643_), .B(new_n18259_), .ZN(new_n19160_));
  NAND2_X1   g18158(.A1(new_n19159_), .A2(new_n19160_), .ZN(new_n19161_));
  AOI22_X1   g18159(.A1(new_n19161_), .A2(new_n19157_), .B1(new_n19148_), .B2(new_n19156_), .ZN(new_n19162_));
  AOI21_X1   g18160(.A1(new_n19149_), .A2(new_n19152_), .B(new_n19155_), .ZN(new_n19163_));
  NOR3_X1    g18161(.A1(new_n19039_), .A2(new_n19044_), .A3(new_n19147_), .ZN(new_n19164_));
  AOI21_X1   g18162(.A1(new_n18629_), .A2(new_n18634_), .B(new_n18638_), .ZN(new_n19165_));
  OAI21_X1   g18163(.A1(new_n18654_), .A2(new_n19165_), .B(new_n19157_), .ZN(new_n19166_));
  NOR3_X1    g18164(.A1(new_n19166_), .A2(new_n19163_), .A3(new_n19164_), .ZN(new_n19167_));
  OAI21_X1   g18165(.A1(new_n19162_), .A2(new_n19167_), .B(new_n18843_), .ZN(new_n19168_));
  NOR3_X1    g18166(.A1(new_n19162_), .A2(new_n19167_), .A3(new_n18843_), .ZN(new_n19169_));
  AOI21_X1   g18167(.A1(new_n18658_), .A2(new_n19168_), .B(new_n19169_), .ZN(new_n19170_));
  NOR2_X1    g18168(.A1(new_n18831_), .A2(new_n18827_), .ZN(new_n19171_));
  NAND2_X1   g18169(.A1(new_n18831_), .A2(new_n18827_), .ZN(new_n19172_));
  AOI21_X1   g18170(.A1(new_n18661_), .A2(new_n19172_), .B(new_n19171_), .ZN(new_n19173_));
  NOR2_X1    g18171(.A1(new_n18754_), .A2(new_n18760_), .ZN(new_n19174_));
  NAND2_X1   g18172(.A1(new_n17848_), .A2(new_n18753_), .ZN(new_n19175_));
  NAND2_X1   g18173(.A1(new_n17795_), .A2(new_n18759_), .ZN(new_n19176_));
  AOI21_X1   g18174(.A1(new_n18750_), .A2(new_n17833_), .B(new_n18756_), .ZN(new_n19177_));
  NAND3_X1   g18175(.A1(new_n19175_), .A2(new_n19176_), .A3(new_n19177_), .ZN(new_n19178_));
  AOI21_X1   g18176(.A1(new_n18776_), .A2(new_n19178_), .B(new_n19174_), .ZN(new_n19179_));
  NOR2_X1    g18177(.A1(new_n18786_), .A2(new_n18792_), .ZN(new_n19180_));
  NAND2_X1   g18178(.A1(new_n17744_), .A2(new_n18785_), .ZN(new_n19181_));
  NAND2_X1   g18179(.A1(new_n17763_), .A2(new_n18791_), .ZN(new_n19182_));
  NOR2_X1    g18180(.A1(new_n18781_), .A2(new_n18787_), .ZN(new_n19183_));
  NAND3_X1   g18181(.A1(new_n19182_), .A2(new_n19181_), .A3(new_n19183_), .ZN(new_n19184_));
  AOI21_X1   g18182(.A1(new_n18818_), .A2(new_n19184_), .B(new_n19180_), .ZN(new_n19185_));
  XNOR2_X1   g18183(.A1(new_n19185_), .A2(new_n19179_), .ZN(new_n19186_));
  NOR2_X1    g18184(.A1(new_n18820_), .A2(new_n18780_), .ZN(new_n19187_));
  AOI21_X1   g18185(.A1(new_n18746_), .A2(new_n18823_), .B(new_n19187_), .ZN(new_n19188_));
  NAND2_X1   g18186(.A1(new_n18823_), .A2(new_n18746_), .ZN(new_n19189_));
  INV_X1     g18187(.I(new_n19187_), .ZN(new_n19190_));
  NOR2_X1    g18188(.A1(new_n18813_), .A2(new_n18811_), .ZN(new_n19191_));
  NOR2_X1    g18189(.A1(new_n18812_), .A2(new_n18814_), .ZN(new_n19192_));
  NOR2_X1    g18190(.A1(new_n18804_), .A2(new_n18797_), .ZN(new_n19193_));
  NOR2_X1    g18191(.A1(new_n18808_), .A2(new_n18798_), .ZN(new_n19194_));
  NOR4_X1    g18192(.A1(new_n19193_), .A2(new_n19191_), .A3(new_n19192_), .A4(new_n19194_), .ZN(new_n19195_));
  AOI21_X1   g18193(.A1(new_n19189_), .A2(new_n19190_), .B(new_n19195_), .ZN(new_n19196_));
  INV_X1     g18194(.I(new_n19179_), .ZN(new_n19197_));
  NAND2_X1   g18195(.A1(new_n19197_), .A2(new_n19185_), .ZN(new_n19198_));
  INV_X1     g18196(.I(new_n19185_), .ZN(new_n19199_));
  NAND2_X1   g18197(.A1(new_n19199_), .A2(new_n19179_), .ZN(new_n19200_));
  INV_X1     g18198(.I(new_n19193_), .ZN(new_n19201_));
  NOR3_X1    g18199(.A1(new_n19191_), .A2(new_n19192_), .A3(new_n19194_), .ZN(new_n19202_));
  NAND2_X1   g18200(.A1(new_n19202_), .A2(new_n19201_), .ZN(new_n19203_));
  NAND3_X1   g18201(.A1(new_n19203_), .A2(new_n19200_), .A3(new_n19198_), .ZN(new_n19204_));
  OAI22_X1   g18202(.A1(new_n19196_), .A2(new_n19186_), .B1(new_n19188_), .B2(new_n19204_), .ZN(new_n19205_));
  NOR2_X1    g18203(.A1(new_n18677_), .A2(new_n18670_), .ZN(new_n19206_));
  INV_X1     g18204(.I(new_n19206_), .ZN(new_n19207_));
  NAND2_X1   g18205(.A1(new_n18003_), .A2(new_n18668_), .ZN(new_n19208_));
  NAND2_X1   g18206(.A1(new_n18011_), .A2(new_n18676_), .ZN(new_n19209_));
  NOR2_X1    g18207(.A1(new_n18672_), .A2(new_n18669_), .ZN(new_n19210_));
  NAND3_X1   g18208(.A1(new_n19209_), .A2(new_n19208_), .A3(new_n19210_), .ZN(new_n19211_));
  INV_X1     g18209(.I(new_n19211_), .ZN(new_n19212_));
  OAI21_X1   g18210(.A1(new_n18692_), .A2(new_n19212_), .B(new_n19207_), .ZN(new_n19213_));
  NOR2_X1    g18211(.A1(new_n18707_), .A2(new_n18702_), .ZN(new_n19214_));
  NAND2_X1   g18212(.A1(new_n17929_), .A2(new_n18700_), .ZN(new_n19215_));
  NAND2_X1   g18213(.A1(new_n17935_), .A2(new_n18706_), .ZN(new_n19216_));
  AOI21_X1   g18214(.A1(new_n17896_), .A2(new_n17898_), .B(new_n18701_), .ZN(new_n19217_));
  NAND3_X1   g18215(.A1(new_n19216_), .A2(new_n19215_), .A3(new_n19217_), .ZN(new_n19218_));
  AOI21_X1   g18216(.A1(new_n18723_), .A2(new_n19218_), .B(new_n19214_), .ZN(new_n19219_));
  NAND2_X1   g18217(.A1(new_n19213_), .A2(new_n19219_), .ZN(new_n19220_));
  OR2_X2     g18218(.A1(new_n19213_), .A2(new_n19219_), .Z(new_n19221_));
  NAND2_X1   g18219(.A1(new_n19221_), .A2(new_n19220_), .ZN(new_n19222_));
  NAND2_X1   g18220(.A1(new_n18696_), .A2(new_n18738_), .ZN(new_n19223_));
  OAI21_X1   g18221(.A1(new_n18741_), .A2(new_n18662_), .B(new_n19223_), .ZN(new_n19224_));
  NOR2_X1    g18222(.A1(new_n18692_), .A2(new_n18681_), .ZN(new_n19225_));
  NOR2_X1    g18223(.A1(new_n18684_), .A2(new_n18695_), .ZN(new_n19226_));
  NOR2_X1    g18224(.A1(new_n18736_), .A2(new_n18734_), .ZN(new_n19227_));
  NOR2_X1    g18225(.A1(new_n18737_), .A2(new_n18735_), .ZN(new_n19228_));
  NOR4_X1    g18226(.A1(new_n19227_), .A2(new_n19225_), .A3(new_n19226_), .A4(new_n19228_), .ZN(new_n19229_));
  INV_X1     g18227(.I(new_n19229_), .ZN(new_n19230_));
  NAND2_X1   g18228(.A1(new_n19224_), .A2(new_n19230_), .ZN(new_n19231_));
  NOR2_X1    g18229(.A1(new_n19222_), .A2(new_n19229_), .ZN(new_n19232_));
  AOI22_X1   g18230(.A1(new_n19231_), .A2(new_n19222_), .B1(new_n19232_), .B2(new_n19224_), .ZN(new_n19233_));
  NAND2_X1   g18231(.A1(new_n19233_), .A2(new_n19205_), .ZN(new_n19234_));
  NOR2_X1    g18232(.A1(new_n19196_), .A2(new_n19186_), .ZN(new_n19235_));
  NOR2_X1    g18233(.A1(new_n19204_), .A2(new_n19188_), .ZN(new_n19236_));
  NOR2_X1    g18234(.A1(new_n19235_), .A2(new_n19236_), .ZN(new_n19237_));
  INV_X1     g18235(.I(new_n19222_), .ZN(new_n19238_));
  INV_X1     g18236(.I(new_n19224_), .ZN(new_n19239_));
  NAND2_X1   g18237(.A1(new_n18664_), .A2(new_n18663_), .ZN(new_n19240_));
  AOI21_X1   g18238(.A1(new_n19240_), .A2(new_n19223_), .B(new_n19229_), .ZN(new_n19241_));
  NAND3_X1   g18239(.A1(new_n19230_), .A2(new_n19221_), .A3(new_n19220_), .ZN(new_n19242_));
  OAI22_X1   g18240(.A1(new_n19239_), .A2(new_n19242_), .B1(new_n19241_), .B2(new_n19238_), .ZN(new_n19243_));
  NAND2_X1   g18241(.A1(new_n19237_), .A2(new_n19243_), .ZN(new_n19244_));
  AOI21_X1   g18242(.A1(new_n19234_), .A2(new_n19244_), .B(new_n19173_), .ZN(new_n19245_));
  NAND2_X1   g18243(.A1(new_n18745_), .A2(new_n18834_), .ZN(new_n19246_));
  AOI22_X1   g18244(.A1(new_n18829_), .A2(new_n18830_), .B1(new_n18822_), .B2(new_n18826_), .ZN(new_n19247_));
  OAI21_X1   g18245(.A1(new_n18839_), .A2(new_n19247_), .B(new_n19246_), .ZN(new_n19248_));
  NOR2_X1    g18246(.A1(new_n19237_), .A2(new_n19243_), .ZN(new_n19249_));
  NOR2_X1    g18247(.A1(new_n19233_), .A2(new_n19205_), .ZN(new_n19250_));
  NOR3_X1    g18248(.A1(new_n19248_), .A2(new_n19249_), .A3(new_n19250_), .ZN(new_n19251_));
  NOR2_X1    g18249(.A1(new_n19245_), .A2(new_n19251_), .ZN(new_n19252_));
  NOR2_X1    g18250(.A1(new_n18939_), .A2(new_n19037_), .ZN(new_n19253_));
  AOI22_X1   g18251(.A1(new_n18927_), .A2(new_n18938_), .B1(new_n19036_), .B2(new_n19035_), .ZN(new_n19254_));
  AOI21_X1   g18252(.A1(new_n18846_), .A2(new_n18844_), .B(new_n19254_), .ZN(new_n19255_));
  NAND2_X1   g18253(.A1(new_n18382_), .A2(new_n18947_), .ZN(new_n19256_));
  INV_X1     g18254(.I(new_n18949_), .ZN(new_n19257_));
  NAND2_X1   g18255(.A1(new_n18405_), .A2(new_n18957_), .ZN(new_n19258_));
  NAND4_X1   g18256(.A1(new_n19258_), .A2(new_n19256_), .A3(new_n19257_), .A4(new_n18952_), .ZN(new_n19259_));
  AOI21_X1   g18257(.A1(new_n18952_), .A2(new_n19258_), .B(new_n18950_), .ZN(new_n19260_));
  AOI21_X1   g18258(.A1(new_n19012_), .A2(new_n19259_), .B(new_n19260_), .ZN(new_n19261_));
  NAND2_X1   g18259(.A1(new_n18330_), .A2(new_n18329_), .ZN(new_n19262_));
  AOI21_X1   g18260(.A1(new_n19262_), .A2(new_n18995_), .B(new_n19006_), .ZN(new_n19263_));
  NAND2_X1   g18261(.A1(new_n18324_), .A2(new_n18981_), .ZN(new_n19264_));
  NAND2_X1   g18262(.A1(new_n18286_), .A2(new_n18989_), .ZN(new_n19265_));
  NAND4_X1   g18263(.A1(new_n19265_), .A2(new_n19264_), .A3(new_n18983_), .A4(new_n18992_), .ZN(new_n19266_));
  INV_X1     g18264(.I(new_n19266_), .ZN(new_n19267_));
  NOR2_X1    g18265(.A1(new_n19004_), .A2(new_n19002_), .ZN(new_n19268_));
  INV_X1     g18266(.I(new_n19268_), .ZN(new_n19269_));
  OAI21_X1   g18267(.A1(new_n19263_), .A2(new_n19267_), .B(new_n19269_), .ZN(new_n19270_));
  XOR2_X1    g18268(.A1(new_n19270_), .A2(new_n19261_), .Z(new_n19271_));
  NAND2_X1   g18269(.A1(new_n19018_), .A2(new_n18976_), .ZN(new_n19272_));
  OAI21_X1   g18270(.A1(new_n19023_), .A2(new_n19021_), .B(new_n19272_), .ZN(new_n19273_));
  NAND2_X1   g18271(.A1(new_n19012_), .A2(new_n19010_), .ZN(new_n19274_));
  NAND2_X1   g18272(.A1(new_n19013_), .A2(new_n19011_), .ZN(new_n19275_));
  NAND4_X1   g18273(.A1(new_n19274_), .A2(new_n19275_), .A3(new_n19015_), .A4(new_n19017_), .ZN(new_n19276_));
  AOI21_X1   g18274(.A1(new_n19273_), .A2(new_n19276_), .B(new_n19271_), .ZN(new_n19277_));
  NOR2_X1    g18275(.A1(new_n19014_), .A2(new_n19008_), .ZN(new_n19278_));
  AOI21_X1   g18276(.A1(new_n18942_), .A2(new_n18940_), .B(new_n19278_), .ZN(new_n19279_));
  INV_X1     g18277(.I(new_n19259_), .ZN(new_n19280_));
  INV_X1     g18278(.I(new_n19260_), .ZN(new_n19281_));
  OAI21_X1   g18279(.A1(new_n18972_), .A2(new_n19280_), .B(new_n19281_), .ZN(new_n19282_));
  NAND2_X1   g18280(.A1(new_n19001_), .A2(new_n19266_), .ZN(new_n19283_));
  NAND3_X1   g18281(.A1(new_n19282_), .A2(new_n19283_), .A3(new_n19269_), .ZN(new_n19284_));
  NAND2_X1   g18282(.A1(new_n19270_), .A2(new_n19261_), .ZN(new_n19285_));
  NAND3_X1   g18283(.A1(new_n19285_), .A2(new_n19284_), .A3(new_n19276_), .ZN(new_n19286_));
  NOR2_X1    g18284(.A1(new_n19279_), .A2(new_n19286_), .ZN(new_n19287_));
  NOR2_X1    g18285(.A1(new_n19277_), .A2(new_n19287_), .ZN(new_n19288_));
  NAND4_X1   g18286(.A1(new_n18866_), .A2(new_n18864_), .A3(new_n18856_), .A4(new_n18858_), .ZN(new_n19289_));
  NAND2_X1   g18287(.A1(new_n18868_), .A2(new_n18857_), .ZN(new_n19290_));
  INV_X1     g18288(.I(new_n19290_), .ZN(new_n19291_));
  AOI21_X1   g18289(.A1(new_n18876_), .A2(new_n19289_), .B(new_n19291_), .ZN(new_n19292_));
  NAND2_X1   g18290(.A1(new_n18444_), .A2(new_n18443_), .ZN(new_n19293_));
  AOI21_X1   g18291(.A1(new_n19293_), .A2(new_n18906_), .B(new_n18921_), .ZN(new_n19294_));
  NAND2_X1   g18292(.A1(new_n18479_), .A2(new_n18887_), .ZN(new_n19295_));
  NAND2_X1   g18293(.A1(new_n18510_), .A2(new_n18897_), .ZN(new_n19296_));
  NAND4_X1   g18294(.A1(new_n19296_), .A2(new_n19295_), .A3(new_n18890_), .A4(new_n18901_), .ZN(new_n19297_));
  INV_X1     g18295(.I(new_n19297_), .ZN(new_n19298_));
  NOR2_X1    g18296(.A1(new_n18898_), .A2(new_n18900_), .ZN(new_n19299_));
  INV_X1     g18297(.I(new_n19299_), .ZN(new_n19300_));
  OAI21_X1   g18298(.A1(new_n19294_), .A2(new_n19298_), .B(new_n19300_), .ZN(new_n19301_));
  NOR2_X1    g18299(.A1(new_n19301_), .A2(new_n19292_), .ZN(new_n19302_));
  NAND2_X1   g18300(.A1(new_n18595_), .A2(new_n18591_), .ZN(new_n19303_));
  AOI21_X1   g18301(.A1(new_n19303_), .A2(new_n18879_), .B(new_n18931_), .ZN(new_n19304_));
  INV_X1     g18302(.I(new_n19289_), .ZN(new_n19305_));
  OAI21_X1   g18303(.A1(new_n19304_), .A2(new_n19305_), .B(new_n19290_), .ZN(new_n19306_));
  AOI21_X1   g18304(.A1(new_n18916_), .A2(new_n19297_), .B(new_n19299_), .ZN(new_n19307_));
  NOR2_X1    g18305(.A1(new_n19306_), .A2(new_n19307_), .ZN(new_n19308_));
  NOR2_X1    g18306(.A1(new_n19302_), .A2(new_n19308_), .ZN(new_n19309_));
  NOR2_X1    g18307(.A1(new_n18933_), .A2(new_n18923_), .ZN(new_n19310_));
  AOI21_X1   g18308(.A1(new_n18928_), .A2(new_n18847_), .B(new_n19310_), .ZN(new_n19311_));
  NAND2_X1   g18309(.A1(new_n18936_), .A2(new_n18882_), .ZN(new_n19312_));
  AOI22_X1   g18310(.A1(new_n18907_), .A2(new_n18915_), .B1(new_n18899_), .B2(new_n18904_), .ZN(new_n19313_));
  NOR2_X1    g18311(.A1(new_n18909_), .A2(new_n18910_), .ZN(new_n19314_));
  NOR3_X1    g18312(.A1(new_n19314_), .A2(new_n18905_), .A3(new_n18921_), .ZN(new_n19315_));
  NOR4_X1    g18313(.A1(new_n19313_), .A2(new_n19315_), .A3(new_n18932_), .A4(new_n18929_), .ZN(new_n19316_));
  AOI21_X1   g18314(.A1(new_n19032_), .A2(new_n19312_), .B(new_n19316_), .ZN(new_n19317_));
  NAND2_X1   g18315(.A1(new_n19306_), .A2(new_n19307_), .ZN(new_n19318_));
  NAND2_X1   g18316(.A1(new_n19301_), .A2(new_n19292_), .ZN(new_n19319_));
  NAND4_X1   g18317(.A1(new_n18877_), .A2(new_n18934_), .A3(new_n18935_), .A4(new_n18881_), .ZN(new_n19320_));
  NAND3_X1   g18318(.A1(new_n19319_), .A2(new_n19318_), .A3(new_n19320_), .ZN(new_n19321_));
  OAI22_X1   g18319(.A1(new_n19317_), .A2(new_n19309_), .B1(new_n19311_), .B2(new_n19321_), .ZN(new_n19322_));
  NOR2_X1    g18320(.A1(new_n19288_), .A2(new_n19322_), .ZN(new_n19323_));
  INV_X1     g18321(.I(new_n18427_), .ZN(new_n19324_));
  AOI21_X1   g18322(.A1(new_n19324_), .A2(new_n11439_), .B(new_n18619_), .ZN(new_n19325_));
  OAI21_X1   g18323(.A1(new_n19325_), .A2(new_n19022_), .B(new_n18940_), .ZN(new_n19326_));
  INV_X1     g18324(.I(new_n19276_), .ZN(new_n19327_));
  AOI21_X1   g18325(.A1(new_n19326_), .A2(new_n19272_), .B(new_n19327_), .ZN(new_n19328_));
  OAI22_X1   g18326(.A1(new_n19328_), .A2(new_n19271_), .B1(new_n19279_), .B2(new_n19286_), .ZN(new_n19329_));
  OAI21_X1   g18327(.A1(new_n18850_), .A2(new_n18848_), .B(new_n19312_), .ZN(new_n19330_));
  AOI21_X1   g18328(.A1(new_n19330_), .A2(new_n19320_), .B(new_n19309_), .ZN(new_n19331_));
  AOI21_X1   g18329(.A1(new_n19032_), .A2(new_n19312_), .B(new_n19321_), .ZN(new_n19332_));
  NOR2_X1    g18330(.A1(new_n19331_), .A2(new_n19332_), .ZN(new_n19333_));
  NOR2_X1    g18331(.A1(new_n19333_), .A2(new_n19329_), .ZN(new_n19334_));
  OAI22_X1   g18332(.A1(new_n19255_), .A2(new_n19253_), .B1(new_n19323_), .B2(new_n19334_), .ZN(new_n19335_));
  NAND2_X1   g18333(.A1(new_n19034_), .A2(new_n19027_), .ZN(new_n19336_));
  AOI21_X1   g18334(.A1(new_n10665_), .A2(new_n10661_), .B(new_n10673_), .ZN(new_n19337_));
  OAI22_X1   g18335(.A1(new_n19337_), .A2(new_n10701_), .B1(new_n11443_), .B2(new_n11447_), .ZN(new_n19338_));
  AOI21_X1   g18336(.A1(new_n19338_), .A2(new_n18640_), .B(new_n19040_), .ZN(new_n19339_));
  OAI22_X1   g18337(.A1(new_n19033_), .A2(new_n19029_), .B1(new_n19020_), .B2(new_n19026_), .ZN(new_n19340_));
  OAI21_X1   g18338(.A1(new_n19339_), .A2(new_n19150_), .B(new_n19340_), .ZN(new_n19341_));
  NAND2_X1   g18339(.A1(new_n19333_), .A2(new_n19329_), .ZN(new_n19342_));
  NAND2_X1   g18340(.A1(new_n19284_), .A2(new_n19285_), .ZN(new_n19343_));
  AOI21_X1   g18341(.A1(new_n18428_), .A2(new_n18941_), .B(new_n19021_), .ZN(new_n19344_));
  OAI21_X1   g18342(.A1(new_n19344_), .A2(new_n19278_), .B(new_n19276_), .ZN(new_n19345_));
  NAND2_X1   g18343(.A1(new_n19345_), .A2(new_n19343_), .ZN(new_n19346_));
  NAND3_X1   g18344(.A1(new_n19273_), .A2(new_n19271_), .A3(new_n19276_), .ZN(new_n19347_));
  NAND3_X1   g18345(.A1(new_n19322_), .A2(new_n19346_), .A3(new_n19347_), .ZN(new_n19348_));
  NAND4_X1   g18346(.A1(new_n19341_), .A2(new_n19336_), .A3(new_n19342_), .A4(new_n19348_), .ZN(new_n19349_));
  OAI21_X1   g18347(.A1(new_n19131_), .A2(new_n19135_), .B(new_n19071_), .ZN(new_n19350_));
  NOR3_X1    g18348(.A1(new_n19131_), .A2(new_n19071_), .A3(new_n19135_), .ZN(new_n19351_));
  AOI21_X1   g18349(.A1(new_n19139_), .A2(new_n19350_), .B(new_n19351_), .ZN(new_n19352_));
  AOI21_X1   g18350(.A1(new_n18238_), .A2(new_n19051_), .B(new_n19049_), .ZN(new_n19353_));
  NAND2_X1   g18351(.A1(new_n18224_), .A2(new_n19057_), .ZN(new_n19354_));
  NAND2_X1   g18352(.A1(new_n18202_), .A2(new_n18206_), .ZN(new_n19355_));
  NAND2_X1   g18353(.A1(new_n18190_), .A2(new_n19059_), .ZN(new_n19356_));
  INV_X1     g18354(.I(new_n19060_), .ZN(new_n19357_));
  NAND4_X1   g18355(.A1(new_n19354_), .A2(new_n19356_), .A3(new_n19355_), .A4(new_n19357_), .ZN(new_n19358_));
  INV_X1     g18356(.I(new_n19358_), .ZN(new_n19359_));
  OAI22_X1   g18357(.A1(new_n19353_), .A2(new_n19359_), .B1(new_n19058_), .B2(new_n19061_), .ZN(new_n19360_));
  INV_X1     g18358(.I(new_n19360_), .ZN(new_n19361_));
  OAI21_X1   g18359(.A1(new_n19092_), .A2(new_n19120_), .B(new_n19112_), .ZN(new_n19362_));
  OAI21_X1   g18360(.A1(new_n19132_), .A2(new_n19129_), .B(new_n19362_), .ZN(new_n19363_));
  AOI21_X1   g18361(.A1(new_n19097_), .A2(new_n19104_), .B(new_n19112_), .ZN(new_n19364_));
  NAND2_X1   g18362(.A1(new_n19364_), .A2(new_n19123_), .ZN(new_n19365_));
  INV_X1     g18363(.I(new_n18095_), .ZN(new_n19366_));
  NAND2_X1   g18364(.A1(new_n18092_), .A2(new_n19366_), .ZN(new_n19367_));
  NAND4_X1   g18365(.A1(new_n19076_), .A2(new_n19367_), .A3(new_n19078_), .A4(new_n19077_), .ZN(new_n19368_));
  NAND2_X1   g18366(.A1(new_n19103_), .A2(new_n19368_), .ZN(new_n19369_));
  NAND2_X1   g18367(.A1(new_n19093_), .A2(new_n19079_), .ZN(new_n19370_));
  NAND2_X1   g18368(.A1(new_n19369_), .A2(new_n19370_), .ZN(new_n19371_));
  AOI21_X1   g18369(.A1(new_n19363_), .A2(new_n19365_), .B(new_n19371_), .ZN(new_n19372_));
  INV_X1     g18370(.I(new_n19371_), .ZN(new_n19373_));
  AOI22_X1   g18371(.A1(new_n19123_), .A2(new_n19364_), .B1(new_n19369_), .B2(new_n19370_), .ZN(new_n19374_));
  NOR2_X1    g18372(.A1(new_n19105_), .A2(new_n19121_), .ZN(new_n19375_));
  OAI21_X1   g18373(.A1(new_n19130_), .A2(new_n19375_), .B(new_n19365_), .ZN(new_n19376_));
  AOI22_X1   g18374(.A1(new_n19376_), .A2(new_n19373_), .B1(new_n19363_), .B2(new_n19374_), .ZN(new_n19377_));
  OAI21_X1   g18375(.A1(new_n19130_), .A2(new_n19375_), .B(new_n19374_), .ZN(new_n19378_));
  NAND2_X1   g18376(.A1(new_n19378_), .A2(new_n19361_), .ZN(new_n19379_));
  OAI22_X1   g18377(.A1(new_n19377_), .A2(new_n19361_), .B1(new_n19379_), .B2(new_n19372_), .ZN(new_n19380_));
  NAND2_X1   g18378(.A1(new_n19352_), .A2(new_n19380_), .ZN(new_n19381_));
  AOI21_X1   g18379(.A1(new_n19117_), .A2(new_n19126_), .B(new_n19128_), .ZN(new_n19382_));
  NAND3_X1   g18380(.A1(new_n19117_), .A2(new_n19126_), .A3(new_n19128_), .ZN(new_n19383_));
  OAI21_X1   g18381(.A1(new_n19145_), .A2(new_n19382_), .B(new_n19383_), .ZN(new_n19384_));
  AOI22_X1   g18382(.A1(new_n19074_), .A2(new_n19362_), .B1(new_n19123_), .B2(new_n19364_), .ZN(new_n19385_));
  OAI21_X1   g18383(.A1(new_n19385_), .A2(new_n19371_), .B(new_n19378_), .ZN(new_n19386_));
  NAND2_X1   g18384(.A1(new_n19386_), .A2(new_n19360_), .ZN(new_n19387_));
  NAND2_X1   g18385(.A1(new_n19376_), .A2(new_n19373_), .ZN(new_n19388_));
  AOI21_X1   g18386(.A1(new_n19363_), .A2(new_n19374_), .B(new_n19360_), .ZN(new_n19389_));
  NAND2_X1   g18387(.A1(new_n19389_), .A2(new_n19388_), .ZN(new_n19390_));
  NAND3_X1   g18388(.A1(new_n19384_), .A2(new_n19387_), .A3(new_n19390_), .ZN(new_n19391_));
  NAND2_X1   g18389(.A1(new_n19381_), .A2(new_n19391_), .ZN(new_n19392_));
  NAND3_X1   g18390(.A1(new_n19335_), .A2(new_n19349_), .A3(new_n19392_), .ZN(new_n19393_));
  AOI22_X1   g18391(.A1(new_n19341_), .A2(new_n19336_), .B1(new_n19342_), .B2(new_n19348_), .ZN(new_n19394_));
  NOR4_X1    g18392(.A1(new_n19255_), .A2(new_n19323_), .A3(new_n19334_), .A4(new_n19253_), .ZN(new_n19395_));
  AOI22_X1   g18393(.A1(new_n19386_), .A2(new_n19360_), .B1(new_n19388_), .B2(new_n19389_), .ZN(new_n19396_));
  NOR2_X1    g18394(.A1(new_n19396_), .A2(new_n19384_), .ZN(new_n19397_));
  NOR2_X1    g18395(.A1(new_n19352_), .A2(new_n19380_), .ZN(new_n19398_));
  NOR2_X1    g18396(.A1(new_n19398_), .A2(new_n19397_), .ZN(new_n19399_));
  OAI21_X1   g18397(.A1(new_n19395_), .A2(new_n19394_), .B(new_n19399_), .ZN(new_n19400_));
  NAND2_X1   g18398(.A1(new_n19400_), .A2(new_n19393_), .ZN(new_n19401_));
  NOR3_X1    g18399(.A1(new_n18639_), .A2(new_n18643_), .A3(new_n18259_), .ZN(new_n19402_));
  AOI21_X1   g18400(.A1(new_n19159_), .A2(new_n19160_), .B(new_n19402_), .ZN(new_n19403_));
  AOI21_X1   g18401(.A1(new_n19149_), .A2(new_n19152_), .B(new_n19147_), .ZN(new_n19404_));
  NAND3_X1   g18402(.A1(new_n19149_), .A2(new_n19152_), .A3(new_n19147_), .ZN(new_n19405_));
  OAI21_X1   g18403(.A1(new_n19403_), .A2(new_n19404_), .B(new_n19405_), .ZN(new_n19406_));
  NAND2_X1   g18404(.A1(new_n19401_), .A2(new_n19406_), .ZN(new_n19407_));
  OAI21_X1   g18405(.A1(new_n19039_), .A2(new_n19044_), .B(new_n19155_), .ZN(new_n19408_));
  NOR3_X1    g18406(.A1(new_n19039_), .A2(new_n19044_), .A3(new_n19155_), .ZN(new_n19409_));
  AOI21_X1   g18407(.A1(new_n19166_), .A2(new_n19408_), .B(new_n19409_), .ZN(new_n19410_));
  NAND3_X1   g18408(.A1(new_n19410_), .A2(new_n19393_), .A3(new_n19400_), .ZN(new_n19411_));
  AOI21_X1   g18409(.A1(new_n19407_), .A2(new_n19411_), .B(new_n19252_), .ZN(new_n19412_));
  NAND3_X1   g18410(.A1(new_n19407_), .A2(new_n19411_), .A3(new_n19252_), .ZN(new_n19413_));
  OAI21_X1   g18411(.A1(new_n19170_), .A2(new_n19412_), .B(new_n19413_), .ZN(new_n19414_));
  NAND2_X1   g18412(.A1(new_n19376_), .A2(new_n19371_), .ZN(new_n19415_));
  NAND2_X1   g18413(.A1(new_n19384_), .A2(new_n19390_), .ZN(new_n19416_));
  AOI21_X1   g18414(.A1(new_n19416_), .A2(new_n19387_), .B(new_n19415_), .ZN(new_n19417_));
  AOI22_X1   g18415(.A1(new_n19386_), .A2(new_n19360_), .B1(new_n19371_), .B2(new_n19376_), .ZN(new_n19418_));
  NAND2_X1   g18416(.A1(new_n19416_), .A2(new_n19418_), .ZN(new_n19419_));
  INV_X1     g18417(.I(new_n19419_), .ZN(new_n19420_));
  NOR2_X1    g18418(.A1(new_n19420_), .A2(new_n19417_), .ZN(new_n19421_));
  NOR2_X1    g18419(.A1(new_n19304_), .A2(new_n19305_), .ZN(new_n19422_));
  NOR2_X1    g18420(.A1(new_n19294_), .A2(new_n19298_), .ZN(new_n19423_));
  NOR4_X1    g18421(.A1(new_n19423_), .A2(new_n19422_), .A3(new_n19291_), .A4(new_n19299_), .ZN(new_n19424_));
  INV_X1     g18422(.I(new_n19424_), .ZN(new_n19425_));
  OAI21_X1   g18423(.A1(new_n19311_), .A2(new_n19316_), .B(new_n19425_), .ZN(new_n19426_));
  NAND2_X1   g18424(.A1(new_n19301_), .A2(new_n19306_), .ZN(new_n19427_));
  NAND2_X1   g18425(.A1(new_n19269_), .A2(new_n19281_), .ZN(new_n19428_));
  AOI21_X1   g18426(.A1(new_n19012_), .A2(new_n19259_), .B(new_n19428_), .ZN(new_n19429_));
  NAND2_X1   g18427(.A1(new_n19429_), .A2(new_n19283_), .ZN(new_n19430_));
  INV_X1     g18428(.I(new_n19430_), .ZN(new_n19431_));
  NAND2_X1   g18429(.A1(new_n19270_), .A2(new_n19282_), .ZN(new_n19432_));
  OAI21_X1   g18430(.A1(new_n19328_), .A2(new_n19431_), .B(new_n19432_), .ZN(new_n19433_));
  AOI21_X1   g18431(.A1(new_n19426_), .A2(new_n19427_), .B(new_n19433_), .ZN(new_n19434_));
  OAI21_X1   g18432(.A1(new_n19317_), .A2(new_n19424_), .B(new_n19427_), .ZN(new_n19435_));
  AOI22_X1   g18433(.A1(new_n19345_), .A2(new_n19430_), .B1(new_n19282_), .B2(new_n19270_), .ZN(new_n19436_));
  NOR2_X1    g18434(.A1(new_n19436_), .A2(new_n19435_), .ZN(new_n19437_));
  NOR2_X1    g18435(.A1(new_n19434_), .A2(new_n19437_), .ZN(new_n19438_));
  OAI21_X1   g18436(.A1(new_n19151_), .A2(new_n19254_), .B(new_n19336_), .ZN(new_n19439_));
  NAND2_X1   g18437(.A1(new_n19329_), .A2(new_n19322_), .ZN(new_n19440_));
  NOR4_X1    g18438(.A1(new_n19277_), .A2(new_n19331_), .A3(new_n19287_), .A4(new_n19332_), .ZN(new_n19441_));
  AOI21_X1   g18439(.A1(new_n19439_), .A2(new_n19440_), .B(new_n19441_), .ZN(new_n19442_));
  NOR2_X1    g18440(.A1(new_n19442_), .A2(new_n19438_), .ZN(new_n19443_));
  INV_X1     g18441(.I(new_n19438_), .ZN(new_n19444_));
  OAI21_X1   g18442(.A1(new_n19255_), .A2(new_n19253_), .B(new_n19440_), .ZN(new_n19445_));
  AOI21_X1   g18443(.A1(new_n19041_), .A2(new_n19340_), .B(new_n19253_), .ZN(new_n19446_));
  INV_X1     g18444(.I(new_n19440_), .ZN(new_n19447_));
  NAND2_X1   g18445(.A1(new_n19319_), .A2(new_n19318_), .ZN(new_n19448_));
  OAI21_X1   g18446(.A1(new_n19311_), .A2(new_n19316_), .B(new_n19448_), .ZN(new_n19449_));
  NOR3_X1    g18447(.A1(new_n19302_), .A2(new_n19308_), .A3(new_n19316_), .ZN(new_n19450_));
  NAND2_X1   g18448(.A1(new_n19330_), .A2(new_n19450_), .ZN(new_n19451_));
  NAND4_X1   g18449(.A1(new_n19346_), .A2(new_n19449_), .A3(new_n19347_), .A4(new_n19451_), .ZN(new_n19452_));
  OAI21_X1   g18450(.A1(new_n19446_), .A2(new_n19447_), .B(new_n19452_), .ZN(new_n19453_));
  NOR3_X1    g18451(.A1(new_n19434_), .A2(new_n19437_), .A3(new_n19441_), .ZN(new_n19454_));
  AOI22_X1   g18452(.A1(new_n19453_), .A2(new_n19444_), .B1(new_n19445_), .B2(new_n19454_), .ZN(new_n19455_));
  INV_X1     g18453(.I(new_n19417_), .ZN(new_n19456_));
  NAND2_X1   g18454(.A1(new_n19445_), .A2(new_n19454_), .ZN(new_n19457_));
  NAND3_X1   g18455(.A1(new_n19457_), .A2(new_n19456_), .A3(new_n19419_), .ZN(new_n19458_));
  OAI22_X1   g18456(.A1(new_n19458_), .A2(new_n19443_), .B1(new_n19455_), .B2(new_n19421_), .ZN(new_n19459_));
  OAI21_X1   g18457(.A1(new_n19395_), .A2(new_n19394_), .B(new_n19392_), .ZN(new_n19460_));
  NOR3_X1    g18458(.A1(new_n19395_), .A2(new_n19394_), .A3(new_n19392_), .ZN(new_n19461_));
  AOI21_X1   g18459(.A1(new_n19406_), .A2(new_n19460_), .B(new_n19461_), .ZN(new_n19462_));
  NAND2_X1   g18460(.A1(new_n19459_), .A2(new_n19462_), .ZN(new_n19463_));
  INV_X1     g18461(.I(new_n19214_), .ZN(new_n19464_));
  NAND2_X1   g18462(.A1(new_n18723_), .A2(new_n19218_), .ZN(new_n19465_));
  NAND2_X1   g18463(.A1(new_n19465_), .A2(new_n19464_), .ZN(new_n19466_));
  NOR2_X1    g18464(.A1(new_n18692_), .A2(new_n19212_), .ZN(new_n19467_));
  INV_X1     g18465(.I(new_n19467_), .ZN(new_n19468_));
  NAND4_X1   g18466(.A1(new_n19468_), .A2(new_n19207_), .A3(new_n19464_), .A4(new_n19465_), .ZN(new_n19469_));
  AOI22_X1   g18467(.A1(new_n19231_), .A2(new_n19469_), .B1(new_n19213_), .B2(new_n19466_), .ZN(new_n19470_));
  NOR2_X1    g18468(.A1(new_n19185_), .A2(new_n19179_), .ZN(new_n19471_));
  INV_X1     g18469(.I(new_n19471_), .ZN(new_n19472_));
  INV_X1     g18470(.I(new_n19174_), .ZN(new_n19473_));
  NAND2_X1   g18471(.A1(new_n18776_), .A2(new_n19178_), .ZN(new_n19474_));
  INV_X1     g18472(.I(new_n19180_), .ZN(new_n19475_));
  NAND2_X1   g18473(.A1(new_n18818_), .A2(new_n19184_), .ZN(new_n19476_));
  NAND4_X1   g18474(.A1(new_n19476_), .A2(new_n19474_), .A3(new_n19473_), .A4(new_n19475_), .ZN(new_n19477_));
  INV_X1     g18475(.I(new_n19477_), .ZN(new_n19478_));
  OAI21_X1   g18476(.A1(new_n19196_), .A2(new_n19478_), .B(new_n19472_), .ZN(new_n19479_));
  NOR2_X1    g18477(.A1(new_n19470_), .A2(new_n19479_), .ZN(new_n19480_));
  NAND2_X1   g18478(.A1(new_n19470_), .A2(new_n19479_), .ZN(new_n19481_));
  INV_X1     g18479(.I(new_n19481_), .ZN(new_n19482_));
  NOR2_X1    g18480(.A1(new_n19482_), .A2(new_n19480_), .ZN(new_n19483_));
  NOR2_X1    g18481(.A1(new_n19237_), .A2(new_n19233_), .ZN(new_n19484_));
  NOR2_X1    g18482(.A1(new_n19173_), .A2(new_n19484_), .ZN(new_n19485_));
  NOR2_X1    g18483(.A1(new_n19241_), .A2(new_n19238_), .ZN(new_n19486_));
  NOR2_X1    g18484(.A1(new_n19239_), .A2(new_n19242_), .ZN(new_n19487_));
  NOR4_X1    g18485(.A1(new_n19486_), .A2(new_n19487_), .A3(new_n19235_), .A4(new_n19236_), .ZN(new_n19488_));
  NOR2_X1    g18486(.A1(new_n19485_), .A2(new_n19488_), .ZN(new_n19489_));
  INV_X1     g18487(.I(new_n19480_), .ZN(new_n19490_));
  INV_X1     g18488(.I(new_n19488_), .ZN(new_n19491_));
  NAND3_X1   g18489(.A1(new_n19490_), .A2(new_n19491_), .A3(new_n19481_), .ZN(new_n19492_));
  OAI22_X1   g18490(.A1(new_n19489_), .A2(new_n19483_), .B1(new_n19485_), .B2(new_n19492_), .ZN(new_n19493_));
  NOR2_X1    g18491(.A1(new_n19459_), .A2(new_n19462_), .ZN(new_n19494_));
  NAND2_X1   g18492(.A1(new_n19456_), .A2(new_n19419_), .ZN(new_n19495_));
  NAND2_X1   g18493(.A1(new_n19453_), .A2(new_n19444_), .ZN(new_n19496_));
  NOR2_X1    g18494(.A1(new_n19446_), .A2(new_n19447_), .ZN(new_n19497_));
  NAND2_X1   g18495(.A1(new_n19436_), .A2(new_n19435_), .ZN(new_n19498_));
  NAND3_X1   g18496(.A1(new_n19433_), .A2(new_n19426_), .A3(new_n19427_), .ZN(new_n19499_));
  NAND3_X1   g18497(.A1(new_n19498_), .A2(new_n19499_), .A3(new_n19452_), .ZN(new_n19500_));
  OAI22_X1   g18498(.A1(new_n19442_), .A2(new_n19438_), .B1(new_n19497_), .B2(new_n19500_), .ZN(new_n19501_));
  AOI21_X1   g18499(.A1(new_n19439_), .A2(new_n19440_), .B(new_n19500_), .ZN(new_n19502_));
  NOR3_X1    g18500(.A1(new_n19502_), .A2(new_n19417_), .A3(new_n19420_), .ZN(new_n19503_));
  AOI22_X1   g18501(.A1(new_n19503_), .A2(new_n19496_), .B1(new_n19501_), .B2(new_n19495_), .ZN(new_n19504_));
  AOI21_X1   g18502(.A1(new_n19335_), .A2(new_n19349_), .B(new_n19399_), .ZN(new_n19505_));
  NAND3_X1   g18503(.A1(new_n19335_), .A2(new_n19399_), .A3(new_n19349_), .ZN(new_n19506_));
  OAI21_X1   g18504(.A1(new_n19410_), .A2(new_n19505_), .B(new_n19506_), .ZN(new_n19507_));
  NOR2_X1    g18505(.A1(new_n19504_), .A2(new_n19507_), .ZN(new_n19508_));
  OAI21_X1   g18506(.A1(new_n19494_), .A2(new_n19508_), .B(new_n19493_), .ZN(new_n19509_));
  NOR2_X1    g18507(.A1(new_n19494_), .A2(new_n19493_), .ZN(new_n19510_));
  AOI22_X1   g18508(.A1(new_n19414_), .A2(new_n19509_), .B1(new_n19463_), .B2(new_n19510_), .ZN(new_n19511_));
  INV_X1     g18509(.I(new_n19470_), .ZN(new_n19512_));
  OAI21_X1   g18510(.A1(new_n17661_), .A2(new_n17655_), .B(new_n16959_), .ZN(new_n19513_));
  AOI22_X1   g18511(.A1(new_n16943_), .A2(new_n19513_), .B1(new_n17633_), .B2(new_n17629_), .ZN(new_n19514_));
  OAI22_X1   g18512(.A1(new_n19514_), .A2(new_n17701_), .B1(new_n18048_), .B2(new_n18042_), .ZN(new_n19515_));
  AOI21_X1   g18513(.A1(new_n19515_), .A2(new_n18659_), .B(new_n19247_), .ZN(new_n19516_));
  OAI22_X1   g18514(.A1(new_n19516_), .A2(new_n19171_), .B1(new_n19237_), .B2(new_n19233_), .ZN(new_n19517_));
  NAND2_X1   g18515(.A1(new_n19517_), .A2(new_n19491_), .ZN(new_n19518_));
  NAND2_X1   g18516(.A1(new_n19466_), .A2(new_n19213_), .ZN(new_n19519_));
  NAND2_X1   g18517(.A1(new_n19231_), .A2(new_n19469_), .ZN(new_n19520_));
  INV_X1     g18518(.I(new_n19196_), .ZN(new_n19521_));
  NAND2_X1   g18519(.A1(new_n19521_), .A2(new_n19477_), .ZN(new_n19522_));
  NAND4_X1   g18520(.A1(new_n19522_), .A2(new_n19520_), .A3(new_n19519_), .A4(new_n19472_), .ZN(new_n19523_));
  AOI22_X1   g18521(.A1(new_n19518_), .A2(new_n19523_), .B1(new_n19512_), .B2(new_n19479_), .ZN(new_n19524_));
  INV_X1     g18522(.I(new_n19524_), .ZN(new_n19525_));
  NAND2_X1   g18523(.A1(new_n19503_), .A2(new_n19496_), .ZN(new_n19526_));
  NAND2_X1   g18524(.A1(new_n19501_), .A2(new_n19495_), .ZN(new_n19527_));
  NAND2_X1   g18525(.A1(new_n19507_), .A2(new_n19527_), .ZN(new_n19528_));
  INV_X1     g18526(.I(new_n19426_), .ZN(new_n19529_));
  NOR2_X1    g18527(.A1(new_n19328_), .A2(new_n19431_), .ZN(new_n19530_));
  NAND2_X1   g18528(.A1(new_n19427_), .A2(new_n19432_), .ZN(new_n19531_));
  NOR3_X1    g18529(.A1(new_n19529_), .A2(new_n19530_), .A3(new_n19531_), .ZN(new_n19532_));
  NAND2_X1   g18530(.A1(new_n19433_), .A2(new_n19435_), .ZN(new_n19533_));
  INV_X1     g18531(.I(new_n19533_), .ZN(new_n19534_));
  NOR2_X1    g18532(.A1(new_n19417_), .A2(new_n19534_), .ZN(new_n19535_));
  OAI21_X1   g18533(.A1(new_n19442_), .A2(new_n19532_), .B(new_n19535_), .ZN(new_n19536_));
  OAI21_X1   g18534(.A1(new_n19442_), .A2(new_n19532_), .B(new_n19533_), .ZN(new_n19537_));
  NAND2_X1   g18535(.A1(new_n19537_), .A2(new_n19417_), .ZN(new_n19538_));
  NAND2_X1   g18536(.A1(new_n19538_), .A2(new_n19536_), .ZN(new_n19539_));
  AOI21_X1   g18537(.A1(new_n19528_), .A2(new_n19526_), .B(new_n19539_), .ZN(new_n19540_));
  INV_X1     g18538(.I(new_n19540_), .ZN(new_n19541_));
  AOI22_X1   g18539(.A1(new_n19538_), .A2(new_n19536_), .B1(new_n19496_), .B2(new_n19503_), .ZN(new_n19542_));
  NAND2_X1   g18540(.A1(new_n19528_), .A2(new_n19542_), .ZN(new_n19543_));
  AOI21_X1   g18541(.A1(new_n19541_), .A2(new_n19543_), .B(new_n19525_), .ZN(new_n19544_));
  NOR2_X1    g18542(.A1(new_n19511_), .A2(new_n19544_), .ZN(new_n19545_));
  NAND2_X1   g18543(.A1(new_n19528_), .A2(new_n19526_), .ZN(new_n19546_));
  NAND2_X1   g18544(.A1(new_n19546_), .A2(new_n19536_), .ZN(new_n19547_));
  NAND2_X1   g18545(.A1(new_n19547_), .A2(new_n19538_), .ZN(new_n19548_));
  NAND3_X1   g18546(.A1(new_n19541_), .A2(new_n19525_), .A3(new_n19543_), .ZN(new_n19549_));
  NAND2_X1   g18547(.A1(new_n19549_), .A2(new_n19548_), .ZN(new_n19550_));
  NAND2_X1   g18548(.A1(new_n19414_), .A2(new_n19509_), .ZN(new_n19551_));
  NAND2_X1   g18549(.A1(new_n19490_), .A2(new_n19481_), .ZN(new_n19552_));
  NOR3_X1    g18550(.A1(new_n19482_), .A2(new_n19488_), .A3(new_n19480_), .ZN(new_n19553_));
  AOI22_X1   g18551(.A1(new_n19518_), .A2(new_n19552_), .B1(new_n19553_), .B2(new_n19517_), .ZN(new_n19554_));
  NAND3_X1   g18552(.A1(new_n19507_), .A2(new_n19526_), .A3(new_n19527_), .ZN(new_n19555_));
  NAND3_X1   g18553(.A1(new_n19463_), .A2(new_n19555_), .A3(new_n19554_), .ZN(new_n19556_));
  NAND2_X1   g18554(.A1(new_n19551_), .A2(new_n19556_), .ZN(new_n19557_));
  INV_X1     g18555(.I(new_n19543_), .ZN(new_n19558_));
  OAI21_X1   g18556(.A1(new_n19558_), .A2(new_n19540_), .B(new_n19524_), .ZN(new_n19559_));
  NOR3_X1    g18557(.A1(new_n19558_), .A2(new_n19524_), .A3(new_n19540_), .ZN(new_n19560_));
  AOI21_X1   g18558(.A1(new_n19557_), .A2(new_n19559_), .B(new_n19560_), .ZN(new_n19561_));
  OAI22_X1   g18559(.A1(new_n19561_), .A2(new_n19548_), .B1(new_n19545_), .B2(new_n19550_), .ZN(new_n19562_));
  INV_X1     g18560(.I(new_n17690_), .ZN(new_n19563_));
  INV_X1     g18561(.I(new_n17676_), .ZN(new_n19564_));
  AOI21_X1   g18562(.A1(new_n19564_), .A2(new_n17677_), .B(new_n10692_), .ZN(new_n19565_));
  NAND3_X1   g18563(.A1(new_n17680_), .A2(new_n17675_), .A3(new_n17681_), .ZN(new_n19566_));
  AOI21_X1   g18564(.A1(new_n19566_), .A2(new_n10687_), .B(new_n10693_), .ZN(new_n19567_));
  NOR3_X1    g18565(.A1(new_n19565_), .A2(new_n19567_), .A3(new_n17674_), .ZN(new_n19568_));
  AOI21_X1   g18566(.A1(new_n17679_), .A2(new_n17683_), .B(new_n17673_), .ZN(new_n19569_));
  OAI21_X1   g18567(.A1(new_n19569_), .A2(new_n19568_), .B(new_n19563_), .ZN(new_n19570_));
  NOR3_X1    g18568(.A1(new_n19565_), .A2(new_n19567_), .A3(new_n17673_), .ZN(new_n19571_));
  OAI21_X1   g18569(.A1(new_n17684_), .A2(new_n19571_), .B(new_n17690_), .ZN(new_n19572_));
  INV_X1     g18570(.I(\A[1000] ), .ZN(new_n19573_));
  NOR3_X1    g18571(.A1(new_n17671_), .A2(new_n17667_), .A3(new_n17669_), .ZN(new_n19574_));
  OAI21_X1   g18572(.A1(new_n17671_), .A2(new_n17669_), .B(new_n17667_), .ZN(new_n19575_));
  INV_X1     g18573(.I(new_n19575_), .ZN(new_n19576_));
  NOR2_X1    g18574(.A1(new_n19576_), .A2(new_n19574_), .ZN(new_n19577_));
  NOR2_X1    g18575(.A1(new_n19577_), .A2(new_n19573_), .ZN(new_n19578_));
  INV_X1     g18576(.I(new_n19578_), .ZN(new_n19579_));
  AOI21_X1   g18577(.A1(new_n19570_), .A2(new_n19572_), .B(new_n19579_), .ZN(new_n19580_));
  OAI21_X1   g18578(.A1(new_n17663_), .A2(new_n17662_), .B(new_n16959_), .ZN(new_n19581_));
  NAND3_X1   g18579(.A1(new_n17656_), .A2(new_n17657_), .A3(new_n16960_), .ZN(new_n19582_));
  NAND2_X1   g18580(.A1(new_n19581_), .A2(new_n19582_), .ZN(new_n19583_));
  NAND3_X1   g18581(.A1(new_n17695_), .A2(new_n17652_), .A3(new_n19583_), .ZN(new_n19584_));
  NOR3_X1    g18582(.A1(new_n17693_), .A2(new_n17694_), .A3(new_n10695_), .ZN(new_n19585_));
  OAI21_X1   g18583(.A1(new_n19585_), .A2(new_n17651_), .B(new_n17665_), .ZN(new_n19586_));
  NAND3_X1   g18584(.A1(new_n19586_), .A2(new_n19584_), .A3(new_n17692_), .ZN(new_n19587_));
  OAI21_X1   g18585(.A1(new_n19565_), .A2(new_n19567_), .B(new_n17673_), .ZN(new_n19588_));
  OAI21_X1   g18586(.A1(new_n19563_), .A2(new_n19571_), .B(new_n19588_), .ZN(new_n19589_));
  NOR3_X1    g18587(.A1(new_n19585_), .A2(new_n17651_), .A3(new_n17665_), .ZN(new_n19590_));
  AOI21_X1   g18588(.A1(new_n17695_), .A2(new_n17652_), .B(new_n19583_), .ZN(new_n19591_));
  OAI21_X1   g18589(.A1(new_n19590_), .A2(new_n19591_), .B(new_n19589_), .ZN(new_n19592_));
  NAND3_X1   g18590(.A1(new_n19592_), .A2(new_n19587_), .A3(new_n19580_), .ZN(new_n19593_));
  NOR2_X1    g18591(.A1(new_n11875_), .A2(new_n11874_), .ZN(new_n19594_));
  OAI22_X1   g18592(.A1(new_n11877_), .A2(new_n11878_), .B1(new_n19594_), .B2(new_n18646_), .ZN(new_n19595_));
  NAND4_X1   g18593(.A1(new_n10700_), .A2(new_n11866_), .A3(new_n11872_), .A4(new_n10677_), .ZN(new_n19596_));
  AOI21_X1   g18594(.A1(new_n19595_), .A2(new_n19596_), .B(new_n17647_), .ZN(new_n19597_));
  AOI22_X1   g18595(.A1(new_n17644_), .A2(new_n17645_), .B1(new_n16943_), .B2(new_n19513_), .ZN(new_n19598_));
  NOR3_X1    g18596(.A1(new_n17637_), .A2(new_n17630_), .A3(new_n16962_), .ZN(new_n19599_));
  NOR2_X1    g18597(.A1(new_n19598_), .A2(new_n19599_), .ZN(new_n19600_));
  NOR3_X1    g18598(.A1(new_n11873_), .A2(new_n11879_), .A3(new_n19600_), .ZN(new_n19601_));
  NOR3_X1    g18599(.A1(new_n17697_), .A2(new_n19597_), .A3(new_n19601_), .ZN(new_n19602_));
  NOR2_X1    g18600(.A1(new_n19585_), .A2(new_n19583_), .ZN(new_n19603_));
  OAI21_X1   g18601(.A1(new_n19585_), .A2(new_n17651_), .B(new_n19583_), .ZN(new_n19604_));
  AOI22_X1   g18602(.A1(new_n19604_), .A2(new_n19589_), .B1(new_n19603_), .B2(new_n17695_), .ZN(new_n19605_));
  OAI21_X1   g18603(.A1(new_n11873_), .A2(new_n11879_), .B(new_n19600_), .ZN(new_n19606_));
  NAND3_X1   g18604(.A1(new_n19595_), .A2(new_n19596_), .A3(new_n17647_), .ZN(new_n19607_));
  AOI21_X1   g18605(.A1(new_n19606_), .A2(new_n19607_), .B(new_n19605_), .ZN(new_n19608_));
  NOR3_X1    g18606(.A1(new_n19608_), .A2(new_n19602_), .A3(new_n19593_), .ZN(new_n19609_));
  OAI21_X1   g18607(.A1(new_n18057_), .A2(new_n18058_), .B(new_n18056_), .ZN(new_n19610_));
  NAND3_X1   g18608(.A1(new_n18043_), .A2(new_n18052_), .A3(new_n17702_), .ZN(new_n19611_));
  NAND2_X1   g18609(.A1(new_n19610_), .A2(new_n19611_), .ZN(new_n19612_));
  NAND3_X1   g18610(.A1(new_n18650_), .A2(new_n18655_), .A3(new_n19612_), .ZN(new_n19613_));
  NAND2_X1   g18611(.A1(new_n11876_), .A2(new_n18653_), .ZN(new_n19614_));
  AOI22_X1   g18612(.A1(new_n19614_), .A2(new_n19158_), .B1(new_n18651_), .B2(new_n18652_), .ZN(new_n19615_));
  NOR3_X1    g18613(.A1(new_n19159_), .A2(new_n18635_), .A3(new_n18644_), .ZN(new_n19616_));
  OAI21_X1   g18614(.A1(new_n19616_), .A2(new_n19615_), .B(new_n18060_), .ZN(new_n19617_));
  NAND3_X1   g18615(.A1(new_n17699_), .A2(new_n19617_), .A3(new_n19613_), .ZN(new_n19618_));
  NAND3_X1   g18616(.A1(new_n19595_), .A2(new_n19596_), .A3(new_n19600_), .ZN(new_n19619_));
  AOI21_X1   g18617(.A1(new_n19595_), .A2(new_n19596_), .B(new_n19600_), .ZN(new_n19620_));
  OAI21_X1   g18618(.A1(new_n19605_), .A2(new_n19620_), .B(new_n19619_), .ZN(new_n19621_));
  NOR3_X1    g18619(.A1(new_n19616_), .A2(new_n19615_), .A3(new_n18060_), .ZN(new_n19622_));
  AOI21_X1   g18620(.A1(new_n18650_), .A2(new_n18655_), .B(new_n19612_), .ZN(new_n19623_));
  OAI21_X1   g18621(.A1(new_n19622_), .A2(new_n19623_), .B(new_n19621_), .ZN(new_n19624_));
  NAND3_X1   g18622(.A1(new_n19624_), .A2(new_n19609_), .A3(new_n19618_), .ZN(new_n19625_));
  OAI21_X1   g18623(.A1(new_n19163_), .A2(new_n19164_), .B(new_n19166_), .ZN(new_n19626_));
  NAND3_X1   g18624(.A1(new_n19403_), .A2(new_n19148_), .A3(new_n19156_), .ZN(new_n19627_));
  AOI21_X1   g18625(.A1(new_n19626_), .A2(new_n19627_), .B(new_n18843_), .ZN(new_n19628_));
  AOI21_X1   g18626(.A1(new_n18840_), .A2(new_n18841_), .B(new_n18839_), .ZN(new_n19629_));
  NOR3_X1    g18627(.A1(new_n18835_), .A2(new_n18828_), .A3(new_n18661_), .ZN(new_n19630_));
  NOR2_X1    g18628(.A1(new_n19629_), .A2(new_n19630_), .ZN(new_n19631_));
  NOR3_X1    g18629(.A1(new_n19162_), .A2(new_n19167_), .A3(new_n19631_), .ZN(new_n19632_));
  NOR3_X1    g18630(.A1(new_n18658_), .A2(new_n19628_), .A3(new_n19632_), .ZN(new_n19633_));
  OAI21_X1   g18631(.A1(new_n19616_), .A2(new_n19615_), .B(new_n19612_), .ZN(new_n19634_));
  NOR3_X1    g18632(.A1(new_n19616_), .A2(new_n19615_), .A3(new_n19612_), .ZN(new_n19635_));
  AOI21_X1   g18633(.A1(new_n19621_), .A2(new_n19634_), .B(new_n19635_), .ZN(new_n19636_));
  OAI21_X1   g18634(.A1(new_n19162_), .A2(new_n19167_), .B(new_n19631_), .ZN(new_n19637_));
  NAND3_X1   g18635(.A1(new_n19626_), .A2(new_n19627_), .A3(new_n18843_), .ZN(new_n19638_));
  AOI21_X1   g18636(.A1(new_n19637_), .A2(new_n19638_), .B(new_n19636_), .ZN(new_n19639_));
  NOR3_X1    g18637(.A1(new_n19639_), .A2(new_n19625_), .A3(new_n19633_), .ZN(new_n19640_));
  OAI22_X1   g18638(.A1(new_n19249_), .A2(new_n19250_), .B1(new_n19516_), .B2(new_n19171_), .ZN(new_n19641_));
  NAND3_X1   g18639(.A1(new_n19173_), .A2(new_n19244_), .A3(new_n19234_), .ZN(new_n19642_));
  NAND2_X1   g18640(.A1(new_n19641_), .A2(new_n19642_), .ZN(new_n19643_));
  NAND3_X1   g18641(.A1(new_n19407_), .A2(new_n19411_), .A3(new_n19643_), .ZN(new_n19644_));
  NAND2_X1   g18642(.A1(new_n19166_), .A2(new_n19408_), .ZN(new_n19645_));
  AOI22_X1   g18643(.A1(new_n19645_), .A2(new_n19405_), .B1(new_n19393_), .B2(new_n19400_), .ZN(new_n19646_));
  NOR2_X1    g18644(.A1(new_n19401_), .A2(new_n19406_), .ZN(new_n19647_));
  OAI21_X1   g18645(.A1(new_n19647_), .A2(new_n19646_), .B(new_n19252_), .ZN(new_n19648_));
  NAND3_X1   g18646(.A1(new_n19170_), .A2(new_n19648_), .A3(new_n19644_), .ZN(new_n19649_));
  AOI21_X1   g18647(.A1(new_n19626_), .A2(new_n19627_), .B(new_n19631_), .ZN(new_n19650_));
  NOR2_X1    g18648(.A1(new_n19636_), .A2(new_n19650_), .ZN(new_n19651_));
  NOR3_X1    g18649(.A1(new_n19647_), .A2(new_n19646_), .A3(new_n19252_), .ZN(new_n19652_));
  AOI21_X1   g18650(.A1(new_n19407_), .A2(new_n19411_), .B(new_n19643_), .ZN(new_n19653_));
  OAI22_X1   g18651(.A1(new_n19651_), .A2(new_n19169_), .B1(new_n19652_), .B2(new_n19653_), .ZN(new_n19654_));
  NAND3_X1   g18652(.A1(new_n19640_), .A2(new_n19654_), .A3(new_n19649_), .ZN(new_n19655_));
  AOI21_X1   g18653(.A1(new_n19463_), .A2(new_n19555_), .B(new_n19493_), .ZN(new_n19656_));
  NOR3_X1    g18654(.A1(new_n19494_), .A2(new_n19508_), .A3(new_n19554_), .ZN(new_n19657_));
  NOR3_X1    g18655(.A1(new_n19414_), .A2(new_n19657_), .A3(new_n19656_), .ZN(new_n19658_));
  NAND3_X1   g18656(.A1(new_n19626_), .A2(new_n19627_), .A3(new_n19631_), .ZN(new_n19659_));
  OAI21_X1   g18657(.A1(new_n19636_), .A2(new_n19650_), .B(new_n19659_), .ZN(new_n19660_));
  OAI21_X1   g18658(.A1(new_n19647_), .A2(new_n19646_), .B(new_n19643_), .ZN(new_n19661_));
  NAND2_X1   g18659(.A1(new_n19660_), .A2(new_n19661_), .ZN(new_n19662_));
  OAI21_X1   g18660(.A1(new_n19494_), .A2(new_n19508_), .B(new_n19554_), .ZN(new_n19663_));
  NAND3_X1   g18661(.A1(new_n19463_), .A2(new_n19555_), .A3(new_n19493_), .ZN(new_n19664_));
  AOI22_X1   g18662(.A1(new_n19662_), .A2(new_n19413_), .B1(new_n19663_), .B2(new_n19664_), .ZN(new_n19665_));
  NOR3_X1    g18663(.A1(new_n19655_), .A2(new_n19665_), .A3(new_n19658_), .ZN(new_n19666_));
  OAI21_X1   g18664(.A1(new_n19558_), .A2(new_n19540_), .B(new_n19525_), .ZN(new_n19667_));
  NAND3_X1   g18665(.A1(new_n19541_), .A2(new_n19524_), .A3(new_n19543_), .ZN(new_n19668_));
  NAND2_X1   g18666(.A1(new_n19668_), .A2(new_n19667_), .ZN(new_n19669_));
  NAND2_X1   g18667(.A1(new_n19669_), .A2(new_n19557_), .ZN(new_n19670_));
  NAND4_X1   g18668(.A1(new_n19668_), .A2(new_n19667_), .A3(new_n19551_), .A4(new_n19556_), .ZN(new_n19671_));
  NAND3_X1   g18669(.A1(new_n19670_), .A2(new_n19666_), .A3(new_n19671_), .ZN(new_n19672_));
  NAND3_X1   g18670(.A1(new_n17679_), .A2(new_n17683_), .A3(new_n17673_), .ZN(new_n19673_));
  OAI21_X1   g18671(.A1(new_n19565_), .A2(new_n19567_), .B(new_n17674_), .ZN(new_n19674_));
  AOI21_X1   g18672(.A1(new_n19674_), .A2(new_n19673_), .B(new_n17690_), .ZN(new_n19675_));
  AOI21_X1   g18673(.A1(new_n19588_), .A2(new_n17691_), .B(new_n19563_), .ZN(new_n19676_));
  OAI21_X1   g18674(.A1(new_n19676_), .A2(new_n19675_), .B(new_n19578_), .ZN(new_n19677_));
  NOR3_X1    g18675(.A1(new_n19590_), .A2(new_n19591_), .A3(new_n19589_), .ZN(new_n19678_));
  AOI21_X1   g18676(.A1(new_n19586_), .A2(new_n19584_), .B(new_n17692_), .ZN(new_n19679_));
  NOR3_X1    g18677(.A1(new_n19678_), .A2(new_n19679_), .A3(new_n19677_), .ZN(new_n19680_));
  NAND3_X1   g18678(.A1(new_n19605_), .A2(new_n19606_), .A3(new_n19607_), .ZN(new_n19681_));
  OAI21_X1   g18679(.A1(new_n19597_), .A2(new_n19601_), .B(new_n17697_), .ZN(new_n19682_));
  NAND3_X1   g18680(.A1(new_n19682_), .A2(new_n19681_), .A3(new_n19680_), .ZN(new_n19683_));
  NOR3_X1    g18681(.A1(new_n19621_), .A2(new_n19622_), .A3(new_n19623_), .ZN(new_n19684_));
  NAND2_X1   g18682(.A1(new_n17697_), .A2(new_n17698_), .ZN(new_n19685_));
  AOI22_X1   g18683(.A1(new_n19617_), .A2(new_n19613_), .B1(new_n19685_), .B2(new_n19619_), .ZN(new_n19686_));
  NOR3_X1    g18684(.A1(new_n19683_), .A2(new_n19686_), .A3(new_n19684_), .ZN(new_n19687_));
  NAND3_X1   g18685(.A1(new_n19636_), .A2(new_n19637_), .A3(new_n19638_), .ZN(new_n19688_));
  OAI21_X1   g18686(.A1(new_n19628_), .A2(new_n19632_), .B(new_n18658_), .ZN(new_n19689_));
  NAND3_X1   g18687(.A1(new_n19687_), .A2(new_n19689_), .A3(new_n19688_), .ZN(new_n19690_));
  NOR3_X1    g18688(.A1(new_n19660_), .A2(new_n19652_), .A3(new_n19653_), .ZN(new_n19691_));
  AOI21_X1   g18689(.A1(new_n19644_), .A2(new_n19648_), .B(new_n19170_), .ZN(new_n19692_));
  NOR2_X1    g18690(.A1(new_n19692_), .A2(new_n19691_), .ZN(new_n19693_));
  OAI21_X1   g18691(.A1(new_n19639_), .A2(new_n19633_), .B(new_n19625_), .ZN(new_n19694_));
  OAI21_X1   g18692(.A1(new_n19608_), .A2(new_n19602_), .B(new_n19593_), .ZN(new_n19695_));
  AOI21_X1   g18693(.A1(new_n19592_), .A2(new_n19587_), .B(new_n19580_), .ZN(new_n19696_));
  NOR3_X1    g18694(.A1(new_n19676_), .A2(new_n19675_), .A3(new_n19579_), .ZN(new_n19697_));
  AOI21_X1   g18695(.A1(new_n19570_), .A2(new_n19572_), .B(new_n19578_), .ZN(new_n19698_));
  NOR2_X1    g18696(.A1(new_n19698_), .A2(new_n19697_), .ZN(new_n19699_));
  OAI21_X1   g18697(.A1(new_n19680_), .A2(new_n19696_), .B(new_n19699_), .ZN(new_n19700_));
  NAND3_X1   g18698(.A1(new_n19695_), .A2(new_n19683_), .A3(new_n19700_), .ZN(new_n19701_));
  AOI21_X1   g18699(.A1(new_n19618_), .A2(new_n19624_), .B(new_n19609_), .ZN(new_n19702_));
  OAI21_X1   g18700(.A1(new_n19702_), .A2(new_n19687_), .B(new_n19701_), .ZN(new_n19703_));
  NAND4_X1   g18701(.A1(new_n19693_), .A2(new_n19690_), .A3(new_n19694_), .A4(new_n19703_), .ZN(new_n19704_));
  NOR3_X1    g18702(.A1(new_n19647_), .A2(new_n19646_), .A3(new_n19643_), .ZN(new_n19705_));
  AOI21_X1   g18703(.A1(new_n19660_), .A2(new_n19661_), .B(new_n19705_), .ZN(new_n19706_));
  NAND3_X1   g18704(.A1(new_n19706_), .A2(new_n19663_), .A3(new_n19664_), .ZN(new_n19707_));
  OAI21_X1   g18705(.A1(new_n19656_), .A2(new_n19657_), .B(new_n19414_), .ZN(new_n19708_));
  AOI22_X1   g18706(.A1(new_n19708_), .A2(new_n19707_), .B1(new_n19693_), .B2(new_n19640_), .ZN(new_n19709_));
  NOR3_X1    g18707(.A1(new_n19709_), .A2(new_n19666_), .A3(new_n19704_), .ZN(new_n19710_));
  NAND2_X1   g18708(.A1(new_n19708_), .A2(new_n19707_), .ZN(new_n19711_));
  AOI21_X1   g18709(.A1(new_n19667_), .A2(new_n19668_), .B(new_n19511_), .ZN(new_n19712_));
  INV_X1     g18710(.I(new_n19509_), .ZN(new_n19713_));
  NOR2_X1    g18711(.A1(new_n19713_), .A2(new_n19706_), .ZN(new_n19714_));
  AOI21_X1   g18712(.A1(new_n19541_), .A2(new_n19543_), .B(new_n19524_), .ZN(new_n19715_));
  NAND2_X1   g18713(.A1(new_n19543_), .A2(new_n19524_), .ZN(new_n19716_));
  OAI21_X1   g18714(.A1(new_n19716_), .A2(new_n19540_), .B(new_n19556_), .ZN(new_n19717_));
  NOR3_X1    g18715(.A1(new_n19714_), .A2(new_n19715_), .A3(new_n19717_), .ZN(new_n19718_));
  OAI22_X1   g18716(.A1(new_n19712_), .A2(new_n19718_), .B1(new_n19655_), .B2(new_n19711_), .ZN(new_n19719_));
  NAND4_X1   g18717(.A1(new_n19562_), .A2(new_n19672_), .A3(new_n19719_), .A4(new_n19710_), .ZN(new_n19720_));
  NAND2_X1   g18718(.A1(new_n19557_), .A2(new_n19559_), .ZN(new_n19721_));
  INV_X1     g18719(.I(new_n19548_), .ZN(new_n19722_));
  NOR4_X1    g18720(.A1(new_n19712_), .A2(new_n19718_), .A3(new_n19655_), .A4(new_n19711_), .ZN(new_n19723_));
  AOI21_X1   g18721(.A1(new_n19721_), .A2(new_n19549_), .B(new_n19722_), .ZN(new_n19724_));
  INV_X1     g18722(.I(new_n19724_), .ZN(new_n19725_));
  OAI21_X1   g18723(.A1(new_n19511_), .A2(new_n19544_), .B(new_n19549_), .ZN(new_n19726_));
  NAND2_X1   g18724(.A1(new_n19726_), .A2(new_n19548_), .ZN(new_n19727_));
  NAND3_X1   g18725(.A1(new_n19562_), .A2(new_n19723_), .A3(new_n19727_), .ZN(new_n19728_));
  NOR3_X1    g18726(.A1(new_n19690_), .A2(new_n19692_), .A3(new_n19691_), .ZN(new_n19729_));
  NAND2_X1   g18727(.A1(new_n19729_), .A2(new_n19548_), .ZN(new_n19730_));
  NOR4_X1    g18728(.A1(new_n19712_), .A2(new_n19718_), .A3(new_n19730_), .A4(new_n19711_), .ZN(new_n19731_));
  NAND3_X1   g18729(.A1(new_n19562_), .A2(new_n19731_), .A3(new_n19726_), .ZN(new_n19732_));
  NAND4_X1   g18730(.A1(new_n19720_), .A2(new_n19728_), .A3(new_n19732_), .A4(new_n19725_), .ZN(new_n19733_));
  INV_X1     g18731(.I(new_n19733_), .ZN(new_n19734_));
  NOR2_X1    g18732(.A1(new_n19665_), .A2(new_n19658_), .ZN(new_n19735_));
  AOI21_X1   g18733(.A1(new_n19688_), .A2(new_n19689_), .B(new_n19687_), .ZN(new_n19736_));
  AOI21_X1   g18734(.A1(new_n19682_), .A2(new_n19681_), .B(new_n19680_), .ZN(new_n19737_));
  OAI21_X1   g18735(.A1(new_n19678_), .A2(new_n19679_), .B(new_n19677_), .ZN(new_n19738_));
  OR2_X2     g18736(.A1(new_n19698_), .A2(new_n19697_), .Z(new_n19739_));
  AOI21_X1   g18737(.A1(new_n19738_), .A2(new_n19593_), .B(new_n19739_), .ZN(new_n19740_));
  NOR3_X1    g18738(.A1(new_n19609_), .A2(new_n19737_), .A3(new_n19740_), .ZN(new_n19741_));
  OAI21_X1   g18739(.A1(new_n19684_), .A2(new_n19686_), .B(new_n19683_), .ZN(new_n19742_));
  AOI21_X1   g18740(.A1(new_n19625_), .A2(new_n19742_), .B(new_n19741_), .ZN(new_n19743_));
  NOR3_X1    g18741(.A1(new_n19736_), .A2(new_n19743_), .A3(new_n19640_), .ZN(new_n19744_));
  OAI21_X1   g18742(.A1(new_n19691_), .A2(new_n19692_), .B(new_n19690_), .ZN(new_n19745_));
  NAND4_X1   g18743(.A1(new_n19735_), .A2(new_n19655_), .A3(new_n19744_), .A4(new_n19745_), .ZN(new_n19746_));
  NAND2_X1   g18744(.A1(new_n19672_), .A2(new_n19719_), .ZN(new_n19747_));
  INV_X1     g18745(.I(new_n19550_), .ZN(new_n19748_));
  AOI22_X1   g18746(.A1(new_n19748_), .A2(new_n19721_), .B1(new_n19722_), .B2(new_n19726_), .ZN(new_n19749_));
  AOI21_X1   g18747(.A1(new_n19670_), .A2(new_n19671_), .B(new_n19666_), .ZN(new_n19750_));
  NOR4_X1    g18748(.A1(new_n19749_), .A2(new_n19750_), .A3(new_n19723_), .A4(new_n19746_), .ZN(new_n19751_));
  NOR2_X1    g18749(.A1(new_n19709_), .A2(new_n19666_), .ZN(new_n19752_));
  NOR2_X1    g18750(.A1(new_n19736_), .A2(new_n19640_), .ZN(new_n19753_));
  NAND2_X1   g18751(.A1(new_n19695_), .A2(new_n19683_), .ZN(new_n19754_));
  NAND2_X1   g18752(.A1(new_n19738_), .A2(new_n19593_), .ZN(new_n19755_));
  INV_X1     g18753(.I(new_n19577_), .ZN(new_n19756_));
  NOR2_X1    g18754(.A1(new_n19574_), .A2(new_n19573_), .ZN(new_n19757_));
  AOI22_X1   g18755(.A1(new_n19756_), .A2(new_n19573_), .B1(new_n19575_), .B2(new_n19757_), .ZN(new_n19758_));
  MUX2_X1    g18756(.I0(new_n19758_), .I1(new_n19755_), .S(new_n19739_), .Z(new_n19759_));
  AOI21_X1   g18757(.A1(new_n19759_), .A2(new_n19700_), .B(new_n19754_), .ZN(new_n19760_));
  AOI21_X1   g18758(.A1(new_n19695_), .A2(new_n19683_), .B(new_n19700_), .ZN(new_n19761_));
  NOR3_X1    g18759(.A1(new_n19759_), .A2(new_n19761_), .A3(new_n19741_), .ZN(new_n19762_));
  OAI21_X1   g18760(.A1(new_n19762_), .A2(new_n19760_), .B(new_n19701_), .ZN(new_n19763_));
  NAND3_X1   g18761(.A1(new_n19625_), .A2(new_n19742_), .A3(new_n19741_), .ZN(new_n19764_));
  NAND3_X1   g18762(.A1(new_n19694_), .A2(new_n19703_), .A3(new_n19690_), .ZN(new_n19765_));
  OAI21_X1   g18763(.A1(new_n19640_), .A2(new_n19736_), .B(new_n19743_), .ZN(new_n19766_));
  NAND2_X1   g18764(.A1(new_n19766_), .A2(new_n19765_), .ZN(new_n19767_));
  NAND3_X1   g18765(.A1(new_n19767_), .A2(new_n19763_), .A3(new_n19764_), .ZN(new_n19768_));
  NAND3_X1   g18766(.A1(new_n19768_), .A2(new_n19753_), .A3(new_n19703_), .ZN(new_n19770_));
  INV_X1     g18767(.I(new_n19745_), .ZN(new_n19771_));
  NOR2_X1    g18768(.A1(new_n19771_), .A2(new_n19729_), .ZN(new_n19772_));
  NAND2_X1   g18769(.A1(new_n19772_), .A2(new_n19765_), .ZN(new_n19773_));
  OAI21_X1   g18770(.A1(new_n19709_), .A2(new_n19666_), .B(new_n19704_), .ZN(new_n19774_));
  NAND2_X1   g18771(.A1(new_n19774_), .A2(new_n19746_), .ZN(new_n19775_));
  NAND3_X1   g18772(.A1(new_n19770_), .A2(new_n19775_), .A3(new_n19773_), .ZN(new_n19776_));
  INV_X1     g18773(.I(new_n19704_), .ZN(new_n19777_));
  NAND4_X1   g18774(.A1(new_n19672_), .A2(new_n19719_), .A3(new_n19777_), .A4(new_n19752_), .ZN(new_n19779_));
  AOI21_X1   g18775(.A1(new_n19776_), .A2(new_n19752_), .B(new_n19779_), .ZN(new_n19780_));
  NOR4_X1    g18776(.A1(new_n19780_), .A2(new_n19746_), .A3(new_n19747_), .A4(new_n19751_), .ZN(new_n19783_));
  XOR2_X1    g18777(.A1(new_n19749_), .A2(new_n19672_), .Z(new_n19787_));
  NAND4_X1   g18778(.A1(new_n19562_), .A2(new_n19672_), .A3(new_n19719_), .A4(new_n19710_), .ZN(new_n19789_));
  NOR2_X1    g18779(.A1(new_n19789_), .A2(new_n19724_), .ZN(new_n19790_));
  NOR2_X1    g18780(.A1(new_n19730_), .A2(new_n19711_), .ZN(new_n19791_));
  NAND2_X1   g18781(.A1(new_n19791_), .A2(new_n19670_), .ZN(new_n19792_));
  NOR4_X1    g18782(.A1(new_n19792_), .A2(new_n19749_), .A3(new_n19561_), .A4(new_n19718_), .ZN(new_n19793_));
  NAND4_X1   g18783(.A1(new_n19727_), .A2(new_n19666_), .A3(new_n19670_), .A4(new_n19671_), .ZN(new_n19794_));
  OAI21_X1   g18784(.A1(new_n19794_), .A2(new_n19749_), .B(new_n19725_), .ZN(new_n19795_));
  OAI21_X1   g18785(.A1(new_n19795_), .A2(new_n19751_), .B(new_n19793_), .ZN(new_n19796_));
  AOI21_X1   g18786(.A1(new_n19796_), .A2(new_n19733_), .B(new_n19790_), .ZN(new_n19797_));
  OAI21_X1   g18787(.A1(new_n19783_), .A2(new_n19787_), .B(new_n19797_), .ZN(new_n19798_));
  NAND2_X1   g18788(.A1(new_n19798_), .A2(new_n19734_), .ZN(maj));
endmodule


