// Benchmark "testing" written by ABC on Fri Feb 25 15:12:55 2022

module g625 ( 
    B9278, B9277, B9276, B9275, B9274, B9245, B9244, B9243, B9242, B9241,
    B9212, B9211, B9210, B9209, B9208, B9179, B9178, B9177, B9176, B9175,
    B9146, B9145, B9144, B9143, B9142, B9113, B9112, B9111, B9110, B9109,
    B9080, B9079, B9078, B9077, B9076, B9047, B9046, B9045, B9044, B9043,
    B9014, B9013, B9012, B9011, B9010, B8981, B8980, B8979, B8978, B8977,
    B8948, B8947, B8946, B8945, B8944, B8915, B8914, B8913, B8912, B8911,
    B8882, B8881, B8880, B8879, B8878, B8849, B8848, B8847, B8846, B8845,
    B8816, B8815, B8814, B8813, B8812, B8783, B8782, B8781, B8780, B8779,
    B8750, B8749, B8748, B8747, B8746, B8717, B8716, B8715, B8714, B8713,
    B8684, B8683, B8682, B8681, B8680, B8651, B8650, B8649, B8648, B8647,
    B8618, B8617, B8616, B8615, B8614, B8585, B8584, B8583, B8582, B8581,
    B8552, B8551, B8550, B8549, B8548, B8519, B8518, B8517, B8516, B8515,
    B8486, B8485, B8484, B8483, B8482, B8453, B8452, B8451, B8450, B8449,
    B8420, B8419, B8418, B8417, B8416, B8387, B8386, B8385, B8384, B8383,
    B8354, B8353, B8352, B8351, B8350, B8321, B8320, B8319, B8318, B8317,
    B8288, B8287, B8286, B8285, B8284, B8255, B8254, B8253, B8252, B8251,
    B8222, B8221, B8220, B8219, B8218, B8189, B8188, B8187, B8186, B8185,
    B8156, B8155, B8154, B8153, B8152, B8123, B8122, B8121, B8120, B8119,
    B8090, B8089, B8088, B8087, B8086, B8057, B8056, B8055, B8054, B8053,
    B8024, B8023, B8022, B8021, B8020, B7991, B7990, B7989, B7988, B7987,
    B7958, B7957, B7956, B7955, B7954, B7925, B7924, B7923, B7922, B7921,
    B7892, B7891, B7890, B7889, B7888, B7859, B7858, B7857, B7856, B7855,
    B7826, B7825, B7824, B7823, B7822, B7793, B7792, B7791, B7790, B7789,
    B7760, B7759, B7758, B7757, B7756, B7727, B7726, B7725, B7724, B7723,
    B7694, B7693, B7692, B7691, B7690, B7661, B7660, B7659, B7658, B7657,
    B7628, B7627, B7626, B7625, B7624, B7595, B7594, B7593, B7592, B7591,
    B7562, B7561, B7560, B7559, B7558, B7529, B7528, B7527, B7526, B7525,
    B7496, B7495, B7494, B7493, B7492, B7463, B7462, B7461, B7460, B7459,
    B7430, B7429, B7428, B7427, B7426, B7397, B7396, B7395, B7394, B7393,
    B7364, B7363, B7362, B7361, B7360, B7331, B7330, B7329, B7328, B7327,
    B7298, B7297, B7296, B7295, B7294, B7265, B7264, B7263, B7262, B7261,
    B7232, B7231, B7230, B7229, B7228, B7199, B7198, B7197, B7196, B7195,
    B7166, B7165, B7164, B7163, B7162, B7133, B7132, B7131, B7130, B7129,
    B7100, B7099, B7098, B7097, B7096, B7067, B7066, B7065, B7064, B7063,
    B7034, B7033, B7032, B7031, B7030, B7001, B7000, B6999, B6998, B6997,
    B6968, B6967, B6966, B6965, B6964, B6935, B6934, B6933, B6932, B6931,
    B6902, B6901, B6900, B6899, B6898, B6869, B6868, B6867, B6866, B6865,
    B6836, B6835, B6834, B6833, B6832, B6803, B6802, B6801, B6800, B6799,
    B6770, B6769, B6768, B6767, B6766, B6737, B6736, B6735, B6734, B6733,
    B6704, B6703, B6702, B6701, B6700, B6671, B6670, B6669, B6668, B6667,
    B6638, B6637, B6636, B6635, B6634, B6605, B6604, B6603, B6602, B6601,
    B6572, B6571, B6570, B6569, B6568, B6539, B6538, B6537, B6536, B6535,
    B6506, B6505, B6504, B6503, B6502, B6473, B6472, B6471, B6470, B6469,
    B6440, B6439, B6438, B6437, B6436, B6407, B6406, B6405, B6404, B6403,
    B6374, B6373, B6372, B6371, B6370, B6341, B6340, B6339, B6338, B6337,
    B6308, B6307, B6306, B6305, B6304, B6275, B6274, B6273, B6272, B6271,
    B6242, B6241, B6240, B6239, B6238, B6209, B6208, B6207, B6206, B6205,
    B6176, B6175, B6174, B6173, B6172, B6143, B6142, B6141, B6140, B6139,
    B6110, B6109, B6108, B6107, B6106, B6077, B6076, B6075, B6074, B6073,
    B6044, B6043, B6042, B6041, B6040, B6011, B6010, B6009, B6008, B6007,
    B5978, B5977, B5976, B5975, B5974, B5945, B5944, B5943, B5942, B5941,
    B5912, B5911, B5910, B5909, B5908, B5879, B5878, B5877, B5876, B5875,
    B5846, B5845, B5844, B5843, B5842, B5813, B5812, B5811, B5810, B5809,
    B5780, B5779, B5778, B5777, B5776, B5747, B5746, B5745, B5744, B5743,
    B5714, B5713, B5712, B5711, B5710, B5681, B5680, B5679, B5678, B5677,
    B5648, B5647, B5646, B5645, B5644, B5615, B5614, B5613, B5612, B5611,
    B5582, B5581, B5580, B5579, B5578, B5549, B5548, B5547, B5546, B5545,
    B5516, B5515, B5514, B5513, B5512, B5483, B5482, B5481, B5480, B5479,
    B5450, B5449, B5448, B5447, B5446, B5417, B5416, B5415, B5414, B5413,
    B5384, B5383, B5382, B5381, B5380, B5351, B5350, B5349, B5348, B5347,
    B5318, B5317, B5316, B5315, B5314, B5285, B5284, B5283, B5282, B5281,
    B5252, B5251, B5250, B5249, B5248, B5219, B5218, B5217, B5216, B5215,
    B5182, B5183, B5184, B5185, B5186,
    A6907, A6906, A6905, A6904, A6903, A6874, A6873, A6872, A6871, A6870,
    A6841, A6840, A6839, A6838, A6837, A6808, A6807, A6806, A6805, A6804,
    A6775, A6774, A6773, A6772, A6771, A6742, A6741, A6740, A6739, A6738,
    A6709, A6708, A6707, A6706, A6705, A6676, A6675, A6674, A6673, A6672,
    A6643, A6642, A6641, A6640, A6639, A6610, A6609, A6608, A6607, A6606,
    A6577, A6576, A6575, A6574, A6573, A6544, A6543, A6542, A6541, A6540,
    A6511, A6510, A6509, A6508, A6507, A6478, A6477, A6476, A6475, A6474,
    A6445, A6444, A6443, A6442, A6441, A6412, A6411, A6410, A6409, A6408,
    A6379, A6378, A6377, A6376, A6375, A6346, A6345, A6344, A6343, A6342,
    A6313, A6312, A6311, A6310, A6309, A6280, A6279, A6278, A6277, A6276,
    A6247, A6246, A6245, A6244, A6243, A6214, A6213, A6212, A6211, A6210,
    A6181, A6180, A6179, A6178, A6177, A6148, A6147, A6146, A6145, A6144,
    A6115, A6114, A6113, A6112, A6111, A6082, A6081, A6080, A6079, A6078,
    A6049, A6048, A6047, A6046, A6045, A6016, A6015, A6014, A6013, A6012,
    A5983, A5982, A5981, A5980, A5979, A5950, A5949, A5948, A5947, A5946,
    A5917, A5916, A5915, A5914, A5913, A5884, A5883, A5882, A5881, A5880,
    A5851, A5850, A5849, A5848, A5847, A5818, A5817, A5816, A5815, A5814,
    A5785, A5784, A5783, A5782, A5781, A5752, A5751, A5750, A5749, A5748,
    A5719, A5718, A5717, A5716, A5715, A5686, A5685, A5684, A5683, A5682,
    A5653, A5652, A5651, A5650, A5649, A5620, A5619, A5618, A5617, A5616,
    A5587, A5586, A5585, A5584, A5583, A5554, A5553, A5552, A5551, A5550,
    A5521, A5520, A5519, A5518, A5517, A5488, A5487, A5486, A5485, A5484,
    A5455, A5454, A5453, A5452, A5451, A5422, A5421, A5420, A5419, A5418,
    A5389, A5388, A5387, A5386, A5385, A5356, A5355, A5354, A5353, A5352,
    A5323, A5322, A5321, A5320, A5319, A5290, A5289, A5288, A5287, A5286,
    A5257, A5256, A5255, A5254, A5253, A5224, A5223, A5222, A5221, A5220,
    A5191, A5190, A5189, A5188, A5187, A5158, A5157, A5156, A5155, A5154,
    A5125, A5124, A5123, A5122, A5121, A5092, A5091, A5090, A5089, A5088,
    A5059, A5058, A5057, A5056, A5055, A5026, A5025, A5024, A5023, A5022,
    A4993, A4992, A4991, A4990, A4989, A4960, A4959, A4958, A4957, A4956,
    A4927, A4926, A4925, A4924, A4923, A4894, A4893, A4892, A4891, A4890,
    A4861, A4860, A4859, A4858, A4857, A4828, A4827, A4826, A4825, A4824,
    A4795, A4794, A4793, A4792, A4791, A4762, A4761, A4760, A4759, A4758,
    A4729, A4728, A4727, A4726, A4725, A4696, A4695, A4694, A4693, A4692,
    A4663, A4662, A4661, A4660, A4659, A4630, A4629, A4628, A4627, A4626,
    A4597, A4596, A4595, A4594, A4593, A4564, A4563, A4562, A4561, A4560,
    A4531, A4530, A4529, A4528, A4527, A4498, A4497, A4496, A4495, A4494,
    A4465, A4464, A4463, A4462, A4461, A4432, A4431, A4430, A4429, A4428,
    A4399, A4398, A4397, A4396, A4395, A4366, A4365, A4364, A4363, A4362,
    A4333, A4332, A4331, A4330, A4329, A4300, A4299, A4298, A4297, A4296,
    A4267, A4266, A4265, A4264, A4263, A4234, A4233, A4232, A4231, A4230,
    A4201, A4200, A4199, A4198, A4197, A4168, A4167, A4166, A4165, A4164,
    A4135, A4134, A4133, A4132, A4131, A4102, A4101, A4100, A4099, A4098,
    A4069, A4068, A4067, A4066, A4065, A4036, A4035, A4034, A4033, A4032,
    A4003, A4002, A4001, A4000, A3999, A3970, A3969, A3968, A3967, A3966,
    A3937, A3936, A3935, A3934, A3933, A3904, A3903, A3902, A3901, A3900,
    A3871, A3870, A3869, A3868, A3867, A3838, A3837, A3836, A3835, A3834,
    A3805, A3804, A3803, A3802, A3801, A3772, A3771, A3770, A3769, A3768,
    A3739, A3738, A3737, A3736, A3735, A3706, A3705, A3704, A3703, A3702,
    A3673, A3672, A3671, A3670, A3669, A3640, A3639, A3638, A3637, A3636,
    A3607, A3606, A3605, A3604, A3603, A3574, A3573, A3572, A3571, A3570,
    A3541, A3540, A3539, A3538, A3537, A3508, A3507, A3506, A3505, A3504,
    A3475, A3474, A3473, A3472, A3471, A3442, A3441, A3440, A3439, A3438,
    A3409, A3408, A3407, A3406, A3405, A3376, A3375, A3374, A3373, A3372,
    A3343, A3342, A3341, A3340, A3339, A3310, A3309, A3308, A3307, A3306,
    A3277, A3276, A3275, A3274, A3273, A3244, A3243, A3242, A3241, A3240,
    A3211, A3210, A3209, A3208, A3207, A3178, A3177, A3176, A3175, A3174,
    A3145, A3144, A3143, A3142, A3141, A3112, A3111, A3110, A3109, A3108,
    A3079, A3078, A3077, A3076, A3075, A3046, A3045, A3044, A3043, A3042,
    A3013, A3012, A3011, A3010, A3009, A2980, A2979, A2978, A2977, A2976,
    A2947, A2946, A2945, A2944, A2943, A2914, A2913, A2912, A2911, A2910,
    A2881, A2880, A2879, A2878, A2877, A2848, A2847, A2846, A2845, A2844,
    A2811, A2812, A2813, A2814, A2815  );
  input  B9278, B9277, B9276, B9275, B9274, B9245, B9244, B9243, B9242,
    B9241, B9212, B9211, B9210, B9209, B9208, B9179, B9178, B9177, B9176,
    B9175, B9146, B9145, B9144, B9143, B9142, B9113, B9112, B9111, B9110,
    B9109, B9080, B9079, B9078, B9077, B9076, B9047, B9046, B9045, B9044,
    B9043, B9014, B9013, B9012, B9011, B9010, B8981, B8980, B8979, B8978,
    B8977, B8948, B8947, B8946, B8945, B8944, B8915, B8914, B8913, B8912,
    B8911, B8882, B8881, B8880, B8879, B8878, B8849, B8848, B8847, B8846,
    B8845, B8816, B8815, B8814, B8813, B8812, B8783, B8782, B8781, B8780,
    B8779, B8750, B8749, B8748, B8747, B8746, B8717, B8716, B8715, B8714,
    B8713, B8684, B8683, B8682, B8681, B8680, B8651, B8650, B8649, B8648,
    B8647, B8618, B8617, B8616, B8615, B8614, B8585, B8584, B8583, B8582,
    B8581, B8552, B8551, B8550, B8549, B8548, B8519, B8518, B8517, B8516,
    B8515, B8486, B8485, B8484, B8483, B8482, B8453, B8452, B8451, B8450,
    B8449, B8420, B8419, B8418, B8417, B8416, B8387, B8386, B8385, B8384,
    B8383, B8354, B8353, B8352, B8351, B8350, B8321, B8320, B8319, B8318,
    B8317, B8288, B8287, B8286, B8285, B8284, B8255, B8254, B8253, B8252,
    B8251, B8222, B8221, B8220, B8219, B8218, B8189, B8188, B8187, B8186,
    B8185, B8156, B8155, B8154, B8153, B8152, B8123, B8122, B8121, B8120,
    B8119, B8090, B8089, B8088, B8087, B8086, B8057, B8056, B8055, B8054,
    B8053, B8024, B8023, B8022, B8021, B8020, B7991, B7990, B7989, B7988,
    B7987, B7958, B7957, B7956, B7955, B7954, B7925, B7924, B7923, B7922,
    B7921, B7892, B7891, B7890, B7889, B7888, B7859, B7858, B7857, B7856,
    B7855, B7826, B7825, B7824, B7823, B7822, B7793, B7792, B7791, B7790,
    B7789, B7760, B7759, B7758, B7757, B7756, B7727, B7726, B7725, B7724,
    B7723, B7694, B7693, B7692, B7691, B7690, B7661, B7660, B7659, B7658,
    B7657, B7628, B7627, B7626, B7625, B7624, B7595, B7594, B7593, B7592,
    B7591, B7562, B7561, B7560, B7559, B7558, B7529, B7528, B7527, B7526,
    B7525, B7496, B7495, B7494, B7493, B7492, B7463, B7462, B7461, B7460,
    B7459, B7430, B7429, B7428, B7427, B7426, B7397, B7396, B7395, B7394,
    B7393, B7364, B7363, B7362, B7361, B7360, B7331, B7330, B7329, B7328,
    B7327, B7298, B7297, B7296, B7295, B7294, B7265, B7264, B7263, B7262,
    B7261, B7232, B7231, B7230, B7229, B7228, B7199, B7198, B7197, B7196,
    B7195, B7166, B7165, B7164, B7163, B7162, B7133, B7132, B7131, B7130,
    B7129, B7100, B7099, B7098, B7097, B7096, B7067, B7066, B7065, B7064,
    B7063, B7034, B7033, B7032, B7031, B7030, B7001, B7000, B6999, B6998,
    B6997, B6968, B6967, B6966, B6965, B6964, B6935, B6934, B6933, B6932,
    B6931, B6902, B6901, B6900, B6899, B6898, B6869, B6868, B6867, B6866,
    B6865, B6836, B6835, B6834, B6833, B6832, B6803, B6802, B6801, B6800,
    B6799, B6770, B6769, B6768, B6767, B6766, B6737, B6736, B6735, B6734,
    B6733, B6704, B6703, B6702, B6701, B6700, B6671, B6670, B6669, B6668,
    B6667, B6638, B6637, B6636, B6635, B6634, B6605, B6604, B6603, B6602,
    B6601, B6572, B6571, B6570, B6569, B6568, B6539, B6538, B6537, B6536,
    B6535, B6506, B6505, B6504, B6503, B6502, B6473, B6472, B6471, B6470,
    B6469, B6440, B6439, B6438, B6437, B6436, B6407, B6406, B6405, B6404,
    B6403, B6374, B6373, B6372, B6371, B6370, B6341, B6340, B6339, B6338,
    B6337, B6308, B6307, B6306, B6305, B6304, B6275, B6274, B6273, B6272,
    B6271, B6242, B6241, B6240, B6239, B6238, B6209, B6208, B6207, B6206,
    B6205, B6176, B6175, B6174, B6173, B6172, B6143, B6142, B6141, B6140,
    B6139, B6110, B6109, B6108, B6107, B6106, B6077, B6076, B6075, B6074,
    B6073, B6044, B6043, B6042, B6041, B6040, B6011, B6010, B6009, B6008,
    B6007, B5978, B5977, B5976, B5975, B5974, B5945, B5944, B5943, B5942,
    B5941, B5912, B5911, B5910, B5909, B5908, B5879, B5878, B5877, B5876,
    B5875, B5846, B5845, B5844, B5843, B5842, B5813, B5812, B5811, B5810,
    B5809, B5780, B5779, B5778, B5777, B5776, B5747, B5746, B5745, B5744,
    B5743, B5714, B5713, B5712, B5711, B5710, B5681, B5680, B5679, B5678,
    B5677, B5648, B5647, B5646, B5645, B5644, B5615, B5614, B5613, B5612,
    B5611, B5582, B5581, B5580, B5579, B5578, B5549, B5548, B5547, B5546,
    B5545, B5516, B5515, B5514, B5513, B5512, B5483, B5482, B5481, B5480,
    B5479, B5450, B5449, B5448, B5447, B5446, B5417, B5416, B5415, B5414,
    B5413, B5384, B5383, B5382, B5381, B5380, B5351, B5350, B5349, B5348,
    B5347, B5318, B5317, B5316, B5315, B5314, B5285, B5284, B5283, B5282,
    B5281, B5252, B5251, B5250, B5249, B5248, B5219, B5218, B5217, B5216,
    B5215, B5182, B5183, B5184, B5185, B5186;
  output A6907, A6906, A6905, A6904, A6903, A6874, A6873, A6872, A6871, A6870,
    A6841, A6840, A6839, A6838, A6837, A6808, A6807, A6806, A6805, A6804,
    A6775, A6774, A6773, A6772, A6771, A6742, A6741, A6740, A6739, A6738,
    A6709, A6708, A6707, A6706, A6705, A6676, A6675, A6674, A6673, A6672,
    A6643, A6642, A6641, A6640, A6639, A6610, A6609, A6608, A6607, A6606,
    A6577, A6576, A6575, A6574, A6573, A6544, A6543, A6542, A6541, A6540,
    A6511, A6510, A6509, A6508, A6507, A6478, A6477, A6476, A6475, A6474,
    A6445, A6444, A6443, A6442, A6441, A6412, A6411, A6410, A6409, A6408,
    A6379, A6378, A6377, A6376, A6375, A6346, A6345, A6344, A6343, A6342,
    A6313, A6312, A6311, A6310, A6309, A6280, A6279, A6278, A6277, A6276,
    A6247, A6246, A6245, A6244, A6243, A6214, A6213, A6212, A6211, A6210,
    A6181, A6180, A6179, A6178, A6177, A6148, A6147, A6146, A6145, A6144,
    A6115, A6114, A6113, A6112, A6111, A6082, A6081, A6080, A6079, A6078,
    A6049, A6048, A6047, A6046, A6045, A6016, A6015, A6014, A6013, A6012,
    A5983, A5982, A5981, A5980, A5979, A5950, A5949, A5948, A5947, A5946,
    A5917, A5916, A5915, A5914, A5913, A5884, A5883, A5882, A5881, A5880,
    A5851, A5850, A5849, A5848, A5847, A5818, A5817, A5816, A5815, A5814,
    A5785, A5784, A5783, A5782, A5781, A5752, A5751, A5750, A5749, A5748,
    A5719, A5718, A5717, A5716, A5715, A5686, A5685, A5684, A5683, A5682,
    A5653, A5652, A5651, A5650, A5649, A5620, A5619, A5618, A5617, A5616,
    A5587, A5586, A5585, A5584, A5583, A5554, A5553, A5552, A5551, A5550,
    A5521, A5520, A5519, A5518, A5517, A5488, A5487, A5486, A5485, A5484,
    A5455, A5454, A5453, A5452, A5451, A5422, A5421, A5420, A5419, A5418,
    A5389, A5388, A5387, A5386, A5385, A5356, A5355, A5354, A5353, A5352,
    A5323, A5322, A5321, A5320, A5319, A5290, A5289, A5288, A5287, A5286,
    A5257, A5256, A5255, A5254, A5253, A5224, A5223, A5222, A5221, A5220,
    A5191, A5190, A5189, A5188, A5187, A5158, A5157, A5156, A5155, A5154,
    A5125, A5124, A5123, A5122, A5121, A5092, A5091, A5090, A5089, A5088,
    A5059, A5058, A5057, A5056, A5055, A5026, A5025, A5024, A5023, A5022,
    A4993, A4992, A4991, A4990, A4989, A4960, A4959, A4958, A4957, A4956,
    A4927, A4926, A4925, A4924, A4923, A4894, A4893, A4892, A4891, A4890,
    A4861, A4860, A4859, A4858, A4857, A4828, A4827, A4826, A4825, A4824,
    A4795, A4794, A4793, A4792, A4791, A4762, A4761, A4760, A4759, A4758,
    A4729, A4728, A4727, A4726, A4725, A4696, A4695, A4694, A4693, A4692,
    A4663, A4662, A4661, A4660, A4659, A4630, A4629, A4628, A4627, A4626,
    A4597, A4596, A4595, A4594, A4593, A4564, A4563, A4562, A4561, A4560,
    A4531, A4530, A4529, A4528, A4527, A4498, A4497, A4496, A4495, A4494,
    A4465, A4464, A4463, A4462, A4461, A4432, A4431, A4430, A4429, A4428,
    A4399, A4398, A4397, A4396, A4395, A4366, A4365, A4364, A4363, A4362,
    A4333, A4332, A4331, A4330, A4329, A4300, A4299, A4298, A4297, A4296,
    A4267, A4266, A4265, A4264, A4263, A4234, A4233, A4232, A4231, A4230,
    A4201, A4200, A4199, A4198, A4197, A4168, A4167, A4166, A4165, A4164,
    A4135, A4134, A4133, A4132, A4131, A4102, A4101, A4100, A4099, A4098,
    A4069, A4068, A4067, A4066, A4065, A4036, A4035, A4034, A4033, A4032,
    A4003, A4002, A4001, A4000, A3999, A3970, A3969, A3968, A3967, A3966,
    A3937, A3936, A3935, A3934, A3933, A3904, A3903, A3902, A3901, A3900,
    A3871, A3870, A3869, A3868, A3867, A3838, A3837, A3836, A3835, A3834,
    A3805, A3804, A3803, A3802, A3801, A3772, A3771, A3770, A3769, A3768,
    A3739, A3738, A3737, A3736, A3735, A3706, A3705, A3704, A3703, A3702,
    A3673, A3672, A3671, A3670, A3669, A3640, A3639, A3638, A3637, A3636,
    A3607, A3606, A3605, A3604, A3603, A3574, A3573, A3572, A3571, A3570,
    A3541, A3540, A3539, A3538, A3537, A3508, A3507, A3506, A3505, A3504,
    A3475, A3474, A3473, A3472, A3471, A3442, A3441, A3440, A3439, A3438,
    A3409, A3408, A3407, A3406, A3405, A3376, A3375, A3374, A3373, A3372,
    A3343, A3342, A3341, A3340, A3339, A3310, A3309, A3308, A3307, A3306,
    A3277, A3276, A3275, A3274, A3273, A3244, A3243, A3242, A3241, A3240,
    A3211, A3210, A3209, A3208, A3207, A3178, A3177, A3176, A3175, A3174,
    A3145, A3144, A3143, A3142, A3141, A3112, A3111, A3110, A3109, A3108,
    A3079, A3078, A3077, A3076, A3075, A3046, A3045, A3044, A3043, A3042,
    A3013, A3012, A3011, A3010, A3009, A2980, A2979, A2978, A2977, A2976,
    A2947, A2946, A2945, A2944, A2943, A2914, A2913, A2912, A2911, A2910,
    A2881, A2880, A2879, A2878, A2877, A2848, A2847, A2846, A2845, A2844,
    A2811, A2812, A2813, A2814, A2815;
  wire new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2815_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2831_,
    new_n2832_, new_n2833_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_,
    new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_,
    new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3400_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3416_, new_n3417_, new_n3418_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4601_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4610_,
    new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4617_,
    new_n4618_, new_n4619_, new_n4621_, new_n4622_, new_n4623_, new_n4624_,
    new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_,
    new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_,
    new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_,
    new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_,
    new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_,
    new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_,
    new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_,
    new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_,
    new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_,
    new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_,
    new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_,
    new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_,
    new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_,
    new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_,
    new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_,
    new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_,
    new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_,
    new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_,
    new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_,
    new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_,
    new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_,
    new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_,
    new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_,
    new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_,
    new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_,
    new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_,
    new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_,
    new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_,
    new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_,
    new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_,
    new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_,
    new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_,
    new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_,
    new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_,
    new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_,
    new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_,
    new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_,
    new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_,
    new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_,
    new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_,
    new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_,
    new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_,
    new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_,
    new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_,
    new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_,
    new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_,
    new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_,
    new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_,
    new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_,
    new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_,
    new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_,
    new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_,
    new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_,
    new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_,
    new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_,
    new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_,
    new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_,
    new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_,
    new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_,
    new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_,
    new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_,
    new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_,
    new_n5802_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_,
    new_n5809_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5818_, new_n5819_, new_n5820_, new_n5822_, new_n5823_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_,
    new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_,
    new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_,
    new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_,
    new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_,
    new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_,
    new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_,
    new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_,
    new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_,
    new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_,
    new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_,
    new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_,
    new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_,
    new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_,
    new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_,
    new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_,
    new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_,
    new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_,
    new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_,
    new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_,
    new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_,
    new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_,
    new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_,
    new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_,
    new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_,
    new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_,
    new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_,
    new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_,
    new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_,
    new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_,
    new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_,
    new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_,
    new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_,
    new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_,
    new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_,
    new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_,
    new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_,
    new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_,
    new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_,
    new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_,
    new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_,
    new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_,
    new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_,
    new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_,
    new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_,
    new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_,
    new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_,
    new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_,
    new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_,
    new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_,
    new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_,
    new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_,
    new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_,
    new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_,
    new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_,
    new_n6635_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_,
    new_n6649_, new_n6651_, new_n6652_, new_n6653_, new_n6655_, new_n6656_,
    new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_,
    new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_,
    new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_,
    new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_,
    new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_,
    new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_,
    new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_,
    new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_,
    new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_,
    new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_,
    new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_,
    new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_,
    new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_,
    new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_,
    new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6765_,
    new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6781_, new_n6782_, new_n6783_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6895_, new_n6897_,
    new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6904_,
    new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6911_,
    new_n6912_, new_n6913_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7025_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7034_, new_n7035_,
    new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7041_, new_n7042_,
    new_n7043_, new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_,
    new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_,
    new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_,
    new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_,
    new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_,
    new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_,
    new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_,
    new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_,
    new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_,
    new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_,
    new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_,
    new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7155_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7171_, new_n7172_, new_n7173_,
    new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_,
    new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_,
    new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_,
    new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_,
    new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_,
    new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_,
    new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_,
    new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_,
    new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_,
    new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_,
    new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_,
    new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_,
    new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_,
    new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_,
    new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_,
    new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_,
    new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_,
    new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_,
    new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_,
    new_n7290_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7306_, new_n7307_, new_n7308_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7545_, new_n7547_,
    new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7554_,
    new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7561_,
    new_n7562_, new_n7563_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7800_, new_n7802_, new_n7803_, new_n7804_,
    new_n7805_, new_n7806_, new_n7807_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7816_, new_n7817_, new_n7818_,
    new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_,
    new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_,
    new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_,
    new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_,
    new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_,
    new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_,
    new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_,
    new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_,
    new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_,
    new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_,
    new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_,
    new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_,
    new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_,
    new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_,
    new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_,
    new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_,
    new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_,
    new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_,
    new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_,
    new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_,
    new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_,
    new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_,
    new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_,
    new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_,
    new_n8055_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8071_, new_n8072_, new_n8073_, new_n8075_, new_n8076_,
    new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_,
    new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_,
    new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_,
    new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_,
    new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_,
    new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_,
    new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_,
    new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_,
    new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_,
    new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_,
    new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_,
    new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_,
    new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_,
    new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_,
    new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_,
    new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_,
    new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_,
    new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_,
    new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_,
    new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_,
    new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_,
    new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_,
    new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_,
    new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_,
    new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_,
    new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_,
    new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_,
    new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_,
    new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_,
    new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_,
    new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_,
    new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_,
    new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8310_, new_n8312_,
    new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8319_,
    new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8326_,
    new_n8327_, new_n8328_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8561_, new_n8563_,
    new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8570_,
    new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8577_,
    new_n8578_, new_n8579_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_,
    new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_,
    new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_,
    new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_,
    new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_,
    new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_,
    new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_,
    new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_,
    new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_,
    new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_,
    new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_,
    new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_,
    new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_,
    new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_,
    new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_,
    new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_,
    new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_,
    new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_,
    new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_,
    new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_,
    new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_,
    new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_,
    new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_,
    new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_,
    new_n8813_, new_n8814_, new_n8816_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8832_, new_n8833_, new_n8834_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_,
    new_n8878_, new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_,
    new_n8884_, new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_,
    new_n8890_, new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_,
    new_n8896_, new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_,
    new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_,
    new_n8908_, new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_,
    new_n8914_, new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_,
    new_n8920_, new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_,
    new_n8926_, new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_,
    new_n8932_, new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_,
    new_n8938_, new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_,
    new_n8944_, new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_,
    new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_,
    new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_,
    new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_,
    new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_,
    new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_,
    new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_,
    new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_,
    new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_,
    new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_,
    new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9071_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9087_, new_n9088_, new_n9089_, new_n9091_, new_n9092_,
    new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_,
    new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_,
    new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_,
    new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_,
    new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_,
    new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_,
    new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_,
    new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_,
    new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_,
    new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_,
    new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_,
    new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_,
    new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_,
    new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_,
    new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_,
    new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_,
    new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_,
    new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_,
    new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_,
    new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_,
    new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_,
    new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_,
    new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_,
    new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9326_, new_n9328_,
    new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9335_,
    new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9342_,
    new_n9343_, new_n9344_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_,
    new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_,
    new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_,
    new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_,
    new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_,
    new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_,
    new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_,
    new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_,
    new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_,
    new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_,
    new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_,
    new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_,
    new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_,
    new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_,
    new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_,
    new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_,
    new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_,
    new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_,
    new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_,
    new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_,
    new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_,
    new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_,
    new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_,
    new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_,
    new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_,
    new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9581_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9590_, new_n9591_, new_n9592_,
    new_n9593_, new_n9594_, new_n9595_, new_n9597_, new_n9598_, new_n9599_,
    new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_,
    new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_,
    new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_,
    new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_,
    new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_,
    new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_,
    new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_,
    new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_,
    new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_,
    new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_,
    new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_,
    new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_,
    new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_,
    new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_,
    new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_,
    new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_,
    new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_,
    new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_,
    new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_,
    new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_,
    new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_,
    new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_,
    new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_,
    new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_,
    new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_,
    new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_,
    new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_,
    new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_,
    new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_,
    new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_,
    new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_,
    new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_,
    new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_,
    new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_,
    new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_,
    new_n9829_, new_n9830_, new_n9832_, new_n9834_, new_n9835_, new_n9836_,
    new_n9837_, new_n9838_, new_n9839_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9848_, new_n9849_, new_n9850_,
    new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_,
    new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_,
    new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_,
    new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_,
    new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_,
    new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_,
    new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_,
    new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_,
    new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_,
    new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10012_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10021_, new_n10022_, new_n10023_,
    new_n10024_, new_n10025_, new_n10026_, new_n10028_, new_n10029_,
    new_n10030_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10192_, new_n10194_, new_n10195_, new_n10196_, new_n10197_,
    new_n10198_, new_n10199_, new_n10201_, new_n10202_, new_n10203_,
    new_n10204_, new_n10205_, new_n10206_, new_n10208_, new_n10209_,
    new_n10210_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10372_, new_n10374_, new_n10375_, new_n10376_, new_n10377_,
    new_n10378_, new_n10379_, new_n10381_, new_n10382_, new_n10383_,
    new_n10384_, new_n10385_, new_n10386_, new_n10388_, new_n10389_,
    new_n10390_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10552_, new_n10554_, new_n10555_, new_n10556_, new_n10557_,
    new_n10558_, new_n10559_, new_n10561_, new_n10562_, new_n10563_,
    new_n10564_, new_n10565_, new_n10566_, new_n10568_, new_n10569_,
    new_n10570_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10735_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10744_, new_n10745_, new_n10746_, new_n10747_, new_n10748_,
    new_n10749_, new_n10751_, new_n10752_, new_n10753_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10775_, new_n10777_,
    new_n10778_, new_n10779_, new_n10780_, new_n10781_, new_n10782_,
    new_n10784_, new_n10785_, new_n10786_, new_n10787_, new_n10788_,
    new_n10789_, new_n10791_, new_n10792_, new_n10793_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10815_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10824_, new_n10825_, new_n10826_, new_n10827_, new_n10828_,
    new_n10829_, new_n10831_, new_n10832_, new_n10833_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10855_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10864_, new_n10865_, new_n10866_, new_n10867_, new_n10868_,
    new_n10869_, new_n10871_, new_n10872_, new_n10873_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10895_, new_n10897_,
    new_n10898_, new_n10899_, new_n10900_, new_n10901_, new_n10902_,
    new_n10904_, new_n10905_, new_n10906_, new_n10907_, new_n10908_,
    new_n10909_, new_n10911_, new_n10912_, new_n10913_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10935_, new_n10937_,
    new_n10938_, new_n10939_, new_n10940_, new_n10941_, new_n10942_,
    new_n10944_, new_n10945_, new_n10946_, new_n10947_, new_n10948_,
    new_n10949_, new_n10951_, new_n10952_, new_n10953_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10975_, new_n10977_,
    new_n10978_, new_n10979_, new_n10980_, new_n10981_, new_n10982_,
    new_n10984_, new_n10985_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10991_, new_n10992_, new_n10993_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11015_, new_n11017_,
    new_n11018_, new_n11019_, new_n11020_, new_n11021_, new_n11022_,
    new_n11024_, new_n11025_, new_n11026_, new_n11027_, new_n11028_,
    new_n11029_, new_n11031_, new_n11032_, new_n11033_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11055_, new_n11057_,
    new_n11058_, new_n11059_, new_n11060_, new_n11061_, new_n11062_,
    new_n11064_, new_n11065_, new_n11066_, new_n11067_, new_n11068_,
    new_n11069_, new_n11071_, new_n11072_, new_n11073_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11095_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11101_, new_n11102_,
    new_n11104_, new_n11105_, new_n11106_, new_n11107_, new_n11108_,
    new_n11109_, new_n11111_, new_n11112_, new_n11113_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11135_, new_n11137_,
    new_n11138_, new_n11139_, new_n11140_, new_n11141_, new_n11142_,
    new_n11144_, new_n11145_, new_n11146_, new_n11147_, new_n11148_,
    new_n11149_, new_n11151_, new_n11152_, new_n11153_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11175_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11184_, new_n11185_, new_n11186_, new_n11187_, new_n11188_,
    new_n11189_, new_n11191_, new_n11192_, new_n11193_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11215_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11224_, new_n11225_, new_n11226_, new_n11227_, new_n11228_,
    new_n11229_, new_n11231_, new_n11232_, new_n11233_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11255_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11262_,
    new_n11264_, new_n11265_, new_n11266_, new_n11267_, new_n11268_,
    new_n11269_, new_n11271_, new_n11272_, new_n11273_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11295_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11304_, new_n11305_, new_n11306_, new_n11307_, new_n11308_,
    new_n11309_, new_n11311_, new_n11312_, new_n11313_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11335_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11344_, new_n11345_, new_n11346_, new_n11347_, new_n11348_,
    new_n11349_, new_n11351_, new_n11352_, new_n11353_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11375_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11384_, new_n11385_, new_n11386_, new_n11387_, new_n11388_,
    new_n11389_, new_n11391_, new_n11392_, new_n11393_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11415_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11424_, new_n11425_, new_n11426_, new_n11427_, new_n11428_,
    new_n11429_, new_n11431_, new_n11432_, new_n11433_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11455_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11464_, new_n11465_, new_n11466_, new_n11467_, new_n11468_,
    new_n11469_, new_n11471_, new_n11472_, new_n11473_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11495_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11504_, new_n11505_, new_n11506_, new_n11507_, new_n11508_,
    new_n11509_, new_n11511_, new_n11512_, new_n11513_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11535_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11544_, new_n11545_, new_n11546_, new_n11547_, new_n11548_,
    new_n11549_, new_n11551_, new_n11552_, new_n11553_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11575_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11584_, new_n11585_, new_n11586_, new_n11587_, new_n11588_,
    new_n11589_, new_n11591_, new_n11592_, new_n11593_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11615_, new_n11617_,
    new_n11618_, new_n11619_, new_n11620_, new_n11621_, new_n11622_,
    new_n11624_, new_n11625_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11631_, new_n11632_, new_n11633_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11655_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11664_, new_n11665_, new_n11666_, new_n11667_, new_n11668_,
    new_n11669_, new_n11671_, new_n11672_, new_n11673_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11695_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11704_, new_n11705_, new_n11706_, new_n11707_, new_n11708_,
    new_n11709_, new_n11711_, new_n11712_, new_n11713_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11740_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11749_, new_n11750_, new_n11751_, new_n11752_, new_n11753_,
    new_n11754_, new_n11756_, new_n11757_, new_n11758_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11805_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11814_, new_n11815_, new_n11816_, new_n11817_, new_n11818_,
    new_n11819_, new_n11821_, new_n11822_, new_n11823_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11870_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11884_, new_n11886_, new_n11887_, new_n11888_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11935_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11951_, new_n11952_, new_n11953_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n12000_, new_n12002_,
    new_n12003_, new_n12004_, new_n12005_, new_n12006_, new_n12007_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12016_, new_n12017_, new_n12018_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12065_, new_n12067_,
    new_n12068_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12081_, new_n12082_, new_n12083_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12130_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12139_, new_n12140_, new_n12141_, new_n12142_, new_n12143_,
    new_n12144_, new_n12146_, new_n12147_, new_n12148_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12195_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12211_, new_n12212_, new_n12213_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12260_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12276_, new_n12277_, new_n12278_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12325_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12334_, new_n12335_, new_n12336_, new_n12337_, new_n12338_,
    new_n12339_, new_n12341_, new_n12342_, new_n12343_, new_n12345_,
    new_n12346_, new_n12347_, new_n12348_, new_n12349_, new_n12350_,
    new_n12351_, new_n12352_, new_n12353_, new_n12354_, new_n12355_,
    new_n12356_, new_n12357_, new_n12358_, new_n12359_, new_n12360_,
    new_n12361_, new_n12362_, new_n12363_, new_n12364_, new_n12365_,
    new_n12366_, new_n12367_, new_n12368_, new_n12369_, new_n12370_,
    new_n12371_, new_n12372_, new_n12373_, new_n12374_, new_n12375_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12384_, new_n12385_,
    new_n12386_, new_n12387_, new_n12388_, new_n12390_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12406_, new_n12407_, new_n12408_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12420_,
    new_n12421_, new_n12422_, new_n12423_, new_n12424_, new_n12425_,
    new_n12426_, new_n12427_, new_n12428_, new_n12429_, new_n12430_,
    new_n12431_, new_n12432_, new_n12433_, new_n12434_, new_n12435_,
    new_n12436_, new_n12437_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12455_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12471_, new_n12472_, new_n12473_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12520_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12529_, new_n12530_, new_n12531_, new_n12532_, new_n12533_,
    new_n12534_, new_n12536_, new_n12537_, new_n12538_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12585_, new_n12587_,
    new_n12588_, new_n12589_, new_n12590_, new_n12591_, new_n12592_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12601_, new_n12602_, new_n12603_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12650_, new_n12652_,
    new_n12653_, new_n12654_, new_n12655_, new_n12656_, new_n12657_,
    new_n12659_, new_n12660_, new_n12661_, new_n12662_, new_n12663_,
    new_n12664_, new_n12666_, new_n12667_, new_n12668_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12715_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12724_, new_n12725_, new_n12726_, new_n12727_, new_n12728_,
    new_n12729_, new_n12731_, new_n12732_, new_n12733_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12780_, new_n12782_,
    new_n12783_, new_n12784_, new_n12785_, new_n12786_, new_n12787_,
    new_n12789_, new_n12790_, new_n12791_, new_n12792_, new_n12793_,
    new_n12794_, new_n12796_, new_n12797_, new_n12798_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12845_, new_n12847_,
    new_n12848_, new_n12849_, new_n12850_, new_n12851_, new_n12852_,
    new_n12854_, new_n12855_, new_n12856_, new_n12857_, new_n12858_,
    new_n12859_, new_n12861_, new_n12862_, new_n12863_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12910_, new_n12912_,
    new_n12913_, new_n12914_, new_n12915_, new_n12916_, new_n12917_,
    new_n12919_, new_n12920_, new_n12921_, new_n12922_, new_n12923_,
    new_n12924_, new_n12926_, new_n12927_, new_n12928_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12975_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12984_, new_n12985_, new_n12986_, new_n12987_, new_n12988_,
    new_n12989_, new_n12991_, new_n12992_, new_n12993_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13040_, new_n13042_,
    new_n13043_, new_n13044_, new_n13045_, new_n13046_, new_n13047_,
    new_n13049_, new_n13050_, new_n13051_, new_n13052_, new_n13053_,
    new_n13054_, new_n13056_, new_n13057_, new_n13058_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13105_, new_n13107_,
    new_n13108_, new_n13109_, new_n13110_, new_n13111_, new_n13112_,
    new_n13114_, new_n13115_, new_n13116_, new_n13117_, new_n13118_,
    new_n13119_, new_n13121_, new_n13122_, new_n13123_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13170_, new_n13172_,
    new_n13173_, new_n13174_, new_n13175_, new_n13176_, new_n13177_,
    new_n13179_, new_n13180_, new_n13181_, new_n13182_, new_n13183_,
    new_n13184_, new_n13186_, new_n13187_, new_n13188_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13235_, new_n13237_,
    new_n13238_, new_n13239_, new_n13240_, new_n13241_, new_n13242_,
    new_n13244_, new_n13245_, new_n13246_, new_n13247_, new_n13248_,
    new_n13249_, new_n13251_, new_n13252_, new_n13253_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13300_, new_n13302_,
    new_n13303_, new_n13304_, new_n13305_, new_n13306_, new_n13307_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13316_, new_n13317_, new_n13318_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13361_,
    new_n13363_, new_n13364_, new_n13365_, new_n13366_, new_n13367_,
    new_n13368_, new_n13370_, new_n13371_, new_n13372_, new_n13373_,
    new_n13374_, new_n13375_, new_n13377_, new_n13378_, new_n13379_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13426_,
    new_n13428_, new_n13429_, new_n13430_, new_n13431_, new_n13432_,
    new_n13433_, new_n13435_, new_n13436_, new_n13437_, new_n13438_,
    new_n13439_, new_n13440_, new_n13442_, new_n13443_, new_n13444_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13491_,
    new_n13493_, new_n13494_, new_n13495_, new_n13496_, new_n13497_,
    new_n13498_, new_n13500_, new_n13501_, new_n13502_, new_n13503_,
    new_n13504_, new_n13505_, new_n13507_, new_n13508_, new_n13509_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13556_,
    new_n13558_, new_n13559_, new_n13560_, new_n13561_, new_n13562_,
    new_n13563_, new_n13565_, new_n13566_, new_n13567_, new_n13568_,
    new_n13569_, new_n13570_, new_n13572_, new_n13573_, new_n13574_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13621_,
    new_n13623_, new_n13624_, new_n13625_, new_n13626_, new_n13627_,
    new_n13628_, new_n13630_, new_n13631_, new_n13632_, new_n13633_,
    new_n13634_, new_n13635_, new_n13637_, new_n13638_, new_n13639_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13686_,
    new_n13688_, new_n13689_, new_n13690_, new_n13691_, new_n13692_,
    new_n13693_, new_n13695_, new_n13696_, new_n13697_, new_n13698_,
    new_n13699_, new_n13700_, new_n13702_, new_n13703_, new_n13704_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13751_,
    new_n13753_, new_n13754_, new_n13755_, new_n13756_, new_n13757_,
    new_n13758_, new_n13760_, new_n13761_, new_n13762_, new_n13763_,
    new_n13764_, new_n13765_, new_n13767_, new_n13768_, new_n13769_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13816_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13822_,
    new_n13823_, new_n13825_, new_n13826_, new_n13827_, new_n13828_,
    new_n13829_, new_n13830_, new_n13832_, new_n13833_, new_n13834_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13881_,
    new_n13883_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13890_, new_n13891_, new_n13892_, new_n13893_,
    new_n13894_, new_n13895_, new_n13897_, new_n13898_, new_n13899_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13946_,
    new_n13948_, new_n13949_, new_n13950_, new_n13951_, new_n13952_,
    new_n13953_, new_n13955_, new_n13956_, new_n13957_, new_n13958_,
    new_n13959_, new_n13960_, new_n13962_, new_n13963_, new_n13964_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14011_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14020_, new_n14021_, new_n14022_, new_n14023_,
    new_n14024_, new_n14025_, new_n14027_, new_n14028_, new_n14029_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14076_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14085_, new_n14086_, new_n14087_, new_n14088_,
    new_n14089_, new_n14090_, new_n14092_, new_n14093_, new_n14094_,
    new_n14096_, new_n14097_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14103_, new_n14104_, new_n14105_,
    new_n14106_, new_n14107_, new_n14108_, new_n14109_, new_n14110_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14117_, new_n14118_, new_n14119_, new_n14120_,
    new_n14121_, new_n14122_, new_n14123_, new_n14124_, new_n14125_,
    new_n14126_, new_n14127_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14133_, new_n14134_, new_n14135_,
    new_n14136_, new_n14137_, new_n14138_, new_n14139_, new_n14141_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14150_, new_n14151_, new_n14152_, new_n14153_,
    new_n14154_, new_n14155_, new_n14157_, new_n14158_, new_n14159_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14206_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14215_, new_n14216_, new_n14217_, new_n14218_,
    new_n14219_, new_n14220_, new_n14222_, new_n14223_, new_n14224_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14241_, new_n14242_, new_n14243_, new_n14244_, new_n14245_,
    new_n14246_, new_n14247_, new_n14248_, new_n14249_, new_n14250_,
    new_n14251_, new_n14252_, new_n14253_, new_n14254_, new_n14255_,
    new_n14256_, new_n14257_, new_n14258_, new_n14259_, new_n14260_,
    new_n14261_, new_n14262_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14268_, new_n14269_, new_n14271_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14280_, new_n14281_, new_n14282_, new_n14283_,
    new_n14284_, new_n14285_, new_n14287_, new_n14288_, new_n14289_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14336_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14345_, new_n14346_, new_n14347_, new_n14348_,
    new_n14349_, new_n14350_, new_n14352_, new_n14353_, new_n14354_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14401_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14410_, new_n14411_, new_n14412_, new_n14413_,
    new_n14414_, new_n14415_, new_n14417_, new_n14418_, new_n14419_,
    new_n14421_, new_n14422_, new_n14423_, new_n14424_, new_n14425_,
    new_n14426_, new_n14427_, new_n14428_, new_n14429_, new_n14430_,
    new_n14431_, new_n14432_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14466_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14475_, new_n14476_, new_n14477_, new_n14478_,
    new_n14479_, new_n14480_, new_n14482_, new_n14483_, new_n14484_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14531_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14540_, new_n14541_, new_n14542_, new_n14543_,
    new_n14544_, new_n14545_, new_n14547_, new_n14548_, new_n14549_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14596_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14605_, new_n14606_, new_n14607_, new_n14608_,
    new_n14609_, new_n14610_, new_n14612_, new_n14613_, new_n14614_,
    new_n14616_, new_n14617_, new_n14618_, new_n14619_, new_n14620_,
    new_n14621_, new_n14622_, new_n14623_, new_n14624_, new_n14625_,
    new_n14626_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14661_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14670_, new_n14671_, new_n14672_, new_n14673_,
    new_n14674_, new_n14675_, new_n14677_, new_n14678_, new_n14679_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14726_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14735_, new_n14736_, new_n14737_, new_n14738_,
    new_n14739_, new_n14740_, new_n14742_, new_n14743_, new_n14744_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14791_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14800_, new_n14801_, new_n14802_, new_n14803_,
    new_n14804_, new_n14805_, new_n14807_, new_n14808_, new_n14809_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14840_,
    new_n14841_, new_n14842_, new_n14843_, new_n14844_, new_n14845_,
    new_n14846_, new_n14847_, new_n14848_, new_n14849_, new_n14850_,
    new_n14851_, new_n14852_, new_n14853_, new_n14854_, new_n14856_,
    new_n14858_, new_n14859_, new_n14860_, new_n14861_, new_n14862_,
    new_n14863_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14869_, new_n14870_, new_n14872_, new_n14873_, new_n14874_,
    new_n14876_, new_n14877_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14887_, new_n14888_, new_n14889_, new_n14890_,
    new_n14891_, new_n14892_, new_n14893_, new_n14894_, new_n14895_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14902_, new_n14903_, new_n14904_, new_n14905_,
    new_n14906_, new_n14907_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14921_,
    new_n14923_, new_n14924_, new_n14925_, new_n14926_, new_n14927_,
    new_n14928_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14937_, new_n14938_, new_n14939_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14982_, new_n14984_, new_n14985_, new_n14986_, new_n14987_,
    new_n14988_, new_n14989_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14998_, new_n14999_,
    new_n15000_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15032_, new_n15034_, new_n15035_, new_n15036_, new_n15037_,
    new_n15038_, new_n15039_, new_n15041_, new_n15042_, new_n15043_,
    new_n15044_, new_n15045_, new_n15046_, new_n15048_, new_n15049_,
    new_n15050_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15082_, new_n15084_, new_n15085_, new_n15086_, new_n15087_,
    new_n15088_, new_n15089_, new_n15091_, new_n15092_, new_n15093_,
    new_n15094_, new_n15095_, new_n15096_, new_n15098_, new_n15099_,
    new_n15100_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15132_, new_n15134_, new_n15135_, new_n15136_, new_n15137_,
    new_n15138_, new_n15139_, new_n15141_, new_n15142_, new_n15143_,
    new_n15144_, new_n15145_, new_n15146_, new_n15148_, new_n15149_,
    new_n15150_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15182_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15188_, new_n15189_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15198_, new_n15199_,
    new_n15200_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15232_, new_n15234_, new_n15235_, new_n15236_, new_n15237_,
    new_n15238_, new_n15239_, new_n15241_, new_n15242_, new_n15243_,
    new_n15244_, new_n15245_, new_n15246_, new_n15248_, new_n15249_,
    new_n15250_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15282_, new_n15284_, new_n15285_, new_n15286_, new_n15287_,
    new_n15288_, new_n15289_, new_n15291_, new_n15292_, new_n15293_,
    new_n15294_, new_n15295_, new_n15296_, new_n15298_, new_n15299_,
    new_n15300_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15328_, new_n15329_, new_n15330_,
    new_n15332_, new_n15334_, new_n15335_, new_n15336_, new_n15337_,
    new_n15338_, new_n15339_, new_n15341_, new_n15342_, new_n15343_,
    new_n15344_, new_n15345_, new_n15346_, new_n15348_, new_n15349_,
    new_n15350_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15382_, new_n15384_, new_n15385_, new_n15386_, new_n15387_,
    new_n15388_, new_n15389_, new_n15391_, new_n15392_, new_n15393_,
    new_n15394_, new_n15395_, new_n15396_, new_n15398_, new_n15399_,
    new_n15400_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15432_, new_n15434_, new_n15435_, new_n15436_, new_n15437_,
    new_n15438_, new_n15439_, new_n15441_, new_n15442_, new_n15443_,
    new_n15444_, new_n15445_, new_n15446_, new_n15448_, new_n15449_,
    new_n15450_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15482_, new_n15484_, new_n15485_, new_n15486_, new_n15487_,
    new_n15488_, new_n15489_, new_n15491_, new_n15492_, new_n15493_,
    new_n15494_, new_n15495_, new_n15496_, new_n15498_, new_n15499_,
    new_n15500_, new_n15502_, new_n15503_, new_n15504_, new_n15505_,
    new_n15506_, new_n15507_, new_n15508_, new_n15509_, new_n15510_,
    new_n15511_, new_n15512_, new_n15513_, new_n15514_, new_n15515_,
    new_n15516_, new_n15517_, new_n15518_, new_n15519_, new_n15520_,
    new_n15521_, new_n15522_, new_n15523_, new_n15524_, new_n15525_,
    new_n15526_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15532_, new_n15534_, new_n15535_, new_n15536_, new_n15537_,
    new_n15538_, new_n15539_, new_n15541_, new_n15542_, new_n15543_,
    new_n15544_, new_n15545_, new_n15546_, new_n15548_, new_n15549_,
    new_n15550_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15582_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15591_, new_n15592_, new_n15593_,
    new_n15594_, new_n15595_, new_n15596_, new_n15598_, new_n15599_,
    new_n15600_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15632_, new_n15634_, new_n15635_, new_n15636_, new_n15637_,
    new_n15638_, new_n15639_, new_n15641_, new_n15642_, new_n15643_,
    new_n15644_, new_n15645_, new_n15646_, new_n15648_, new_n15649_,
    new_n15650_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15682_, new_n15684_, new_n15685_, new_n15686_, new_n15687_,
    new_n15688_, new_n15689_, new_n15691_, new_n15692_, new_n15693_,
    new_n15694_, new_n15695_, new_n15696_, new_n15698_, new_n15699_,
    new_n15700_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15732_, new_n15734_, new_n15735_, new_n15736_, new_n15737_,
    new_n15738_, new_n15739_, new_n15741_, new_n15742_, new_n15743_,
    new_n15744_, new_n15745_, new_n15746_, new_n15748_, new_n15749_,
    new_n15750_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15782_, new_n15784_, new_n15785_, new_n15786_, new_n15787_,
    new_n15788_, new_n15789_, new_n15791_, new_n15792_, new_n15793_,
    new_n15794_, new_n15795_, new_n15796_, new_n15798_, new_n15799_,
    new_n15800_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15832_, new_n15834_, new_n15835_, new_n15836_, new_n15837_,
    new_n15838_, new_n15839_, new_n15841_, new_n15842_, new_n15843_,
    new_n15844_, new_n15845_, new_n15846_, new_n15848_, new_n15849_,
    new_n15850_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15882_, new_n15884_, new_n15885_, new_n15886_, new_n15887_,
    new_n15888_, new_n15889_, new_n15891_, new_n15892_, new_n15893_,
    new_n15894_, new_n15895_, new_n15896_, new_n15898_, new_n15899_,
    new_n15900_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15932_, new_n15934_, new_n15935_, new_n15936_, new_n15937_,
    new_n15938_, new_n15939_, new_n15941_, new_n15942_, new_n15943_,
    new_n15944_, new_n15945_, new_n15946_, new_n15948_, new_n15949_,
    new_n15950_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15982_, new_n15984_, new_n15985_, new_n15986_, new_n15987_,
    new_n15988_, new_n15989_, new_n15991_, new_n15992_, new_n15993_,
    new_n15994_, new_n15995_, new_n15996_, new_n15998_, new_n15999_,
    new_n16000_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16032_, new_n16034_, new_n16035_, new_n16036_, new_n16037_,
    new_n16038_, new_n16039_, new_n16041_, new_n16042_, new_n16043_,
    new_n16044_, new_n16045_, new_n16046_, new_n16048_, new_n16049_,
    new_n16050_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16082_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16091_, new_n16092_, new_n16093_,
    new_n16094_, new_n16095_, new_n16096_, new_n16098_, new_n16099_,
    new_n16100_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16132_, new_n16134_, new_n16135_, new_n16136_, new_n16137_,
    new_n16138_, new_n16139_, new_n16141_, new_n16142_, new_n16143_,
    new_n16144_, new_n16145_, new_n16146_, new_n16148_, new_n16149_,
    new_n16150_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16182_, new_n16184_, new_n16185_, new_n16186_, new_n16187_,
    new_n16188_, new_n16189_, new_n16191_, new_n16192_, new_n16193_,
    new_n16194_, new_n16195_, new_n16196_, new_n16198_, new_n16199_,
    new_n16200_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16242_,
    new_n16243_, new_n16245_, new_n16246_, new_n16248_, new_n16249_;
  assign new_n1251_ = B5185 & B5186;
  assign new_n1252_ = ~B5185 & ~B5186;
  assign new_n1253_ = ~new_n1251_ & ~new_n1252_;
  assign new_n1254_ = ~B5182 & B5183;
  assign new_n1255_ = B5182 & ~B5183;
  assign new_n1256_ = ~new_n1254_ & ~new_n1255_;
  assign new_n1257_ = ~B5185 & ~new_n1256_;
  assign new_n1258_ = B5185 & new_n1256_;
  assign new_n1259_ = ~new_n1257_ & ~new_n1258_;
  assign new_n1260_ = new_n1253_ & ~new_n1259_;
  assign new_n1261_ = B5184 & ~new_n1260_;
  assign new_n1262_ = ~B5184 & new_n1260_;
  assign new_n1263_ = ~new_n1261_ & ~new_n1262_;
  assign new_n1264_ = ~new_n1256_ & ~new_n1263_;
  assign new_n1265_ = B5216 & ~B5215;
  assign new_n1266_ = ~B5216 & B5215;
  assign new_n1267_ = ~new_n1265_ & ~new_n1266_;
  assign new_n1268_ = ~B5218 & new_n1267_;
  assign new_n1269_ = ~B5219 & ~B5218;
  assign new_n1270_ = ~new_n1268_ & ~new_n1269_;
  assign new_n1271_ = B5217 & new_n1270_;
  assign new_n1272_ = ~B5217 & ~new_n1270_;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1274_ = ~new_n1267_ & ~new_n1273_;
  assign new_n1275_ = ~new_n1264_ & new_n1274_;
  assign new_n1276_ = new_n1264_ & ~new_n1274_;
  assign new_n1277_ = ~new_n1275_ & ~new_n1276_;
  assign new_n1278_ = B5249 & ~B5248;
  assign new_n1279_ = ~B5249 & B5248;
  assign new_n1280_ = ~new_n1278_ & ~new_n1279_;
  assign new_n1281_ = ~B5251 & new_n1280_;
  assign new_n1282_ = ~B5252 & ~B5251;
  assign new_n1283_ = ~new_n1281_ & ~new_n1282_;
  assign new_n1284_ = B5250 & new_n1283_;
  assign new_n1285_ = ~B5250 & ~new_n1283_;
  assign new_n1286_ = ~new_n1284_ & ~new_n1285_;
  assign new_n1287_ = ~new_n1280_ & ~new_n1286_;
  assign new_n1288_ = B5282 & ~B5281;
  assign new_n1289_ = ~B5282 & B5281;
  assign new_n1290_ = ~new_n1288_ & ~new_n1289_;
  assign new_n1291_ = ~B5284 & new_n1290_;
  assign new_n1292_ = ~B5285 & ~B5284;
  assign new_n1293_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1294_ = B5283 & new_n1293_;
  assign new_n1295_ = ~B5283 & ~new_n1293_;
  assign new_n1296_ = ~new_n1294_ & ~new_n1295_;
  assign new_n1297_ = ~new_n1290_ & ~new_n1296_;
  assign new_n1298_ = new_n1277_ & ~new_n1297_;
  assign new_n1299_ = B5315 & ~B5314;
  assign new_n1300_ = ~B5315 & B5314;
  assign new_n1301_ = ~new_n1299_ & ~new_n1300_;
  assign new_n1302_ = ~B5317 & new_n1301_;
  assign new_n1303_ = ~B5318 & ~B5317;
  assign new_n1304_ = ~new_n1302_ & ~new_n1303_;
  assign new_n1305_ = B5316 & new_n1304_;
  assign new_n1306_ = ~B5316 & ~new_n1304_;
  assign new_n1307_ = ~new_n1305_ & ~new_n1306_;
  assign new_n1308_ = ~new_n1301_ & ~new_n1307_;
  assign new_n1309_ = ~new_n1297_ & ~new_n1308_;
  assign new_n1310_ = ~new_n1298_ & ~new_n1309_;
  assign new_n1311_ = new_n1287_ & new_n1310_;
  assign new_n1312_ = ~new_n1287_ & ~new_n1310_;
  assign new_n1313_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1314_ = ~new_n1277_ & ~new_n1313_;
  assign new_n1315_ = B5348 & ~B5347;
  assign new_n1316_ = ~B5348 & B5347;
  assign new_n1317_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1318_ = ~B5350 & new_n1317_;
  assign new_n1319_ = ~B5351 & ~B5350;
  assign new_n1320_ = ~new_n1318_ & ~new_n1319_;
  assign new_n1321_ = B5349 & new_n1320_;
  assign new_n1322_ = ~B5349 & ~new_n1320_;
  assign new_n1323_ = ~new_n1321_ & ~new_n1322_;
  assign new_n1324_ = ~new_n1317_ & ~new_n1323_;
  assign new_n1325_ = B5381 & ~B5380;
  assign new_n1326_ = ~B5381 & B5380;
  assign new_n1327_ = ~new_n1325_ & ~new_n1326_;
  assign new_n1328_ = ~B5383 & new_n1327_;
  assign new_n1329_ = ~B5384 & ~B5383;
  assign new_n1330_ = ~new_n1328_ & ~new_n1329_;
  assign new_n1331_ = B5382 & new_n1330_;
  assign new_n1332_ = ~B5382 & ~new_n1330_;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = ~new_n1327_ & ~new_n1333_;
  assign new_n1335_ = ~new_n1324_ & new_n1334_;
  assign new_n1336_ = new_n1324_ & ~new_n1334_;
  assign new_n1337_ = ~new_n1335_ & ~new_n1336_;
  assign new_n1338_ = B5414 & ~B5413;
  assign new_n1339_ = ~B5414 & B5413;
  assign new_n1340_ = ~new_n1338_ & ~new_n1339_;
  assign new_n1341_ = ~B5416 & new_n1340_;
  assign new_n1342_ = ~B5417 & ~B5416;
  assign new_n1343_ = ~new_n1341_ & ~new_n1342_;
  assign new_n1344_ = B5415 & new_n1343_;
  assign new_n1345_ = ~B5415 & ~new_n1343_;
  assign new_n1346_ = ~new_n1344_ & ~new_n1345_;
  assign new_n1347_ = ~new_n1340_ & ~new_n1346_;
  assign new_n1348_ = B5447 & ~B5446;
  assign new_n1349_ = ~B5447 & B5446;
  assign new_n1350_ = ~new_n1348_ & ~new_n1349_;
  assign new_n1351_ = ~B5449 & new_n1350_;
  assign new_n1352_ = ~B5450 & ~B5449;
  assign new_n1353_ = ~new_n1351_ & ~new_n1352_;
  assign new_n1354_ = B5448 & new_n1353_;
  assign new_n1355_ = ~B5448 & ~new_n1353_;
  assign new_n1356_ = ~new_n1354_ & ~new_n1355_;
  assign new_n1357_ = ~new_n1350_ & ~new_n1356_;
  assign new_n1358_ = new_n1337_ & ~new_n1357_;
  assign new_n1359_ = B5480 & ~B5479;
  assign new_n1360_ = ~B5480 & B5479;
  assign new_n1361_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1362_ = ~B5482 & new_n1361_;
  assign new_n1363_ = ~B5483 & ~B5482;
  assign new_n1364_ = ~new_n1362_ & ~new_n1363_;
  assign new_n1365_ = B5481 & new_n1364_;
  assign new_n1366_ = ~B5481 & ~new_n1364_;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign new_n1368_ = ~new_n1361_ & ~new_n1367_;
  assign new_n1369_ = ~new_n1357_ & ~new_n1368_;
  assign new_n1370_ = ~new_n1358_ & ~new_n1369_;
  assign new_n1371_ = new_n1347_ & new_n1370_;
  assign new_n1372_ = ~new_n1347_ & ~new_n1370_;
  assign new_n1373_ = ~new_n1371_ & ~new_n1372_;
  assign new_n1374_ = ~new_n1337_ & ~new_n1373_;
  assign new_n1375_ = ~new_n1314_ & new_n1374_;
  assign new_n1376_ = new_n1314_ & ~new_n1374_;
  assign new_n1377_ = ~new_n1375_ & ~new_n1376_;
  assign new_n1378_ = B5513 & ~B5512;
  assign new_n1379_ = ~B5513 & B5512;
  assign new_n1380_ = ~new_n1378_ & ~new_n1379_;
  assign new_n1381_ = ~B5515 & new_n1380_;
  assign new_n1382_ = ~B5516 & ~B5515;
  assign new_n1383_ = ~new_n1381_ & ~new_n1382_;
  assign new_n1384_ = B5514 & new_n1383_;
  assign new_n1385_ = ~B5514 & ~new_n1383_;
  assign new_n1386_ = ~new_n1384_ & ~new_n1385_;
  assign new_n1387_ = ~new_n1380_ & ~new_n1386_;
  assign new_n1388_ = B5546 & ~B5545;
  assign new_n1389_ = ~B5546 & B5545;
  assign new_n1390_ = ~new_n1388_ & ~new_n1389_;
  assign new_n1391_ = ~B5548 & new_n1390_;
  assign new_n1392_ = ~B5549 & ~B5548;
  assign new_n1393_ = ~new_n1391_ & ~new_n1392_;
  assign new_n1394_ = B5547 & new_n1393_;
  assign new_n1395_ = ~B5547 & ~new_n1393_;
  assign new_n1396_ = ~new_n1394_ & ~new_n1395_;
  assign new_n1397_ = ~new_n1390_ & ~new_n1396_;
  assign new_n1398_ = ~new_n1387_ & new_n1397_;
  assign new_n1399_ = new_n1387_ & ~new_n1397_;
  assign new_n1400_ = ~new_n1398_ & ~new_n1399_;
  assign new_n1401_ = B5579 & ~B5578;
  assign new_n1402_ = ~B5579 & B5578;
  assign new_n1403_ = ~new_n1401_ & ~new_n1402_;
  assign new_n1404_ = ~B5581 & new_n1403_;
  assign new_n1405_ = ~B5582 & ~B5581;
  assign new_n1406_ = ~new_n1404_ & ~new_n1405_;
  assign new_n1407_ = B5580 & new_n1406_;
  assign new_n1408_ = ~B5580 & ~new_n1406_;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1410_ = ~new_n1403_ & ~new_n1409_;
  assign new_n1411_ = B5612 & ~B5611;
  assign new_n1412_ = ~B5612 & B5611;
  assign new_n1413_ = ~new_n1411_ & ~new_n1412_;
  assign new_n1414_ = ~B5614 & new_n1413_;
  assign new_n1415_ = ~B5615 & ~B5614;
  assign new_n1416_ = ~new_n1414_ & ~new_n1415_;
  assign new_n1417_ = B5613 & new_n1416_;
  assign new_n1418_ = ~B5613 & ~new_n1416_;
  assign new_n1419_ = ~new_n1417_ & ~new_n1418_;
  assign new_n1420_ = ~new_n1413_ & ~new_n1419_;
  assign new_n1421_ = new_n1400_ & ~new_n1420_;
  assign new_n1422_ = B5645 & ~B5644;
  assign new_n1423_ = ~B5645 & B5644;
  assign new_n1424_ = ~new_n1422_ & ~new_n1423_;
  assign new_n1425_ = ~B5647 & new_n1424_;
  assign new_n1426_ = ~B5648 & ~B5647;
  assign new_n1427_ = ~new_n1425_ & ~new_n1426_;
  assign new_n1428_ = B5646 & new_n1427_;
  assign new_n1429_ = ~B5646 & ~new_n1427_;
  assign new_n1430_ = ~new_n1428_ & ~new_n1429_;
  assign new_n1431_ = ~new_n1424_ & ~new_n1430_;
  assign new_n1432_ = ~new_n1420_ & ~new_n1431_;
  assign new_n1433_ = ~new_n1421_ & ~new_n1432_;
  assign new_n1434_ = new_n1410_ & new_n1433_;
  assign new_n1435_ = ~new_n1410_ & ~new_n1433_;
  assign new_n1436_ = ~new_n1434_ & ~new_n1435_;
  assign new_n1437_ = ~new_n1400_ & ~new_n1436_;
  assign new_n1438_ = B5678 & ~B5677;
  assign new_n1439_ = ~B5678 & B5677;
  assign new_n1440_ = ~new_n1438_ & ~new_n1439_;
  assign new_n1441_ = ~B5680 & new_n1440_;
  assign new_n1442_ = ~B5681 & ~B5680;
  assign new_n1443_ = ~new_n1441_ & ~new_n1442_;
  assign new_n1444_ = B5679 & new_n1443_;
  assign new_n1445_ = ~B5679 & ~new_n1443_;
  assign new_n1446_ = ~new_n1444_ & ~new_n1445_;
  assign new_n1447_ = ~new_n1440_ & ~new_n1446_;
  assign new_n1448_ = B5711 & ~B5710;
  assign new_n1449_ = ~B5711 & B5710;
  assign new_n1450_ = ~new_n1448_ & ~new_n1449_;
  assign new_n1451_ = ~B5713 & new_n1450_;
  assign new_n1452_ = ~B5714 & ~B5713;
  assign new_n1453_ = ~new_n1451_ & ~new_n1452_;
  assign new_n1454_ = B5712 & new_n1453_;
  assign new_n1455_ = ~B5712 & ~new_n1453_;
  assign new_n1456_ = ~new_n1454_ & ~new_n1455_;
  assign new_n1457_ = ~new_n1450_ & ~new_n1456_;
  assign new_n1458_ = ~new_n1447_ & new_n1457_;
  assign new_n1459_ = new_n1447_ & ~new_n1457_;
  assign new_n1460_ = ~new_n1458_ & ~new_n1459_;
  assign new_n1461_ = B5744 & ~B5743;
  assign new_n1462_ = ~B5744 & B5743;
  assign new_n1463_ = ~new_n1461_ & ~new_n1462_;
  assign new_n1464_ = ~B5746 & new_n1463_;
  assign new_n1465_ = ~B5747 & ~B5746;
  assign new_n1466_ = ~new_n1464_ & ~new_n1465_;
  assign new_n1467_ = B5745 & new_n1466_;
  assign new_n1468_ = ~B5745 & ~new_n1466_;
  assign new_n1469_ = ~new_n1467_ & ~new_n1468_;
  assign new_n1470_ = ~new_n1463_ & ~new_n1469_;
  assign new_n1471_ = B5777 & ~B5776;
  assign new_n1472_ = ~B5777 & B5776;
  assign new_n1473_ = ~new_n1471_ & ~new_n1472_;
  assign new_n1474_ = ~B5779 & new_n1473_;
  assign new_n1475_ = ~B5780 & ~B5779;
  assign new_n1476_ = ~new_n1474_ & ~new_n1475_;
  assign new_n1477_ = B5778 & new_n1476_;
  assign new_n1478_ = ~B5778 & ~new_n1476_;
  assign new_n1479_ = ~new_n1477_ & ~new_n1478_;
  assign new_n1480_ = ~new_n1473_ & ~new_n1479_;
  assign new_n1481_ = new_n1460_ & ~new_n1480_;
  assign new_n1482_ = B5810 & ~B5809;
  assign new_n1483_ = ~B5810 & B5809;
  assign new_n1484_ = ~new_n1482_ & ~new_n1483_;
  assign new_n1485_ = ~B5812 & new_n1484_;
  assign new_n1486_ = ~B5813 & ~B5812;
  assign new_n1487_ = ~new_n1485_ & ~new_n1486_;
  assign new_n1488_ = B5811 & new_n1487_;
  assign new_n1489_ = ~B5811 & ~new_n1487_;
  assign new_n1490_ = ~new_n1488_ & ~new_n1489_;
  assign new_n1491_ = ~new_n1484_ & ~new_n1490_;
  assign new_n1492_ = ~new_n1480_ & ~new_n1491_;
  assign new_n1493_ = ~new_n1481_ & ~new_n1492_;
  assign new_n1494_ = new_n1470_ & new_n1493_;
  assign new_n1495_ = ~new_n1470_ & ~new_n1493_;
  assign new_n1496_ = ~new_n1494_ & ~new_n1495_;
  assign new_n1497_ = ~new_n1460_ & ~new_n1496_;
  assign new_n1498_ = new_n1377_ & ~new_n1497_;
  assign new_n1499_ = B5843 & ~B5842;
  assign new_n1500_ = ~B5843 & B5842;
  assign new_n1501_ = ~new_n1499_ & ~new_n1500_;
  assign new_n1502_ = ~B5845 & new_n1501_;
  assign new_n1503_ = ~B5846 & ~B5845;
  assign new_n1504_ = ~new_n1502_ & ~new_n1503_;
  assign new_n1505_ = B5844 & new_n1504_;
  assign new_n1506_ = ~B5844 & ~new_n1504_;
  assign new_n1507_ = ~new_n1505_ & ~new_n1506_;
  assign new_n1508_ = ~new_n1501_ & ~new_n1507_;
  assign new_n1509_ = B5876 & ~B5875;
  assign new_n1510_ = ~B5876 & B5875;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign new_n1512_ = ~B5878 & new_n1511_;
  assign new_n1513_ = ~B5879 & ~B5878;
  assign new_n1514_ = ~new_n1512_ & ~new_n1513_;
  assign new_n1515_ = B5877 & new_n1514_;
  assign new_n1516_ = ~B5877 & ~new_n1514_;
  assign new_n1517_ = ~new_n1515_ & ~new_n1516_;
  assign new_n1518_ = ~new_n1511_ & ~new_n1517_;
  assign new_n1519_ = ~new_n1508_ & new_n1518_;
  assign new_n1520_ = new_n1508_ & ~new_n1518_;
  assign new_n1521_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1522_ = B5909 & ~B5908;
  assign new_n1523_ = ~B5909 & B5908;
  assign new_n1524_ = ~new_n1522_ & ~new_n1523_;
  assign new_n1525_ = ~B5911 & new_n1524_;
  assign new_n1526_ = ~B5912 & ~B5911;
  assign new_n1527_ = ~new_n1525_ & ~new_n1526_;
  assign new_n1528_ = B5910 & new_n1527_;
  assign new_n1529_ = ~B5910 & ~new_n1527_;
  assign new_n1530_ = ~new_n1528_ & ~new_n1529_;
  assign new_n1531_ = ~new_n1524_ & ~new_n1530_;
  assign new_n1532_ = B5942 & ~B5941;
  assign new_n1533_ = ~B5942 & B5941;
  assign new_n1534_ = ~new_n1532_ & ~new_n1533_;
  assign new_n1535_ = ~B5944 & new_n1534_;
  assign new_n1536_ = ~B5945 & ~B5944;
  assign new_n1537_ = ~new_n1535_ & ~new_n1536_;
  assign new_n1538_ = B5943 & new_n1537_;
  assign new_n1539_ = ~B5943 & ~new_n1537_;
  assign new_n1540_ = ~new_n1538_ & ~new_n1539_;
  assign new_n1541_ = ~new_n1534_ & ~new_n1540_;
  assign new_n1542_ = new_n1521_ & ~new_n1541_;
  assign new_n1543_ = B5975 & ~B5974;
  assign new_n1544_ = ~B5975 & B5974;
  assign new_n1545_ = ~new_n1543_ & ~new_n1544_;
  assign new_n1546_ = ~B5977 & new_n1545_;
  assign new_n1547_ = ~B5978 & ~B5977;
  assign new_n1548_ = ~new_n1546_ & ~new_n1547_;
  assign new_n1549_ = B5976 & new_n1548_;
  assign new_n1550_ = ~B5976 & ~new_n1548_;
  assign new_n1551_ = ~new_n1549_ & ~new_n1550_;
  assign new_n1552_ = ~new_n1545_ & ~new_n1551_;
  assign new_n1553_ = ~new_n1541_ & ~new_n1552_;
  assign new_n1554_ = ~new_n1542_ & ~new_n1553_;
  assign new_n1555_ = new_n1531_ & new_n1554_;
  assign new_n1556_ = ~new_n1531_ & ~new_n1554_;
  assign new_n1557_ = ~new_n1555_ & ~new_n1556_;
  assign new_n1558_ = ~new_n1521_ & ~new_n1557_;
  assign new_n1559_ = ~new_n1497_ & ~new_n1558_;
  assign new_n1560_ = ~new_n1498_ & ~new_n1559_;
  assign new_n1561_ = new_n1437_ & new_n1560_;
  assign new_n1562_ = ~new_n1437_ & ~new_n1560_;
  assign new_n1563_ = ~new_n1561_ & ~new_n1562_;
  assign new_n1564_ = ~new_n1377_ & ~new_n1563_;
  assign new_n1565_ = B6008 & ~B6007;
  assign new_n1566_ = ~B6008 & B6007;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = ~B6010 & new_n1567_;
  assign new_n1569_ = ~B6011 & ~B6010;
  assign new_n1570_ = ~new_n1568_ & ~new_n1569_;
  assign new_n1571_ = B6009 & new_n1570_;
  assign new_n1572_ = ~B6009 & ~new_n1570_;
  assign new_n1573_ = ~new_n1571_ & ~new_n1572_;
  assign new_n1574_ = ~new_n1567_ & ~new_n1573_;
  assign new_n1575_ = B6041 & ~B6040;
  assign new_n1576_ = ~B6041 & B6040;
  assign new_n1577_ = ~new_n1575_ & ~new_n1576_;
  assign new_n1578_ = ~B6043 & new_n1577_;
  assign new_n1579_ = ~B6044 & ~B6043;
  assign new_n1580_ = ~new_n1578_ & ~new_n1579_;
  assign new_n1581_ = B6042 & new_n1580_;
  assign new_n1582_ = ~B6042 & ~new_n1580_;
  assign new_n1583_ = ~new_n1581_ & ~new_n1582_;
  assign new_n1584_ = ~new_n1577_ & ~new_n1583_;
  assign new_n1585_ = ~new_n1574_ & new_n1584_;
  assign new_n1586_ = new_n1574_ & ~new_n1584_;
  assign new_n1587_ = ~new_n1585_ & ~new_n1586_;
  assign new_n1588_ = B6074 & ~B6073;
  assign new_n1589_ = ~B6074 & B6073;
  assign new_n1590_ = ~new_n1588_ & ~new_n1589_;
  assign new_n1591_ = ~B6076 & new_n1590_;
  assign new_n1592_ = ~B6077 & ~B6076;
  assign new_n1593_ = ~new_n1591_ & ~new_n1592_;
  assign new_n1594_ = B6075 & new_n1593_;
  assign new_n1595_ = ~B6075 & ~new_n1593_;
  assign new_n1596_ = ~new_n1594_ & ~new_n1595_;
  assign new_n1597_ = ~new_n1590_ & ~new_n1596_;
  assign new_n1598_ = B6107 & ~B6106;
  assign new_n1599_ = ~B6107 & B6106;
  assign new_n1600_ = ~new_n1598_ & ~new_n1599_;
  assign new_n1601_ = ~B6109 & new_n1600_;
  assign new_n1602_ = ~B6110 & ~B6109;
  assign new_n1603_ = ~new_n1601_ & ~new_n1602_;
  assign new_n1604_ = B6108 & new_n1603_;
  assign new_n1605_ = ~B6108 & ~new_n1603_;
  assign new_n1606_ = ~new_n1604_ & ~new_n1605_;
  assign new_n1607_ = ~new_n1600_ & ~new_n1606_;
  assign new_n1608_ = new_n1587_ & ~new_n1607_;
  assign new_n1609_ = B6140 & ~B6139;
  assign new_n1610_ = ~B6140 & B6139;
  assign new_n1611_ = ~new_n1609_ & ~new_n1610_;
  assign new_n1612_ = ~B6142 & new_n1611_;
  assign new_n1613_ = ~B6143 & ~B6142;
  assign new_n1614_ = ~new_n1612_ & ~new_n1613_;
  assign new_n1615_ = B6141 & new_n1614_;
  assign new_n1616_ = ~B6141 & ~new_n1614_;
  assign new_n1617_ = ~new_n1615_ & ~new_n1616_;
  assign new_n1618_ = ~new_n1611_ & ~new_n1617_;
  assign new_n1619_ = ~new_n1607_ & ~new_n1618_;
  assign new_n1620_ = ~new_n1608_ & ~new_n1619_;
  assign new_n1621_ = new_n1597_ & new_n1620_;
  assign new_n1622_ = ~new_n1597_ & ~new_n1620_;
  assign new_n1623_ = ~new_n1621_ & ~new_n1622_;
  assign new_n1624_ = ~new_n1587_ & ~new_n1623_;
  assign new_n1625_ = B6173 & ~B6172;
  assign new_n1626_ = ~B6173 & B6172;
  assign new_n1627_ = ~new_n1625_ & ~new_n1626_;
  assign new_n1628_ = ~B6175 & new_n1627_;
  assign new_n1629_ = ~B6176 & ~B6175;
  assign new_n1630_ = ~new_n1628_ & ~new_n1629_;
  assign new_n1631_ = B6174 & new_n1630_;
  assign new_n1632_ = ~B6174 & ~new_n1630_;
  assign new_n1633_ = ~new_n1631_ & ~new_n1632_;
  assign new_n1634_ = ~new_n1627_ & ~new_n1633_;
  assign new_n1635_ = B6206 & ~B6205;
  assign new_n1636_ = ~B6206 & B6205;
  assign new_n1637_ = ~new_n1635_ & ~new_n1636_;
  assign new_n1638_ = ~B6208 & new_n1637_;
  assign new_n1639_ = ~B6209 & ~B6208;
  assign new_n1640_ = ~new_n1638_ & ~new_n1639_;
  assign new_n1641_ = B6207 & new_n1640_;
  assign new_n1642_ = ~B6207 & ~new_n1640_;
  assign new_n1643_ = ~new_n1641_ & ~new_n1642_;
  assign new_n1644_ = ~new_n1637_ & ~new_n1643_;
  assign new_n1645_ = ~new_n1634_ & new_n1644_;
  assign new_n1646_ = new_n1634_ & ~new_n1644_;
  assign new_n1647_ = ~new_n1645_ & ~new_n1646_;
  assign new_n1648_ = B6239 & ~B6238;
  assign new_n1649_ = ~B6239 & B6238;
  assign new_n1650_ = ~new_n1648_ & ~new_n1649_;
  assign new_n1651_ = ~B6241 & new_n1650_;
  assign new_n1652_ = ~B6242 & ~B6241;
  assign new_n1653_ = ~new_n1651_ & ~new_n1652_;
  assign new_n1654_ = B6240 & new_n1653_;
  assign new_n1655_ = ~B6240 & ~new_n1653_;
  assign new_n1656_ = ~new_n1654_ & ~new_n1655_;
  assign new_n1657_ = ~new_n1650_ & ~new_n1656_;
  assign new_n1658_ = B6272 & ~B6271;
  assign new_n1659_ = ~B6272 & B6271;
  assign new_n1660_ = ~new_n1658_ & ~new_n1659_;
  assign new_n1661_ = ~B6274 & new_n1660_;
  assign new_n1662_ = ~B6275 & ~B6274;
  assign new_n1663_ = ~new_n1661_ & ~new_n1662_;
  assign new_n1664_ = B6273 & new_n1663_;
  assign new_n1665_ = ~B6273 & ~new_n1663_;
  assign new_n1666_ = ~new_n1664_ & ~new_n1665_;
  assign new_n1667_ = ~new_n1660_ & ~new_n1666_;
  assign new_n1668_ = new_n1647_ & ~new_n1667_;
  assign new_n1669_ = B6305 & ~B6304;
  assign new_n1670_ = ~B6305 & B6304;
  assign new_n1671_ = ~new_n1669_ & ~new_n1670_;
  assign new_n1672_ = ~B6307 & new_n1671_;
  assign new_n1673_ = ~B6308 & ~B6307;
  assign new_n1674_ = ~new_n1672_ & ~new_n1673_;
  assign new_n1675_ = B6306 & new_n1674_;
  assign new_n1676_ = ~B6306 & ~new_n1674_;
  assign new_n1677_ = ~new_n1675_ & ~new_n1676_;
  assign new_n1678_ = ~new_n1671_ & ~new_n1677_;
  assign new_n1679_ = ~new_n1667_ & ~new_n1678_;
  assign new_n1680_ = ~new_n1668_ & ~new_n1679_;
  assign new_n1681_ = new_n1657_ & new_n1680_;
  assign new_n1682_ = ~new_n1657_ & ~new_n1680_;
  assign new_n1683_ = ~new_n1681_ & ~new_n1682_;
  assign new_n1684_ = ~new_n1647_ & ~new_n1683_;
  assign new_n1685_ = ~new_n1624_ & new_n1684_;
  assign new_n1686_ = new_n1624_ & ~new_n1684_;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = B6338 & ~B6337;
  assign new_n1689_ = ~B6338 & B6337;
  assign new_n1690_ = ~new_n1688_ & ~new_n1689_;
  assign new_n1691_ = ~B6340 & new_n1690_;
  assign new_n1692_ = ~B6341 & ~B6340;
  assign new_n1693_ = ~new_n1691_ & ~new_n1692_;
  assign new_n1694_ = B6339 & new_n1693_;
  assign new_n1695_ = ~B6339 & ~new_n1693_;
  assign new_n1696_ = ~new_n1694_ & ~new_n1695_;
  assign new_n1697_ = ~new_n1690_ & ~new_n1696_;
  assign new_n1698_ = B6371 & ~B6370;
  assign new_n1699_ = ~B6371 & B6370;
  assign new_n1700_ = ~new_n1698_ & ~new_n1699_;
  assign new_n1701_ = ~B6373 & new_n1700_;
  assign new_n1702_ = ~B6374 & ~B6373;
  assign new_n1703_ = ~new_n1701_ & ~new_n1702_;
  assign new_n1704_ = B6372 & new_n1703_;
  assign new_n1705_ = ~B6372 & ~new_n1703_;
  assign new_n1706_ = ~new_n1704_ & ~new_n1705_;
  assign new_n1707_ = ~new_n1700_ & ~new_n1706_;
  assign new_n1708_ = ~new_n1697_ & new_n1707_;
  assign new_n1709_ = new_n1697_ & ~new_n1707_;
  assign new_n1710_ = ~new_n1708_ & ~new_n1709_;
  assign new_n1711_ = B6404 & ~B6403;
  assign new_n1712_ = ~B6404 & B6403;
  assign new_n1713_ = ~new_n1711_ & ~new_n1712_;
  assign new_n1714_ = ~B6406 & new_n1713_;
  assign new_n1715_ = ~B6407 & ~B6406;
  assign new_n1716_ = ~new_n1714_ & ~new_n1715_;
  assign new_n1717_ = B6405 & new_n1716_;
  assign new_n1718_ = ~B6405 & ~new_n1716_;
  assign new_n1719_ = ~new_n1717_ & ~new_n1718_;
  assign new_n1720_ = ~new_n1713_ & ~new_n1719_;
  assign new_n1721_ = B6437 & ~B6436;
  assign new_n1722_ = ~B6437 & B6436;
  assign new_n1723_ = ~new_n1721_ & ~new_n1722_;
  assign new_n1724_ = ~B6439 & new_n1723_;
  assign new_n1725_ = ~B6440 & ~B6439;
  assign new_n1726_ = ~new_n1724_ & ~new_n1725_;
  assign new_n1727_ = B6438 & new_n1726_;
  assign new_n1728_ = ~B6438 & ~new_n1726_;
  assign new_n1729_ = ~new_n1727_ & ~new_n1728_;
  assign new_n1730_ = ~new_n1723_ & ~new_n1729_;
  assign new_n1731_ = new_n1710_ & ~new_n1730_;
  assign new_n1732_ = B6470 & ~B6469;
  assign new_n1733_ = ~B6470 & B6469;
  assign new_n1734_ = ~new_n1732_ & ~new_n1733_;
  assign new_n1735_ = ~B6472 & new_n1734_;
  assign new_n1736_ = ~B6473 & ~B6472;
  assign new_n1737_ = ~new_n1735_ & ~new_n1736_;
  assign new_n1738_ = B6471 & new_n1737_;
  assign new_n1739_ = ~B6471 & ~new_n1737_;
  assign new_n1740_ = ~new_n1738_ & ~new_n1739_;
  assign new_n1741_ = ~new_n1734_ & ~new_n1740_;
  assign new_n1742_ = ~new_n1730_ & ~new_n1741_;
  assign new_n1743_ = ~new_n1731_ & ~new_n1742_;
  assign new_n1744_ = new_n1720_ & new_n1743_;
  assign new_n1745_ = ~new_n1720_ & ~new_n1743_;
  assign new_n1746_ = ~new_n1744_ & ~new_n1745_;
  assign new_n1747_ = ~new_n1710_ & ~new_n1746_;
  assign new_n1748_ = B6503 & ~B6502;
  assign new_n1749_ = ~B6503 & B6502;
  assign new_n1750_ = ~new_n1748_ & ~new_n1749_;
  assign new_n1751_ = ~B6505 & new_n1750_;
  assign new_n1752_ = ~B6506 & ~B6505;
  assign new_n1753_ = ~new_n1751_ & ~new_n1752_;
  assign new_n1754_ = B6504 & new_n1753_;
  assign new_n1755_ = ~B6504 & ~new_n1753_;
  assign new_n1756_ = ~new_n1754_ & ~new_n1755_;
  assign new_n1757_ = ~new_n1750_ & ~new_n1756_;
  assign new_n1758_ = B6536 & ~B6535;
  assign new_n1759_ = ~B6536 & B6535;
  assign new_n1760_ = ~new_n1758_ & ~new_n1759_;
  assign new_n1761_ = ~B6538 & new_n1760_;
  assign new_n1762_ = ~B6539 & ~B6538;
  assign new_n1763_ = ~new_n1761_ & ~new_n1762_;
  assign new_n1764_ = B6537 & new_n1763_;
  assign new_n1765_ = ~B6537 & ~new_n1763_;
  assign new_n1766_ = ~new_n1764_ & ~new_n1765_;
  assign new_n1767_ = ~new_n1760_ & ~new_n1766_;
  assign new_n1768_ = ~new_n1757_ & new_n1767_;
  assign new_n1769_ = new_n1757_ & ~new_n1767_;
  assign new_n1770_ = ~new_n1768_ & ~new_n1769_;
  assign new_n1771_ = B6569 & ~B6568;
  assign new_n1772_ = ~B6569 & B6568;
  assign new_n1773_ = ~new_n1771_ & ~new_n1772_;
  assign new_n1774_ = ~B6571 & new_n1773_;
  assign new_n1775_ = ~B6572 & ~B6571;
  assign new_n1776_ = ~new_n1774_ & ~new_n1775_;
  assign new_n1777_ = B6570 & new_n1776_;
  assign new_n1778_ = ~B6570 & ~new_n1776_;
  assign new_n1779_ = ~new_n1777_ & ~new_n1778_;
  assign new_n1780_ = ~new_n1773_ & ~new_n1779_;
  assign new_n1781_ = B6602 & ~B6601;
  assign new_n1782_ = ~B6602 & B6601;
  assign new_n1783_ = ~new_n1781_ & ~new_n1782_;
  assign new_n1784_ = ~B6604 & new_n1783_;
  assign new_n1785_ = ~B6605 & ~B6604;
  assign new_n1786_ = ~new_n1784_ & ~new_n1785_;
  assign new_n1787_ = B6603 & new_n1786_;
  assign new_n1788_ = ~B6603 & ~new_n1786_;
  assign new_n1789_ = ~new_n1787_ & ~new_n1788_;
  assign new_n1790_ = ~new_n1783_ & ~new_n1789_;
  assign new_n1791_ = new_n1770_ & ~new_n1790_;
  assign new_n1792_ = B6635 & ~B6634;
  assign new_n1793_ = ~B6635 & B6634;
  assign new_n1794_ = ~new_n1792_ & ~new_n1793_;
  assign new_n1795_ = ~B6637 & new_n1794_;
  assign new_n1796_ = ~B6638 & ~B6637;
  assign new_n1797_ = ~new_n1795_ & ~new_n1796_;
  assign new_n1798_ = B6636 & new_n1797_;
  assign new_n1799_ = ~B6636 & ~new_n1797_;
  assign new_n1800_ = ~new_n1798_ & ~new_n1799_;
  assign new_n1801_ = ~new_n1794_ & ~new_n1800_;
  assign new_n1802_ = ~new_n1790_ & ~new_n1801_;
  assign new_n1803_ = ~new_n1791_ & ~new_n1802_;
  assign new_n1804_ = new_n1780_ & new_n1803_;
  assign new_n1805_ = ~new_n1780_ & ~new_n1803_;
  assign new_n1806_ = ~new_n1804_ & ~new_n1805_;
  assign new_n1807_ = ~new_n1770_ & ~new_n1806_;
  assign new_n1808_ = new_n1687_ & ~new_n1807_;
  assign new_n1809_ = B6668 & ~B6667;
  assign new_n1810_ = ~B6668 & B6667;
  assign new_n1811_ = ~new_n1809_ & ~new_n1810_;
  assign new_n1812_ = ~B6670 & new_n1811_;
  assign new_n1813_ = ~B6671 & ~B6670;
  assign new_n1814_ = ~new_n1812_ & ~new_n1813_;
  assign new_n1815_ = B6669 & new_n1814_;
  assign new_n1816_ = ~B6669 & ~new_n1814_;
  assign new_n1817_ = ~new_n1815_ & ~new_n1816_;
  assign new_n1818_ = ~new_n1811_ & ~new_n1817_;
  assign new_n1819_ = B6701 & ~B6700;
  assign new_n1820_ = ~B6701 & B6700;
  assign new_n1821_ = ~new_n1819_ & ~new_n1820_;
  assign new_n1822_ = ~B6703 & new_n1821_;
  assign new_n1823_ = ~B6704 & ~B6703;
  assign new_n1824_ = ~new_n1822_ & ~new_n1823_;
  assign new_n1825_ = B6702 & new_n1824_;
  assign new_n1826_ = ~B6702 & ~new_n1824_;
  assign new_n1827_ = ~new_n1825_ & ~new_n1826_;
  assign new_n1828_ = ~new_n1821_ & ~new_n1827_;
  assign new_n1829_ = ~new_n1818_ & new_n1828_;
  assign new_n1830_ = new_n1818_ & ~new_n1828_;
  assign new_n1831_ = ~new_n1829_ & ~new_n1830_;
  assign new_n1832_ = B6734 & ~B6733;
  assign new_n1833_ = ~B6734 & B6733;
  assign new_n1834_ = ~new_n1832_ & ~new_n1833_;
  assign new_n1835_ = ~B6736 & new_n1834_;
  assign new_n1836_ = ~B6737 & ~B6736;
  assign new_n1837_ = ~new_n1835_ & ~new_n1836_;
  assign new_n1838_ = B6735 & new_n1837_;
  assign new_n1839_ = ~B6735 & ~new_n1837_;
  assign new_n1840_ = ~new_n1838_ & ~new_n1839_;
  assign new_n1841_ = ~new_n1834_ & ~new_n1840_;
  assign new_n1842_ = B6767 & ~B6766;
  assign new_n1843_ = ~B6767 & B6766;
  assign new_n1844_ = ~new_n1842_ & ~new_n1843_;
  assign new_n1845_ = ~B6769 & new_n1844_;
  assign new_n1846_ = ~B6770 & ~B6769;
  assign new_n1847_ = ~new_n1845_ & ~new_n1846_;
  assign new_n1848_ = B6768 & new_n1847_;
  assign new_n1849_ = ~B6768 & ~new_n1847_;
  assign new_n1850_ = ~new_n1848_ & ~new_n1849_;
  assign new_n1851_ = ~new_n1844_ & ~new_n1850_;
  assign new_n1852_ = new_n1831_ & ~new_n1851_;
  assign new_n1853_ = B6800 & ~B6799;
  assign new_n1854_ = ~B6800 & B6799;
  assign new_n1855_ = ~new_n1853_ & ~new_n1854_;
  assign new_n1856_ = ~B6802 & new_n1855_;
  assign new_n1857_ = ~B6803 & ~B6802;
  assign new_n1858_ = ~new_n1856_ & ~new_n1857_;
  assign new_n1859_ = B6801 & new_n1858_;
  assign new_n1860_ = ~B6801 & ~new_n1858_;
  assign new_n1861_ = ~new_n1859_ & ~new_n1860_;
  assign new_n1862_ = ~new_n1855_ & ~new_n1861_;
  assign new_n1863_ = ~new_n1851_ & ~new_n1862_;
  assign new_n1864_ = ~new_n1852_ & ~new_n1863_;
  assign new_n1865_ = new_n1841_ & new_n1864_;
  assign new_n1866_ = ~new_n1841_ & ~new_n1864_;
  assign new_n1867_ = ~new_n1865_ & ~new_n1866_;
  assign new_n1868_ = ~new_n1831_ & ~new_n1867_;
  assign new_n1869_ = ~new_n1807_ & ~new_n1868_;
  assign new_n1870_ = ~new_n1808_ & ~new_n1869_;
  assign new_n1871_ = new_n1747_ & new_n1870_;
  assign new_n1872_ = ~new_n1747_ & ~new_n1870_;
  assign new_n1873_ = ~new_n1871_ & ~new_n1872_;
  assign new_n1874_ = ~new_n1687_ & ~new_n1873_;
  assign new_n1875_ = ~new_n1564_ & new_n1874_;
  assign new_n1876_ = new_n1564_ & ~new_n1874_;
  assign new_n1877_ = ~new_n1875_ & ~new_n1876_;
  assign new_n1878_ = B6833 & ~B6832;
  assign new_n1879_ = ~B6833 & B6832;
  assign new_n1880_ = ~new_n1878_ & ~new_n1879_;
  assign new_n1881_ = ~B6835 & new_n1880_;
  assign new_n1882_ = ~B6836 & ~B6835;
  assign new_n1883_ = ~new_n1881_ & ~new_n1882_;
  assign new_n1884_ = B6834 & new_n1883_;
  assign new_n1885_ = ~B6834 & ~new_n1883_;
  assign new_n1886_ = ~new_n1884_ & ~new_n1885_;
  assign new_n1887_ = ~new_n1880_ & ~new_n1886_;
  assign new_n1888_ = B6866 & ~B6865;
  assign new_n1889_ = ~B6866 & B6865;
  assign new_n1890_ = ~new_n1888_ & ~new_n1889_;
  assign new_n1891_ = ~B6868 & new_n1890_;
  assign new_n1892_ = ~B6869 & ~B6868;
  assign new_n1893_ = ~new_n1891_ & ~new_n1892_;
  assign new_n1894_ = B6867 & new_n1893_;
  assign new_n1895_ = ~B6867 & ~new_n1893_;
  assign new_n1896_ = ~new_n1894_ & ~new_n1895_;
  assign new_n1897_ = ~new_n1890_ & ~new_n1896_;
  assign new_n1898_ = ~new_n1887_ & new_n1897_;
  assign new_n1899_ = new_n1887_ & ~new_n1897_;
  assign new_n1900_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1901_ = B6899 & ~B6898;
  assign new_n1902_ = ~B6899 & B6898;
  assign new_n1903_ = ~new_n1901_ & ~new_n1902_;
  assign new_n1904_ = ~B6901 & new_n1903_;
  assign new_n1905_ = ~B6902 & ~B6901;
  assign new_n1906_ = ~new_n1904_ & ~new_n1905_;
  assign new_n1907_ = B6900 & new_n1906_;
  assign new_n1908_ = ~B6900 & ~new_n1906_;
  assign new_n1909_ = ~new_n1907_ & ~new_n1908_;
  assign new_n1910_ = ~new_n1903_ & ~new_n1909_;
  assign new_n1911_ = B6932 & ~B6931;
  assign new_n1912_ = ~B6932 & B6931;
  assign new_n1913_ = ~new_n1911_ & ~new_n1912_;
  assign new_n1914_ = ~B6934 & new_n1913_;
  assign new_n1915_ = ~B6935 & ~B6934;
  assign new_n1916_ = ~new_n1914_ & ~new_n1915_;
  assign new_n1917_ = B6933 & new_n1916_;
  assign new_n1918_ = ~B6933 & ~new_n1916_;
  assign new_n1919_ = ~new_n1917_ & ~new_n1918_;
  assign new_n1920_ = ~new_n1913_ & ~new_n1919_;
  assign new_n1921_ = new_n1900_ & ~new_n1920_;
  assign new_n1922_ = B6965 & ~B6964;
  assign new_n1923_ = ~B6965 & B6964;
  assign new_n1924_ = ~new_n1922_ & ~new_n1923_;
  assign new_n1925_ = ~B6967 & new_n1924_;
  assign new_n1926_ = ~B6968 & ~B6967;
  assign new_n1927_ = ~new_n1925_ & ~new_n1926_;
  assign new_n1928_ = B6966 & new_n1927_;
  assign new_n1929_ = ~B6966 & ~new_n1927_;
  assign new_n1930_ = ~new_n1928_ & ~new_n1929_;
  assign new_n1931_ = ~new_n1924_ & ~new_n1930_;
  assign new_n1932_ = ~new_n1920_ & ~new_n1931_;
  assign new_n1933_ = ~new_n1921_ & ~new_n1932_;
  assign new_n1934_ = new_n1910_ & new_n1933_;
  assign new_n1935_ = ~new_n1910_ & ~new_n1933_;
  assign new_n1936_ = ~new_n1934_ & ~new_n1935_;
  assign new_n1937_ = ~new_n1900_ & ~new_n1936_;
  assign new_n1938_ = B6998 & ~B6997;
  assign new_n1939_ = ~B6998 & B6997;
  assign new_n1940_ = ~new_n1938_ & ~new_n1939_;
  assign new_n1941_ = ~B7000 & new_n1940_;
  assign new_n1942_ = ~B7001 & ~B7000;
  assign new_n1943_ = ~new_n1941_ & ~new_n1942_;
  assign new_n1944_ = B6999 & new_n1943_;
  assign new_n1945_ = ~B6999 & ~new_n1943_;
  assign new_n1946_ = ~new_n1944_ & ~new_n1945_;
  assign new_n1947_ = ~new_n1940_ & ~new_n1946_;
  assign new_n1948_ = B7031 & ~B7030;
  assign new_n1949_ = ~B7031 & B7030;
  assign new_n1950_ = ~new_n1948_ & ~new_n1949_;
  assign new_n1951_ = ~B7033 & new_n1950_;
  assign new_n1952_ = ~B7034 & ~B7033;
  assign new_n1953_ = ~new_n1951_ & ~new_n1952_;
  assign new_n1954_ = B7032 & new_n1953_;
  assign new_n1955_ = ~B7032 & ~new_n1953_;
  assign new_n1956_ = ~new_n1954_ & ~new_n1955_;
  assign new_n1957_ = ~new_n1950_ & ~new_n1956_;
  assign new_n1958_ = ~new_n1947_ & new_n1957_;
  assign new_n1959_ = new_n1947_ & ~new_n1957_;
  assign new_n1960_ = ~new_n1958_ & ~new_n1959_;
  assign new_n1961_ = B7064 & ~B7063;
  assign new_n1962_ = ~B7064 & B7063;
  assign new_n1963_ = ~new_n1961_ & ~new_n1962_;
  assign new_n1964_ = ~B7066 & new_n1963_;
  assign new_n1965_ = ~B7067 & ~B7066;
  assign new_n1966_ = ~new_n1964_ & ~new_n1965_;
  assign new_n1967_ = B7065 & new_n1966_;
  assign new_n1968_ = ~B7065 & ~new_n1966_;
  assign new_n1969_ = ~new_n1967_ & ~new_n1968_;
  assign new_n1970_ = ~new_n1963_ & ~new_n1969_;
  assign new_n1971_ = B7097 & ~B7096;
  assign new_n1972_ = ~B7097 & B7096;
  assign new_n1973_ = ~new_n1971_ & ~new_n1972_;
  assign new_n1974_ = ~B7099 & new_n1973_;
  assign new_n1975_ = ~B7100 & ~B7099;
  assign new_n1976_ = ~new_n1974_ & ~new_n1975_;
  assign new_n1977_ = B7098 & new_n1976_;
  assign new_n1978_ = ~B7098 & ~new_n1976_;
  assign new_n1979_ = ~new_n1977_ & ~new_n1978_;
  assign new_n1980_ = ~new_n1973_ & ~new_n1979_;
  assign new_n1981_ = new_n1960_ & ~new_n1980_;
  assign new_n1982_ = B7130 & ~B7129;
  assign new_n1983_ = ~B7130 & B7129;
  assign new_n1984_ = ~new_n1982_ & ~new_n1983_;
  assign new_n1985_ = ~B7132 & new_n1984_;
  assign new_n1986_ = ~B7133 & ~B7132;
  assign new_n1987_ = ~new_n1985_ & ~new_n1986_;
  assign new_n1988_ = B7131 & new_n1987_;
  assign new_n1989_ = ~B7131 & ~new_n1987_;
  assign new_n1990_ = ~new_n1988_ & ~new_n1989_;
  assign new_n1991_ = ~new_n1984_ & ~new_n1990_;
  assign new_n1992_ = ~new_n1980_ & ~new_n1991_;
  assign new_n1993_ = ~new_n1981_ & ~new_n1992_;
  assign new_n1994_ = new_n1970_ & new_n1993_;
  assign new_n1995_ = ~new_n1970_ & ~new_n1993_;
  assign new_n1996_ = ~new_n1994_ & ~new_n1995_;
  assign new_n1997_ = ~new_n1960_ & ~new_n1996_;
  assign new_n1998_ = ~new_n1937_ & new_n1997_;
  assign new_n1999_ = new_n1937_ & ~new_n1997_;
  assign new_n2000_ = ~new_n1998_ & ~new_n1999_;
  assign new_n2001_ = B7163 & ~B7162;
  assign new_n2002_ = ~B7163 & B7162;
  assign new_n2003_ = ~new_n2001_ & ~new_n2002_;
  assign new_n2004_ = ~B7165 & new_n2003_;
  assign new_n2005_ = ~B7166 & ~B7165;
  assign new_n2006_ = ~new_n2004_ & ~new_n2005_;
  assign new_n2007_ = B7164 & new_n2006_;
  assign new_n2008_ = ~B7164 & ~new_n2006_;
  assign new_n2009_ = ~new_n2007_ & ~new_n2008_;
  assign new_n2010_ = ~new_n2003_ & ~new_n2009_;
  assign new_n2011_ = B7196 & ~B7195;
  assign new_n2012_ = ~B7196 & B7195;
  assign new_n2013_ = ~new_n2011_ & ~new_n2012_;
  assign new_n2014_ = ~B7198 & new_n2013_;
  assign new_n2015_ = ~B7199 & ~B7198;
  assign new_n2016_ = ~new_n2014_ & ~new_n2015_;
  assign new_n2017_ = B7197 & new_n2016_;
  assign new_n2018_ = ~B7197 & ~new_n2016_;
  assign new_n2019_ = ~new_n2017_ & ~new_n2018_;
  assign new_n2020_ = ~new_n2013_ & ~new_n2019_;
  assign new_n2021_ = ~new_n2010_ & new_n2020_;
  assign new_n2022_ = new_n2010_ & ~new_n2020_;
  assign new_n2023_ = ~new_n2021_ & ~new_n2022_;
  assign new_n2024_ = B7229 & ~B7228;
  assign new_n2025_ = ~B7229 & B7228;
  assign new_n2026_ = ~new_n2024_ & ~new_n2025_;
  assign new_n2027_ = ~B7231 & new_n2026_;
  assign new_n2028_ = ~B7232 & ~B7231;
  assign new_n2029_ = ~new_n2027_ & ~new_n2028_;
  assign new_n2030_ = B7230 & new_n2029_;
  assign new_n2031_ = ~B7230 & ~new_n2029_;
  assign new_n2032_ = ~new_n2030_ & ~new_n2031_;
  assign new_n2033_ = ~new_n2026_ & ~new_n2032_;
  assign new_n2034_ = B7262 & ~B7261;
  assign new_n2035_ = ~B7262 & B7261;
  assign new_n2036_ = ~new_n2034_ & ~new_n2035_;
  assign new_n2037_ = ~B7264 & new_n2036_;
  assign new_n2038_ = ~B7265 & ~B7264;
  assign new_n2039_ = ~new_n2037_ & ~new_n2038_;
  assign new_n2040_ = B7263 & new_n2039_;
  assign new_n2041_ = ~B7263 & ~new_n2039_;
  assign new_n2042_ = ~new_n2040_ & ~new_n2041_;
  assign new_n2043_ = ~new_n2036_ & ~new_n2042_;
  assign new_n2044_ = new_n2023_ & ~new_n2043_;
  assign new_n2045_ = B7295 & ~B7294;
  assign new_n2046_ = ~B7295 & B7294;
  assign new_n2047_ = ~new_n2045_ & ~new_n2046_;
  assign new_n2048_ = ~B7297 & new_n2047_;
  assign new_n2049_ = ~B7298 & ~B7297;
  assign new_n2050_ = ~new_n2048_ & ~new_n2049_;
  assign new_n2051_ = B7296 & new_n2050_;
  assign new_n2052_ = ~B7296 & ~new_n2050_;
  assign new_n2053_ = ~new_n2051_ & ~new_n2052_;
  assign new_n2054_ = ~new_n2047_ & ~new_n2053_;
  assign new_n2055_ = ~new_n2043_ & ~new_n2054_;
  assign new_n2056_ = ~new_n2044_ & ~new_n2055_;
  assign new_n2057_ = new_n2033_ & new_n2056_;
  assign new_n2058_ = ~new_n2033_ & ~new_n2056_;
  assign new_n2059_ = ~new_n2057_ & ~new_n2058_;
  assign new_n2060_ = ~new_n2023_ & ~new_n2059_;
  assign new_n2061_ = B7328 & ~B7327;
  assign new_n2062_ = ~B7328 & B7327;
  assign new_n2063_ = ~new_n2061_ & ~new_n2062_;
  assign new_n2064_ = ~B7330 & new_n2063_;
  assign new_n2065_ = ~B7331 & ~B7330;
  assign new_n2066_ = ~new_n2064_ & ~new_n2065_;
  assign new_n2067_ = B7329 & new_n2066_;
  assign new_n2068_ = ~B7329 & ~new_n2066_;
  assign new_n2069_ = ~new_n2067_ & ~new_n2068_;
  assign new_n2070_ = ~new_n2063_ & ~new_n2069_;
  assign new_n2071_ = B7361 & ~B7360;
  assign new_n2072_ = ~B7361 & B7360;
  assign new_n2073_ = ~new_n2071_ & ~new_n2072_;
  assign new_n2074_ = ~B7363 & new_n2073_;
  assign new_n2075_ = ~B7364 & ~B7363;
  assign new_n2076_ = ~new_n2074_ & ~new_n2075_;
  assign new_n2077_ = B7362 & new_n2076_;
  assign new_n2078_ = ~B7362 & ~new_n2076_;
  assign new_n2079_ = ~new_n2077_ & ~new_n2078_;
  assign new_n2080_ = ~new_n2073_ & ~new_n2079_;
  assign new_n2081_ = ~new_n2070_ & new_n2080_;
  assign new_n2082_ = new_n2070_ & ~new_n2080_;
  assign new_n2083_ = ~new_n2081_ & ~new_n2082_;
  assign new_n2084_ = B7394 & ~B7393;
  assign new_n2085_ = ~B7394 & B7393;
  assign new_n2086_ = ~new_n2084_ & ~new_n2085_;
  assign new_n2087_ = ~B7396 & new_n2086_;
  assign new_n2088_ = ~B7397 & ~B7396;
  assign new_n2089_ = ~new_n2087_ & ~new_n2088_;
  assign new_n2090_ = B7395 & new_n2089_;
  assign new_n2091_ = ~B7395 & ~new_n2089_;
  assign new_n2092_ = ~new_n2090_ & ~new_n2091_;
  assign new_n2093_ = ~new_n2086_ & ~new_n2092_;
  assign new_n2094_ = B7427 & ~B7426;
  assign new_n2095_ = ~B7427 & B7426;
  assign new_n2096_ = ~new_n2094_ & ~new_n2095_;
  assign new_n2097_ = ~B7429 & new_n2096_;
  assign new_n2098_ = ~B7430 & ~B7429;
  assign new_n2099_ = ~new_n2097_ & ~new_n2098_;
  assign new_n2100_ = B7428 & new_n2099_;
  assign new_n2101_ = ~B7428 & ~new_n2099_;
  assign new_n2102_ = ~new_n2100_ & ~new_n2101_;
  assign new_n2103_ = ~new_n2096_ & ~new_n2102_;
  assign new_n2104_ = new_n2083_ & ~new_n2103_;
  assign new_n2105_ = B7460 & ~B7459;
  assign new_n2106_ = ~B7460 & B7459;
  assign new_n2107_ = ~new_n2105_ & ~new_n2106_;
  assign new_n2108_ = ~B7462 & new_n2107_;
  assign new_n2109_ = ~B7463 & ~B7462;
  assign new_n2110_ = ~new_n2108_ & ~new_n2109_;
  assign new_n2111_ = B7461 & new_n2110_;
  assign new_n2112_ = ~B7461 & ~new_n2110_;
  assign new_n2113_ = ~new_n2111_ & ~new_n2112_;
  assign new_n2114_ = ~new_n2107_ & ~new_n2113_;
  assign new_n2115_ = ~new_n2103_ & ~new_n2114_;
  assign new_n2116_ = ~new_n2104_ & ~new_n2115_;
  assign new_n2117_ = new_n2093_ & new_n2116_;
  assign new_n2118_ = ~new_n2093_ & ~new_n2116_;
  assign new_n2119_ = ~new_n2117_ & ~new_n2118_;
  assign new_n2120_ = ~new_n2083_ & ~new_n2119_;
  assign new_n2121_ = new_n2000_ & ~new_n2120_;
  assign new_n2122_ = B7493 & ~B7492;
  assign new_n2123_ = ~B7493 & B7492;
  assign new_n2124_ = ~new_n2122_ & ~new_n2123_;
  assign new_n2125_ = ~B7495 & new_n2124_;
  assign new_n2126_ = ~B7496 & ~B7495;
  assign new_n2127_ = ~new_n2125_ & ~new_n2126_;
  assign new_n2128_ = B7494 & new_n2127_;
  assign new_n2129_ = ~B7494 & ~new_n2127_;
  assign new_n2130_ = ~new_n2128_ & ~new_n2129_;
  assign new_n2131_ = ~new_n2124_ & ~new_n2130_;
  assign new_n2132_ = B7526 & ~B7525;
  assign new_n2133_ = ~B7526 & B7525;
  assign new_n2134_ = ~new_n2132_ & ~new_n2133_;
  assign new_n2135_ = ~B7528 & new_n2134_;
  assign new_n2136_ = ~B7529 & ~B7528;
  assign new_n2137_ = ~new_n2135_ & ~new_n2136_;
  assign new_n2138_ = B7527 & new_n2137_;
  assign new_n2139_ = ~B7527 & ~new_n2137_;
  assign new_n2140_ = ~new_n2138_ & ~new_n2139_;
  assign new_n2141_ = ~new_n2134_ & ~new_n2140_;
  assign new_n2142_ = ~new_n2131_ & new_n2141_;
  assign new_n2143_ = new_n2131_ & ~new_n2141_;
  assign new_n2144_ = ~new_n2142_ & ~new_n2143_;
  assign new_n2145_ = B7559 & ~B7558;
  assign new_n2146_ = ~B7559 & B7558;
  assign new_n2147_ = ~new_n2145_ & ~new_n2146_;
  assign new_n2148_ = ~B7561 & new_n2147_;
  assign new_n2149_ = ~B7562 & ~B7561;
  assign new_n2150_ = ~new_n2148_ & ~new_n2149_;
  assign new_n2151_ = B7560 & new_n2150_;
  assign new_n2152_ = ~B7560 & ~new_n2150_;
  assign new_n2153_ = ~new_n2151_ & ~new_n2152_;
  assign new_n2154_ = ~new_n2147_ & ~new_n2153_;
  assign new_n2155_ = B7592 & ~B7591;
  assign new_n2156_ = ~B7592 & B7591;
  assign new_n2157_ = ~new_n2155_ & ~new_n2156_;
  assign new_n2158_ = ~B7594 & new_n2157_;
  assign new_n2159_ = ~B7595 & ~B7594;
  assign new_n2160_ = ~new_n2158_ & ~new_n2159_;
  assign new_n2161_ = B7593 & new_n2160_;
  assign new_n2162_ = ~B7593 & ~new_n2160_;
  assign new_n2163_ = ~new_n2161_ & ~new_n2162_;
  assign new_n2164_ = ~new_n2157_ & ~new_n2163_;
  assign new_n2165_ = new_n2144_ & ~new_n2164_;
  assign new_n2166_ = B7625 & ~B7624;
  assign new_n2167_ = ~B7625 & B7624;
  assign new_n2168_ = ~new_n2166_ & ~new_n2167_;
  assign new_n2169_ = ~B7627 & new_n2168_;
  assign new_n2170_ = ~B7628 & ~B7627;
  assign new_n2171_ = ~new_n2169_ & ~new_n2170_;
  assign new_n2172_ = B7626 & new_n2171_;
  assign new_n2173_ = ~B7626 & ~new_n2171_;
  assign new_n2174_ = ~new_n2172_ & ~new_n2173_;
  assign new_n2175_ = ~new_n2168_ & ~new_n2174_;
  assign new_n2176_ = ~new_n2164_ & ~new_n2175_;
  assign new_n2177_ = ~new_n2165_ & ~new_n2176_;
  assign new_n2178_ = new_n2154_ & new_n2177_;
  assign new_n2179_ = ~new_n2154_ & ~new_n2177_;
  assign new_n2180_ = ~new_n2178_ & ~new_n2179_;
  assign new_n2181_ = ~new_n2144_ & ~new_n2180_;
  assign new_n2182_ = ~new_n2120_ & ~new_n2181_;
  assign new_n2183_ = ~new_n2121_ & ~new_n2182_;
  assign new_n2184_ = new_n2060_ & new_n2183_;
  assign new_n2185_ = ~new_n2060_ & ~new_n2183_;
  assign new_n2186_ = ~new_n2184_ & ~new_n2185_;
  assign new_n2187_ = ~new_n2000_ & ~new_n2186_;
  assign new_n2188_ = B7658 & ~B7657;
  assign new_n2189_ = ~B7658 & B7657;
  assign new_n2190_ = ~new_n2188_ & ~new_n2189_;
  assign new_n2191_ = ~B7660 & new_n2190_;
  assign new_n2192_ = ~B7661 & ~B7660;
  assign new_n2193_ = ~new_n2191_ & ~new_n2192_;
  assign new_n2194_ = B7659 & new_n2193_;
  assign new_n2195_ = ~B7659 & ~new_n2193_;
  assign new_n2196_ = ~new_n2194_ & ~new_n2195_;
  assign new_n2197_ = ~new_n2190_ & ~new_n2196_;
  assign new_n2198_ = B7691 & ~B7690;
  assign new_n2199_ = ~B7691 & B7690;
  assign new_n2200_ = ~new_n2198_ & ~new_n2199_;
  assign new_n2201_ = ~B7693 & new_n2200_;
  assign new_n2202_ = ~B7694 & ~B7693;
  assign new_n2203_ = ~new_n2201_ & ~new_n2202_;
  assign new_n2204_ = B7692 & new_n2203_;
  assign new_n2205_ = ~B7692 & ~new_n2203_;
  assign new_n2206_ = ~new_n2204_ & ~new_n2205_;
  assign new_n2207_ = ~new_n2200_ & ~new_n2206_;
  assign new_n2208_ = ~new_n2197_ & new_n2207_;
  assign new_n2209_ = new_n2197_ & ~new_n2207_;
  assign new_n2210_ = ~new_n2208_ & ~new_n2209_;
  assign new_n2211_ = B7724 & ~B7723;
  assign new_n2212_ = ~B7724 & B7723;
  assign new_n2213_ = ~new_n2211_ & ~new_n2212_;
  assign new_n2214_ = ~B7726 & new_n2213_;
  assign new_n2215_ = ~B7727 & ~B7726;
  assign new_n2216_ = ~new_n2214_ & ~new_n2215_;
  assign new_n2217_ = B7725 & new_n2216_;
  assign new_n2218_ = ~B7725 & ~new_n2216_;
  assign new_n2219_ = ~new_n2217_ & ~new_n2218_;
  assign new_n2220_ = ~new_n2213_ & ~new_n2219_;
  assign new_n2221_ = B7757 & ~B7756;
  assign new_n2222_ = ~B7757 & B7756;
  assign new_n2223_ = ~new_n2221_ & ~new_n2222_;
  assign new_n2224_ = ~B7759 & new_n2223_;
  assign new_n2225_ = ~B7760 & ~B7759;
  assign new_n2226_ = ~new_n2224_ & ~new_n2225_;
  assign new_n2227_ = B7758 & new_n2226_;
  assign new_n2228_ = ~B7758 & ~new_n2226_;
  assign new_n2229_ = ~new_n2227_ & ~new_n2228_;
  assign new_n2230_ = ~new_n2223_ & ~new_n2229_;
  assign new_n2231_ = new_n2210_ & ~new_n2230_;
  assign new_n2232_ = B7790 & ~B7789;
  assign new_n2233_ = ~B7790 & B7789;
  assign new_n2234_ = ~new_n2232_ & ~new_n2233_;
  assign new_n2235_ = ~B7792 & new_n2234_;
  assign new_n2236_ = ~B7793 & ~B7792;
  assign new_n2237_ = ~new_n2235_ & ~new_n2236_;
  assign new_n2238_ = B7791 & new_n2237_;
  assign new_n2239_ = ~B7791 & ~new_n2237_;
  assign new_n2240_ = ~new_n2238_ & ~new_n2239_;
  assign new_n2241_ = ~new_n2234_ & ~new_n2240_;
  assign new_n2242_ = ~new_n2230_ & ~new_n2241_;
  assign new_n2243_ = ~new_n2231_ & ~new_n2242_;
  assign new_n2244_ = new_n2220_ & new_n2243_;
  assign new_n2245_ = ~new_n2220_ & ~new_n2243_;
  assign new_n2246_ = ~new_n2244_ & ~new_n2245_;
  assign new_n2247_ = ~new_n2210_ & ~new_n2246_;
  assign new_n2248_ = B7823 & ~B7822;
  assign new_n2249_ = ~B7823 & B7822;
  assign new_n2250_ = ~new_n2248_ & ~new_n2249_;
  assign new_n2251_ = ~B7825 & new_n2250_;
  assign new_n2252_ = ~B7826 & ~B7825;
  assign new_n2253_ = ~new_n2251_ & ~new_n2252_;
  assign new_n2254_ = B7824 & new_n2253_;
  assign new_n2255_ = ~B7824 & ~new_n2253_;
  assign new_n2256_ = ~new_n2254_ & ~new_n2255_;
  assign new_n2257_ = ~new_n2250_ & ~new_n2256_;
  assign new_n2258_ = B7856 & ~B7855;
  assign new_n2259_ = ~B7856 & B7855;
  assign new_n2260_ = ~new_n2258_ & ~new_n2259_;
  assign new_n2261_ = ~B7858 & new_n2260_;
  assign new_n2262_ = ~B7859 & ~B7858;
  assign new_n2263_ = ~new_n2261_ & ~new_n2262_;
  assign new_n2264_ = B7857 & new_n2263_;
  assign new_n2265_ = ~B7857 & ~new_n2263_;
  assign new_n2266_ = ~new_n2264_ & ~new_n2265_;
  assign new_n2267_ = ~new_n2260_ & ~new_n2266_;
  assign new_n2268_ = ~new_n2257_ & new_n2267_;
  assign new_n2269_ = new_n2257_ & ~new_n2267_;
  assign new_n2270_ = ~new_n2268_ & ~new_n2269_;
  assign new_n2271_ = B7889 & ~B7888;
  assign new_n2272_ = ~B7889 & B7888;
  assign new_n2273_ = ~new_n2271_ & ~new_n2272_;
  assign new_n2274_ = ~B7891 & new_n2273_;
  assign new_n2275_ = ~B7892 & ~B7891;
  assign new_n2276_ = ~new_n2274_ & ~new_n2275_;
  assign new_n2277_ = B7890 & new_n2276_;
  assign new_n2278_ = ~B7890 & ~new_n2276_;
  assign new_n2279_ = ~new_n2277_ & ~new_n2278_;
  assign new_n2280_ = ~new_n2273_ & ~new_n2279_;
  assign new_n2281_ = B7922 & ~B7921;
  assign new_n2282_ = ~B7922 & B7921;
  assign new_n2283_ = ~new_n2281_ & ~new_n2282_;
  assign new_n2284_ = ~B7924 & new_n2283_;
  assign new_n2285_ = ~B7925 & ~B7924;
  assign new_n2286_ = ~new_n2284_ & ~new_n2285_;
  assign new_n2287_ = B7923 & new_n2286_;
  assign new_n2288_ = ~B7923 & ~new_n2286_;
  assign new_n2289_ = ~new_n2287_ & ~new_n2288_;
  assign new_n2290_ = ~new_n2283_ & ~new_n2289_;
  assign new_n2291_ = new_n2270_ & ~new_n2290_;
  assign new_n2292_ = B7955 & ~B7954;
  assign new_n2293_ = ~B7955 & B7954;
  assign new_n2294_ = ~new_n2292_ & ~new_n2293_;
  assign new_n2295_ = ~B7957 & new_n2294_;
  assign new_n2296_ = ~B7958 & ~B7957;
  assign new_n2297_ = ~new_n2295_ & ~new_n2296_;
  assign new_n2298_ = B7956 & new_n2297_;
  assign new_n2299_ = ~B7956 & ~new_n2297_;
  assign new_n2300_ = ~new_n2298_ & ~new_n2299_;
  assign new_n2301_ = ~new_n2294_ & ~new_n2300_;
  assign new_n2302_ = ~new_n2290_ & ~new_n2301_;
  assign new_n2303_ = ~new_n2291_ & ~new_n2302_;
  assign new_n2304_ = new_n2280_ & new_n2303_;
  assign new_n2305_ = ~new_n2280_ & ~new_n2303_;
  assign new_n2306_ = ~new_n2304_ & ~new_n2305_;
  assign new_n2307_ = ~new_n2270_ & ~new_n2306_;
  assign new_n2308_ = ~new_n2247_ & new_n2307_;
  assign new_n2309_ = new_n2247_ & ~new_n2307_;
  assign new_n2310_ = ~new_n2308_ & ~new_n2309_;
  assign new_n2311_ = B7988 & ~B7987;
  assign new_n2312_ = ~B7988 & B7987;
  assign new_n2313_ = ~new_n2311_ & ~new_n2312_;
  assign new_n2314_ = ~B7990 & new_n2313_;
  assign new_n2315_ = ~B7991 & ~B7990;
  assign new_n2316_ = ~new_n2314_ & ~new_n2315_;
  assign new_n2317_ = B7989 & new_n2316_;
  assign new_n2318_ = ~B7989 & ~new_n2316_;
  assign new_n2319_ = ~new_n2317_ & ~new_n2318_;
  assign new_n2320_ = ~new_n2313_ & ~new_n2319_;
  assign new_n2321_ = B8021 & ~B8020;
  assign new_n2322_ = ~B8021 & B8020;
  assign new_n2323_ = ~new_n2321_ & ~new_n2322_;
  assign new_n2324_ = ~B8023 & new_n2323_;
  assign new_n2325_ = ~B8024 & ~B8023;
  assign new_n2326_ = ~new_n2324_ & ~new_n2325_;
  assign new_n2327_ = B8022 & new_n2326_;
  assign new_n2328_ = ~B8022 & ~new_n2326_;
  assign new_n2329_ = ~new_n2327_ & ~new_n2328_;
  assign new_n2330_ = ~new_n2323_ & ~new_n2329_;
  assign new_n2331_ = ~new_n2320_ & new_n2330_;
  assign new_n2332_ = new_n2320_ & ~new_n2330_;
  assign new_n2333_ = ~new_n2331_ & ~new_n2332_;
  assign new_n2334_ = B8054 & ~B8053;
  assign new_n2335_ = ~B8054 & B8053;
  assign new_n2336_ = ~new_n2334_ & ~new_n2335_;
  assign new_n2337_ = ~B8056 & new_n2336_;
  assign new_n2338_ = ~B8057 & ~B8056;
  assign new_n2339_ = ~new_n2337_ & ~new_n2338_;
  assign new_n2340_ = B8055 & new_n2339_;
  assign new_n2341_ = ~B8055 & ~new_n2339_;
  assign new_n2342_ = ~new_n2340_ & ~new_n2341_;
  assign new_n2343_ = ~new_n2336_ & ~new_n2342_;
  assign new_n2344_ = B8087 & ~B8086;
  assign new_n2345_ = ~B8087 & B8086;
  assign new_n2346_ = ~new_n2344_ & ~new_n2345_;
  assign new_n2347_ = ~B8089 & new_n2346_;
  assign new_n2348_ = ~B8090 & ~B8089;
  assign new_n2349_ = ~new_n2347_ & ~new_n2348_;
  assign new_n2350_ = B8088 & new_n2349_;
  assign new_n2351_ = ~B8088 & ~new_n2349_;
  assign new_n2352_ = ~new_n2350_ & ~new_n2351_;
  assign new_n2353_ = ~new_n2346_ & ~new_n2352_;
  assign new_n2354_ = new_n2333_ & ~new_n2353_;
  assign new_n2355_ = B8120 & ~B8119;
  assign new_n2356_ = ~B8120 & B8119;
  assign new_n2357_ = ~new_n2355_ & ~new_n2356_;
  assign new_n2358_ = ~B8122 & new_n2357_;
  assign new_n2359_ = ~B8123 & ~B8122;
  assign new_n2360_ = ~new_n2358_ & ~new_n2359_;
  assign new_n2361_ = B8121 & new_n2360_;
  assign new_n2362_ = ~B8121 & ~new_n2360_;
  assign new_n2363_ = ~new_n2361_ & ~new_n2362_;
  assign new_n2364_ = ~new_n2357_ & ~new_n2363_;
  assign new_n2365_ = ~new_n2353_ & ~new_n2364_;
  assign new_n2366_ = ~new_n2354_ & ~new_n2365_;
  assign new_n2367_ = new_n2343_ & new_n2366_;
  assign new_n2368_ = ~new_n2343_ & ~new_n2366_;
  assign new_n2369_ = ~new_n2367_ & ~new_n2368_;
  assign new_n2370_ = ~new_n2333_ & ~new_n2369_;
  assign new_n2371_ = B8153 & ~B8152;
  assign new_n2372_ = ~B8153 & B8152;
  assign new_n2373_ = ~new_n2371_ & ~new_n2372_;
  assign new_n2374_ = ~B8155 & new_n2373_;
  assign new_n2375_ = ~B8156 & ~B8155;
  assign new_n2376_ = ~new_n2374_ & ~new_n2375_;
  assign new_n2377_ = B8154 & new_n2376_;
  assign new_n2378_ = ~B8154 & ~new_n2376_;
  assign new_n2379_ = ~new_n2377_ & ~new_n2378_;
  assign new_n2380_ = ~new_n2373_ & ~new_n2379_;
  assign new_n2381_ = B8186 & ~B8185;
  assign new_n2382_ = ~B8186 & B8185;
  assign new_n2383_ = ~new_n2381_ & ~new_n2382_;
  assign new_n2384_ = ~B8188 & new_n2383_;
  assign new_n2385_ = ~B8189 & ~B8188;
  assign new_n2386_ = ~new_n2384_ & ~new_n2385_;
  assign new_n2387_ = B8187 & new_n2386_;
  assign new_n2388_ = ~B8187 & ~new_n2386_;
  assign new_n2389_ = ~new_n2387_ & ~new_n2388_;
  assign new_n2390_ = ~new_n2383_ & ~new_n2389_;
  assign new_n2391_ = ~new_n2380_ & new_n2390_;
  assign new_n2392_ = new_n2380_ & ~new_n2390_;
  assign new_n2393_ = ~new_n2391_ & ~new_n2392_;
  assign new_n2394_ = B8219 & ~B8218;
  assign new_n2395_ = ~B8219 & B8218;
  assign new_n2396_ = ~new_n2394_ & ~new_n2395_;
  assign new_n2397_ = ~B8221 & new_n2396_;
  assign new_n2398_ = ~B8222 & ~B8221;
  assign new_n2399_ = ~new_n2397_ & ~new_n2398_;
  assign new_n2400_ = B8220 & new_n2399_;
  assign new_n2401_ = ~B8220 & ~new_n2399_;
  assign new_n2402_ = ~new_n2400_ & ~new_n2401_;
  assign new_n2403_ = ~new_n2396_ & ~new_n2402_;
  assign new_n2404_ = B8252 & ~B8251;
  assign new_n2405_ = ~B8252 & B8251;
  assign new_n2406_ = ~new_n2404_ & ~new_n2405_;
  assign new_n2407_ = ~B8254 & new_n2406_;
  assign new_n2408_ = ~B8255 & ~B8254;
  assign new_n2409_ = ~new_n2407_ & ~new_n2408_;
  assign new_n2410_ = B8253 & new_n2409_;
  assign new_n2411_ = ~B8253 & ~new_n2409_;
  assign new_n2412_ = ~new_n2410_ & ~new_n2411_;
  assign new_n2413_ = ~new_n2406_ & ~new_n2412_;
  assign new_n2414_ = new_n2393_ & ~new_n2413_;
  assign new_n2415_ = B8285 & ~B8284;
  assign new_n2416_ = ~B8285 & B8284;
  assign new_n2417_ = ~new_n2415_ & ~new_n2416_;
  assign new_n2418_ = ~B8287 & new_n2417_;
  assign new_n2419_ = ~B8288 & ~B8287;
  assign new_n2420_ = ~new_n2418_ & ~new_n2419_;
  assign new_n2421_ = B8286 & new_n2420_;
  assign new_n2422_ = ~B8286 & ~new_n2420_;
  assign new_n2423_ = ~new_n2421_ & ~new_n2422_;
  assign new_n2424_ = ~new_n2417_ & ~new_n2423_;
  assign new_n2425_ = ~new_n2413_ & ~new_n2424_;
  assign new_n2426_ = ~new_n2414_ & ~new_n2425_;
  assign new_n2427_ = new_n2403_ & new_n2426_;
  assign new_n2428_ = ~new_n2403_ & ~new_n2426_;
  assign new_n2429_ = ~new_n2427_ & ~new_n2428_;
  assign new_n2430_ = ~new_n2393_ & ~new_n2429_;
  assign new_n2431_ = new_n2310_ & ~new_n2430_;
  assign new_n2432_ = B8318 & ~B8317;
  assign new_n2433_ = ~B8318 & B8317;
  assign new_n2434_ = ~new_n2432_ & ~new_n2433_;
  assign new_n2435_ = ~B8320 & new_n2434_;
  assign new_n2436_ = ~B8321 & ~B8320;
  assign new_n2437_ = ~new_n2435_ & ~new_n2436_;
  assign new_n2438_ = B8319 & new_n2437_;
  assign new_n2439_ = ~B8319 & ~new_n2437_;
  assign new_n2440_ = ~new_n2438_ & ~new_n2439_;
  assign new_n2441_ = ~new_n2434_ & ~new_n2440_;
  assign new_n2442_ = B8351 & ~B8350;
  assign new_n2443_ = ~B8351 & B8350;
  assign new_n2444_ = ~new_n2442_ & ~new_n2443_;
  assign new_n2445_ = ~B8353 & new_n2444_;
  assign new_n2446_ = ~B8354 & ~B8353;
  assign new_n2447_ = ~new_n2445_ & ~new_n2446_;
  assign new_n2448_ = B8352 & new_n2447_;
  assign new_n2449_ = ~B8352 & ~new_n2447_;
  assign new_n2450_ = ~new_n2448_ & ~new_n2449_;
  assign new_n2451_ = ~new_n2444_ & ~new_n2450_;
  assign new_n2452_ = ~new_n2441_ & new_n2451_;
  assign new_n2453_ = new_n2441_ & ~new_n2451_;
  assign new_n2454_ = ~new_n2452_ & ~new_n2453_;
  assign new_n2455_ = B8384 & ~B8383;
  assign new_n2456_ = ~B8384 & B8383;
  assign new_n2457_ = ~new_n2455_ & ~new_n2456_;
  assign new_n2458_ = ~B8386 & new_n2457_;
  assign new_n2459_ = ~B8387 & ~B8386;
  assign new_n2460_ = ~new_n2458_ & ~new_n2459_;
  assign new_n2461_ = B8385 & new_n2460_;
  assign new_n2462_ = ~B8385 & ~new_n2460_;
  assign new_n2463_ = ~new_n2461_ & ~new_n2462_;
  assign new_n2464_ = ~new_n2457_ & ~new_n2463_;
  assign new_n2465_ = B8417 & ~B8416;
  assign new_n2466_ = ~B8417 & B8416;
  assign new_n2467_ = ~new_n2465_ & ~new_n2466_;
  assign new_n2468_ = ~B8419 & new_n2467_;
  assign new_n2469_ = ~B8420 & ~B8419;
  assign new_n2470_ = ~new_n2468_ & ~new_n2469_;
  assign new_n2471_ = B8418 & new_n2470_;
  assign new_n2472_ = ~B8418 & ~new_n2470_;
  assign new_n2473_ = ~new_n2471_ & ~new_n2472_;
  assign new_n2474_ = ~new_n2467_ & ~new_n2473_;
  assign new_n2475_ = new_n2454_ & ~new_n2474_;
  assign new_n2476_ = B8450 & ~B8449;
  assign new_n2477_ = ~B8450 & B8449;
  assign new_n2478_ = ~new_n2476_ & ~new_n2477_;
  assign new_n2479_ = ~B8452 & new_n2478_;
  assign new_n2480_ = ~B8453 & ~B8452;
  assign new_n2481_ = ~new_n2479_ & ~new_n2480_;
  assign new_n2482_ = B8451 & new_n2481_;
  assign new_n2483_ = ~B8451 & ~new_n2481_;
  assign new_n2484_ = ~new_n2482_ & ~new_n2483_;
  assign new_n2485_ = ~new_n2478_ & ~new_n2484_;
  assign new_n2486_ = ~new_n2474_ & ~new_n2485_;
  assign new_n2487_ = ~new_n2475_ & ~new_n2486_;
  assign new_n2488_ = new_n2464_ & new_n2487_;
  assign new_n2489_ = ~new_n2464_ & ~new_n2487_;
  assign new_n2490_ = ~new_n2488_ & ~new_n2489_;
  assign new_n2491_ = ~new_n2454_ & ~new_n2490_;
  assign new_n2492_ = ~new_n2430_ & ~new_n2491_;
  assign new_n2493_ = ~new_n2431_ & ~new_n2492_;
  assign new_n2494_ = new_n2370_ & new_n2493_;
  assign new_n2495_ = ~new_n2370_ & ~new_n2493_;
  assign new_n2496_ = ~new_n2494_ & ~new_n2495_;
  assign new_n2497_ = ~new_n2310_ & ~new_n2496_;
  assign new_n2498_ = new_n1877_ & ~new_n2497_;
  assign new_n2499_ = B8483 & ~B8482;
  assign new_n2500_ = ~B8483 & B8482;
  assign new_n2501_ = ~new_n2499_ & ~new_n2500_;
  assign new_n2502_ = ~B8485 & new_n2501_;
  assign new_n2503_ = ~B8486 & ~B8485;
  assign new_n2504_ = ~new_n2502_ & ~new_n2503_;
  assign new_n2505_ = B8484 & new_n2504_;
  assign new_n2506_ = ~B8484 & ~new_n2504_;
  assign new_n2507_ = ~new_n2505_ & ~new_n2506_;
  assign new_n2508_ = ~new_n2501_ & ~new_n2507_;
  assign new_n2509_ = B8516 & ~B8515;
  assign new_n2510_ = ~B8516 & B8515;
  assign new_n2511_ = ~new_n2509_ & ~new_n2510_;
  assign new_n2512_ = ~B8518 & new_n2511_;
  assign new_n2513_ = ~B8519 & ~B8518;
  assign new_n2514_ = ~new_n2512_ & ~new_n2513_;
  assign new_n2515_ = B8517 & new_n2514_;
  assign new_n2516_ = ~B8517 & ~new_n2514_;
  assign new_n2517_ = ~new_n2515_ & ~new_n2516_;
  assign new_n2518_ = ~new_n2511_ & ~new_n2517_;
  assign new_n2519_ = ~new_n2508_ & new_n2518_;
  assign new_n2520_ = new_n2508_ & ~new_n2518_;
  assign new_n2521_ = ~new_n2519_ & ~new_n2520_;
  assign new_n2522_ = B8549 & ~B8548;
  assign new_n2523_ = ~B8549 & B8548;
  assign new_n2524_ = ~new_n2522_ & ~new_n2523_;
  assign new_n2525_ = ~B8551 & new_n2524_;
  assign new_n2526_ = ~B8552 & ~B8551;
  assign new_n2527_ = ~new_n2525_ & ~new_n2526_;
  assign new_n2528_ = B8550 & new_n2527_;
  assign new_n2529_ = ~B8550 & ~new_n2527_;
  assign new_n2530_ = ~new_n2528_ & ~new_n2529_;
  assign new_n2531_ = ~new_n2524_ & ~new_n2530_;
  assign new_n2532_ = B8582 & ~B8581;
  assign new_n2533_ = ~B8582 & B8581;
  assign new_n2534_ = ~new_n2532_ & ~new_n2533_;
  assign new_n2535_ = ~B8584 & new_n2534_;
  assign new_n2536_ = ~B8585 & ~B8584;
  assign new_n2537_ = ~new_n2535_ & ~new_n2536_;
  assign new_n2538_ = B8583 & new_n2537_;
  assign new_n2539_ = ~B8583 & ~new_n2537_;
  assign new_n2540_ = ~new_n2538_ & ~new_n2539_;
  assign new_n2541_ = ~new_n2534_ & ~new_n2540_;
  assign new_n2542_ = new_n2521_ & ~new_n2541_;
  assign new_n2543_ = B8615 & ~B8614;
  assign new_n2544_ = ~B8615 & B8614;
  assign new_n2545_ = ~new_n2543_ & ~new_n2544_;
  assign new_n2546_ = ~B8617 & new_n2545_;
  assign new_n2547_ = ~B8618 & ~B8617;
  assign new_n2548_ = ~new_n2546_ & ~new_n2547_;
  assign new_n2549_ = B8616 & new_n2548_;
  assign new_n2550_ = ~B8616 & ~new_n2548_;
  assign new_n2551_ = ~new_n2549_ & ~new_n2550_;
  assign new_n2552_ = ~new_n2545_ & ~new_n2551_;
  assign new_n2553_ = ~new_n2541_ & ~new_n2552_;
  assign new_n2554_ = ~new_n2542_ & ~new_n2553_;
  assign new_n2555_ = new_n2531_ & new_n2554_;
  assign new_n2556_ = ~new_n2531_ & ~new_n2554_;
  assign new_n2557_ = ~new_n2555_ & ~new_n2556_;
  assign new_n2558_ = ~new_n2521_ & ~new_n2557_;
  assign new_n2559_ = B8648 & ~B8647;
  assign new_n2560_ = ~B8648 & B8647;
  assign new_n2561_ = ~new_n2559_ & ~new_n2560_;
  assign new_n2562_ = ~B8650 & new_n2561_;
  assign new_n2563_ = ~B8651 & ~B8650;
  assign new_n2564_ = ~new_n2562_ & ~new_n2563_;
  assign new_n2565_ = B8649 & new_n2564_;
  assign new_n2566_ = ~B8649 & ~new_n2564_;
  assign new_n2567_ = ~new_n2565_ & ~new_n2566_;
  assign new_n2568_ = ~new_n2561_ & ~new_n2567_;
  assign new_n2569_ = B8681 & ~B8680;
  assign new_n2570_ = ~B8681 & B8680;
  assign new_n2571_ = ~new_n2569_ & ~new_n2570_;
  assign new_n2572_ = ~B8683 & new_n2571_;
  assign new_n2573_ = ~B8684 & ~B8683;
  assign new_n2574_ = ~new_n2572_ & ~new_n2573_;
  assign new_n2575_ = B8682 & new_n2574_;
  assign new_n2576_ = ~B8682 & ~new_n2574_;
  assign new_n2577_ = ~new_n2575_ & ~new_n2576_;
  assign new_n2578_ = ~new_n2571_ & ~new_n2577_;
  assign new_n2579_ = ~new_n2568_ & new_n2578_;
  assign new_n2580_ = new_n2568_ & ~new_n2578_;
  assign new_n2581_ = ~new_n2579_ & ~new_n2580_;
  assign new_n2582_ = B8714 & ~B8713;
  assign new_n2583_ = ~B8714 & B8713;
  assign new_n2584_ = ~new_n2582_ & ~new_n2583_;
  assign new_n2585_ = ~B8716 & new_n2584_;
  assign new_n2586_ = ~B8717 & ~B8716;
  assign new_n2587_ = ~new_n2585_ & ~new_n2586_;
  assign new_n2588_ = B8715 & new_n2587_;
  assign new_n2589_ = ~B8715 & ~new_n2587_;
  assign new_n2590_ = ~new_n2588_ & ~new_n2589_;
  assign new_n2591_ = ~new_n2584_ & ~new_n2590_;
  assign new_n2592_ = B8747 & ~B8746;
  assign new_n2593_ = ~B8747 & B8746;
  assign new_n2594_ = ~new_n2592_ & ~new_n2593_;
  assign new_n2595_ = ~B8749 & new_n2594_;
  assign new_n2596_ = ~B8750 & ~B8749;
  assign new_n2597_ = ~new_n2595_ & ~new_n2596_;
  assign new_n2598_ = B8748 & new_n2597_;
  assign new_n2599_ = ~B8748 & ~new_n2597_;
  assign new_n2600_ = ~new_n2598_ & ~new_n2599_;
  assign new_n2601_ = ~new_n2594_ & ~new_n2600_;
  assign new_n2602_ = new_n2581_ & ~new_n2601_;
  assign new_n2603_ = B8780 & ~B8779;
  assign new_n2604_ = ~B8780 & B8779;
  assign new_n2605_ = ~new_n2603_ & ~new_n2604_;
  assign new_n2606_ = ~B8782 & new_n2605_;
  assign new_n2607_ = ~B8783 & ~B8782;
  assign new_n2608_ = ~new_n2606_ & ~new_n2607_;
  assign new_n2609_ = B8781 & new_n2608_;
  assign new_n2610_ = ~B8781 & ~new_n2608_;
  assign new_n2611_ = ~new_n2609_ & ~new_n2610_;
  assign new_n2612_ = ~new_n2605_ & ~new_n2611_;
  assign new_n2613_ = ~new_n2601_ & ~new_n2612_;
  assign new_n2614_ = ~new_n2602_ & ~new_n2613_;
  assign new_n2615_ = new_n2591_ & new_n2614_;
  assign new_n2616_ = ~new_n2591_ & ~new_n2614_;
  assign new_n2617_ = ~new_n2615_ & ~new_n2616_;
  assign new_n2618_ = ~new_n2581_ & ~new_n2617_;
  assign new_n2619_ = ~new_n2558_ & new_n2618_;
  assign new_n2620_ = new_n2558_ & ~new_n2618_;
  assign new_n2621_ = ~new_n2619_ & ~new_n2620_;
  assign new_n2622_ = B8813 & ~B8812;
  assign new_n2623_ = ~B8813 & B8812;
  assign new_n2624_ = ~new_n2622_ & ~new_n2623_;
  assign new_n2625_ = ~B8815 & new_n2624_;
  assign new_n2626_ = ~B8816 & ~B8815;
  assign new_n2627_ = ~new_n2625_ & ~new_n2626_;
  assign new_n2628_ = B8814 & new_n2627_;
  assign new_n2629_ = ~B8814 & ~new_n2627_;
  assign new_n2630_ = ~new_n2628_ & ~new_n2629_;
  assign new_n2631_ = ~new_n2624_ & ~new_n2630_;
  assign new_n2632_ = B8846 & ~B8845;
  assign new_n2633_ = ~B8846 & B8845;
  assign new_n2634_ = ~new_n2632_ & ~new_n2633_;
  assign new_n2635_ = ~B8848 & new_n2634_;
  assign new_n2636_ = ~B8849 & ~B8848;
  assign new_n2637_ = ~new_n2635_ & ~new_n2636_;
  assign new_n2638_ = B8847 & new_n2637_;
  assign new_n2639_ = ~B8847 & ~new_n2637_;
  assign new_n2640_ = ~new_n2638_ & ~new_n2639_;
  assign new_n2641_ = ~new_n2634_ & ~new_n2640_;
  assign new_n2642_ = ~new_n2631_ & new_n2641_;
  assign new_n2643_ = new_n2631_ & ~new_n2641_;
  assign new_n2644_ = ~new_n2642_ & ~new_n2643_;
  assign new_n2645_ = B8879 & ~B8878;
  assign new_n2646_ = ~B8879 & B8878;
  assign new_n2647_ = ~new_n2645_ & ~new_n2646_;
  assign new_n2648_ = ~B8881 & new_n2647_;
  assign new_n2649_ = ~B8882 & ~B8881;
  assign new_n2650_ = ~new_n2648_ & ~new_n2649_;
  assign new_n2651_ = B8880 & new_n2650_;
  assign new_n2652_ = ~B8880 & ~new_n2650_;
  assign new_n2653_ = ~new_n2651_ & ~new_n2652_;
  assign new_n2654_ = ~new_n2647_ & ~new_n2653_;
  assign new_n2655_ = B8912 & ~B8911;
  assign new_n2656_ = ~B8912 & B8911;
  assign new_n2657_ = ~new_n2655_ & ~new_n2656_;
  assign new_n2658_ = ~B8914 & new_n2657_;
  assign new_n2659_ = ~B8915 & ~B8914;
  assign new_n2660_ = ~new_n2658_ & ~new_n2659_;
  assign new_n2661_ = B8913 & new_n2660_;
  assign new_n2662_ = ~B8913 & ~new_n2660_;
  assign new_n2663_ = ~new_n2661_ & ~new_n2662_;
  assign new_n2664_ = ~new_n2657_ & ~new_n2663_;
  assign new_n2665_ = new_n2644_ & ~new_n2664_;
  assign new_n2666_ = B8945 & ~B8944;
  assign new_n2667_ = ~B8945 & B8944;
  assign new_n2668_ = ~new_n2666_ & ~new_n2667_;
  assign new_n2669_ = ~B8947 & new_n2668_;
  assign new_n2670_ = ~B8948 & ~B8947;
  assign new_n2671_ = ~new_n2669_ & ~new_n2670_;
  assign new_n2672_ = B8946 & new_n2671_;
  assign new_n2673_ = ~B8946 & ~new_n2671_;
  assign new_n2674_ = ~new_n2672_ & ~new_n2673_;
  assign new_n2675_ = ~new_n2668_ & ~new_n2674_;
  assign new_n2676_ = ~new_n2664_ & ~new_n2675_;
  assign new_n2677_ = ~new_n2665_ & ~new_n2676_;
  assign new_n2678_ = new_n2654_ & new_n2677_;
  assign new_n2679_ = ~new_n2654_ & ~new_n2677_;
  assign new_n2680_ = ~new_n2678_ & ~new_n2679_;
  assign new_n2681_ = ~new_n2644_ & ~new_n2680_;
  assign new_n2682_ = B8978 & ~B8977;
  assign new_n2683_ = ~B8978 & B8977;
  assign new_n2684_ = ~new_n2682_ & ~new_n2683_;
  assign new_n2685_ = ~B8980 & new_n2684_;
  assign new_n2686_ = ~B8981 & ~B8980;
  assign new_n2687_ = ~new_n2685_ & ~new_n2686_;
  assign new_n2688_ = B8979 & new_n2687_;
  assign new_n2689_ = ~B8979 & ~new_n2687_;
  assign new_n2690_ = ~new_n2688_ & ~new_n2689_;
  assign new_n2691_ = ~new_n2684_ & ~new_n2690_;
  assign new_n2692_ = B9011 & ~B9010;
  assign new_n2693_ = ~B9011 & B9010;
  assign new_n2694_ = ~new_n2692_ & ~new_n2693_;
  assign new_n2695_ = ~B9013 & new_n2694_;
  assign new_n2696_ = ~B9014 & ~B9013;
  assign new_n2697_ = ~new_n2695_ & ~new_n2696_;
  assign new_n2698_ = B9012 & new_n2697_;
  assign new_n2699_ = ~B9012 & ~new_n2697_;
  assign new_n2700_ = ~new_n2698_ & ~new_n2699_;
  assign new_n2701_ = ~new_n2694_ & ~new_n2700_;
  assign new_n2702_ = ~new_n2691_ & new_n2701_;
  assign new_n2703_ = new_n2691_ & ~new_n2701_;
  assign new_n2704_ = ~new_n2702_ & ~new_n2703_;
  assign new_n2705_ = B9044 & ~B9043;
  assign new_n2706_ = ~B9044 & B9043;
  assign new_n2707_ = ~new_n2705_ & ~new_n2706_;
  assign new_n2708_ = ~B9046 & new_n2707_;
  assign new_n2709_ = ~B9047 & ~B9046;
  assign new_n2710_ = ~new_n2708_ & ~new_n2709_;
  assign new_n2711_ = B9045 & new_n2710_;
  assign new_n2712_ = ~B9045 & ~new_n2710_;
  assign new_n2713_ = ~new_n2711_ & ~new_n2712_;
  assign new_n2714_ = ~new_n2707_ & ~new_n2713_;
  assign new_n2715_ = B9077 & ~B9076;
  assign new_n2716_ = ~B9077 & B9076;
  assign new_n2717_ = ~new_n2715_ & ~new_n2716_;
  assign new_n2718_ = ~B9079 & new_n2717_;
  assign new_n2719_ = ~B9080 & ~B9079;
  assign new_n2720_ = ~new_n2718_ & ~new_n2719_;
  assign new_n2721_ = B9078 & new_n2720_;
  assign new_n2722_ = ~B9078 & ~new_n2720_;
  assign new_n2723_ = ~new_n2721_ & ~new_n2722_;
  assign new_n2724_ = ~new_n2717_ & ~new_n2723_;
  assign new_n2725_ = new_n2704_ & ~new_n2724_;
  assign new_n2726_ = B9110 & ~B9109;
  assign new_n2727_ = ~B9110 & B9109;
  assign new_n2728_ = ~new_n2726_ & ~new_n2727_;
  assign new_n2729_ = ~B9112 & new_n2728_;
  assign new_n2730_ = ~B9113 & ~B9112;
  assign new_n2731_ = ~new_n2729_ & ~new_n2730_;
  assign new_n2732_ = B9111 & new_n2731_;
  assign new_n2733_ = ~B9111 & ~new_n2731_;
  assign new_n2734_ = ~new_n2732_ & ~new_n2733_;
  assign new_n2735_ = ~new_n2728_ & ~new_n2734_;
  assign new_n2736_ = ~new_n2724_ & ~new_n2735_;
  assign new_n2737_ = ~new_n2725_ & ~new_n2736_;
  assign new_n2738_ = new_n2714_ & new_n2737_;
  assign new_n2739_ = ~new_n2714_ & ~new_n2737_;
  assign new_n2740_ = ~new_n2738_ & ~new_n2739_;
  assign new_n2741_ = ~new_n2704_ & ~new_n2740_;
  assign new_n2742_ = new_n2621_ & ~new_n2741_;
  assign new_n2743_ = B9143 & ~B9142;
  assign new_n2744_ = ~B9143 & B9142;
  assign new_n2745_ = ~new_n2743_ & ~new_n2744_;
  assign new_n2746_ = ~B9145 & new_n2745_;
  assign new_n2747_ = ~B9146 & ~B9145;
  assign new_n2748_ = ~new_n2746_ & ~new_n2747_;
  assign new_n2749_ = B9144 & new_n2748_;
  assign new_n2750_ = ~B9144 & ~new_n2748_;
  assign new_n2751_ = ~new_n2749_ & ~new_n2750_;
  assign new_n2752_ = ~new_n2745_ & ~new_n2751_;
  assign new_n2753_ = B9176 & ~B9175;
  assign new_n2754_ = ~B9176 & B9175;
  assign new_n2755_ = ~new_n2753_ & ~new_n2754_;
  assign new_n2756_ = ~B9178 & new_n2755_;
  assign new_n2757_ = ~B9179 & ~B9178;
  assign new_n2758_ = ~new_n2756_ & ~new_n2757_;
  assign new_n2759_ = B9177 & new_n2758_;
  assign new_n2760_ = ~B9177 & ~new_n2758_;
  assign new_n2761_ = ~new_n2759_ & ~new_n2760_;
  assign new_n2762_ = ~new_n2755_ & ~new_n2761_;
  assign new_n2763_ = ~new_n2752_ & new_n2762_;
  assign new_n2764_ = new_n2752_ & ~new_n2762_;
  assign new_n2765_ = ~new_n2763_ & ~new_n2764_;
  assign new_n2766_ = B9209 & ~B9208;
  assign new_n2767_ = ~B9209 & B9208;
  assign new_n2768_ = ~new_n2766_ & ~new_n2767_;
  assign new_n2769_ = ~B9211 & new_n2768_;
  assign new_n2770_ = ~B9212 & ~B9211;
  assign new_n2771_ = ~new_n2769_ & ~new_n2770_;
  assign new_n2772_ = B9210 & new_n2771_;
  assign new_n2773_ = ~B9210 & ~new_n2771_;
  assign new_n2774_ = ~new_n2772_ & ~new_n2773_;
  assign new_n2775_ = ~new_n2768_ & ~new_n2774_;
  assign new_n2776_ = B9242 & ~B9241;
  assign new_n2777_ = ~B9242 & B9241;
  assign new_n2778_ = ~new_n2776_ & ~new_n2777_;
  assign new_n2779_ = ~B9244 & new_n2778_;
  assign new_n2780_ = ~B9245 & ~B9244;
  assign new_n2781_ = ~new_n2779_ & ~new_n2780_;
  assign new_n2782_ = B9243 & new_n2781_;
  assign new_n2783_ = ~B9243 & ~new_n2781_;
  assign new_n2784_ = ~new_n2782_ & ~new_n2783_;
  assign new_n2785_ = ~new_n2778_ & ~new_n2784_;
  assign new_n2786_ = new_n2765_ & ~new_n2785_;
  assign new_n2787_ = B9275 & ~B9274;
  assign new_n2788_ = ~B9275 & B9274;
  assign new_n2789_ = ~new_n2787_ & ~new_n2788_;
  assign new_n2790_ = ~B9277 & new_n2789_;
  assign new_n2791_ = ~B9278 & ~B9277;
  assign new_n2792_ = ~new_n2790_ & ~new_n2791_;
  assign new_n2793_ = B9276 & new_n2792_;
  assign new_n2794_ = ~B9276 & ~new_n2792_;
  assign new_n2795_ = ~new_n2793_ & ~new_n2794_;
  assign new_n2796_ = ~new_n2789_ & ~new_n2795_;
  assign new_n2797_ = ~new_n2785_ & ~new_n2796_;
  assign new_n2798_ = ~new_n2786_ & ~new_n2797_;
  assign new_n2799_ = new_n2775_ & new_n2798_;
  assign new_n2800_ = ~new_n2775_ & ~new_n2798_;
  assign new_n2801_ = ~new_n2799_ & ~new_n2800_;
  assign new_n2802_ = ~new_n2765_ & ~new_n2801_;
  assign new_n2803_ = ~new_n2741_ & ~new_n2802_;
  assign new_n2804_ = ~new_n2742_ & ~new_n2803_;
  assign new_n2805_ = new_n2681_ & new_n2804_;
  assign new_n2806_ = ~new_n2681_ & ~new_n2804_;
  assign new_n2807_ = ~new_n2805_ & ~new_n2806_;
  assign new_n2808_ = ~new_n2621_ & ~new_n2807_;
  assign new_n2809_ = ~new_n2497_ & ~new_n2808_;
  assign new_n2810_ = ~new_n2498_ & ~new_n2809_;
  assign new_n2811_ = new_n2187_ & new_n2810_;
  assign new_n2812_ = ~new_n2187_ & ~new_n2810_;
  assign new_n2813_ = ~new_n2811_ & ~new_n2812_;
  assign A6907 = ~new_n1877_ & ~new_n2813_;
  assign new_n2815_ = ~new_n1874_ & ~new_n2811_;
  assign A6906 = ~new_n1877_ & ~new_n2815_;
  assign new_n2817_ = new_n1874_ & new_n2187_;
  assign new_n2818_ = ~new_n1877_ & ~new_n2817_;
  assign new_n2819_ = new_n1877_ & ~new_n2818_;
  assign new_n2820_ = new_n1877_ & new_n2817_;
  assign new_n2821_ = new_n2819_ & ~new_n2820_;
  assign new_n2822_ = new_n2187_ & ~new_n2821_;
  assign A6905 = new_n2810_ | new_n2822_;
  assign new_n2824_ = new_n2497_ & new_n2808_;
  assign new_n2825_ = ~new_n2809_ & ~new_n2824_;
  assign new_n2826_ = ~new_n1877_ & ~new_n2497_;
  assign new_n2827_ = new_n1877_ & new_n2497_;
  assign new_n2828_ = ~new_n2826_ & ~new_n2827_;
  assign new_n2829_ = new_n2825_ & ~new_n2828_;
  assign A6904 = new_n2822_ | new_n2829_;
  assign new_n2831_ = new_n2187_ & ~new_n2829_;
  assign new_n2832_ = ~new_n2187_ & new_n2829_;
  assign new_n2833_ = ~new_n2831_ & ~new_n2832_;
  assign A6903 = ~new_n1877_ & ~new_n2833_;
  assign new_n2835_ = B5183 & B5184;
  assign new_n2836_ = ~new_n1256_ & ~new_n2835_;
  assign new_n2837_ = new_n1256_ & ~new_n2836_;
  assign new_n2838_ = new_n1256_ & new_n2835_;
  assign new_n2839_ = new_n2837_ & ~new_n2838_;
  assign new_n2840_ = B5184 & ~new_n2839_;
  assign new_n2841_ = ~new_n1260_ & ~new_n2840_;
  assign new_n2842_ = ~B5216 & ~new_n1271_;
  assign new_n2843_ = ~new_n1267_ & ~new_n2842_;
  assign new_n2844_ = new_n2841_ & new_n2843_;
  assign new_n2845_ = ~new_n2841_ & ~new_n2843_;
  assign new_n2846_ = ~new_n2844_ & ~new_n2845_;
  assign new_n2847_ = ~B5249 & ~new_n1284_;
  assign new_n2848_ = ~new_n1280_ & ~new_n2847_;
  assign new_n2849_ = ~B5282 & ~new_n1294_;
  assign new_n2850_ = ~new_n1290_ & ~new_n2849_;
  assign new_n2851_ = new_n2846_ & ~new_n2850_;
  assign new_n2852_ = ~B5315 & ~new_n1305_;
  assign new_n2853_ = ~new_n1301_ & ~new_n2852_;
  assign new_n2854_ = ~new_n2850_ & ~new_n2853_;
  assign new_n2855_ = ~new_n2851_ & ~new_n2854_;
  assign new_n2856_ = new_n2848_ & new_n2855_;
  assign new_n2857_ = ~new_n2848_ & ~new_n2855_;
  assign new_n2858_ = ~new_n2856_ & ~new_n2857_;
  assign new_n2859_ = ~new_n2846_ & ~new_n2858_;
  assign new_n2860_ = ~B5348 & ~new_n1321_;
  assign new_n2861_ = ~new_n1317_ & ~new_n2860_;
  assign new_n2862_ = ~B5381 & ~new_n1331_;
  assign new_n2863_ = ~new_n1327_ & ~new_n2862_;
  assign new_n2864_ = ~new_n2861_ & new_n2863_;
  assign new_n2865_ = new_n2861_ & ~new_n2863_;
  assign new_n2866_ = ~new_n2864_ & ~new_n2865_;
  assign new_n2867_ = ~B5414 & ~new_n1344_;
  assign new_n2868_ = ~new_n1340_ & ~new_n2867_;
  assign new_n2869_ = ~B5447 & ~new_n1354_;
  assign new_n2870_ = ~new_n1350_ & ~new_n2869_;
  assign new_n2871_ = new_n2866_ & ~new_n2870_;
  assign new_n2872_ = ~B5480 & ~new_n1365_;
  assign new_n2873_ = ~new_n1361_ & ~new_n2872_;
  assign new_n2874_ = ~new_n2870_ & ~new_n2873_;
  assign new_n2875_ = ~new_n2871_ & ~new_n2874_;
  assign new_n2876_ = new_n2868_ & new_n2875_;
  assign new_n2877_ = ~new_n2868_ & ~new_n2875_;
  assign new_n2878_ = ~new_n2876_ & ~new_n2877_;
  assign new_n2879_ = ~new_n2866_ & ~new_n2878_;
  assign new_n2880_ = ~new_n2859_ & new_n2879_;
  assign new_n2881_ = new_n2859_ & ~new_n2879_;
  assign new_n2882_ = ~new_n2880_ & ~new_n2881_;
  assign new_n2883_ = ~B5513 & ~new_n1384_;
  assign new_n2884_ = ~new_n1380_ & ~new_n2883_;
  assign new_n2885_ = ~B5546 & ~new_n1394_;
  assign new_n2886_ = ~new_n1390_ & ~new_n2885_;
  assign new_n2887_ = ~new_n2884_ & new_n2886_;
  assign new_n2888_ = new_n2884_ & ~new_n2886_;
  assign new_n2889_ = ~new_n2887_ & ~new_n2888_;
  assign new_n2890_ = ~B5579 & ~new_n1407_;
  assign new_n2891_ = ~new_n1403_ & ~new_n2890_;
  assign new_n2892_ = ~B5612 & ~new_n1417_;
  assign new_n2893_ = ~new_n1413_ & ~new_n2892_;
  assign new_n2894_ = new_n2889_ & ~new_n2893_;
  assign new_n2895_ = ~B5645 & ~new_n1428_;
  assign new_n2896_ = ~new_n1424_ & ~new_n2895_;
  assign new_n2897_ = ~new_n2893_ & ~new_n2896_;
  assign new_n2898_ = ~new_n2894_ & ~new_n2897_;
  assign new_n2899_ = new_n2891_ & new_n2898_;
  assign new_n2900_ = ~new_n2891_ & ~new_n2898_;
  assign new_n2901_ = ~new_n2899_ & ~new_n2900_;
  assign new_n2902_ = ~new_n2889_ & ~new_n2901_;
  assign new_n2903_ = ~B5678 & ~new_n1444_;
  assign new_n2904_ = ~new_n1440_ & ~new_n2903_;
  assign new_n2905_ = ~B5711 & ~new_n1454_;
  assign new_n2906_ = ~new_n1450_ & ~new_n2905_;
  assign new_n2907_ = ~new_n2904_ & new_n2906_;
  assign new_n2908_ = new_n2904_ & ~new_n2906_;
  assign new_n2909_ = ~new_n2907_ & ~new_n2908_;
  assign new_n2910_ = ~B5744 & ~new_n1467_;
  assign new_n2911_ = ~new_n1463_ & ~new_n2910_;
  assign new_n2912_ = ~B5777 & ~new_n1477_;
  assign new_n2913_ = ~new_n1473_ & ~new_n2912_;
  assign new_n2914_ = new_n2909_ & ~new_n2913_;
  assign new_n2915_ = ~B5810 & ~new_n1488_;
  assign new_n2916_ = ~new_n1484_ & ~new_n2915_;
  assign new_n2917_ = ~new_n2913_ & ~new_n2916_;
  assign new_n2918_ = ~new_n2914_ & ~new_n2917_;
  assign new_n2919_ = new_n2911_ & new_n2918_;
  assign new_n2920_ = ~new_n2911_ & ~new_n2918_;
  assign new_n2921_ = ~new_n2919_ & ~new_n2920_;
  assign new_n2922_ = ~new_n2909_ & ~new_n2921_;
  assign new_n2923_ = new_n2882_ & ~new_n2922_;
  assign new_n2924_ = ~B5843 & ~new_n1505_;
  assign new_n2925_ = ~new_n1501_ & ~new_n2924_;
  assign new_n2926_ = ~B5876 & ~new_n1515_;
  assign new_n2927_ = ~new_n1511_ & ~new_n2926_;
  assign new_n2928_ = ~new_n2925_ & new_n2927_;
  assign new_n2929_ = new_n2925_ & ~new_n2927_;
  assign new_n2930_ = ~new_n2928_ & ~new_n2929_;
  assign new_n2931_ = ~B5909 & ~new_n1528_;
  assign new_n2932_ = ~new_n1524_ & ~new_n2931_;
  assign new_n2933_ = ~B5942 & ~new_n1538_;
  assign new_n2934_ = ~new_n1534_ & ~new_n2933_;
  assign new_n2935_ = new_n2930_ & ~new_n2934_;
  assign new_n2936_ = ~B5975 & ~new_n1549_;
  assign new_n2937_ = ~new_n1545_ & ~new_n2936_;
  assign new_n2938_ = ~new_n2934_ & ~new_n2937_;
  assign new_n2939_ = ~new_n2935_ & ~new_n2938_;
  assign new_n2940_ = new_n2932_ & new_n2939_;
  assign new_n2941_ = ~new_n2932_ & ~new_n2939_;
  assign new_n2942_ = ~new_n2940_ & ~new_n2941_;
  assign new_n2943_ = ~new_n2930_ & ~new_n2942_;
  assign new_n2944_ = ~new_n2922_ & ~new_n2943_;
  assign new_n2945_ = ~new_n2923_ & ~new_n2944_;
  assign new_n2946_ = new_n2902_ & new_n2945_;
  assign new_n2947_ = ~new_n2902_ & ~new_n2945_;
  assign new_n2948_ = ~new_n2946_ & ~new_n2947_;
  assign new_n2949_ = ~new_n2882_ & ~new_n2948_;
  assign new_n2950_ = ~B6008 & ~new_n1571_;
  assign new_n2951_ = ~new_n1567_ & ~new_n2950_;
  assign new_n2952_ = ~B6041 & ~new_n1581_;
  assign new_n2953_ = ~new_n1577_ & ~new_n2952_;
  assign new_n2954_ = ~new_n2951_ & new_n2953_;
  assign new_n2955_ = new_n2951_ & ~new_n2953_;
  assign new_n2956_ = ~new_n2954_ & ~new_n2955_;
  assign new_n2957_ = ~B6074 & ~new_n1594_;
  assign new_n2958_ = ~new_n1590_ & ~new_n2957_;
  assign new_n2959_ = ~B6107 & ~new_n1604_;
  assign new_n2960_ = ~new_n1600_ & ~new_n2959_;
  assign new_n2961_ = new_n2956_ & ~new_n2960_;
  assign new_n2962_ = ~B6140 & ~new_n1615_;
  assign new_n2963_ = ~new_n1611_ & ~new_n2962_;
  assign new_n2964_ = ~new_n2960_ & ~new_n2963_;
  assign new_n2965_ = ~new_n2961_ & ~new_n2964_;
  assign new_n2966_ = new_n2958_ & new_n2965_;
  assign new_n2967_ = ~new_n2958_ & ~new_n2965_;
  assign new_n2968_ = ~new_n2966_ & ~new_n2967_;
  assign new_n2969_ = ~new_n2956_ & ~new_n2968_;
  assign new_n2970_ = ~B6173 & ~new_n1631_;
  assign new_n2971_ = ~new_n1627_ & ~new_n2970_;
  assign new_n2972_ = ~B6206 & ~new_n1641_;
  assign new_n2973_ = ~new_n1637_ & ~new_n2972_;
  assign new_n2974_ = ~new_n2971_ & new_n2973_;
  assign new_n2975_ = new_n2971_ & ~new_n2973_;
  assign new_n2976_ = ~new_n2974_ & ~new_n2975_;
  assign new_n2977_ = ~B6239 & ~new_n1654_;
  assign new_n2978_ = ~new_n1650_ & ~new_n2977_;
  assign new_n2979_ = ~B6272 & ~new_n1664_;
  assign new_n2980_ = ~new_n1660_ & ~new_n2979_;
  assign new_n2981_ = new_n2976_ & ~new_n2980_;
  assign new_n2982_ = ~B6305 & ~new_n1675_;
  assign new_n2983_ = ~new_n1671_ & ~new_n2982_;
  assign new_n2984_ = ~new_n2980_ & ~new_n2983_;
  assign new_n2985_ = ~new_n2981_ & ~new_n2984_;
  assign new_n2986_ = new_n2978_ & new_n2985_;
  assign new_n2987_ = ~new_n2978_ & ~new_n2985_;
  assign new_n2988_ = ~new_n2986_ & ~new_n2987_;
  assign new_n2989_ = ~new_n2976_ & ~new_n2988_;
  assign new_n2990_ = ~new_n2969_ & new_n2989_;
  assign new_n2991_ = new_n2969_ & ~new_n2989_;
  assign new_n2992_ = ~new_n2990_ & ~new_n2991_;
  assign new_n2993_ = ~B6338 & ~new_n1694_;
  assign new_n2994_ = ~new_n1690_ & ~new_n2993_;
  assign new_n2995_ = ~B6371 & ~new_n1704_;
  assign new_n2996_ = ~new_n1700_ & ~new_n2995_;
  assign new_n2997_ = ~new_n2994_ & new_n2996_;
  assign new_n2998_ = new_n2994_ & ~new_n2996_;
  assign new_n2999_ = ~new_n2997_ & ~new_n2998_;
  assign new_n3000_ = ~B6404 & ~new_n1717_;
  assign new_n3001_ = ~new_n1713_ & ~new_n3000_;
  assign new_n3002_ = ~B6437 & ~new_n1727_;
  assign new_n3003_ = ~new_n1723_ & ~new_n3002_;
  assign new_n3004_ = new_n2999_ & ~new_n3003_;
  assign new_n3005_ = ~B6470 & ~new_n1738_;
  assign new_n3006_ = ~new_n1734_ & ~new_n3005_;
  assign new_n3007_ = ~new_n3003_ & ~new_n3006_;
  assign new_n3008_ = ~new_n3004_ & ~new_n3007_;
  assign new_n3009_ = new_n3001_ & new_n3008_;
  assign new_n3010_ = ~new_n3001_ & ~new_n3008_;
  assign new_n3011_ = ~new_n3009_ & ~new_n3010_;
  assign new_n3012_ = ~new_n2999_ & ~new_n3011_;
  assign new_n3013_ = ~B6503 & ~new_n1754_;
  assign new_n3014_ = ~new_n1750_ & ~new_n3013_;
  assign new_n3015_ = ~B6536 & ~new_n1764_;
  assign new_n3016_ = ~new_n1760_ & ~new_n3015_;
  assign new_n3017_ = ~new_n3014_ & new_n3016_;
  assign new_n3018_ = new_n3014_ & ~new_n3016_;
  assign new_n3019_ = ~new_n3017_ & ~new_n3018_;
  assign new_n3020_ = ~B6569 & ~new_n1777_;
  assign new_n3021_ = ~new_n1773_ & ~new_n3020_;
  assign new_n3022_ = ~B6602 & ~new_n1787_;
  assign new_n3023_ = ~new_n1783_ & ~new_n3022_;
  assign new_n3024_ = new_n3019_ & ~new_n3023_;
  assign new_n3025_ = ~B6635 & ~new_n1798_;
  assign new_n3026_ = ~new_n1794_ & ~new_n3025_;
  assign new_n3027_ = ~new_n3023_ & ~new_n3026_;
  assign new_n3028_ = ~new_n3024_ & ~new_n3027_;
  assign new_n3029_ = new_n3021_ & new_n3028_;
  assign new_n3030_ = ~new_n3021_ & ~new_n3028_;
  assign new_n3031_ = ~new_n3029_ & ~new_n3030_;
  assign new_n3032_ = ~new_n3019_ & ~new_n3031_;
  assign new_n3033_ = new_n2992_ & ~new_n3032_;
  assign new_n3034_ = ~B6668 & ~new_n1815_;
  assign new_n3035_ = ~new_n1811_ & ~new_n3034_;
  assign new_n3036_ = ~B6701 & ~new_n1825_;
  assign new_n3037_ = ~new_n1821_ & ~new_n3036_;
  assign new_n3038_ = ~new_n3035_ & new_n3037_;
  assign new_n3039_ = new_n3035_ & ~new_n3037_;
  assign new_n3040_ = ~new_n3038_ & ~new_n3039_;
  assign new_n3041_ = ~B6734 & ~new_n1838_;
  assign new_n3042_ = ~new_n1834_ & ~new_n3041_;
  assign new_n3043_ = ~B6767 & ~new_n1848_;
  assign new_n3044_ = ~new_n1844_ & ~new_n3043_;
  assign new_n3045_ = new_n3040_ & ~new_n3044_;
  assign new_n3046_ = ~B6800 & ~new_n1859_;
  assign new_n3047_ = ~new_n1855_ & ~new_n3046_;
  assign new_n3048_ = ~new_n3044_ & ~new_n3047_;
  assign new_n3049_ = ~new_n3045_ & ~new_n3048_;
  assign new_n3050_ = new_n3042_ & new_n3049_;
  assign new_n3051_ = ~new_n3042_ & ~new_n3049_;
  assign new_n3052_ = ~new_n3050_ & ~new_n3051_;
  assign new_n3053_ = ~new_n3040_ & ~new_n3052_;
  assign new_n3054_ = ~new_n3032_ & ~new_n3053_;
  assign new_n3055_ = ~new_n3033_ & ~new_n3054_;
  assign new_n3056_ = new_n3012_ & new_n3055_;
  assign new_n3057_ = ~new_n3012_ & ~new_n3055_;
  assign new_n3058_ = ~new_n3056_ & ~new_n3057_;
  assign new_n3059_ = ~new_n2992_ & ~new_n3058_;
  assign new_n3060_ = ~new_n2949_ & new_n3059_;
  assign new_n3061_ = new_n2949_ & ~new_n3059_;
  assign new_n3062_ = ~new_n3060_ & ~new_n3061_;
  assign new_n3063_ = ~B6833 & ~new_n1884_;
  assign new_n3064_ = ~new_n1880_ & ~new_n3063_;
  assign new_n3065_ = ~B6866 & ~new_n1894_;
  assign new_n3066_ = ~new_n1890_ & ~new_n3065_;
  assign new_n3067_ = ~new_n3064_ & new_n3066_;
  assign new_n3068_ = new_n3064_ & ~new_n3066_;
  assign new_n3069_ = ~new_n3067_ & ~new_n3068_;
  assign new_n3070_ = ~B6899 & ~new_n1907_;
  assign new_n3071_ = ~new_n1903_ & ~new_n3070_;
  assign new_n3072_ = ~B6932 & ~new_n1917_;
  assign new_n3073_ = ~new_n1913_ & ~new_n3072_;
  assign new_n3074_ = new_n3069_ & ~new_n3073_;
  assign new_n3075_ = ~B6965 & ~new_n1928_;
  assign new_n3076_ = ~new_n1924_ & ~new_n3075_;
  assign new_n3077_ = ~new_n3073_ & ~new_n3076_;
  assign new_n3078_ = ~new_n3074_ & ~new_n3077_;
  assign new_n3079_ = new_n3071_ & new_n3078_;
  assign new_n3080_ = ~new_n3071_ & ~new_n3078_;
  assign new_n3081_ = ~new_n3079_ & ~new_n3080_;
  assign new_n3082_ = ~new_n3069_ & ~new_n3081_;
  assign new_n3083_ = ~B6998 & ~new_n1944_;
  assign new_n3084_ = ~new_n1940_ & ~new_n3083_;
  assign new_n3085_ = ~B7031 & ~new_n1954_;
  assign new_n3086_ = ~new_n1950_ & ~new_n3085_;
  assign new_n3087_ = ~new_n3084_ & new_n3086_;
  assign new_n3088_ = new_n3084_ & ~new_n3086_;
  assign new_n3089_ = ~new_n3087_ & ~new_n3088_;
  assign new_n3090_ = ~B7064 & ~new_n1967_;
  assign new_n3091_ = ~new_n1963_ & ~new_n3090_;
  assign new_n3092_ = ~B7097 & ~new_n1977_;
  assign new_n3093_ = ~new_n1973_ & ~new_n3092_;
  assign new_n3094_ = new_n3089_ & ~new_n3093_;
  assign new_n3095_ = ~B7130 & ~new_n1988_;
  assign new_n3096_ = ~new_n1984_ & ~new_n3095_;
  assign new_n3097_ = ~new_n3093_ & ~new_n3096_;
  assign new_n3098_ = ~new_n3094_ & ~new_n3097_;
  assign new_n3099_ = new_n3091_ & new_n3098_;
  assign new_n3100_ = ~new_n3091_ & ~new_n3098_;
  assign new_n3101_ = ~new_n3099_ & ~new_n3100_;
  assign new_n3102_ = ~new_n3089_ & ~new_n3101_;
  assign new_n3103_ = ~new_n3082_ & new_n3102_;
  assign new_n3104_ = new_n3082_ & ~new_n3102_;
  assign new_n3105_ = ~new_n3103_ & ~new_n3104_;
  assign new_n3106_ = ~B7163 & ~new_n2007_;
  assign new_n3107_ = ~new_n2003_ & ~new_n3106_;
  assign new_n3108_ = ~B7196 & ~new_n2017_;
  assign new_n3109_ = ~new_n2013_ & ~new_n3108_;
  assign new_n3110_ = ~new_n3107_ & new_n3109_;
  assign new_n3111_ = new_n3107_ & ~new_n3109_;
  assign new_n3112_ = ~new_n3110_ & ~new_n3111_;
  assign new_n3113_ = ~B7229 & ~new_n2030_;
  assign new_n3114_ = ~new_n2026_ & ~new_n3113_;
  assign new_n3115_ = ~B7262 & ~new_n2040_;
  assign new_n3116_ = ~new_n2036_ & ~new_n3115_;
  assign new_n3117_ = new_n3112_ & ~new_n3116_;
  assign new_n3118_ = ~B7295 & ~new_n2051_;
  assign new_n3119_ = ~new_n2047_ & ~new_n3118_;
  assign new_n3120_ = ~new_n3116_ & ~new_n3119_;
  assign new_n3121_ = ~new_n3117_ & ~new_n3120_;
  assign new_n3122_ = new_n3114_ & new_n3121_;
  assign new_n3123_ = ~new_n3114_ & ~new_n3121_;
  assign new_n3124_ = ~new_n3122_ & ~new_n3123_;
  assign new_n3125_ = ~new_n3112_ & ~new_n3124_;
  assign new_n3126_ = ~B7328 & ~new_n2067_;
  assign new_n3127_ = ~new_n2063_ & ~new_n3126_;
  assign new_n3128_ = ~B7361 & ~new_n2077_;
  assign new_n3129_ = ~new_n2073_ & ~new_n3128_;
  assign new_n3130_ = ~new_n3127_ & new_n3129_;
  assign new_n3131_ = new_n3127_ & ~new_n3129_;
  assign new_n3132_ = ~new_n3130_ & ~new_n3131_;
  assign new_n3133_ = ~B7394 & ~new_n2090_;
  assign new_n3134_ = ~new_n2086_ & ~new_n3133_;
  assign new_n3135_ = ~B7427 & ~new_n2100_;
  assign new_n3136_ = ~new_n2096_ & ~new_n3135_;
  assign new_n3137_ = new_n3132_ & ~new_n3136_;
  assign new_n3138_ = ~B7460 & ~new_n2111_;
  assign new_n3139_ = ~new_n2107_ & ~new_n3138_;
  assign new_n3140_ = ~new_n3136_ & ~new_n3139_;
  assign new_n3141_ = ~new_n3137_ & ~new_n3140_;
  assign new_n3142_ = new_n3134_ & new_n3141_;
  assign new_n3143_ = ~new_n3134_ & ~new_n3141_;
  assign new_n3144_ = ~new_n3142_ & ~new_n3143_;
  assign new_n3145_ = ~new_n3132_ & ~new_n3144_;
  assign new_n3146_ = new_n3105_ & ~new_n3145_;
  assign new_n3147_ = ~B7493 & ~new_n2128_;
  assign new_n3148_ = ~new_n2124_ & ~new_n3147_;
  assign new_n3149_ = ~B7526 & ~new_n2138_;
  assign new_n3150_ = ~new_n2134_ & ~new_n3149_;
  assign new_n3151_ = ~new_n3148_ & new_n3150_;
  assign new_n3152_ = new_n3148_ & ~new_n3150_;
  assign new_n3153_ = ~new_n3151_ & ~new_n3152_;
  assign new_n3154_ = ~B7559 & ~new_n2151_;
  assign new_n3155_ = ~new_n2147_ & ~new_n3154_;
  assign new_n3156_ = ~B7592 & ~new_n2161_;
  assign new_n3157_ = ~new_n2157_ & ~new_n3156_;
  assign new_n3158_ = new_n3153_ & ~new_n3157_;
  assign new_n3159_ = ~B7625 & ~new_n2172_;
  assign new_n3160_ = ~new_n2168_ & ~new_n3159_;
  assign new_n3161_ = ~new_n3157_ & ~new_n3160_;
  assign new_n3162_ = ~new_n3158_ & ~new_n3161_;
  assign new_n3163_ = new_n3155_ & new_n3162_;
  assign new_n3164_ = ~new_n3155_ & ~new_n3162_;
  assign new_n3165_ = ~new_n3163_ & ~new_n3164_;
  assign new_n3166_ = ~new_n3153_ & ~new_n3165_;
  assign new_n3167_ = ~new_n3145_ & ~new_n3166_;
  assign new_n3168_ = ~new_n3146_ & ~new_n3167_;
  assign new_n3169_ = new_n3125_ & new_n3168_;
  assign new_n3170_ = ~new_n3125_ & ~new_n3168_;
  assign new_n3171_ = ~new_n3169_ & ~new_n3170_;
  assign new_n3172_ = ~new_n3105_ & ~new_n3171_;
  assign new_n3173_ = ~B7658 & ~new_n2194_;
  assign new_n3174_ = ~new_n2190_ & ~new_n3173_;
  assign new_n3175_ = ~B7691 & ~new_n2204_;
  assign new_n3176_ = ~new_n2200_ & ~new_n3175_;
  assign new_n3177_ = ~new_n3174_ & new_n3176_;
  assign new_n3178_ = new_n3174_ & ~new_n3176_;
  assign new_n3179_ = ~new_n3177_ & ~new_n3178_;
  assign new_n3180_ = ~B7724 & ~new_n2217_;
  assign new_n3181_ = ~new_n2213_ & ~new_n3180_;
  assign new_n3182_ = ~B7757 & ~new_n2227_;
  assign new_n3183_ = ~new_n2223_ & ~new_n3182_;
  assign new_n3184_ = new_n3179_ & ~new_n3183_;
  assign new_n3185_ = ~B7790 & ~new_n2238_;
  assign new_n3186_ = ~new_n2234_ & ~new_n3185_;
  assign new_n3187_ = ~new_n3183_ & ~new_n3186_;
  assign new_n3188_ = ~new_n3184_ & ~new_n3187_;
  assign new_n3189_ = new_n3181_ & new_n3188_;
  assign new_n3190_ = ~new_n3181_ & ~new_n3188_;
  assign new_n3191_ = ~new_n3189_ & ~new_n3190_;
  assign new_n3192_ = ~new_n3179_ & ~new_n3191_;
  assign new_n3193_ = ~B7823 & ~new_n2254_;
  assign new_n3194_ = ~new_n2250_ & ~new_n3193_;
  assign new_n3195_ = ~B7856 & ~new_n2264_;
  assign new_n3196_ = ~new_n2260_ & ~new_n3195_;
  assign new_n3197_ = ~new_n3194_ & new_n3196_;
  assign new_n3198_ = new_n3194_ & ~new_n3196_;
  assign new_n3199_ = ~new_n3197_ & ~new_n3198_;
  assign new_n3200_ = ~B7889 & ~new_n2277_;
  assign new_n3201_ = ~new_n2273_ & ~new_n3200_;
  assign new_n3202_ = ~B7922 & ~new_n2287_;
  assign new_n3203_ = ~new_n2283_ & ~new_n3202_;
  assign new_n3204_ = new_n3199_ & ~new_n3203_;
  assign new_n3205_ = ~B7955 & ~new_n2298_;
  assign new_n3206_ = ~new_n2294_ & ~new_n3205_;
  assign new_n3207_ = ~new_n3203_ & ~new_n3206_;
  assign new_n3208_ = ~new_n3204_ & ~new_n3207_;
  assign new_n3209_ = new_n3201_ & new_n3208_;
  assign new_n3210_ = ~new_n3201_ & ~new_n3208_;
  assign new_n3211_ = ~new_n3209_ & ~new_n3210_;
  assign new_n3212_ = ~new_n3199_ & ~new_n3211_;
  assign new_n3213_ = ~new_n3192_ & new_n3212_;
  assign new_n3214_ = new_n3192_ & ~new_n3212_;
  assign new_n3215_ = ~new_n3213_ & ~new_n3214_;
  assign new_n3216_ = ~B7988 & ~new_n2317_;
  assign new_n3217_ = ~new_n2313_ & ~new_n3216_;
  assign new_n3218_ = ~B8021 & ~new_n2327_;
  assign new_n3219_ = ~new_n2323_ & ~new_n3218_;
  assign new_n3220_ = ~new_n3217_ & new_n3219_;
  assign new_n3221_ = new_n3217_ & ~new_n3219_;
  assign new_n3222_ = ~new_n3220_ & ~new_n3221_;
  assign new_n3223_ = ~B8054 & ~new_n2340_;
  assign new_n3224_ = ~new_n2336_ & ~new_n3223_;
  assign new_n3225_ = ~B8087 & ~new_n2350_;
  assign new_n3226_ = ~new_n2346_ & ~new_n3225_;
  assign new_n3227_ = new_n3222_ & ~new_n3226_;
  assign new_n3228_ = ~B8120 & ~new_n2361_;
  assign new_n3229_ = ~new_n2357_ & ~new_n3228_;
  assign new_n3230_ = ~new_n3226_ & ~new_n3229_;
  assign new_n3231_ = ~new_n3227_ & ~new_n3230_;
  assign new_n3232_ = new_n3224_ & new_n3231_;
  assign new_n3233_ = ~new_n3224_ & ~new_n3231_;
  assign new_n3234_ = ~new_n3232_ & ~new_n3233_;
  assign new_n3235_ = ~new_n3222_ & ~new_n3234_;
  assign new_n3236_ = ~B8153 & ~new_n2377_;
  assign new_n3237_ = ~new_n2373_ & ~new_n3236_;
  assign new_n3238_ = ~B8186 & ~new_n2387_;
  assign new_n3239_ = ~new_n2383_ & ~new_n3238_;
  assign new_n3240_ = ~new_n3237_ & new_n3239_;
  assign new_n3241_ = new_n3237_ & ~new_n3239_;
  assign new_n3242_ = ~new_n3240_ & ~new_n3241_;
  assign new_n3243_ = ~B8219 & ~new_n2400_;
  assign new_n3244_ = ~new_n2396_ & ~new_n3243_;
  assign new_n3245_ = ~B8252 & ~new_n2410_;
  assign new_n3246_ = ~new_n2406_ & ~new_n3245_;
  assign new_n3247_ = new_n3242_ & ~new_n3246_;
  assign new_n3248_ = ~B8285 & ~new_n2421_;
  assign new_n3249_ = ~new_n2417_ & ~new_n3248_;
  assign new_n3250_ = ~new_n3246_ & ~new_n3249_;
  assign new_n3251_ = ~new_n3247_ & ~new_n3250_;
  assign new_n3252_ = new_n3244_ & new_n3251_;
  assign new_n3253_ = ~new_n3244_ & ~new_n3251_;
  assign new_n3254_ = ~new_n3252_ & ~new_n3253_;
  assign new_n3255_ = ~new_n3242_ & ~new_n3254_;
  assign new_n3256_ = new_n3215_ & ~new_n3255_;
  assign new_n3257_ = ~B8318 & ~new_n2438_;
  assign new_n3258_ = ~new_n2434_ & ~new_n3257_;
  assign new_n3259_ = ~B8351 & ~new_n2448_;
  assign new_n3260_ = ~new_n2444_ & ~new_n3259_;
  assign new_n3261_ = ~new_n3258_ & new_n3260_;
  assign new_n3262_ = new_n3258_ & ~new_n3260_;
  assign new_n3263_ = ~new_n3261_ & ~new_n3262_;
  assign new_n3264_ = ~B8384 & ~new_n2461_;
  assign new_n3265_ = ~new_n2457_ & ~new_n3264_;
  assign new_n3266_ = ~B8417 & ~new_n2471_;
  assign new_n3267_ = ~new_n2467_ & ~new_n3266_;
  assign new_n3268_ = new_n3263_ & ~new_n3267_;
  assign new_n3269_ = ~B8450 & ~new_n2482_;
  assign new_n3270_ = ~new_n2478_ & ~new_n3269_;
  assign new_n3271_ = ~new_n3267_ & ~new_n3270_;
  assign new_n3272_ = ~new_n3268_ & ~new_n3271_;
  assign new_n3273_ = new_n3265_ & new_n3272_;
  assign new_n3274_ = ~new_n3265_ & ~new_n3272_;
  assign new_n3275_ = ~new_n3273_ & ~new_n3274_;
  assign new_n3276_ = ~new_n3263_ & ~new_n3275_;
  assign new_n3277_ = ~new_n3255_ & ~new_n3276_;
  assign new_n3278_ = ~new_n3256_ & ~new_n3277_;
  assign new_n3279_ = new_n3235_ & new_n3278_;
  assign new_n3280_ = ~new_n3235_ & ~new_n3278_;
  assign new_n3281_ = ~new_n3279_ & ~new_n3280_;
  assign new_n3282_ = ~new_n3215_ & ~new_n3281_;
  assign new_n3283_ = new_n3062_ & ~new_n3282_;
  assign new_n3284_ = ~B8483 & ~new_n2505_;
  assign new_n3285_ = ~new_n2501_ & ~new_n3284_;
  assign new_n3286_ = ~B8516 & ~new_n2515_;
  assign new_n3287_ = ~new_n2511_ & ~new_n3286_;
  assign new_n3288_ = ~new_n3285_ & new_n3287_;
  assign new_n3289_ = new_n3285_ & ~new_n3287_;
  assign new_n3290_ = ~new_n3288_ & ~new_n3289_;
  assign new_n3291_ = ~B8549 & ~new_n2528_;
  assign new_n3292_ = ~new_n2524_ & ~new_n3291_;
  assign new_n3293_ = ~B8582 & ~new_n2538_;
  assign new_n3294_ = ~new_n2534_ & ~new_n3293_;
  assign new_n3295_ = new_n3290_ & ~new_n3294_;
  assign new_n3296_ = ~B8615 & ~new_n2549_;
  assign new_n3297_ = ~new_n2545_ & ~new_n3296_;
  assign new_n3298_ = ~new_n3294_ & ~new_n3297_;
  assign new_n3299_ = ~new_n3295_ & ~new_n3298_;
  assign new_n3300_ = new_n3292_ & new_n3299_;
  assign new_n3301_ = ~new_n3292_ & ~new_n3299_;
  assign new_n3302_ = ~new_n3300_ & ~new_n3301_;
  assign new_n3303_ = ~new_n3290_ & ~new_n3302_;
  assign new_n3304_ = ~B8648 & ~new_n2565_;
  assign new_n3305_ = ~new_n2561_ & ~new_n3304_;
  assign new_n3306_ = ~B8681 & ~new_n2575_;
  assign new_n3307_ = ~new_n2571_ & ~new_n3306_;
  assign new_n3308_ = ~new_n3305_ & new_n3307_;
  assign new_n3309_ = new_n3305_ & ~new_n3307_;
  assign new_n3310_ = ~new_n3308_ & ~new_n3309_;
  assign new_n3311_ = ~B8714 & ~new_n2588_;
  assign new_n3312_ = ~new_n2584_ & ~new_n3311_;
  assign new_n3313_ = ~B8747 & ~new_n2598_;
  assign new_n3314_ = ~new_n2594_ & ~new_n3313_;
  assign new_n3315_ = new_n3310_ & ~new_n3314_;
  assign new_n3316_ = ~B8780 & ~new_n2609_;
  assign new_n3317_ = ~new_n2605_ & ~new_n3316_;
  assign new_n3318_ = ~new_n3314_ & ~new_n3317_;
  assign new_n3319_ = ~new_n3315_ & ~new_n3318_;
  assign new_n3320_ = new_n3312_ & new_n3319_;
  assign new_n3321_ = ~new_n3312_ & ~new_n3319_;
  assign new_n3322_ = ~new_n3320_ & ~new_n3321_;
  assign new_n3323_ = ~new_n3310_ & ~new_n3322_;
  assign new_n3324_ = ~new_n3303_ & new_n3323_;
  assign new_n3325_ = new_n3303_ & ~new_n3323_;
  assign new_n3326_ = ~new_n3324_ & ~new_n3325_;
  assign new_n3327_ = ~B8813 & ~new_n2628_;
  assign new_n3328_ = ~new_n2624_ & ~new_n3327_;
  assign new_n3329_ = ~B8846 & ~new_n2638_;
  assign new_n3330_ = ~new_n2634_ & ~new_n3329_;
  assign new_n3331_ = ~new_n3328_ & new_n3330_;
  assign new_n3332_ = new_n3328_ & ~new_n3330_;
  assign new_n3333_ = ~new_n3331_ & ~new_n3332_;
  assign new_n3334_ = ~B8879 & ~new_n2651_;
  assign new_n3335_ = ~new_n2647_ & ~new_n3334_;
  assign new_n3336_ = ~B8912 & ~new_n2661_;
  assign new_n3337_ = ~new_n2657_ & ~new_n3336_;
  assign new_n3338_ = new_n3333_ & ~new_n3337_;
  assign new_n3339_ = ~B8945 & ~new_n2672_;
  assign new_n3340_ = ~new_n2668_ & ~new_n3339_;
  assign new_n3341_ = ~new_n3337_ & ~new_n3340_;
  assign new_n3342_ = ~new_n3338_ & ~new_n3341_;
  assign new_n3343_ = new_n3335_ & new_n3342_;
  assign new_n3344_ = ~new_n3335_ & ~new_n3342_;
  assign new_n3345_ = ~new_n3343_ & ~new_n3344_;
  assign new_n3346_ = ~new_n3333_ & ~new_n3345_;
  assign new_n3347_ = ~B8978 & ~new_n2688_;
  assign new_n3348_ = ~new_n2684_ & ~new_n3347_;
  assign new_n3349_ = ~B9011 & ~new_n2698_;
  assign new_n3350_ = ~new_n2694_ & ~new_n3349_;
  assign new_n3351_ = ~new_n3348_ & new_n3350_;
  assign new_n3352_ = new_n3348_ & ~new_n3350_;
  assign new_n3353_ = ~new_n3351_ & ~new_n3352_;
  assign new_n3354_ = ~B9044 & ~new_n2711_;
  assign new_n3355_ = ~new_n2707_ & ~new_n3354_;
  assign new_n3356_ = ~B9077 & ~new_n2721_;
  assign new_n3357_ = ~new_n2717_ & ~new_n3356_;
  assign new_n3358_ = new_n3353_ & ~new_n3357_;
  assign new_n3359_ = ~B9110 & ~new_n2732_;
  assign new_n3360_ = ~new_n2728_ & ~new_n3359_;
  assign new_n3361_ = ~new_n3357_ & ~new_n3360_;
  assign new_n3362_ = ~new_n3358_ & ~new_n3361_;
  assign new_n3363_ = new_n3355_ & new_n3362_;
  assign new_n3364_ = ~new_n3355_ & ~new_n3362_;
  assign new_n3365_ = ~new_n3363_ & ~new_n3364_;
  assign new_n3366_ = ~new_n3353_ & ~new_n3365_;
  assign new_n3367_ = new_n3326_ & ~new_n3366_;
  assign new_n3368_ = ~B9143 & ~new_n2749_;
  assign new_n3369_ = ~new_n2745_ & ~new_n3368_;
  assign new_n3370_ = ~B9176 & ~new_n2759_;
  assign new_n3371_ = ~new_n2755_ & ~new_n3370_;
  assign new_n3372_ = ~new_n3369_ & new_n3371_;
  assign new_n3373_ = new_n3369_ & ~new_n3371_;
  assign new_n3374_ = ~new_n3372_ & ~new_n3373_;
  assign new_n3375_ = ~B9209 & ~new_n2772_;
  assign new_n3376_ = ~new_n2768_ & ~new_n3375_;
  assign new_n3377_ = ~B9242 & ~new_n2782_;
  assign new_n3378_ = ~new_n2778_ & ~new_n3377_;
  assign new_n3379_ = new_n3374_ & ~new_n3378_;
  assign new_n3380_ = ~B9275 & ~new_n2793_;
  assign new_n3381_ = ~new_n2789_ & ~new_n3380_;
  assign new_n3382_ = ~new_n3378_ & ~new_n3381_;
  assign new_n3383_ = ~new_n3379_ & ~new_n3382_;
  assign new_n3384_ = new_n3376_ & new_n3383_;
  assign new_n3385_ = ~new_n3376_ & ~new_n3383_;
  assign new_n3386_ = ~new_n3384_ & ~new_n3385_;
  assign new_n3387_ = ~new_n3374_ & ~new_n3386_;
  assign new_n3388_ = ~new_n3366_ & ~new_n3387_;
  assign new_n3389_ = ~new_n3367_ & ~new_n3388_;
  assign new_n3390_ = new_n3346_ & new_n3389_;
  assign new_n3391_ = ~new_n3346_ & ~new_n3389_;
  assign new_n3392_ = ~new_n3390_ & ~new_n3391_;
  assign new_n3393_ = ~new_n3326_ & ~new_n3392_;
  assign new_n3394_ = ~new_n3282_ & ~new_n3393_;
  assign new_n3395_ = ~new_n3283_ & ~new_n3394_;
  assign new_n3396_ = new_n3172_ & new_n3395_;
  assign new_n3397_ = ~new_n3172_ & ~new_n3395_;
  assign new_n3398_ = ~new_n3396_ & ~new_n3397_;
  assign A6874 = ~new_n3062_ & ~new_n3398_;
  assign new_n3400_ = ~new_n3059_ & ~new_n3396_;
  assign A6873 = ~new_n3062_ & ~new_n3400_;
  assign new_n3402_ = new_n3059_ & new_n3172_;
  assign new_n3403_ = ~new_n3062_ & ~new_n3402_;
  assign new_n3404_ = new_n3062_ & ~new_n3403_;
  assign new_n3405_ = new_n3062_ & new_n3402_;
  assign new_n3406_ = new_n3404_ & ~new_n3405_;
  assign new_n3407_ = new_n3172_ & ~new_n3406_;
  assign A6872 = new_n3395_ | new_n3407_;
  assign new_n3409_ = new_n3282_ & new_n3393_;
  assign new_n3410_ = ~new_n3394_ & ~new_n3409_;
  assign new_n3411_ = ~new_n3062_ & ~new_n3282_;
  assign new_n3412_ = new_n3062_ & new_n3282_;
  assign new_n3413_ = ~new_n3411_ & ~new_n3412_;
  assign new_n3414_ = new_n3410_ & ~new_n3413_;
  assign A6871 = new_n3407_ | new_n3414_;
  assign new_n3416_ = new_n3172_ & ~new_n3414_;
  assign new_n3417_ = ~new_n3172_ & new_n3414_;
  assign new_n3418_ = ~new_n3416_ & ~new_n3417_;
  assign A6870 = ~new_n3062_ & ~new_n3418_;
  assign new_n3420_ = ~B5185 & new_n1256_;
  assign new_n3421_ = ~new_n1252_ & ~new_n3420_;
  assign new_n3422_ = ~new_n2840_ & ~new_n3421_;
  assign new_n3423_ = B5217 & B5216;
  assign new_n3424_ = ~new_n1267_ & ~new_n3423_;
  assign new_n3425_ = new_n1267_ & ~new_n3424_;
  assign new_n3426_ = new_n1267_ & new_n3423_;
  assign new_n3427_ = new_n3425_ & ~new_n3426_;
  assign new_n3428_ = B5217 & ~new_n3427_;
  assign new_n3429_ = ~new_n1270_ & ~new_n3428_;
  assign new_n3430_ = new_n3422_ & ~new_n3429_;
  assign new_n3431_ = ~new_n3422_ & new_n3429_;
  assign new_n3432_ = ~new_n3430_ & ~new_n3431_;
  assign new_n3433_ = B5250 & B5249;
  assign new_n3434_ = ~new_n1280_ & ~new_n3433_;
  assign new_n3435_ = new_n1280_ & ~new_n3434_;
  assign new_n3436_ = new_n1280_ & new_n3433_;
  assign new_n3437_ = new_n3435_ & ~new_n3436_;
  assign new_n3438_ = B5250 & ~new_n3437_;
  assign new_n3439_ = ~new_n1283_ & ~new_n3438_;
  assign new_n3440_ = B5283 & B5282;
  assign new_n3441_ = ~new_n1290_ & ~new_n3440_;
  assign new_n3442_ = new_n1290_ & ~new_n3441_;
  assign new_n3443_ = new_n1290_ & new_n3440_;
  assign new_n3444_ = new_n3442_ & ~new_n3443_;
  assign new_n3445_ = B5283 & ~new_n3444_;
  assign new_n3446_ = ~new_n1293_ & ~new_n3445_;
  assign new_n3447_ = new_n3432_ & new_n3446_;
  assign new_n3448_ = B5316 & B5315;
  assign new_n3449_ = ~new_n1301_ & ~new_n3448_;
  assign new_n3450_ = new_n1301_ & ~new_n3449_;
  assign new_n3451_ = new_n1301_ & new_n3448_;
  assign new_n3452_ = new_n3450_ & ~new_n3451_;
  assign new_n3453_ = B5316 & ~new_n3452_;
  assign new_n3454_ = ~new_n1304_ & ~new_n3453_;
  assign new_n3455_ = new_n3446_ & new_n3454_;
  assign new_n3456_ = ~new_n3447_ & ~new_n3455_;
  assign new_n3457_ = ~new_n3439_ & new_n3456_;
  assign new_n3458_ = new_n3439_ & ~new_n3456_;
  assign new_n3459_ = ~new_n3457_ & ~new_n3458_;
  assign new_n3460_ = ~new_n3432_ & ~new_n3459_;
  assign new_n3461_ = B5349 & B5348;
  assign new_n3462_ = ~new_n1317_ & ~new_n3461_;
  assign new_n3463_ = new_n1317_ & ~new_n3462_;
  assign new_n3464_ = new_n1317_ & new_n3461_;
  assign new_n3465_ = new_n3463_ & ~new_n3464_;
  assign new_n3466_ = B5349 & ~new_n3465_;
  assign new_n3467_ = ~new_n1320_ & ~new_n3466_;
  assign new_n3468_ = B5382 & B5381;
  assign new_n3469_ = ~new_n1327_ & ~new_n3468_;
  assign new_n3470_ = new_n1327_ & ~new_n3469_;
  assign new_n3471_ = new_n1327_ & new_n3468_;
  assign new_n3472_ = new_n3470_ & ~new_n3471_;
  assign new_n3473_ = B5382 & ~new_n3472_;
  assign new_n3474_ = ~new_n1330_ & ~new_n3473_;
  assign new_n3475_ = new_n3467_ & ~new_n3474_;
  assign new_n3476_ = ~new_n3467_ & new_n3474_;
  assign new_n3477_ = ~new_n3475_ & ~new_n3476_;
  assign new_n3478_ = B5415 & B5414;
  assign new_n3479_ = ~new_n1340_ & ~new_n3478_;
  assign new_n3480_ = new_n1340_ & ~new_n3479_;
  assign new_n3481_ = new_n1340_ & new_n3478_;
  assign new_n3482_ = new_n3480_ & ~new_n3481_;
  assign new_n3483_ = B5415 & ~new_n3482_;
  assign new_n3484_ = ~new_n1343_ & ~new_n3483_;
  assign new_n3485_ = B5448 & B5447;
  assign new_n3486_ = ~new_n1350_ & ~new_n3485_;
  assign new_n3487_ = new_n1350_ & ~new_n3486_;
  assign new_n3488_ = new_n1350_ & new_n3485_;
  assign new_n3489_ = new_n3487_ & ~new_n3488_;
  assign new_n3490_ = B5448 & ~new_n3489_;
  assign new_n3491_ = ~new_n1353_ & ~new_n3490_;
  assign new_n3492_ = new_n3477_ & new_n3491_;
  assign new_n3493_ = B5481 & B5480;
  assign new_n3494_ = ~new_n1361_ & ~new_n3493_;
  assign new_n3495_ = new_n1361_ & ~new_n3494_;
  assign new_n3496_ = new_n1361_ & new_n3493_;
  assign new_n3497_ = new_n3495_ & ~new_n3496_;
  assign new_n3498_ = B5481 & ~new_n3497_;
  assign new_n3499_ = ~new_n1364_ & ~new_n3498_;
  assign new_n3500_ = new_n3491_ & new_n3499_;
  assign new_n3501_ = ~new_n3492_ & ~new_n3500_;
  assign new_n3502_ = ~new_n3484_ & new_n3501_;
  assign new_n3503_ = new_n3484_ & ~new_n3501_;
  assign new_n3504_ = ~new_n3502_ & ~new_n3503_;
  assign new_n3505_ = ~new_n3477_ & ~new_n3504_;
  assign new_n3506_ = ~new_n3460_ & new_n3505_;
  assign new_n3507_ = new_n3460_ & ~new_n3505_;
  assign new_n3508_ = ~new_n3506_ & ~new_n3507_;
  assign new_n3509_ = B5514 & B5513;
  assign new_n3510_ = ~new_n1380_ & ~new_n3509_;
  assign new_n3511_ = new_n1380_ & ~new_n3510_;
  assign new_n3512_ = new_n1380_ & new_n3509_;
  assign new_n3513_ = new_n3511_ & ~new_n3512_;
  assign new_n3514_ = B5514 & ~new_n3513_;
  assign new_n3515_ = ~new_n1383_ & ~new_n3514_;
  assign new_n3516_ = B5547 & B5546;
  assign new_n3517_ = ~new_n1390_ & ~new_n3516_;
  assign new_n3518_ = new_n1390_ & ~new_n3517_;
  assign new_n3519_ = new_n1390_ & new_n3516_;
  assign new_n3520_ = new_n3518_ & ~new_n3519_;
  assign new_n3521_ = B5547 & ~new_n3520_;
  assign new_n3522_ = ~new_n1393_ & ~new_n3521_;
  assign new_n3523_ = new_n3515_ & ~new_n3522_;
  assign new_n3524_ = ~new_n3515_ & new_n3522_;
  assign new_n3525_ = ~new_n3523_ & ~new_n3524_;
  assign new_n3526_ = B5580 & B5579;
  assign new_n3527_ = ~new_n1403_ & ~new_n3526_;
  assign new_n3528_ = new_n1403_ & ~new_n3527_;
  assign new_n3529_ = new_n1403_ & new_n3526_;
  assign new_n3530_ = new_n3528_ & ~new_n3529_;
  assign new_n3531_ = B5580 & ~new_n3530_;
  assign new_n3532_ = ~new_n1406_ & ~new_n3531_;
  assign new_n3533_ = B5613 & B5612;
  assign new_n3534_ = ~new_n1413_ & ~new_n3533_;
  assign new_n3535_ = new_n1413_ & ~new_n3534_;
  assign new_n3536_ = new_n1413_ & new_n3533_;
  assign new_n3537_ = new_n3535_ & ~new_n3536_;
  assign new_n3538_ = B5613 & ~new_n3537_;
  assign new_n3539_ = ~new_n1416_ & ~new_n3538_;
  assign new_n3540_ = new_n3525_ & new_n3539_;
  assign new_n3541_ = B5646 & B5645;
  assign new_n3542_ = ~new_n1424_ & ~new_n3541_;
  assign new_n3543_ = new_n1424_ & ~new_n3542_;
  assign new_n3544_ = new_n1424_ & new_n3541_;
  assign new_n3545_ = new_n3543_ & ~new_n3544_;
  assign new_n3546_ = B5646 & ~new_n3545_;
  assign new_n3547_ = ~new_n1427_ & ~new_n3546_;
  assign new_n3548_ = new_n3539_ & new_n3547_;
  assign new_n3549_ = ~new_n3540_ & ~new_n3548_;
  assign new_n3550_ = ~new_n3532_ & new_n3549_;
  assign new_n3551_ = new_n3532_ & ~new_n3549_;
  assign new_n3552_ = ~new_n3550_ & ~new_n3551_;
  assign new_n3553_ = ~new_n3525_ & ~new_n3552_;
  assign new_n3554_ = B5679 & B5678;
  assign new_n3555_ = ~new_n1440_ & ~new_n3554_;
  assign new_n3556_ = new_n1440_ & ~new_n3555_;
  assign new_n3557_ = new_n1440_ & new_n3554_;
  assign new_n3558_ = new_n3556_ & ~new_n3557_;
  assign new_n3559_ = B5679 & ~new_n3558_;
  assign new_n3560_ = ~new_n1443_ & ~new_n3559_;
  assign new_n3561_ = B5712 & B5711;
  assign new_n3562_ = ~new_n1450_ & ~new_n3561_;
  assign new_n3563_ = new_n1450_ & ~new_n3562_;
  assign new_n3564_ = new_n1450_ & new_n3561_;
  assign new_n3565_ = new_n3563_ & ~new_n3564_;
  assign new_n3566_ = B5712 & ~new_n3565_;
  assign new_n3567_ = ~new_n1453_ & ~new_n3566_;
  assign new_n3568_ = new_n3560_ & ~new_n3567_;
  assign new_n3569_ = ~new_n3560_ & new_n3567_;
  assign new_n3570_ = ~new_n3568_ & ~new_n3569_;
  assign new_n3571_ = B5745 & B5744;
  assign new_n3572_ = ~new_n1463_ & ~new_n3571_;
  assign new_n3573_ = new_n1463_ & ~new_n3572_;
  assign new_n3574_ = new_n1463_ & new_n3571_;
  assign new_n3575_ = new_n3573_ & ~new_n3574_;
  assign new_n3576_ = B5745 & ~new_n3575_;
  assign new_n3577_ = ~new_n1466_ & ~new_n3576_;
  assign new_n3578_ = B5778 & B5777;
  assign new_n3579_ = ~new_n1473_ & ~new_n3578_;
  assign new_n3580_ = new_n1473_ & ~new_n3579_;
  assign new_n3581_ = new_n1473_ & new_n3578_;
  assign new_n3582_ = new_n3580_ & ~new_n3581_;
  assign new_n3583_ = B5778 & ~new_n3582_;
  assign new_n3584_ = ~new_n1476_ & ~new_n3583_;
  assign new_n3585_ = new_n3570_ & new_n3584_;
  assign new_n3586_ = B5811 & B5810;
  assign new_n3587_ = ~new_n1484_ & ~new_n3586_;
  assign new_n3588_ = new_n1484_ & ~new_n3587_;
  assign new_n3589_ = new_n1484_ & new_n3586_;
  assign new_n3590_ = new_n3588_ & ~new_n3589_;
  assign new_n3591_ = B5811 & ~new_n3590_;
  assign new_n3592_ = ~new_n1487_ & ~new_n3591_;
  assign new_n3593_ = new_n3584_ & new_n3592_;
  assign new_n3594_ = ~new_n3585_ & ~new_n3593_;
  assign new_n3595_ = ~new_n3577_ & new_n3594_;
  assign new_n3596_ = new_n3577_ & ~new_n3594_;
  assign new_n3597_ = ~new_n3595_ & ~new_n3596_;
  assign new_n3598_ = ~new_n3570_ & ~new_n3597_;
  assign new_n3599_ = new_n3508_ & ~new_n3598_;
  assign new_n3600_ = B5844 & B5843;
  assign new_n3601_ = ~new_n1501_ & ~new_n3600_;
  assign new_n3602_ = new_n1501_ & ~new_n3601_;
  assign new_n3603_ = new_n1501_ & new_n3600_;
  assign new_n3604_ = new_n3602_ & ~new_n3603_;
  assign new_n3605_ = B5844 & ~new_n3604_;
  assign new_n3606_ = ~new_n1504_ & ~new_n3605_;
  assign new_n3607_ = B5877 & B5876;
  assign new_n3608_ = ~new_n1511_ & ~new_n3607_;
  assign new_n3609_ = new_n1511_ & ~new_n3608_;
  assign new_n3610_ = new_n1511_ & new_n3607_;
  assign new_n3611_ = new_n3609_ & ~new_n3610_;
  assign new_n3612_ = B5877 & ~new_n3611_;
  assign new_n3613_ = ~new_n1514_ & ~new_n3612_;
  assign new_n3614_ = new_n3606_ & ~new_n3613_;
  assign new_n3615_ = ~new_n3606_ & new_n3613_;
  assign new_n3616_ = ~new_n3614_ & ~new_n3615_;
  assign new_n3617_ = B5910 & B5909;
  assign new_n3618_ = ~new_n1524_ & ~new_n3617_;
  assign new_n3619_ = new_n1524_ & ~new_n3618_;
  assign new_n3620_ = new_n1524_ & new_n3617_;
  assign new_n3621_ = new_n3619_ & ~new_n3620_;
  assign new_n3622_ = B5910 & ~new_n3621_;
  assign new_n3623_ = ~new_n1527_ & ~new_n3622_;
  assign new_n3624_ = B5943 & B5942;
  assign new_n3625_ = ~new_n1534_ & ~new_n3624_;
  assign new_n3626_ = new_n1534_ & ~new_n3625_;
  assign new_n3627_ = new_n1534_ & new_n3624_;
  assign new_n3628_ = new_n3626_ & ~new_n3627_;
  assign new_n3629_ = B5943 & ~new_n3628_;
  assign new_n3630_ = ~new_n1537_ & ~new_n3629_;
  assign new_n3631_ = new_n3616_ & new_n3630_;
  assign new_n3632_ = B5976 & B5975;
  assign new_n3633_ = ~new_n1545_ & ~new_n3632_;
  assign new_n3634_ = new_n1545_ & ~new_n3633_;
  assign new_n3635_ = new_n1545_ & new_n3632_;
  assign new_n3636_ = new_n3634_ & ~new_n3635_;
  assign new_n3637_ = B5976 & ~new_n3636_;
  assign new_n3638_ = ~new_n1548_ & ~new_n3637_;
  assign new_n3639_ = new_n3630_ & new_n3638_;
  assign new_n3640_ = ~new_n3631_ & ~new_n3639_;
  assign new_n3641_ = ~new_n3623_ & new_n3640_;
  assign new_n3642_ = new_n3623_ & ~new_n3640_;
  assign new_n3643_ = ~new_n3641_ & ~new_n3642_;
  assign new_n3644_ = ~new_n3616_ & ~new_n3643_;
  assign new_n3645_ = ~new_n3598_ & ~new_n3644_;
  assign new_n3646_ = ~new_n3599_ & ~new_n3645_;
  assign new_n3647_ = new_n3553_ & new_n3646_;
  assign new_n3648_ = ~new_n3553_ & ~new_n3646_;
  assign new_n3649_ = ~new_n3647_ & ~new_n3648_;
  assign new_n3650_ = ~new_n3508_ & ~new_n3649_;
  assign new_n3651_ = B6009 & B6008;
  assign new_n3652_ = ~new_n1567_ & ~new_n3651_;
  assign new_n3653_ = new_n1567_ & ~new_n3652_;
  assign new_n3654_ = new_n1567_ & new_n3651_;
  assign new_n3655_ = new_n3653_ & ~new_n3654_;
  assign new_n3656_ = B6009 & ~new_n3655_;
  assign new_n3657_ = ~new_n1570_ & ~new_n3656_;
  assign new_n3658_ = B6042 & B6041;
  assign new_n3659_ = ~new_n1577_ & ~new_n3658_;
  assign new_n3660_ = new_n1577_ & ~new_n3659_;
  assign new_n3661_ = new_n1577_ & new_n3658_;
  assign new_n3662_ = new_n3660_ & ~new_n3661_;
  assign new_n3663_ = B6042 & ~new_n3662_;
  assign new_n3664_ = ~new_n1580_ & ~new_n3663_;
  assign new_n3665_ = new_n3657_ & ~new_n3664_;
  assign new_n3666_ = ~new_n3657_ & new_n3664_;
  assign new_n3667_ = ~new_n3665_ & ~new_n3666_;
  assign new_n3668_ = B6075 & B6074;
  assign new_n3669_ = ~new_n1590_ & ~new_n3668_;
  assign new_n3670_ = new_n1590_ & ~new_n3669_;
  assign new_n3671_ = new_n1590_ & new_n3668_;
  assign new_n3672_ = new_n3670_ & ~new_n3671_;
  assign new_n3673_ = B6075 & ~new_n3672_;
  assign new_n3674_ = ~new_n1593_ & ~new_n3673_;
  assign new_n3675_ = B6108 & B6107;
  assign new_n3676_ = ~new_n1600_ & ~new_n3675_;
  assign new_n3677_ = new_n1600_ & ~new_n3676_;
  assign new_n3678_ = new_n1600_ & new_n3675_;
  assign new_n3679_ = new_n3677_ & ~new_n3678_;
  assign new_n3680_ = B6108 & ~new_n3679_;
  assign new_n3681_ = ~new_n1603_ & ~new_n3680_;
  assign new_n3682_ = new_n3667_ & new_n3681_;
  assign new_n3683_ = B6141 & B6140;
  assign new_n3684_ = ~new_n1611_ & ~new_n3683_;
  assign new_n3685_ = new_n1611_ & ~new_n3684_;
  assign new_n3686_ = new_n1611_ & new_n3683_;
  assign new_n3687_ = new_n3685_ & ~new_n3686_;
  assign new_n3688_ = B6141 & ~new_n3687_;
  assign new_n3689_ = ~new_n1614_ & ~new_n3688_;
  assign new_n3690_ = new_n3681_ & new_n3689_;
  assign new_n3691_ = ~new_n3682_ & ~new_n3690_;
  assign new_n3692_ = ~new_n3674_ & new_n3691_;
  assign new_n3693_ = new_n3674_ & ~new_n3691_;
  assign new_n3694_ = ~new_n3692_ & ~new_n3693_;
  assign new_n3695_ = ~new_n3667_ & ~new_n3694_;
  assign new_n3696_ = B6174 & B6173;
  assign new_n3697_ = ~new_n1627_ & ~new_n3696_;
  assign new_n3698_ = new_n1627_ & ~new_n3697_;
  assign new_n3699_ = new_n1627_ & new_n3696_;
  assign new_n3700_ = new_n3698_ & ~new_n3699_;
  assign new_n3701_ = B6174 & ~new_n3700_;
  assign new_n3702_ = ~new_n1630_ & ~new_n3701_;
  assign new_n3703_ = B6207 & B6206;
  assign new_n3704_ = ~new_n1637_ & ~new_n3703_;
  assign new_n3705_ = new_n1637_ & ~new_n3704_;
  assign new_n3706_ = new_n1637_ & new_n3703_;
  assign new_n3707_ = new_n3705_ & ~new_n3706_;
  assign new_n3708_ = B6207 & ~new_n3707_;
  assign new_n3709_ = ~new_n1640_ & ~new_n3708_;
  assign new_n3710_ = new_n3702_ & ~new_n3709_;
  assign new_n3711_ = ~new_n3702_ & new_n3709_;
  assign new_n3712_ = ~new_n3710_ & ~new_n3711_;
  assign new_n3713_ = B6240 & B6239;
  assign new_n3714_ = ~new_n1650_ & ~new_n3713_;
  assign new_n3715_ = new_n1650_ & ~new_n3714_;
  assign new_n3716_ = new_n1650_ & new_n3713_;
  assign new_n3717_ = new_n3715_ & ~new_n3716_;
  assign new_n3718_ = B6240 & ~new_n3717_;
  assign new_n3719_ = ~new_n1653_ & ~new_n3718_;
  assign new_n3720_ = B6273 & B6272;
  assign new_n3721_ = ~new_n1660_ & ~new_n3720_;
  assign new_n3722_ = new_n1660_ & ~new_n3721_;
  assign new_n3723_ = new_n1660_ & new_n3720_;
  assign new_n3724_ = new_n3722_ & ~new_n3723_;
  assign new_n3725_ = B6273 & ~new_n3724_;
  assign new_n3726_ = ~new_n1663_ & ~new_n3725_;
  assign new_n3727_ = new_n3712_ & new_n3726_;
  assign new_n3728_ = B6306 & B6305;
  assign new_n3729_ = ~new_n1671_ & ~new_n3728_;
  assign new_n3730_ = new_n1671_ & ~new_n3729_;
  assign new_n3731_ = new_n1671_ & new_n3728_;
  assign new_n3732_ = new_n3730_ & ~new_n3731_;
  assign new_n3733_ = B6306 & ~new_n3732_;
  assign new_n3734_ = ~new_n1674_ & ~new_n3733_;
  assign new_n3735_ = new_n3726_ & new_n3734_;
  assign new_n3736_ = ~new_n3727_ & ~new_n3735_;
  assign new_n3737_ = ~new_n3719_ & new_n3736_;
  assign new_n3738_ = new_n3719_ & ~new_n3736_;
  assign new_n3739_ = ~new_n3737_ & ~new_n3738_;
  assign new_n3740_ = ~new_n3712_ & ~new_n3739_;
  assign new_n3741_ = ~new_n3695_ & new_n3740_;
  assign new_n3742_ = new_n3695_ & ~new_n3740_;
  assign new_n3743_ = ~new_n3741_ & ~new_n3742_;
  assign new_n3744_ = B6339 & B6338;
  assign new_n3745_ = ~new_n1690_ & ~new_n3744_;
  assign new_n3746_ = new_n1690_ & ~new_n3745_;
  assign new_n3747_ = new_n1690_ & new_n3744_;
  assign new_n3748_ = new_n3746_ & ~new_n3747_;
  assign new_n3749_ = B6339 & ~new_n3748_;
  assign new_n3750_ = ~new_n1693_ & ~new_n3749_;
  assign new_n3751_ = B6372 & B6371;
  assign new_n3752_ = ~new_n1700_ & ~new_n3751_;
  assign new_n3753_ = new_n1700_ & ~new_n3752_;
  assign new_n3754_ = new_n1700_ & new_n3751_;
  assign new_n3755_ = new_n3753_ & ~new_n3754_;
  assign new_n3756_ = B6372 & ~new_n3755_;
  assign new_n3757_ = ~new_n1703_ & ~new_n3756_;
  assign new_n3758_ = new_n3750_ & ~new_n3757_;
  assign new_n3759_ = ~new_n3750_ & new_n3757_;
  assign new_n3760_ = ~new_n3758_ & ~new_n3759_;
  assign new_n3761_ = B6405 & B6404;
  assign new_n3762_ = ~new_n1713_ & ~new_n3761_;
  assign new_n3763_ = new_n1713_ & ~new_n3762_;
  assign new_n3764_ = new_n1713_ & new_n3761_;
  assign new_n3765_ = new_n3763_ & ~new_n3764_;
  assign new_n3766_ = B6405 & ~new_n3765_;
  assign new_n3767_ = ~new_n1716_ & ~new_n3766_;
  assign new_n3768_ = B6438 & B6437;
  assign new_n3769_ = ~new_n1723_ & ~new_n3768_;
  assign new_n3770_ = new_n1723_ & ~new_n3769_;
  assign new_n3771_ = new_n1723_ & new_n3768_;
  assign new_n3772_ = new_n3770_ & ~new_n3771_;
  assign new_n3773_ = B6438 & ~new_n3772_;
  assign new_n3774_ = ~new_n1726_ & ~new_n3773_;
  assign new_n3775_ = new_n3760_ & new_n3774_;
  assign new_n3776_ = B6471 & B6470;
  assign new_n3777_ = ~new_n1734_ & ~new_n3776_;
  assign new_n3778_ = new_n1734_ & ~new_n3777_;
  assign new_n3779_ = new_n1734_ & new_n3776_;
  assign new_n3780_ = new_n3778_ & ~new_n3779_;
  assign new_n3781_ = B6471 & ~new_n3780_;
  assign new_n3782_ = ~new_n1737_ & ~new_n3781_;
  assign new_n3783_ = new_n3774_ & new_n3782_;
  assign new_n3784_ = ~new_n3775_ & ~new_n3783_;
  assign new_n3785_ = ~new_n3767_ & new_n3784_;
  assign new_n3786_ = new_n3767_ & ~new_n3784_;
  assign new_n3787_ = ~new_n3785_ & ~new_n3786_;
  assign new_n3788_ = ~new_n3760_ & ~new_n3787_;
  assign new_n3789_ = B6504 & B6503;
  assign new_n3790_ = ~new_n1750_ & ~new_n3789_;
  assign new_n3791_ = new_n1750_ & ~new_n3790_;
  assign new_n3792_ = new_n1750_ & new_n3789_;
  assign new_n3793_ = new_n3791_ & ~new_n3792_;
  assign new_n3794_ = B6504 & ~new_n3793_;
  assign new_n3795_ = ~new_n1753_ & ~new_n3794_;
  assign new_n3796_ = B6537 & B6536;
  assign new_n3797_ = ~new_n1760_ & ~new_n3796_;
  assign new_n3798_ = new_n1760_ & ~new_n3797_;
  assign new_n3799_ = new_n1760_ & new_n3796_;
  assign new_n3800_ = new_n3798_ & ~new_n3799_;
  assign new_n3801_ = B6537 & ~new_n3800_;
  assign new_n3802_ = ~new_n1763_ & ~new_n3801_;
  assign new_n3803_ = new_n3795_ & ~new_n3802_;
  assign new_n3804_ = ~new_n3795_ & new_n3802_;
  assign new_n3805_ = ~new_n3803_ & ~new_n3804_;
  assign new_n3806_ = B6570 & B6569;
  assign new_n3807_ = ~new_n1773_ & ~new_n3806_;
  assign new_n3808_ = new_n1773_ & ~new_n3807_;
  assign new_n3809_ = new_n1773_ & new_n3806_;
  assign new_n3810_ = new_n3808_ & ~new_n3809_;
  assign new_n3811_ = B6570 & ~new_n3810_;
  assign new_n3812_ = ~new_n1776_ & ~new_n3811_;
  assign new_n3813_ = B6603 & B6602;
  assign new_n3814_ = ~new_n1783_ & ~new_n3813_;
  assign new_n3815_ = new_n1783_ & ~new_n3814_;
  assign new_n3816_ = new_n1783_ & new_n3813_;
  assign new_n3817_ = new_n3815_ & ~new_n3816_;
  assign new_n3818_ = B6603 & ~new_n3817_;
  assign new_n3819_ = ~new_n1786_ & ~new_n3818_;
  assign new_n3820_ = new_n3805_ & new_n3819_;
  assign new_n3821_ = B6636 & B6635;
  assign new_n3822_ = ~new_n1794_ & ~new_n3821_;
  assign new_n3823_ = new_n1794_ & ~new_n3822_;
  assign new_n3824_ = new_n1794_ & new_n3821_;
  assign new_n3825_ = new_n3823_ & ~new_n3824_;
  assign new_n3826_ = B6636 & ~new_n3825_;
  assign new_n3827_ = ~new_n1797_ & ~new_n3826_;
  assign new_n3828_ = new_n3819_ & new_n3827_;
  assign new_n3829_ = ~new_n3820_ & ~new_n3828_;
  assign new_n3830_ = ~new_n3812_ & new_n3829_;
  assign new_n3831_ = new_n3812_ & ~new_n3829_;
  assign new_n3832_ = ~new_n3830_ & ~new_n3831_;
  assign new_n3833_ = ~new_n3805_ & ~new_n3832_;
  assign new_n3834_ = new_n3743_ & ~new_n3833_;
  assign new_n3835_ = B6669 & B6668;
  assign new_n3836_ = ~new_n1811_ & ~new_n3835_;
  assign new_n3837_ = new_n1811_ & ~new_n3836_;
  assign new_n3838_ = new_n1811_ & new_n3835_;
  assign new_n3839_ = new_n3837_ & ~new_n3838_;
  assign new_n3840_ = B6669 & ~new_n3839_;
  assign new_n3841_ = ~new_n1814_ & ~new_n3840_;
  assign new_n3842_ = B6702 & B6701;
  assign new_n3843_ = ~new_n1821_ & ~new_n3842_;
  assign new_n3844_ = new_n1821_ & ~new_n3843_;
  assign new_n3845_ = new_n1821_ & new_n3842_;
  assign new_n3846_ = new_n3844_ & ~new_n3845_;
  assign new_n3847_ = B6702 & ~new_n3846_;
  assign new_n3848_ = ~new_n1824_ & ~new_n3847_;
  assign new_n3849_ = new_n3841_ & ~new_n3848_;
  assign new_n3850_ = ~new_n3841_ & new_n3848_;
  assign new_n3851_ = ~new_n3849_ & ~new_n3850_;
  assign new_n3852_ = B6735 & B6734;
  assign new_n3853_ = ~new_n1834_ & ~new_n3852_;
  assign new_n3854_ = new_n1834_ & ~new_n3853_;
  assign new_n3855_ = new_n1834_ & new_n3852_;
  assign new_n3856_ = new_n3854_ & ~new_n3855_;
  assign new_n3857_ = B6735 & ~new_n3856_;
  assign new_n3858_ = ~new_n1837_ & ~new_n3857_;
  assign new_n3859_ = B6768 & B6767;
  assign new_n3860_ = ~new_n1844_ & ~new_n3859_;
  assign new_n3861_ = new_n1844_ & ~new_n3860_;
  assign new_n3862_ = new_n1844_ & new_n3859_;
  assign new_n3863_ = new_n3861_ & ~new_n3862_;
  assign new_n3864_ = B6768 & ~new_n3863_;
  assign new_n3865_ = ~new_n1847_ & ~new_n3864_;
  assign new_n3866_ = new_n3851_ & new_n3865_;
  assign new_n3867_ = B6801 & B6800;
  assign new_n3868_ = ~new_n1855_ & ~new_n3867_;
  assign new_n3869_ = new_n1855_ & ~new_n3868_;
  assign new_n3870_ = new_n1855_ & new_n3867_;
  assign new_n3871_ = new_n3869_ & ~new_n3870_;
  assign new_n3872_ = B6801 & ~new_n3871_;
  assign new_n3873_ = ~new_n1858_ & ~new_n3872_;
  assign new_n3874_ = new_n3865_ & new_n3873_;
  assign new_n3875_ = ~new_n3866_ & ~new_n3874_;
  assign new_n3876_ = ~new_n3858_ & new_n3875_;
  assign new_n3877_ = new_n3858_ & ~new_n3875_;
  assign new_n3878_ = ~new_n3876_ & ~new_n3877_;
  assign new_n3879_ = ~new_n3851_ & ~new_n3878_;
  assign new_n3880_ = ~new_n3833_ & ~new_n3879_;
  assign new_n3881_ = ~new_n3834_ & ~new_n3880_;
  assign new_n3882_ = new_n3788_ & new_n3881_;
  assign new_n3883_ = ~new_n3788_ & ~new_n3881_;
  assign new_n3884_ = ~new_n3882_ & ~new_n3883_;
  assign new_n3885_ = ~new_n3743_ & ~new_n3884_;
  assign new_n3886_ = ~new_n3650_ & new_n3885_;
  assign new_n3887_ = new_n3650_ & ~new_n3885_;
  assign new_n3888_ = ~new_n3886_ & ~new_n3887_;
  assign new_n3889_ = B6834 & B6833;
  assign new_n3890_ = ~new_n1880_ & ~new_n3889_;
  assign new_n3891_ = new_n1880_ & ~new_n3890_;
  assign new_n3892_ = new_n1880_ & new_n3889_;
  assign new_n3893_ = new_n3891_ & ~new_n3892_;
  assign new_n3894_ = B6834 & ~new_n3893_;
  assign new_n3895_ = ~new_n1883_ & ~new_n3894_;
  assign new_n3896_ = B6867 & B6866;
  assign new_n3897_ = ~new_n1890_ & ~new_n3896_;
  assign new_n3898_ = new_n1890_ & ~new_n3897_;
  assign new_n3899_ = new_n1890_ & new_n3896_;
  assign new_n3900_ = new_n3898_ & ~new_n3899_;
  assign new_n3901_ = B6867 & ~new_n3900_;
  assign new_n3902_ = ~new_n1893_ & ~new_n3901_;
  assign new_n3903_ = new_n3895_ & ~new_n3902_;
  assign new_n3904_ = ~new_n3895_ & new_n3902_;
  assign new_n3905_ = ~new_n3903_ & ~new_n3904_;
  assign new_n3906_ = B6900 & B6899;
  assign new_n3907_ = ~new_n1903_ & ~new_n3906_;
  assign new_n3908_ = new_n1903_ & ~new_n3907_;
  assign new_n3909_ = new_n1903_ & new_n3906_;
  assign new_n3910_ = new_n3908_ & ~new_n3909_;
  assign new_n3911_ = B6900 & ~new_n3910_;
  assign new_n3912_ = ~new_n1906_ & ~new_n3911_;
  assign new_n3913_ = B6933 & B6932;
  assign new_n3914_ = ~new_n1913_ & ~new_n3913_;
  assign new_n3915_ = new_n1913_ & ~new_n3914_;
  assign new_n3916_ = new_n1913_ & new_n3913_;
  assign new_n3917_ = new_n3915_ & ~new_n3916_;
  assign new_n3918_ = B6933 & ~new_n3917_;
  assign new_n3919_ = ~new_n1916_ & ~new_n3918_;
  assign new_n3920_ = new_n3905_ & new_n3919_;
  assign new_n3921_ = B6966 & B6965;
  assign new_n3922_ = ~new_n1924_ & ~new_n3921_;
  assign new_n3923_ = new_n1924_ & ~new_n3922_;
  assign new_n3924_ = new_n1924_ & new_n3921_;
  assign new_n3925_ = new_n3923_ & ~new_n3924_;
  assign new_n3926_ = B6966 & ~new_n3925_;
  assign new_n3927_ = ~new_n1927_ & ~new_n3926_;
  assign new_n3928_ = new_n3919_ & new_n3927_;
  assign new_n3929_ = ~new_n3920_ & ~new_n3928_;
  assign new_n3930_ = ~new_n3912_ & new_n3929_;
  assign new_n3931_ = new_n3912_ & ~new_n3929_;
  assign new_n3932_ = ~new_n3930_ & ~new_n3931_;
  assign new_n3933_ = ~new_n3905_ & ~new_n3932_;
  assign new_n3934_ = B6999 & B6998;
  assign new_n3935_ = ~new_n1940_ & ~new_n3934_;
  assign new_n3936_ = new_n1940_ & ~new_n3935_;
  assign new_n3937_ = new_n1940_ & new_n3934_;
  assign new_n3938_ = new_n3936_ & ~new_n3937_;
  assign new_n3939_ = B6999 & ~new_n3938_;
  assign new_n3940_ = ~new_n1943_ & ~new_n3939_;
  assign new_n3941_ = B7032 & B7031;
  assign new_n3942_ = ~new_n1950_ & ~new_n3941_;
  assign new_n3943_ = new_n1950_ & ~new_n3942_;
  assign new_n3944_ = new_n1950_ & new_n3941_;
  assign new_n3945_ = new_n3943_ & ~new_n3944_;
  assign new_n3946_ = B7032 & ~new_n3945_;
  assign new_n3947_ = ~new_n1953_ & ~new_n3946_;
  assign new_n3948_ = new_n3940_ & ~new_n3947_;
  assign new_n3949_ = ~new_n3940_ & new_n3947_;
  assign new_n3950_ = ~new_n3948_ & ~new_n3949_;
  assign new_n3951_ = B7065 & B7064;
  assign new_n3952_ = ~new_n1963_ & ~new_n3951_;
  assign new_n3953_ = new_n1963_ & ~new_n3952_;
  assign new_n3954_ = new_n1963_ & new_n3951_;
  assign new_n3955_ = new_n3953_ & ~new_n3954_;
  assign new_n3956_ = B7065 & ~new_n3955_;
  assign new_n3957_ = ~new_n1966_ & ~new_n3956_;
  assign new_n3958_ = B7098 & B7097;
  assign new_n3959_ = ~new_n1973_ & ~new_n3958_;
  assign new_n3960_ = new_n1973_ & ~new_n3959_;
  assign new_n3961_ = new_n1973_ & new_n3958_;
  assign new_n3962_ = new_n3960_ & ~new_n3961_;
  assign new_n3963_ = B7098 & ~new_n3962_;
  assign new_n3964_ = ~new_n1976_ & ~new_n3963_;
  assign new_n3965_ = new_n3950_ & new_n3964_;
  assign new_n3966_ = B7131 & B7130;
  assign new_n3967_ = ~new_n1984_ & ~new_n3966_;
  assign new_n3968_ = new_n1984_ & ~new_n3967_;
  assign new_n3969_ = new_n1984_ & new_n3966_;
  assign new_n3970_ = new_n3968_ & ~new_n3969_;
  assign new_n3971_ = B7131 & ~new_n3970_;
  assign new_n3972_ = ~new_n1987_ & ~new_n3971_;
  assign new_n3973_ = new_n3964_ & new_n3972_;
  assign new_n3974_ = ~new_n3965_ & ~new_n3973_;
  assign new_n3975_ = ~new_n3957_ & new_n3974_;
  assign new_n3976_ = new_n3957_ & ~new_n3974_;
  assign new_n3977_ = ~new_n3975_ & ~new_n3976_;
  assign new_n3978_ = ~new_n3950_ & ~new_n3977_;
  assign new_n3979_ = ~new_n3933_ & new_n3978_;
  assign new_n3980_ = new_n3933_ & ~new_n3978_;
  assign new_n3981_ = ~new_n3979_ & ~new_n3980_;
  assign new_n3982_ = B7164 & B7163;
  assign new_n3983_ = ~new_n2003_ & ~new_n3982_;
  assign new_n3984_ = new_n2003_ & ~new_n3983_;
  assign new_n3985_ = new_n2003_ & new_n3982_;
  assign new_n3986_ = new_n3984_ & ~new_n3985_;
  assign new_n3987_ = B7164 & ~new_n3986_;
  assign new_n3988_ = ~new_n2006_ & ~new_n3987_;
  assign new_n3989_ = B7197 & B7196;
  assign new_n3990_ = ~new_n2013_ & ~new_n3989_;
  assign new_n3991_ = new_n2013_ & ~new_n3990_;
  assign new_n3992_ = new_n2013_ & new_n3989_;
  assign new_n3993_ = new_n3991_ & ~new_n3992_;
  assign new_n3994_ = B7197 & ~new_n3993_;
  assign new_n3995_ = ~new_n2016_ & ~new_n3994_;
  assign new_n3996_ = new_n3988_ & ~new_n3995_;
  assign new_n3997_ = ~new_n3988_ & new_n3995_;
  assign new_n3998_ = ~new_n3996_ & ~new_n3997_;
  assign new_n3999_ = B7230 & B7229;
  assign new_n4000_ = ~new_n2026_ & ~new_n3999_;
  assign new_n4001_ = new_n2026_ & ~new_n4000_;
  assign new_n4002_ = new_n2026_ & new_n3999_;
  assign new_n4003_ = new_n4001_ & ~new_n4002_;
  assign new_n4004_ = B7230 & ~new_n4003_;
  assign new_n4005_ = ~new_n2029_ & ~new_n4004_;
  assign new_n4006_ = B7263 & B7262;
  assign new_n4007_ = ~new_n2036_ & ~new_n4006_;
  assign new_n4008_ = new_n2036_ & ~new_n4007_;
  assign new_n4009_ = new_n2036_ & new_n4006_;
  assign new_n4010_ = new_n4008_ & ~new_n4009_;
  assign new_n4011_ = B7263 & ~new_n4010_;
  assign new_n4012_ = ~new_n2039_ & ~new_n4011_;
  assign new_n4013_ = new_n3998_ & new_n4012_;
  assign new_n4014_ = B7296 & B7295;
  assign new_n4015_ = ~new_n2047_ & ~new_n4014_;
  assign new_n4016_ = new_n2047_ & ~new_n4015_;
  assign new_n4017_ = new_n2047_ & new_n4014_;
  assign new_n4018_ = new_n4016_ & ~new_n4017_;
  assign new_n4019_ = B7296 & ~new_n4018_;
  assign new_n4020_ = ~new_n2050_ & ~new_n4019_;
  assign new_n4021_ = new_n4012_ & new_n4020_;
  assign new_n4022_ = ~new_n4013_ & ~new_n4021_;
  assign new_n4023_ = ~new_n4005_ & new_n4022_;
  assign new_n4024_ = new_n4005_ & ~new_n4022_;
  assign new_n4025_ = ~new_n4023_ & ~new_n4024_;
  assign new_n4026_ = ~new_n3998_ & ~new_n4025_;
  assign new_n4027_ = B7329 & B7328;
  assign new_n4028_ = ~new_n2063_ & ~new_n4027_;
  assign new_n4029_ = new_n2063_ & ~new_n4028_;
  assign new_n4030_ = new_n2063_ & new_n4027_;
  assign new_n4031_ = new_n4029_ & ~new_n4030_;
  assign new_n4032_ = B7329 & ~new_n4031_;
  assign new_n4033_ = ~new_n2066_ & ~new_n4032_;
  assign new_n4034_ = B7362 & B7361;
  assign new_n4035_ = ~new_n2073_ & ~new_n4034_;
  assign new_n4036_ = new_n2073_ & ~new_n4035_;
  assign new_n4037_ = new_n2073_ & new_n4034_;
  assign new_n4038_ = new_n4036_ & ~new_n4037_;
  assign new_n4039_ = B7362 & ~new_n4038_;
  assign new_n4040_ = ~new_n2076_ & ~new_n4039_;
  assign new_n4041_ = new_n4033_ & ~new_n4040_;
  assign new_n4042_ = ~new_n4033_ & new_n4040_;
  assign new_n4043_ = ~new_n4041_ & ~new_n4042_;
  assign new_n4044_ = B7395 & B7394;
  assign new_n4045_ = ~new_n2086_ & ~new_n4044_;
  assign new_n4046_ = new_n2086_ & ~new_n4045_;
  assign new_n4047_ = new_n2086_ & new_n4044_;
  assign new_n4048_ = new_n4046_ & ~new_n4047_;
  assign new_n4049_ = B7395 & ~new_n4048_;
  assign new_n4050_ = ~new_n2089_ & ~new_n4049_;
  assign new_n4051_ = B7428 & B7427;
  assign new_n4052_ = ~new_n2096_ & ~new_n4051_;
  assign new_n4053_ = new_n2096_ & ~new_n4052_;
  assign new_n4054_ = new_n2096_ & new_n4051_;
  assign new_n4055_ = new_n4053_ & ~new_n4054_;
  assign new_n4056_ = B7428 & ~new_n4055_;
  assign new_n4057_ = ~new_n2099_ & ~new_n4056_;
  assign new_n4058_ = new_n4043_ & new_n4057_;
  assign new_n4059_ = B7461 & B7460;
  assign new_n4060_ = ~new_n2107_ & ~new_n4059_;
  assign new_n4061_ = new_n2107_ & ~new_n4060_;
  assign new_n4062_ = new_n2107_ & new_n4059_;
  assign new_n4063_ = new_n4061_ & ~new_n4062_;
  assign new_n4064_ = B7461 & ~new_n4063_;
  assign new_n4065_ = ~new_n2110_ & ~new_n4064_;
  assign new_n4066_ = new_n4057_ & new_n4065_;
  assign new_n4067_ = ~new_n4058_ & ~new_n4066_;
  assign new_n4068_ = ~new_n4050_ & new_n4067_;
  assign new_n4069_ = new_n4050_ & ~new_n4067_;
  assign new_n4070_ = ~new_n4068_ & ~new_n4069_;
  assign new_n4071_ = ~new_n4043_ & ~new_n4070_;
  assign new_n4072_ = new_n3981_ & ~new_n4071_;
  assign new_n4073_ = B7494 & B7493;
  assign new_n4074_ = ~new_n2124_ & ~new_n4073_;
  assign new_n4075_ = new_n2124_ & ~new_n4074_;
  assign new_n4076_ = new_n2124_ & new_n4073_;
  assign new_n4077_ = new_n4075_ & ~new_n4076_;
  assign new_n4078_ = B7494 & ~new_n4077_;
  assign new_n4079_ = ~new_n2127_ & ~new_n4078_;
  assign new_n4080_ = B7527 & B7526;
  assign new_n4081_ = ~new_n2134_ & ~new_n4080_;
  assign new_n4082_ = new_n2134_ & ~new_n4081_;
  assign new_n4083_ = new_n2134_ & new_n4080_;
  assign new_n4084_ = new_n4082_ & ~new_n4083_;
  assign new_n4085_ = B7527 & ~new_n4084_;
  assign new_n4086_ = ~new_n2137_ & ~new_n4085_;
  assign new_n4087_ = new_n4079_ & ~new_n4086_;
  assign new_n4088_ = ~new_n4079_ & new_n4086_;
  assign new_n4089_ = ~new_n4087_ & ~new_n4088_;
  assign new_n4090_ = B7560 & B7559;
  assign new_n4091_ = ~new_n2147_ & ~new_n4090_;
  assign new_n4092_ = new_n2147_ & ~new_n4091_;
  assign new_n4093_ = new_n2147_ & new_n4090_;
  assign new_n4094_ = new_n4092_ & ~new_n4093_;
  assign new_n4095_ = B7560 & ~new_n4094_;
  assign new_n4096_ = ~new_n2150_ & ~new_n4095_;
  assign new_n4097_ = B7593 & B7592;
  assign new_n4098_ = ~new_n2157_ & ~new_n4097_;
  assign new_n4099_ = new_n2157_ & ~new_n4098_;
  assign new_n4100_ = new_n2157_ & new_n4097_;
  assign new_n4101_ = new_n4099_ & ~new_n4100_;
  assign new_n4102_ = B7593 & ~new_n4101_;
  assign new_n4103_ = ~new_n2160_ & ~new_n4102_;
  assign new_n4104_ = new_n4089_ & new_n4103_;
  assign new_n4105_ = B7626 & B7625;
  assign new_n4106_ = ~new_n2168_ & ~new_n4105_;
  assign new_n4107_ = new_n2168_ & ~new_n4106_;
  assign new_n4108_ = new_n2168_ & new_n4105_;
  assign new_n4109_ = new_n4107_ & ~new_n4108_;
  assign new_n4110_ = B7626 & ~new_n4109_;
  assign new_n4111_ = ~new_n2171_ & ~new_n4110_;
  assign new_n4112_ = new_n4103_ & new_n4111_;
  assign new_n4113_ = ~new_n4104_ & ~new_n4112_;
  assign new_n4114_ = ~new_n4096_ & new_n4113_;
  assign new_n4115_ = new_n4096_ & ~new_n4113_;
  assign new_n4116_ = ~new_n4114_ & ~new_n4115_;
  assign new_n4117_ = ~new_n4089_ & ~new_n4116_;
  assign new_n4118_ = ~new_n4071_ & ~new_n4117_;
  assign new_n4119_ = ~new_n4072_ & ~new_n4118_;
  assign new_n4120_ = new_n4026_ & new_n4119_;
  assign new_n4121_ = ~new_n4026_ & ~new_n4119_;
  assign new_n4122_ = ~new_n4120_ & ~new_n4121_;
  assign new_n4123_ = ~new_n3981_ & ~new_n4122_;
  assign new_n4124_ = B7659 & B7658;
  assign new_n4125_ = ~new_n2190_ & ~new_n4124_;
  assign new_n4126_ = new_n2190_ & ~new_n4125_;
  assign new_n4127_ = new_n2190_ & new_n4124_;
  assign new_n4128_ = new_n4126_ & ~new_n4127_;
  assign new_n4129_ = B7659 & ~new_n4128_;
  assign new_n4130_ = ~new_n2193_ & ~new_n4129_;
  assign new_n4131_ = B7692 & B7691;
  assign new_n4132_ = ~new_n2200_ & ~new_n4131_;
  assign new_n4133_ = new_n2200_ & ~new_n4132_;
  assign new_n4134_ = new_n2200_ & new_n4131_;
  assign new_n4135_ = new_n4133_ & ~new_n4134_;
  assign new_n4136_ = B7692 & ~new_n4135_;
  assign new_n4137_ = ~new_n2203_ & ~new_n4136_;
  assign new_n4138_ = new_n4130_ & ~new_n4137_;
  assign new_n4139_ = ~new_n4130_ & new_n4137_;
  assign new_n4140_ = ~new_n4138_ & ~new_n4139_;
  assign new_n4141_ = B7725 & B7724;
  assign new_n4142_ = ~new_n2213_ & ~new_n4141_;
  assign new_n4143_ = new_n2213_ & ~new_n4142_;
  assign new_n4144_ = new_n2213_ & new_n4141_;
  assign new_n4145_ = new_n4143_ & ~new_n4144_;
  assign new_n4146_ = B7725 & ~new_n4145_;
  assign new_n4147_ = ~new_n2216_ & ~new_n4146_;
  assign new_n4148_ = B7758 & B7757;
  assign new_n4149_ = ~new_n2223_ & ~new_n4148_;
  assign new_n4150_ = new_n2223_ & ~new_n4149_;
  assign new_n4151_ = new_n2223_ & new_n4148_;
  assign new_n4152_ = new_n4150_ & ~new_n4151_;
  assign new_n4153_ = B7758 & ~new_n4152_;
  assign new_n4154_ = ~new_n2226_ & ~new_n4153_;
  assign new_n4155_ = new_n4140_ & new_n4154_;
  assign new_n4156_ = B7791 & B7790;
  assign new_n4157_ = ~new_n2234_ & ~new_n4156_;
  assign new_n4158_ = new_n2234_ & ~new_n4157_;
  assign new_n4159_ = new_n2234_ & new_n4156_;
  assign new_n4160_ = new_n4158_ & ~new_n4159_;
  assign new_n4161_ = B7791 & ~new_n4160_;
  assign new_n4162_ = ~new_n2237_ & ~new_n4161_;
  assign new_n4163_ = new_n4154_ & new_n4162_;
  assign new_n4164_ = ~new_n4155_ & ~new_n4163_;
  assign new_n4165_ = ~new_n4147_ & new_n4164_;
  assign new_n4166_ = new_n4147_ & ~new_n4164_;
  assign new_n4167_ = ~new_n4165_ & ~new_n4166_;
  assign new_n4168_ = ~new_n4140_ & ~new_n4167_;
  assign new_n4169_ = B7824 & B7823;
  assign new_n4170_ = ~new_n2250_ & ~new_n4169_;
  assign new_n4171_ = new_n2250_ & ~new_n4170_;
  assign new_n4172_ = new_n2250_ & new_n4169_;
  assign new_n4173_ = new_n4171_ & ~new_n4172_;
  assign new_n4174_ = B7824 & ~new_n4173_;
  assign new_n4175_ = ~new_n2253_ & ~new_n4174_;
  assign new_n4176_ = B7857 & B7856;
  assign new_n4177_ = ~new_n2260_ & ~new_n4176_;
  assign new_n4178_ = new_n2260_ & ~new_n4177_;
  assign new_n4179_ = new_n2260_ & new_n4176_;
  assign new_n4180_ = new_n4178_ & ~new_n4179_;
  assign new_n4181_ = B7857 & ~new_n4180_;
  assign new_n4182_ = ~new_n2263_ & ~new_n4181_;
  assign new_n4183_ = new_n4175_ & ~new_n4182_;
  assign new_n4184_ = ~new_n4175_ & new_n4182_;
  assign new_n4185_ = ~new_n4183_ & ~new_n4184_;
  assign new_n4186_ = B7890 & B7889;
  assign new_n4187_ = ~new_n2273_ & ~new_n4186_;
  assign new_n4188_ = new_n2273_ & ~new_n4187_;
  assign new_n4189_ = new_n2273_ & new_n4186_;
  assign new_n4190_ = new_n4188_ & ~new_n4189_;
  assign new_n4191_ = B7890 & ~new_n4190_;
  assign new_n4192_ = ~new_n2276_ & ~new_n4191_;
  assign new_n4193_ = B7923 & B7922;
  assign new_n4194_ = ~new_n2283_ & ~new_n4193_;
  assign new_n4195_ = new_n2283_ & ~new_n4194_;
  assign new_n4196_ = new_n2283_ & new_n4193_;
  assign new_n4197_ = new_n4195_ & ~new_n4196_;
  assign new_n4198_ = B7923 & ~new_n4197_;
  assign new_n4199_ = ~new_n2286_ & ~new_n4198_;
  assign new_n4200_ = new_n4185_ & new_n4199_;
  assign new_n4201_ = B7956 & B7955;
  assign new_n4202_ = ~new_n2294_ & ~new_n4201_;
  assign new_n4203_ = new_n2294_ & ~new_n4202_;
  assign new_n4204_ = new_n2294_ & new_n4201_;
  assign new_n4205_ = new_n4203_ & ~new_n4204_;
  assign new_n4206_ = B7956 & ~new_n4205_;
  assign new_n4207_ = ~new_n2297_ & ~new_n4206_;
  assign new_n4208_ = new_n4199_ & new_n4207_;
  assign new_n4209_ = ~new_n4200_ & ~new_n4208_;
  assign new_n4210_ = ~new_n4192_ & new_n4209_;
  assign new_n4211_ = new_n4192_ & ~new_n4209_;
  assign new_n4212_ = ~new_n4210_ & ~new_n4211_;
  assign new_n4213_ = ~new_n4185_ & ~new_n4212_;
  assign new_n4214_ = ~new_n4168_ & new_n4213_;
  assign new_n4215_ = new_n4168_ & ~new_n4213_;
  assign new_n4216_ = ~new_n4214_ & ~new_n4215_;
  assign new_n4217_ = B7989 & B7988;
  assign new_n4218_ = ~new_n2313_ & ~new_n4217_;
  assign new_n4219_ = new_n2313_ & ~new_n4218_;
  assign new_n4220_ = new_n2313_ & new_n4217_;
  assign new_n4221_ = new_n4219_ & ~new_n4220_;
  assign new_n4222_ = B7989 & ~new_n4221_;
  assign new_n4223_ = ~new_n2316_ & ~new_n4222_;
  assign new_n4224_ = B8022 & B8021;
  assign new_n4225_ = ~new_n2323_ & ~new_n4224_;
  assign new_n4226_ = new_n2323_ & ~new_n4225_;
  assign new_n4227_ = new_n2323_ & new_n4224_;
  assign new_n4228_ = new_n4226_ & ~new_n4227_;
  assign new_n4229_ = B8022 & ~new_n4228_;
  assign new_n4230_ = ~new_n2326_ & ~new_n4229_;
  assign new_n4231_ = new_n4223_ & ~new_n4230_;
  assign new_n4232_ = ~new_n4223_ & new_n4230_;
  assign new_n4233_ = ~new_n4231_ & ~new_n4232_;
  assign new_n4234_ = B8055 & B8054;
  assign new_n4235_ = ~new_n2336_ & ~new_n4234_;
  assign new_n4236_ = new_n2336_ & ~new_n4235_;
  assign new_n4237_ = new_n2336_ & new_n4234_;
  assign new_n4238_ = new_n4236_ & ~new_n4237_;
  assign new_n4239_ = B8055 & ~new_n4238_;
  assign new_n4240_ = ~new_n2339_ & ~new_n4239_;
  assign new_n4241_ = B8088 & B8087;
  assign new_n4242_ = ~new_n2346_ & ~new_n4241_;
  assign new_n4243_ = new_n2346_ & ~new_n4242_;
  assign new_n4244_ = new_n2346_ & new_n4241_;
  assign new_n4245_ = new_n4243_ & ~new_n4244_;
  assign new_n4246_ = B8088 & ~new_n4245_;
  assign new_n4247_ = ~new_n2349_ & ~new_n4246_;
  assign new_n4248_ = new_n4233_ & new_n4247_;
  assign new_n4249_ = B8121 & B8120;
  assign new_n4250_ = ~new_n2357_ & ~new_n4249_;
  assign new_n4251_ = new_n2357_ & ~new_n4250_;
  assign new_n4252_ = new_n2357_ & new_n4249_;
  assign new_n4253_ = new_n4251_ & ~new_n4252_;
  assign new_n4254_ = B8121 & ~new_n4253_;
  assign new_n4255_ = ~new_n2360_ & ~new_n4254_;
  assign new_n4256_ = new_n4247_ & new_n4255_;
  assign new_n4257_ = ~new_n4248_ & ~new_n4256_;
  assign new_n4258_ = ~new_n4240_ & new_n4257_;
  assign new_n4259_ = new_n4240_ & ~new_n4257_;
  assign new_n4260_ = ~new_n4258_ & ~new_n4259_;
  assign new_n4261_ = ~new_n4233_ & ~new_n4260_;
  assign new_n4262_ = B8154 & B8153;
  assign new_n4263_ = ~new_n2373_ & ~new_n4262_;
  assign new_n4264_ = new_n2373_ & ~new_n4263_;
  assign new_n4265_ = new_n2373_ & new_n4262_;
  assign new_n4266_ = new_n4264_ & ~new_n4265_;
  assign new_n4267_ = B8154 & ~new_n4266_;
  assign new_n4268_ = ~new_n2376_ & ~new_n4267_;
  assign new_n4269_ = B8187 & B8186;
  assign new_n4270_ = ~new_n2383_ & ~new_n4269_;
  assign new_n4271_ = new_n2383_ & ~new_n4270_;
  assign new_n4272_ = new_n2383_ & new_n4269_;
  assign new_n4273_ = new_n4271_ & ~new_n4272_;
  assign new_n4274_ = B8187 & ~new_n4273_;
  assign new_n4275_ = ~new_n2386_ & ~new_n4274_;
  assign new_n4276_ = new_n4268_ & ~new_n4275_;
  assign new_n4277_ = ~new_n4268_ & new_n4275_;
  assign new_n4278_ = ~new_n4276_ & ~new_n4277_;
  assign new_n4279_ = B8220 & B8219;
  assign new_n4280_ = ~new_n2396_ & ~new_n4279_;
  assign new_n4281_ = new_n2396_ & ~new_n4280_;
  assign new_n4282_ = new_n2396_ & new_n4279_;
  assign new_n4283_ = new_n4281_ & ~new_n4282_;
  assign new_n4284_ = B8220 & ~new_n4283_;
  assign new_n4285_ = ~new_n2399_ & ~new_n4284_;
  assign new_n4286_ = B8253 & B8252;
  assign new_n4287_ = ~new_n2406_ & ~new_n4286_;
  assign new_n4288_ = new_n2406_ & ~new_n4287_;
  assign new_n4289_ = new_n2406_ & new_n4286_;
  assign new_n4290_ = new_n4288_ & ~new_n4289_;
  assign new_n4291_ = B8253 & ~new_n4290_;
  assign new_n4292_ = ~new_n2409_ & ~new_n4291_;
  assign new_n4293_ = new_n4278_ & new_n4292_;
  assign new_n4294_ = B8286 & B8285;
  assign new_n4295_ = ~new_n2417_ & ~new_n4294_;
  assign new_n4296_ = new_n2417_ & ~new_n4295_;
  assign new_n4297_ = new_n2417_ & new_n4294_;
  assign new_n4298_ = new_n4296_ & ~new_n4297_;
  assign new_n4299_ = B8286 & ~new_n4298_;
  assign new_n4300_ = ~new_n2420_ & ~new_n4299_;
  assign new_n4301_ = new_n4292_ & new_n4300_;
  assign new_n4302_ = ~new_n4293_ & ~new_n4301_;
  assign new_n4303_ = ~new_n4285_ & new_n4302_;
  assign new_n4304_ = new_n4285_ & ~new_n4302_;
  assign new_n4305_ = ~new_n4303_ & ~new_n4304_;
  assign new_n4306_ = ~new_n4278_ & ~new_n4305_;
  assign new_n4307_ = new_n4216_ & ~new_n4306_;
  assign new_n4308_ = B8319 & B8318;
  assign new_n4309_ = ~new_n2434_ & ~new_n4308_;
  assign new_n4310_ = new_n2434_ & ~new_n4309_;
  assign new_n4311_ = new_n2434_ & new_n4308_;
  assign new_n4312_ = new_n4310_ & ~new_n4311_;
  assign new_n4313_ = B8319 & ~new_n4312_;
  assign new_n4314_ = ~new_n2437_ & ~new_n4313_;
  assign new_n4315_ = B8352 & B8351;
  assign new_n4316_ = ~new_n2444_ & ~new_n4315_;
  assign new_n4317_ = new_n2444_ & ~new_n4316_;
  assign new_n4318_ = new_n2444_ & new_n4315_;
  assign new_n4319_ = new_n4317_ & ~new_n4318_;
  assign new_n4320_ = B8352 & ~new_n4319_;
  assign new_n4321_ = ~new_n2447_ & ~new_n4320_;
  assign new_n4322_ = new_n4314_ & ~new_n4321_;
  assign new_n4323_ = ~new_n4314_ & new_n4321_;
  assign new_n4324_ = ~new_n4322_ & ~new_n4323_;
  assign new_n4325_ = B8385 & B8384;
  assign new_n4326_ = ~new_n2457_ & ~new_n4325_;
  assign new_n4327_ = new_n2457_ & ~new_n4326_;
  assign new_n4328_ = new_n2457_ & new_n4325_;
  assign new_n4329_ = new_n4327_ & ~new_n4328_;
  assign new_n4330_ = B8385 & ~new_n4329_;
  assign new_n4331_ = ~new_n2460_ & ~new_n4330_;
  assign new_n4332_ = B8418 & B8417;
  assign new_n4333_ = ~new_n2467_ & ~new_n4332_;
  assign new_n4334_ = new_n2467_ & ~new_n4333_;
  assign new_n4335_ = new_n2467_ & new_n4332_;
  assign new_n4336_ = new_n4334_ & ~new_n4335_;
  assign new_n4337_ = B8418 & ~new_n4336_;
  assign new_n4338_ = ~new_n2470_ & ~new_n4337_;
  assign new_n4339_ = new_n4324_ & new_n4338_;
  assign new_n4340_ = B8451 & B8450;
  assign new_n4341_ = ~new_n2478_ & ~new_n4340_;
  assign new_n4342_ = new_n2478_ & ~new_n4341_;
  assign new_n4343_ = new_n2478_ & new_n4340_;
  assign new_n4344_ = new_n4342_ & ~new_n4343_;
  assign new_n4345_ = B8451 & ~new_n4344_;
  assign new_n4346_ = ~new_n2481_ & ~new_n4345_;
  assign new_n4347_ = new_n4338_ & new_n4346_;
  assign new_n4348_ = ~new_n4339_ & ~new_n4347_;
  assign new_n4349_ = ~new_n4331_ & new_n4348_;
  assign new_n4350_ = new_n4331_ & ~new_n4348_;
  assign new_n4351_ = ~new_n4349_ & ~new_n4350_;
  assign new_n4352_ = ~new_n4324_ & ~new_n4351_;
  assign new_n4353_ = ~new_n4306_ & ~new_n4352_;
  assign new_n4354_ = ~new_n4307_ & ~new_n4353_;
  assign new_n4355_ = new_n4261_ & new_n4354_;
  assign new_n4356_ = ~new_n4261_ & ~new_n4354_;
  assign new_n4357_ = ~new_n4355_ & ~new_n4356_;
  assign new_n4358_ = ~new_n4216_ & ~new_n4357_;
  assign new_n4359_ = new_n3888_ & ~new_n4358_;
  assign new_n4360_ = B8484 & B8483;
  assign new_n4361_ = ~new_n2501_ & ~new_n4360_;
  assign new_n4362_ = new_n2501_ & ~new_n4361_;
  assign new_n4363_ = new_n2501_ & new_n4360_;
  assign new_n4364_ = new_n4362_ & ~new_n4363_;
  assign new_n4365_ = B8484 & ~new_n4364_;
  assign new_n4366_ = ~new_n2504_ & ~new_n4365_;
  assign new_n4367_ = B8517 & B8516;
  assign new_n4368_ = ~new_n2511_ & ~new_n4367_;
  assign new_n4369_ = new_n2511_ & ~new_n4368_;
  assign new_n4370_ = new_n2511_ & new_n4367_;
  assign new_n4371_ = new_n4369_ & ~new_n4370_;
  assign new_n4372_ = B8517 & ~new_n4371_;
  assign new_n4373_ = ~new_n2514_ & ~new_n4372_;
  assign new_n4374_ = new_n4366_ & ~new_n4373_;
  assign new_n4375_ = ~new_n4366_ & new_n4373_;
  assign new_n4376_ = ~new_n4374_ & ~new_n4375_;
  assign new_n4377_ = B8550 & B8549;
  assign new_n4378_ = ~new_n2524_ & ~new_n4377_;
  assign new_n4379_ = new_n2524_ & ~new_n4378_;
  assign new_n4380_ = new_n2524_ & new_n4377_;
  assign new_n4381_ = new_n4379_ & ~new_n4380_;
  assign new_n4382_ = B8550 & ~new_n4381_;
  assign new_n4383_ = ~new_n2527_ & ~new_n4382_;
  assign new_n4384_ = B8583 & B8582;
  assign new_n4385_ = ~new_n2534_ & ~new_n4384_;
  assign new_n4386_ = new_n2534_ & ~new_n4385_;
  assign new_n4387_ = new_n2534_ & new_n4384_;
  assign new_n4388_ = new_n4386_ & ~new_n4387_;
  assign new_n4389_ = B8583 & ~new_n4388_;
  assign new_n4390_ = ~new_n2537_ & ~new_n4389_;
  assign new_n4391_ = new_n4376_ & new_n4390_;
  assign new_n4392_ = B8616 & B8615;
  assign new_n4393_ = ~new_n2545_ & ~new_n4392_;
  assign new_n4394_ = new_n2545_ & ~new_n4393_;
  assign new_n4395_ = new_n2545_ & new_n4392_;
  assign new_n4396_ = new_n4394_ & ~new_n4395_;
  assign new_n4397_ = B8616 & ~new_n4396_;
  assign new_n4398_ = ~new_n2548_ & ~new_n4397_;
  assign new_n4399_ = new_n4390_ & new_n4398_;
  assign new_n4400_ = ~new_n4391_ & ~new_n4399_;
  assign new_n4401_ = ~new_n4383_ & new_n4400_;
  assign new_n4402_ = new_n4383_ & ~new_n4400_;
  assign new_n4403_ = ~new_n4401_ & ~new_n4402_;
  assign new_n4404_ = ~new_n4376_ & ~new_n4403_;
  assign new_n4405_ = B8649 & B8648;
  assign new_n4406_ = ~new_n2561_ & ~new_n4405_;
  assign new_n4407_ = new_n2561_ & ~new_n4406_;
  assign new_n4408_ = new_n2561_ & new_n4405_;
  assign new_n4409_ = new_n4407_ & ~new_n4408_;
  assign new_n4410_ = B8649 & ~new_n4409_;
  assign new_n4411_ = ~new_n2564_ & ~new_n4410_;
  assign new_n4412_ = B8682 & B8681;
  assign new_n4413_ = ~new_n2571_ & ~new_n4412_;
  assign new_n4414_ = new_n2571_ & ~new_n4413_;
  assign new_n4415_ = new_n2571_ & new_n4412_;
  assign new_n4416_ = new_n4414_ & ~new_n4415_;
  assign new_n4417_ = B8682 & ~new_n4416_;
  assign new_n4418_ = ~new_n2574_ & ~new_n4417_;
  assign new_n4419_ = new_n4411_ & ~new_n4418_;
  assign new_n4420_ = ~new_n4411_ & new_n4418_;
  assign new_n4421_ = ~new_n4419_ & ~new_n4420_;
  assign new_n4422_ = B8715 & B8714;
  assign new_n4423_ = ~new_n2584_ & ~new_n4422_;
  assign new_n4424_ = new_n2584_ & ~new_n4423_;
  assign new_n4425_ = new_n2584_ & new_n4422_;
  assign new_n4426_ = new_n4424_ & ~new_n4425_;
  assign new_n4427_ = B8715 & ~new_n4426_;
  assign new_n4428_ = ~new_n2587_ & ~new_n4427_;
  assign new_n4429_ = B8748 & B8747;
  assign new_n4430_ = ~new_n2594_ & ~new_n4429_;
  assign new_n4431_ = new_n2594_ & ~new_n4430_;
  assign new_n4432_ = new_n2594_ & new_n4429_;
  assign new_n4433_ = new_n4431_ & ~new_n4432_;
  assign new_n4434_ = B8748 & ~new_n4433_;
  assign new_n4435_ = ~new_n2597_ & ~new_n4434_;
  assign new_n4436_ = new_n4421_ & new_n4435_;
  assign new_n4437_ = B8781 & B8780;
  assign new_n4438_ = ~new_n2605_ & ~new_n4437_;
  assign new_n4439_ = new_n2605_ & ~new_n4438_;
  assign new_n4440_ = new_n2605_ & new_n4437_;
  assign new_n4441_ = new_n4439_ & ~new_n4440_;
  assign new_n4442_ = B8781 & ~new_n4441_;
  assign new_n4443_ = ~new_n2608_ & ~new_n4442_;
  assign new_n4444_ = new_n4435_ & new_n4443_;
  assign new_n4445_ = ~new_n4436_ & ~new_n4444_;
  assign new_n4446_ = ~new_n4428_ & new_n4445_;
  assign new_n4447_ = new_n4428_ & ~new_n4445_;
  assign new_n4448_ = ~new_n4446_ & ~new_n4447_;
  assign new_n4449_ = ~new_n4421_ & ~new_n4448_;
  assign new_n4450_ = ~new_n4404_ & new_n4449_;
  assign new_n4451_ = new_n4404_ & ~new_n4449_;
  assign new_n4452_ = ~new_n4450_ & ~new_n4451_;
  assign new_n4453_ = B8814 & B8813;
  assign new_n4454_ = ~new_n2624_ & ~new_n4453_;
  assign new_n4455_ = new_n2624_ & ~new_n4454_;
  assign new_n4456_ = new_n2624_ & new_n4453_;
  assign new_n4457_ = new_n4455_ & ~new_n4456_;
  assign new_n4458_ = B8814 & ~new_n4457_;
  assign new_n4459_ = ~new_n2627_ & ~new_n4458_;
  assign new_n4460_ = B8847 & B8846;
  assign new_n4461_ = ~new_n2634_ & ~new_n4460_;
  assign new_n4462_ = new_n2634_ & ~new_n4461_;
  assign new_n4463_ = new_n2634_ & new_n4460_;
  assign new_n4464_ = new_n4462_ & ~new_n4463_;
  assign new_n4465_ = B8847 & ~new_n4464_;
  assign new_n4466_ = ~new_n2637_ & ~new_n4465_;
  assign new_n4467_ = new_n4459_ & ~new_n4466_;
  assign new_n4468_ = ~new_n4459_ & new_n4466_;
  assign new_n4469_ = ~new_n4467_ & ~new_n4468_;
  assign new_n4470_ = B8880 & B8879;
  assign new_n4471_ = ~new_n2647_ & ~new_n4470_;
  assign new_n4472_ = new_n2647_ & ~new_n4471_;
  assign new_n4473_ = new_n2647_ & new_n4470_;
  assign new_n4474_ = new_n4472_ & ~new_n4473_;
  assign new_n4475_ = B8880 & ~new_n4474_;
  assign new_n4476_ = ~new_n2650_ & ~new_n4475_;
  assign new_n4477_ = B8913 & B8912;
  assign new_n4478_ = ~new_n2657_ & ~new_n4477_;
  assign new_n4479_ = new_n2657_ & ~new_n4478_;
  assign new_n4480_ = new_n2657_ & new_n4477_;
  assign new_n4481_ = new_n4479_ & ~new_n4480_;
  assign new_n4482_ = B8913 & ~new_n4481_;
  assign new_n4483_ = ~new_n2660_ & ~new_n4482_;
  assign new_n4484_ = new_n4469_ & new_n4483_;
  assign new_n4485_ = B8946 & B8945;
  assign new_n4486_ = ~new_n2668_ & ~new_n4485_;
  assign new_n4487_ = new_n2668_ & ~new_n4486_;
  assign new_n4488_ = new_n2668_ & new_n4485_;
  assign new_n4489_ = new_n4487_ & ~new_n4488_;
  assign new_n4490_ = B8946 & ~new_n4489_;
  assign new_n4491_ = ~new_n2671_ & ~new_n4490_;
  assign new_n4492_ = new_n4483_ & new_n4491_;
  assign new_n4493_ = ~new_n4484_ & ~new_n4492_;
  assign new_n4494_ = ~new_n4476_ & new_n4493_;
  assign new_n4495_ = new_n4476_ & ~new_n4493_;
  assign new_n4496_ = ~new_n4494_ & ~new_n4495_;
  assign new_n4497_ = ~new_n4469_ & ~new_n4496_;
  assign new_n4498_ = B8979 & B8978;
  assign new_n4499_ = ~new_n2684_ & ~new_n4498_;
  assign new_n4500_ = new_n2684_ & ~new_n4499_;
  assign new_n4501_ = new_n2684_ & new_n4498_;
  assign new_n4502_ = new_n4500_ & ~new_n4501_;
  assign new_n4503_ = B8979 & ~new_n4502_;
  assign new_n4504_ = ~new_n2687_ & ~new_n4503_;
  assign new_n4505_ = B9012 & B9011;
  assign new_n4506_ = ~new_n2694_ & ~new_n4505_;
  assign new_n4507_ = new_n2694_ & ~new_n4506_;
  assign new_n4508_ = new_n2694_ & new_n4505_;
  assign new_n4509_ = new_n4507_ & ~new_n4508_;
  assign new_n4510_ = B9012 & ~new_n4509_;
  assign new_n4511_ = ~new_n2697_ & ~new_n4510_;
  assign new_n4512_ = new_n4504_ & ~new_n4511_;
  assign new_n4513_ = ~new_n4504_ & new_n4511_;
  assign new_n4514_ = ~new_n4512_ & ~new_n4513_;
  assign new_n4515_ = B9045 & B9044;
  assign new_n4516_ = ~new_n2707_ & ~new_n4515_;
  assign new_n4517_ = new_n2707_ & ~new_n4516_;
  assign new_n4518_ = new_n2707_ & new_n4515_;
  assign new_n4519_ = new_n4517_ & ~new_n4518_;
  assign new_n4520_ = B9045 & ~new_n4519_;
  assign new_n4521_ = ~new_n2710_ & ~new_n4520_;
  assign new_n4522_ = B9078 & B9077;
  assign new_n4523_ = ~new_n2717_ & ~new_n4522_;
  assign new_n4524_ = new_n2717_ & ~new_n4523_;
  assign new_n4525_ = new_n2717_ & new_n4522_;
  assign new_n4526_ = new_n4524_ & ~new_n4525_;
  assign new_n4527_ = B9078 & ~new_n4526_;
  assign new_n4528_ = ~new_n2720_ & ~new_n4527_;
  assign new_n4529_ = new_n4514_ & new_n4528_;
  assign new_n4530_ = B9111 & B9110;
  assign new_n4531_ = ~new_n2728_ & ~new_n4530_;
  assign new_n4532_ = new_n2728_ & ~new_n4531_;
  assign new_n4533_ = new_n2728_ & new_n4530_;
  assign new_n4534_ = new_n4532_ & ~new_n4533_;
  assign new_n4535_ = B9111 & ~new_n4534_;
  assign new_n4536_ = ~new_n2731_ & ~new_n4535_;
  assign new_n4537_ = new_n4528_ & new_n4536_;
  assign new_n4538_ = ~new_n4529_ & ~new_n4537_;
  assign new_n4539_ = ~new_n4521_ & new_n4538_;
  assign new_n4540_ = new_n4521_ & ~new_n4538_;
  assign new_n4541_ = ~new_n4539_ & ~new_n4540_;
  assign new_n4542_ = ~new_n4514_ & ~new_n4541_;
  assign new_n4543_ = new_n4452_ & ~new_n4542_;
  assign new_n4544_ = B9144 & B9143;
  assign new_n4545_ = ~new_n2745_ & ~new_n4544_;
  assign new_n4546_ = new_n2745_ & ~new_n4545_;
  assign new_n4547_ = new_n2745_ & new_n4544_;
  assign new_n4548_ = new_n4546_ & ~new_n4547_;
  assign new_n4549_ = B9144 & ~new_n4548_;
  assign new_n4550_ = ~new_n2748_ & ~new_n4549_;
  assign new_n4551_ = B9177 & B9176;
  assign new_n4552_ = ~new_n2755_ & ~new_n4551_;
  assign new_n4553_ = new_n2755_ & ~new_n4552_;
  assign new_n4554_ = new_n2755_ & new_n4551_;
  assign new_n4555_ = new_n4553_ & ~new_n4554_;
  assign new_n4556_ = B9177 & ~new_n4555_;
  assign new_n4557_ = ~new_n2758_ & ~new_n4556_;
  assign new_n4558_ = new_n4550_ & ~new_n4557_;
  assign new_n4559_ = ~new_n4550_ & new_n4557_;
  assign new_n4560_ = ~new_n4558_ & ~new_n4559_;
  assign new_n4561_ = B9210 & B9209;
  assign new_n4562_ = ~new_n2768_ & ~new_n4561_;
  assign new_n4563_ = new_n2768_ & ~new_n4562_;
  assign new_n4564_ = new_n2768_ & new_n4561_;
  assign new_n4565_ = new_n4563_ & ~new_n4564_;
  assign new_n4566_ = B9210 & ~new_n4565_;
  assign new_n4567_ = ~new_n2771_ & ~new_n4566_;
  assign new_n4568_ = B9243 & B9242;
  assign new_n4569_ = ~new_n2778_ & ~new_n4568_;
  assign new_n4570_ = new_n2778_ & ~new_n4569_;
  assign new_n4571_ = new_n2778_ & new_n4568_;
  assign new_n4572_ = new_n4570_ & ~new_n4571_;
  assign new_n4573_ = B9243 & ~new_n4572_;
  assign new_n4574_ = ~new_n2781_ & ~new_n4573_;
  assign new_n4575_ = new_n4560_ & new_n4574_;
  assign new_n4576_ = B9276 & B9275;
  assign new_n4577_ = ~new_n2789_ & ~new_n4576_;
  assign new_n4578_ = new_n2789_ & ~new_n4577_;
  assign new_n4579_ = new_n2789_ & new_n4576_;
  assign new_n4580_ = new_n4578_ & ~new_n4579_;
  assign new_n4581_ = B9276 & ~new_n4580_;
  assign new_n4582_ = ~new_n2792_ & ~new_n4581_;
  assign new_n4583_ = new_n4574_ & new_n4582_;
  assign new_n4584_ = ~new_n4575_ & ~new_n4583_;
  assign new_n4585_ = ~new_n4567_ & new_n4584_;
  assign new_n4586_ = new_n4567_ & ~new_n4584_;
  assign new_n4587_ = ~new_n4585_ & ~new_n4586_;
  assign new_n4588_ = ~new_n4560_ & ~new_n4587_;
  assign new_n4589_ = ~new_n4542_ & ~new_n4588_;
  assign new_n4590_ = ~new_n4543_ & ~new_n4589_;
  assign new_n4591_ = new_n4497_ & new_n4590_;
  assign new_n4592_ = ~new_n4497_ & ~new_n4590_;
  assign new_n4593_ = ~new_n4591_ & ~new_n4592_;
  assign new_n4594_ = ~new_n4452_ & ~new_n4593_;
  assign new_n4595_ = ~new_n4358_ & ~new_n4594_;
  assign new_n4596_ = ~new_n4359_ & ~new_n4595_;
  assign new_n4597_ = new_n4123_ & new_n4596_;
  assign new_n4598_ = ~new_n4123_ & ~new_n4596_;
  assign new_n4599_ = ~new_n4597_ & ~new_n4598_;
  assign A6841 = ~new_n3888_ & ~new_n4599_;
  assign new_n4601_ = ~new_n3885_ & ~new_n4597_;
  assign A6840 = ~new_n3888_ & ~new_n4601_;
  assign new_n4603_ = new_n3885_ & new_n4123_;
  assign new_n4604_ = ~new_n3888_ & ~new_n4603_;
  assign new_n4605_ = new_n3888_ & ~new_n4604_;
  assign new_n4606_ = new_n3888_ & new_n4603_;
  assign new_n4607_ = new_n4605_ & ~new_n4606_;
  assign new_n4608_ = new_n4123_ & ~new_n4607_;
  assign A6839 = new_n4596_ | new_n4608_;
  assign new_n4610_ = new_n4358_ & new_n4594_;
  assign new_n4611_ = ~new_n4595_ & ~new_n4610_;
  assign new_n4612_ = ~new_n3888_ & ~new_n4358_;
  assign new_n4613_ = new_n3888_ & new_n4358_;
  assign new_n4614_ = ~new_n4612_ & ~new_n4613_;
  assign new_n4615_ = new_n4611_ & ~new_n4614_;
  assign A6838 = new_n4608_ | new_n4615_;
  assign new_n4617_ = new_n4123_ & ~new_n4615_;
  assign new_n4618_ = ~new_n4123_ & new_n4615_;
  assign new_n4619_ = ~new_n4617_ & ~new_n4618_;
  assign A6837 = ~new_n3888_ & ~new_n4619_;
  assign new_n4621_ = B5184 & new_n3421_;
  assign new_n4622_ = ~B5183 & ~new_n4621_;
  assign new_n4623_ = ~new_n1256_ & ~new_n4622_;
  assign new_n4624_ = B5219 & B5218;
  assign new_n4625_ = ~new_n1269_ & ~new_n4624_;
  assign new_n4626_ = ~B5218 & ~new_n1267_;
  assign new_n4627_ = B5218 & new_n1267_;
  assign new_n4628_ = ~new_n4626_ & ~new_n4627_;
  assign new_n4629_ = new_n4625_ & ~new_n4628_;
  assign new_n4630_ = ~new_n3428_ & ~new_n4629_;
  assign new_n4631_ = ~new_n4623_ & ~new_n4630_;
  assign new_n4632_ = new_n4623_ & new_n4630_;
  assign new_n4633_ = ~new_n4631_ & ~new_n4632_;
  assign new_n4634_ = B5252 & B5251;
  assign new_n4635_ = ~new_n1282_ & ~new_n4634_;
  assign new_n4636_ = ~B5251 & ~new_n1280_;
  assign new_n4637_ = B5251 & new_n1280_;
  assign new_n4638_ = ~new_n4636_ & ~new_n4637_;
  assign new_n4639_ = new_n4635_ & ~new_n4638_;
  assign new_n4640_ = ~new_n3438_ & ~new_n4639_;
  assign new_n4641_ = B5285 & B5284;
  assign new_n4642_ = ~new_n1292_ & ~new_n4641_;
  assign new_n4643_ = ~B5284 & ~new_n1290_;
  assign new_n4644_ = B5284 & new_n1290_;
  assign new_n4645_ = ~new_n4643_ & ~new_n4644_;
  assign new_n4646_ = new_n4642_ & ~new_n4645_;
  assign new_n4647_ = ~new_n3445_ & ~new_n4646_;
  assign new_n4648_ = new_n4633_ & new_n4647_;
  assign new_n4649_ = B5318 & B5317;
  assign new_n4650_ = ~new_n1303_ & ~new_n4649_;
  assign new_n4651_ = ~B5317 & ~new_n1301_;
  assign new_n4652_ = B5317 & new_n1301_;
  assign new_n4653_ = ~new_n4651_ & ~new_n4652_;
  assign new_n4654_ = new_n4650_ & ~new_n4653_;
  assign new_n4655_ = ~new_n3453_ & ~new_n4654_;
  assign new_n4656_ = new_n4647_ & new_n4655_;
  assign new_n4657_ = ~new_n4648_ & ~new_n4656_;
  assign new_n4658_ = ~new_n4640_ & new_n4657_;
  assign new_n4659_ = new_n4640_ & ~new_n4657_;
  assign new_n4660_ = ~new_n4658_ & ~new_n4659_;
  assign new_n4661_ = ~new_n4633_ & ~new_n4660_;
  assign new_n4662_ = B5351 & B5350;
  assign new_n4663_ = ~new_n1319_ & ~new_n4662_;
  assign new_n4664_ = ~B5350 & ~new_n1317_;
  assign new_n4665_ = B5350 & new_n1317_;
  assign new_n4666_ = ~new_n4664_ & ~new_n4665_;
  assign new_n4667_ = new_n4663_ & ~new_n4666_;
  assign new_n4668_ = ~new_n3466_ & ~new_n4667_;
  assign new_n4669_ = B5384 & B5383;
  assign new_n4670_ = ~new_n1329_ & ~new_n4669_;
  assign new_n4671_ = ~B5383 & ~new_n1327_;
  assign new_n4672_ = B5383 & new_n1327_;
  assign new_n4673_ = ~new_n4671_ & ~new_n4672_;
  assign new_n4674_ = new_n4670_ & ~new_n4673_;
  assign new_n4675_ = ~new_n3473_ & ~new_n4674_;
  assign new_n4676_ = new_n4668_ & ~new_n4675_;
  assign new_n4677_ = ~new_n4668_ & new_n4675_;
  assign new_n4678_ = ~new_n4676_ & ~new_n4677_;
  assign new_n4679_ = B5417 & B5416;
  assign new_n4680_ = ~new_n1342_ & ~new_n4679_;
  assign new_n4681_ = ~B5416 & ~new_n1340_;
  assign new_n4682_ = B5416 & new_n1340_;
  assign new_n4683_ = ~new_n4681_ & ~new_n4682_;
  assign new_n4684_ = new_n4680_ & ~new_n4683_;
  assign new_n4685_ = ~new_n3483_ & ~new_n4684_;
  assign new_n4686_ = B5450 & B5449;
  assign new_n4687_ = ~new_n1352_ & ~new_n4686_;
  assign new_n4688_ = ~B5449 & ~new_n1350_;
  assign new_n4689_ = B5449 & new_n1350_;
  assign new_n4690_ = ~new_n4688_ & ~new_n4689_;
  assign new_n4691_ = new_n4687_ & ~new_n4690_;
  assign new_n4692_ = ~new_n3490_ & ~new_n4691_;
  assign new_n4693_ = new_n4678_ & new_n4692_;
  assign new_n4694_ = B5483 & B5482;
  assign new_n4695_ = ~new_n1363_ & ~new_n4694_;
  assign new_n4696_ = ~B5482 & ~new_n1361_;
  assign new_n4697_ = B5482 & new_n1361_;
  assign new_n4698_ = ~new_n4696_ & ~new_n4697_;
  assign new_n4699_ = new_n4695_ & ~new_n4698_;
  assign new_n4700_ = ~new_n3498_ & ~new_n4699_;
  assign new_n4701_ = new_n4692_ & new_n4700_;
  assign new_n4702_ = ~new_n4693_ & ~new_n4701_;
  assign new_n4703_ = ~new_n4685_ & new_n4702_;
  assign new_n4704_ = new_n4685_ & ~new_n4702_;
  assign new_n4705_ = ~new_n4703_ & ~new_n4704_;
  assign new_n4706_ = ~new_n4678_ & ~new_n4705_;
  assign new_n4707_ = ~new_n4661_ & new_n4706_;
  assign new_n4708_ = new_n4661_ & ~new_n4706_;
  assign new_n4709_ = ~new_n4707_ & ~new_n4708_;
  assign new_n4710_ = B5516 & B5515;
  assign new_n4711_ = ~new_n1382_ & ~new_n4710_;
  assign new_n4712_ = ~B5515 & ~new_n1380_;
  assign new_n4713_ = B5515 & new_n1380_;
  assign new_n4714_ = ~new_n4712_ & ~new_n4713_;
  assign new_n4715_ = new_n4711_ & ~new_n4714_;
  assign new_n4716_ = ~new_n3514_ & ~new_n4715_;
  assign new_n4717_ = B5549 & B5548;
  assign new_n4718_ = ~new_n1392_ & ~new_n4717_;
  assign new_n4719_ = ~B5548 & ~new_n1390_;
  assign new_n4720_ = B5548 & new_n1390_;
  assign new_n4721_ = ~new_n4719_ & ~new_n4720_;
  assign new_n4722_ = new_n4718_ & ~new_n4721_;
  assign new_n4723_ = ~new_n3521_ & ~new_n4722_;
  assign new_n4724_ = new_n4716_ & ~new_n4723_;
  assign new_n4725_ = ~new_n4716_ & new_n4723_;
  assign new_n4726_ = ~new_n4724_ & ~new_n4725_;
  assign new_n4727_ = B5582 & B5581;
  assign new_n4728_ = ~new_n1405_ & ~new_n4727_;
  assign new_n4729_ = ~B5581 & ~new_n1403_;
  assign new_n4730_ = B5581 & new_n1403_;
  assign new_n4731_ = ~new_n4729_ & ~new_n4730_;
  assign new_n4732_ = new_n4728_ & ~new_n4731_;
  assign new_n4733_ = ~new_n3531_ & ~new_n4732_;
  assign new_n4734_ = B5615 & B5614;
  assign new_n4735_ = ~new_n1415_ & ~new_n4734_;
  assign new_n4736_ = ~B5614 & ~new_n1413_;
  assign new_n4737_ = B5614 & new_n1413_;
  assign new_n4738_ = ~new_n4736_ & ~new_n4737_;
  assign new_n4739_ = new_n4735_ & ~new_n4738_;
  assign new_n4740_ = ~new_n3538_ & ~new_n4739_;
  assign new_n4741_ = new_n4726_ & new_n4740_;
  assign new_n4742_ = B5648 & B5647;
  assign new_n4743_ = ~new_n1426_ & ~new_n4742_;
  assign new_n4744_ = ~B5647 & ~new_n1424_;
  assign new_n4745_ = B5647 & new_n1424_;
  assign new_n4746_ = ~new_n4744_ & ~new_n4745_;
  assign new_n4747_ = new_n4743_ & ~new_n4746_;
  assign new_n4748_ = ~new_n3546_ & ~new_n4747_;
  assign new_n4749_ = new_n4740_ & new_n4748_;
  assign new_n4750_ = ~new_n4741_ & ~new_n4749_;
  assign new_n4751_ = ~new_n4733_ & new_n4750_;
  assign new_n4752_ = new_n4733_ & ~new_n4750_;
  assign new_n4753_ = ~new_n4751_ & ~new_n4752_;
  assign new_n4754_ = ~new_n4726_ & ~new_n4753_;
  assign new_n4755_ = B5681 & B5680;
  assign new_n4756_ = ~new_n1442_ & ~new_n4755_;
  assign new_n4757_ = ~B5680 & ~new_n1440_;
  assign new_n4758_ = B5680 & new_n1440_;
  assign new_n4759_ = ~new_n4757_ & ~new_n4758_;
  assign new_n4760_ = new_n4756_ & ~new_n4759_;
  assign new_n4761_ = ~new_n3559_ & ~new_n4760_;
  assign new_n4762_ = B5714 & B5713;
  assign new_n4763_ = ~new_n1452_ & ~new_n4762_;
  assign new_n4764_ = ~B5713 & ~new_n1450_;
  assign new_n4765_ = B5713 & new_n1450_;
  assign new_n4766_ = ~new_n4764_ & ~new_n4765_;
  assign new_n4767_ = new_n4763_ & ~new_n4766_;
  assign new_n4768_ = ~new_n3566_ & ~new_n4767_;
  assign new_n4769_ = new_n4761_ & ~new_n4768_;
  assign new_n4770_ = ~new_n4761_ & new_n4768_;
  assign new_n4771_ = ~new_n4769_ & ~new_n4770_;
  assign new_n4772_ = B5747 & B5746;
  assign new_n4773_ = ~new_n1465_ & ~new_n4772_;
  assign new_n4774_ = ~B5746 & ~new_n1463_;
  assign new_n4775_ = B5746 & new_n1463_;
  assign new_n4776_ = ~new_n4774_ & ~new_n4775_;
  assign new_n4777_ = new_n4773_ & ~new_n4776_;
  assign new_n4778_ = ~new_n3576_ & ~new_n4777_;
  assign new_n4779_ = B5780 & B5779;
  assign new_n4780_ = ~new_n1475_ & ~new_n4779_;
  assign new_n4781_ = ~B5779 & ~new_n1473_;
  assign new_n4782_ = B5779 & new_n1473_;
  assign new_n4783_ = ~new_n4781_ & ~new_n4782_;
  assign new_n4784_ = new_n4780_ & ~new_n4783_;
  assign new_n4785_ = ~new_n3583_ & ~new_n4784_;
  assign new_n4786_ = new_n4771_ & new_n4785_;
  assign new_n4787_ = B5813 & B5812;
  assign new_n4788_ = ~new_n1486_ & ~new_n4787_;
  assign new_n4789_ = ~B5812 & ~new_n1484_;
  assign new_n4790_ = B5812 & new_n1484_;
  assign new_n4791_ = ~new_n4789_ & ~new_n4790_;
  assign new_n4792_ = new_n4788_ & ~new_n4791_;
  assign new_n4793_ = ~new_n3591_ & ~new_n4792_;
  assign new_n4794_ = new_n4785_ & new_n4793_;
  assign new_n4795_ = ~new_n4786_ & ~new_n4794_;
  assign new_n4796_ = ~new_n4778_ & new_n4795_;
  assign new_n4797_ = new_n4778_ & ~new_n4795_;
  assign new_n4798_ = ~new_n4796_ & ~new_n4797_;
  assign new_n4799_ = ~new_n4771_ & ~new_n4798_;
  assign new_n4800_ = new_n4709_ & ~new_n4799_;
  assign new_n4801_ = B5846 & B5845;
  assign new_n4802_ = ~new_n1503_ & ~new_n4801_;
  assign new_n4803_ = ~B5845 & ~new_n1501_;
  assign new_n4804_ = B5845 & new_n1501_;
  assign new_n4805_ = ~new_n4803_ & ~new_n4804_;
  assign new_n4806_ = new_n4802_ & ~new_n4805_;
  assign new_n4807_ = ~new_n3605_ & ~new_n4806_;
  assign new_n4808_ = B5879 & B5878;
  assign new_n4809_ = ~new_n1513_ & ~new_n4808_;
  assign new_n4810_ = ~B5878 & ~new_n1511_;
  assign new_n4811_ = B5878 & new_n1511_;
  assign new_n4812_ = ~new_n4810_ & ~new_n4811_;
  assign new_n4813_ = new_n4809_ & ~new_n4812_;
  assign new_n4814_ = ~new_n3612_ & ~new_n4813_;
  assign new_n4815_ = new_n4807_ & ~new_n4814_;
  assign new_n4816_ = ~new_n4807_ & new_n4814_;
  assign new_n4817_ = ~new_n4815_ & ~new_n4816_;
  assign new_n4818_ = B5912 & B5911;
  assign new_n4819_ = ~new_n1526_ & ~new_n4818_;
  assign new_n4820_ = ~B5911 & ~new_n1524_;
  assign new_n4821_ = B5911 & new_n1524_;
  assign new_n4822_ = ~new_n4820_ & ~new_n4821_;
  assign new_n4823_ = new_n4819_ & ~new_n4822_;
  assign new_n4824_ = ~new_n3622_ & ~new_n4823_;
  assign new_n4825_ = B5945 & B5944;
  assign new_n4826_ = ~new_n1536_ & ~new_n4825_;
  assign new_n4827_ = ~B5944 & ~new_n1534_;
  assign new_n4828_ = B5944 & new_n1534_;
  assign new_n4829_ = ~new_n4827_ & ~new_n4828_;
  assign new_n4830_ = new_n4826_ & ~new_n4829_;
  assign new_n4831_ = ~new_n3629_ & ~new_n4830_;
  assign new_n4832_ = new_n4817_ & new_n4831_;
  assign new_n4833_ = B5978 & B5977;
  assign new_n4834_ = ~new_n1547_ & ~new_n4833_;
  assign new_n4835_ = ~B5977 & ~new_n1545_;
  assign new_n4836_ = B5977 & new_n1545_;
  assign new_n4837_ = ~new_n4835_ & ~new_n4836_;
  assign new_n4838_ = new_n4834_ & ~new_n4837_;
  assign new_n4839_ = ~new_n3637_ & ~new_n4838_;
  assign new_n4840_ = new_n4831_ & new_n4839_;
  assign new_n4841_ = ~new_n4832_ & ~new_n4840_;
  assign new_n4842_ = ~new_n4824_ & new_n4841_;
  assign new_n4843_ = new_n4824_ & ~new_n4841_;
  assign new_n4844_ = ~new_n4842_ & ~new_n4843_;
  assign new_n4845_ = ~new_n4817_ & ~new_n4844_;
  assign new_n4846_ = ~new_n4799_ & ~new_n4845_;
  assign new_n4847_ = ~new_n4800_ & ~new_n4846_;
  assign new_n4848_ = new_n4754_ & new_n4847_;
  assign new_n4849_ = ~new_n4754_ & ~new_n4847_;
  assign new_n4850_ = ~new_n4848_ & ~new_n4849_;
  assign new_n4851_ = ~new_n4709_ & ~new_n4850_;
  assign new_n4852_ = B6011 & B6010;
  assign new_n4853_ = ~new_n1569_ & ~new_n4852_;
  assign new_n4854_ = ~B6010 & ~new_n1567_;
  assign new_n4855_ = B6010 & new_n1567_;
  assign new_n4856_ = ~new_n4854_ & ~new_n4855_;
  assign new_n4857_ = new_n4853_ & ~new_n4856_;
  assign new_n4858_ = ~new_n3656_ & ~new_n4857_;
  assign new_n4859_ = B6044 & B6043;
  assign new_n4860_ = ~new_n1579_ & ~new_n4859_;
  assign new_n4861_ = ~B6043 & ~new_n1577_;
  assign new_n4862_ = B6043 & new_n1577_;
  assign new_n4863_ = ~new_n4861_ & ~new_n4862_;
  assign new_n4864_ = new_n4860_ & ~new_n4863_;
  assign new_n4865_ = ~new_n3663_ & ~new_n4864_;
  assign new_n4866_ = new_n4858_ & ~new_n4865_;
  assign new_n4867_ = ~new_n4858_ & new_n4865_;
  assign new_n4868_ = ~new_n4866_ & ~new_n4867_;
  assign new_n4869_ = B6077 & B6076;
  assign new_n4870_ = ~new_n1592_ & ~new_n4869_;
  assign new_n4871_ = ~B6076 & ~new_n1590_;
  assign new_n4872_ = B6076 & new_n1590_;
  assign new_n4873_ = ~new_n4871_ & ~new_n4872_;
  assign new_n4874_ = new_n4870_ & ~new_n4873_;
  assign new_n4875_ = ~new_n3673_ & ~new_n4874_;
  assign new_n4876_ = B6110 & B6109;
  assign new_n4877_ = ~new_n1602_ & ~new_n4876_;
  assign new_n4878_ = ~B6109 & ~new_n1600_;
  assign new_n4879_ = B6109 & new_n1600_;
  assign new_n4880_ = ~new_n4878_ & ~new_n4879_;
  assign new_n4881_ = new_n4877_ & ~new_n4880_;
  assign new_n4882_ = ~new_n3680_ & ~new_n4881_;
  assign new_n4883_ = new_n4868_ & new_n4882_;
  assign new_n4884_ = B6143 & B6142;
  assign new_n4885_ = ~new_n1613_ & ~new_n4884_;
  assign new_n4886_ = ~B6142 & ~new_n1611_;
  assign new_n4887_ = B6142 & new_n1611_;
  assign new_n4888_ = ~new_n4886_ & ~new_n4887_;
  assign new_n4889_ = new_n4885_ & ~new_n4888_;
  assign new_n4890_ = ~new_n3688_ & ~new_n4889_;
  assign new_n4891_ = new_n4882_ & new_n4890_;
  assign new_n4892_ = ~new_n4883_ & ~new_n4891_;
  assign new_n4893_ = ~new_n4875_ & new_n4892_;
  assign new_n4894_ = new_n4875_ & ~new_n4892_;
  assign new_n4895_ = ~new_n4893_ & ~new_n4894_;
  assign new_n4896_ = ~new_n4868_ & ~new_n4895_;
  assign new_n4897_ = B6176 & B6175;
  assign new_n4898_ = ~new_n1629_ & ~new_n4897_;
  assign new_n4899_ = ~B6175 & ~new_n1627_;
  assign new_n4900_ = B6175 & new_n1627_;
  assign new_n4901_ = ~new_n4899_ & ~new_n4900_;
  assign new_n4902_ = new_n4898_ & ~new_n4901_;
  assign new_n4903_ = ~new_n3701_ & ~new_n4902_;
  assign new_n4904_ = B6209 & B6208;
  assign new_n4905_ = ~new_n1639_ & ~new_n4904_;
  assign new_n4906_ = ~B6208 & ~new_n1637_;
  assign new_n4907_ = B6208 & new_n1637_;
  assign new_n4908_ = ~new_n4906_ & ~new_n4907_;
  assign new_n4909_ = new_n4905_ & ~new_n4908_;
  assign new_n4910_ = ~new_n3708_ & ~new_n4909_;
  assign new_n4911_ = new_n4903_ & ~new_n4910_;
  assign new_n4912_ = ~new_n4903_ & new_n4910_;
  assign new_n4913_ = ~new_n4911_ & ~new_n4912_;
  assign new_n4914_ = B6242 & B6241;
  assign new_n4915_ = ~new_n1652_ & ~new_n4914_;
  assign new_n4916_ = ~B6241 & ~new_n1650_;
  assign new_n4917_ = B6241 & new_n1650_;
  assign new_n4918_ = ~new_n4916_ & ~new_n4917_;
  assign new_n4919_ = new_n4915_ & ~new_n4918_;
  assign new_n4920_ = ~new_n3718_ & ~new_n4919_;
  assign new_n4921_ = B6275 & B6274;
  assign new_n4922_ = ~new_n1662_ & ~new_n4921_;
  assign new_n4923_ = ~B6274 & ~new_n1660_;
  assign new_n4924_ = B6274 & new_n1660_;
  assign new_n4925_ = ~new_n4923_ & ~new_n4924_;
  assign new_n4926_ = new_n4922_ & ~new_n4925_;
  assign new_n4927_ = ~new_n3725_ & ~new_n4926_;
  assign new_n4928_ = new_n4913_ & new_n4927_;
  assign new_n4929_ = B6308 & B6307;
  assign new_n4930_ = ~new_n1673_ & ~new_n4929_;
  assign new_n4931_ = ~B6307 & ~new_n1671_;
  assign new_n4932_ = B6307 & new_n1671_;
  assign new_n4933_ = ~new_n4931_ & ~new_n4932_;
  assign new_n4934_ = new_n4930_ & ~new_n4933_;
  assign new_n4935_ = ~new_n3733_ & ~new_n4934_;
  assign new_n4936_ = new_n4927_ & new_n4935_;
  assign new_n4937_ = ~new_n4928_ & ~new_n4936_;
  assign new_n4938_ = ~new_n4920_ & new_n4937_;
  assign new_n4939_ = new_n4920_ & ~new_n4937_;
  assign new_n4940_ = ~new_n4938_ & ~new_n4939_;
  assign new_n4941_ = ~new_n4913_ & ~new_n4940_;
  assign new_n4942_ = ~new_n4896_ & new_n4941_;
  assign new_n4943_ = new_n4896_ & ~new_n4941_;
  assign new_n4944_ = ~new_n4942_ & ~new_n4943_;
  assign new_n4945_ = B6341 & B6340;
  assign new_n4946_ = ~new_n1692_ & ~new_n4945_;
  assign new_n4947_ = ~B6340 & ~new_n1690_;
  assign new_n4948_ = B6340 & new_n1690_;
  assign new_n4949_ = ~new_n4947_ & ~new_n4948_;
  assign new_n4950_ = new_n4946_ & ~new_n4949_;
  assign new_n4951_ = ~new_n3749_ & ~new_n4950_;
  assign new_n4952_ = B6374 & B6373;
  assign new_n4953_ = ~new_n1702_ & ~new_n4952_;
  assign new_n4954_ = ~B6373 & ~new_n1700_;
  assign new_n4955_ = B6373 & new_n1700_;
  assign new_n4956_ = ~new_n4954_ & ~new_n4955_;
  assign new_n4957_ = new_n4953_ & ~new_n4956_;
  assign new_n4958_ = ~new_n3756_ & ~new_n4957_;
  assign new_n4959_ = new_n4951_ & ~new_n4958_;
  assign new_n4960_ = ~new_n4951_ & new_n4958_;
  assign new_n4961_ = ~new_n4959_ & ~new_n4960_;
  assign new_n4962_ = B6407 & B6406;
  assign new_n4963_ = ~new_n1715_ & ~new_n4962_;
  assign new_n4964_ = ~B6406 & ~new_n1713_;
  assign new_n4965_ = B6406 & new_n1713_;
  assign new_n4966_ = ~new_n4964_ & ~new_n4965_;
  assign new_n4967_ = new_n4963_ & ~new_n4966_;
  assign new_n4968_ = ~new_n3766_ & ~new_n4967_;
  assign new_n4969_ = B6440 & B6439;
  assign new_n4970_ = ~new_n1725_ & ~new_n4969_;
  assign new_n4971_ = ~B6439 & ~new_n1723_;
  assign new_n4972_ = B6439 & new_n1723_;
  assign new_n4973_ = ~new_n4971_ & ~new_n4972_;
  assign new_n4974_ = new_n4970_ & ~new_n4973_;
  assign new_n4975_ = ~new_n3773_ & ~new_n4974_;
  assign new_n4976_ = new_n4961_ & new_n4975_;
  assign new_n4977_ = B6473 & B6472;
  assign new_n4978_ = ~new_n1736_ & ~new_n4977_;
  assign new_n4979_ = ~B6472 & ~new_n1734_;
  assign new_n4980_ = B6472 & new_n1734_;
  assign new_n4981_ = ~new_n4979_ & ~new_n4980_;
  assign new_n4982_ = new_n4978_ & ~new_n4981_;
  assign new_n4983_ = ~new_n3781_ & ~new_n4982_;
  assign new_n4984_ = new_n4975_ & new_n4983_;
  assign new_n4985_ = ~new_n4976_ & ~new_n4984_;
  assign new_n4986_ = ~new_n4968_ & new_n4985_;
  assign new_n4987_ = new_n4968_ & ~new_n4985_;
  assign new_n4988_ = ~new_n4986_ & ~new_n4987_;
  assign new_n4989_ = ~new_n4961_ & ~new_n4988_;
  assign new_n4990_ = B6506 & B6505;
  assign new_n4991_ = ~new_n1752_ & ~new_n4990_;
  assign new_n4992_ = ~B6505 & ~new_n1750_;
  assign new_n4993_ = B6505 & new_n1750_;
  assign new_n4994_ = ~new_n4992_ & ~new_n4993_;
  assign new_n4995_ = new_n4991_ & ~new_n4994_;
  assign new_n4996_ = ~new_n3794_ & ~new_n4995_;
  assign new_n4997_ = B6539 & B6538;
  assign new_n4998_ = ~new_n1762_ & ~new_n4997_;
  assign new_n4999_ = ~B6538 & ~new_n1760_;
  assign new_n5000_ = B6538 & new_n1760_;
  assign new_n5001_ = ~new_n4999_ & ~new_n5000_;
  assign new_n5002_ = new_n4998_ & ~new_n5001_;
  assign new_n5003_ = ~new_n3801_ & ~new_n5002_;
  assign new_n5004_ = new_n4996_ & ~new_n5003_;
  assign new_n5005_ = ~new_n4996_ & new_n5003_;
  assign new_n5006_ = ~new_n5004_ & ~new_n5005_;
  assign new_n5007_ = B6572 & B6571;
  assign new_n5008_ = ~new_n1775_ & ~new_n5007_;
  assign new_n5009_ = ~B6571 & ~new_n1773_;
  assign new_n5010_ = B6571 & new_n1773_;
  assign new_n5011_ = ~new_n5009_ & ~new_n5010_;
  assign new_n5012_ = new_n5008_ & ~new_n5011_;
  assign new_n5013_ = ~new_n3811_ & ~new_n5012_;
  assign new_n5014_ = B6605 & B6604;
  assign new_n5015_ = ~new_n1785_ & ~new_n5014_;
  assign new_n5016_ = ~B6604 & ~new_n1783_;
  assign new_n5017_ = B6604 & new_n1783_;
  assign new_n5018_ = ~new_n5016_ & ~new_n5017_;
  assign new_n5019_ = new_n5015_ & ~new_n5018_;
  assign new_n5020_ = ~new_n3818_ & ~new_n5019_;
  assign new_n5021_ = new_n5006_ & new_n5020_;
  assign new_n5022_ = B6638 & B6637;
  assign new_n5023_ = ~new_n1796_ & ~new_n5022_;
  assign new_n5024_ = ~B6637 & ~new_n1794_;
  assign new_n5025_ = B6637 & new_n1794_;
  assign new_n5026_ = ~new_n5024_ & ~new_n5025_;
  assign new_n5027_ = new_n5023_ & ~new_n5026_;
  assign new_n5028_ = ~new_n3826_ & ~new_n5027_;
  assign new_n5029_ = new_n5020_ & new_n5028_;
  assign new_n5030_ = ~new_n5021_ & ~new_n5029_;
  assign new_n5031_ = ~new_n5013_ & new_n5030_;
  assign new_n5032_ = new_n5013_ & ~new_n5030_;
  assign new_n5033_ = ~new_n5031_ & ~new_n5032_;
  assign new_n5034_ = ~new_n5006_ & ~new_n5033_;
  assign new_n5035_ = new_n4944_ & ~new_n5034_;
  assign new_n5036_ = B6671 & B6670;
  assign new_n5037_ = ~new_n1813_ & ~new_n5036_;
  assign new_n5038_ = ~B6670 & ~new_n1811_;
  assign new_n5039_ = B6670 & new_n1811_;
  assign new_n5040_ = ~new_n5038_ & ~new_n5039_;
  assign new_n5041_ = new_n5037_ & ~new_n5040_;
  assign new_n5042_ = ~new_n3840_ & ~new_n5041_;
  assign new_n5043_ = B6704 & B6703;
  assign new_n5044_ = ~new_n1823_ & ~new_n5043_;
  assign new_n5045_ = ~B6703 & ~new_n1821_;
  assign new_n5046_ = B6703 & new_n1821_;
  assign new_n5047_ = ~new_n5045_ & ~new_n5046_;
  assign new_n5048_ = new_n5044_ & ~new_n5047_;
  assign new_n5049_ = ~new_n3847_ & ~new_n5048_;
  assign new_n5050_ = new_n5042_ & ~new_n5049_;
  assign new_n5051_ = ~new_n5042_ & new_n5049_;
  assign new_n5052_ = ~new_n5050_ & ~new_n5051_;
  assign new_n5053_ = B6737 & B6736;
  assign new_n5054_ = ~new_n1836_ & ~new_n5053_;
  assign new_n5055_ = ~B6736 & ~new_n1834_;
  assign new_n5056_ = B6736 & new_n1834_;
  assign new_n5057_ = ~new_n5055_ & ~new_n5056_;
  assign new_n5058_ = new_n5054_ & ~new_n5057_;
  assign new_n5059_ = ~new_n3857_ & ~new_n5058_;
  assign new_n5060_ = B6770 & B6769;
  assign new_n5061_ = ~new_n1846_ & ~new_n5060_;
  assign new_n5062_ = ~B6769 & ~new_n1844_;
  assign new_n5063_ = B6769 & new_n1844_;
  assign new_n5064_ = ~new_n5062_ & ~new_n5063_;
  assign new_n5065_ = new_n5061_ & ~new_n5064_;
  assign new_n5066_ = ~new_n3864_ & ~new_n5065_;
  assign new_n5067_ = new_n5052_ & new_n5066_;
  assign new_n5068_ = B6803 & B6802;
  assign new_n5069_ = ~new_n1857_ & ~new_n5068_;
  assign new_n5070_ = ~B6802 & ~new_n1855_;
  assign new_n5071_ = B6802 & new_n1855_;
  assign new_n5072_ = ~new_n5070_ & ~new_n5071_;
  assign new_n5073_ = new_n5069_ & ~new_n5072_;
  assign new_n5074_ = ~new_n3872_ & ~new_n5073_;
  assign new_n5075_ = new_n5066_ & new_n5074_;
  assign new_n5076_ = ~new_n5067_ & ~new_n5075_;
  assign new_n5077_ = ~new_n5059_ & new_n5076_;
  assign new_n5078_ = new_n5059_ & ~new_n5076_;
  assign new_n5079_ = ~new_n5077_ & ~new_n5078_;
  assign new_n5080_ = ~new_n5052_ & ~new_n5079_;
  assign new_n5081_ = ~new_n5034_ & ~new_n5080_;
  assign new_n5082_ = ~new_n5035_ & ~new_n5081_;
  assign new_n5083_ = new_n4989_ & new_n5082_;
  assign new_n5084_ = ~new_n4989_ & ~new_n5082_;
  assign new_n5085_ = ~new_n5083_ & ~new_n5084_;
  assign new_n5086_ = ~new_n4944_ & ~new_n5085_;
  assign new_n5087_ = ~new_n4851_ & new_n5086_;
  assign new_n5088_ = new_n4851_ & ~new_n5086_;
  assign new_n5089_ = ~new_n5087_ & ~new_n5088_;
  assign new_n5090_ = B6836 & B6835;
  assign new_n5091_ = ~new_n1882_ & ~new_n5090_;
  assign new_n5092_ = ~B6835 & ~new_n1880_;
  assign new_n5093_ = B6835 & new_n1880_;
  assign new_n5094_ = ~new_n5092_ & ~new_n5093_;
  assign new_n5095_ = new_n5091_ & ~new_n5094_;
  assign new_n5096_ = ~new_n3894_ & ~new_n5095_;
  assign new_n5097_ = B6869 & B6868;
  assign new_n5098_ = ~new_n1892_ & ~new_n5097_;
  assign new_n5099_ = ~B6868 & ~new_n1890_;
  assign new_n5100_ = B6868 & new_n1890_;
  assign new_n5101_ = ~new_n5099_ & ~new_n5100_;
  assign new_n5102_ = new_n5098_ & ~new_n5101_;
  assign new_n5103_ = ~new_n3901_ & ~new_n5102_;
  assign new_n5104_ = new_n5096_ & ~new_n5103_;
  assign new_n5105_ = ~new_n5096_ & new_n5103_;
  assign new_n5106_ = ~new_n5104_ & ~new_n5105_;
  assign new_n5107_ = B6902 & B6901;
  assign new_n5108_ = ~new_n1905_ & ~new_n5107_;
  assign new_n5109_ = ~B6901 & ~new_n1903_;
  assign new_n5110_ = B6901 & new_n1903_;
  assign new_n5111_ = ~new_n5109_ & ~new_n5110_;
  assign new_n5112_ = new_n5108_ & ~new_n5111_;
  assign new_n5113_ = ~new_n3911_ & ~new_n5112_;
  assign new_n5114_ = B6935 & B6934;
  assign new_n5115_ = ~new_n1915_ & ~new_n5114_;
  assign new_n5116_ = ~B6934 & ~new_n1913_;
  assign new_n5117_ = B6934 & new_n1913_;
  assign new_n5118_ = ~new_n5116_ & ~new_n5117_;
  assign new_n5119_ = new_n5115_ & ~new_n5118_;
  assign new_n5120_ = ~new_n3918_ & ~new_n5119_;
  assign new_n5121_ = new_n5106_ & new_n5120_;
  assign new_n5122_ = B6968 & B6967;
  assign new_n5123_ = ~new_n1926_ & ~new_n5122_;
  assign new_n5124_ = ~B6967 & ~new_n1924_;
  assign new_n5125_ = B6967 & new_n1924_;
  assign new_n5126_ = ~new_n5124_ & ~new_n5125_;
  assign new_n5127_ = new_n5123_ & ~new_n5126_;
  assign new_n5128_ = ~new_n3926_ & ~new_n5127_;
  assign new_n5129_ = new_n5120_ & new_n5128_;
  assign new_n5130_ = ~new_n5121_ & ~new_n5129_;
  assign new_n5131_ = ~new_n5113_ & new_n5130_;
  assign new_n5132_ = new_n5113_ & ~new_n5130_;
  assign new_n5133_ = ~new_n5131_ & ~new_n5132_;
  assign new_n5134_ = ~new_n5106_ & ~new_n5133_;
  assign new_n5135_ = B7001 & B7000;
  assign new_n5136_ = ~new_n1942_ & ~new_n5135_;
  assign new_n5137_ = ~B7000 & ~new_n1940_;
  assign new_n5138_ = B7000 & new_n1940_;
  assign new_n5139_ = ~new_n5137_ & ~new_n5138_;
  assign new_n5140_ = new_n5136_ & ~new_n5139_;
  assign new_n5141_ = ~new_n3939_ & ~new_n5140_;
  assign new_n5142_ = B7034 & B7033;
  assign new_n5143_ = ~new_n1952_ & ~new_n5142_;
  assign new_n5144_ = ~B7033 & ~new_n1950_;
  assign new_n5145_ = B7033 & new_n1950_;
  assign new_n5146_ = ~new_n5144_ & ~new_n5145_;
  assign new_n5147_ = new_n5143_ & ~new_n5146_;
  assign new_n5148_ = ~new_n3946_ & ~new_n5147_;
  assign new_n5149_ = new_n5141_ & ~new_n5148_;
  assign new_n5150_ = ~new_n5141_ & new_n5148_;
  assign new_n5151_ = ~new_n5149_ & ~new_n5150_;
  assign new_n5152_ = B7067 & B7066;
  assign new_n5153_ = ~new_n1965_ & ~new_n5152_;
  assign new_n5154_ = ~B7066 & ~new_n1963_;
  assign new_n5155_ = B7066 & new_n1963_;
  assign new_n5156_ = ~new_n5154_ & ~new_n5155_;
  assign new_n5157_ = new_n5153_ & ~new_n5156_;
  assign new_n5158_ = ~new_n3956_ & ~new_n5157_;
  assign new_n5159_ = B7100 & B7099;
  assign new_n5160_ = ~new_n1975_ & ~new_n5159_;
  assign new_n5161_ = ~B7099 & ~new_n1973_;
  assign new_n5162_ = B7099 & new_n1973_;
  assign new_n5163_ = ~new_n5161_ & ~new_n5162_;
  assign new_n5164_ = new_n5160_ & ~new_n5163_;
  assign new_n5165_ = ~new_n3963_ & ~new_n5164_;
  assign new_n5166_ = new_n5151_ & new_n5165_;
  assign new_n5167_ = B7133 & B7132;
  assign new_n5168_ = ~new_n1986_ & ~new_n5167_;
  assign new_n5169_ = ~B7132 & ~new_n1984_;
  assign new_n5170_ = B7132 & new_n1984_;
  assign new_n5171_ = ~new_n5169_ & ~new_n5170_;
  assign new_n5172_ = new_n5168_ & ~new_n5171_;
  assign new_n5173_ = ~new_n3971_ & ~new_n5172_;
  assign new_n5174_ = new_n5165_ & new_n5173_;
  assign new_n5175_ = ~new_n5166_ & ~new_n5174_;
  assign new_n5176_ = ~new_n5158_ & new_n5175_;
  assign new_n5177_ = new_n5158_ & ~new_n5175_;
  assign new_n5178_ = ~new_n5176_ & ~new_n5177_;
  assign new_n5179_ = ~new_n5151_ & ~new_n5178_;
  assign new_n5180_ = ~new_n5134_ & new_n5179_;
  assign new_n5181_ = new_n5134_ & ~new_n5179_;
  assign new_n5182_ = ~new_n5180_ & ~new_n5181_;
  assign new_n5183_ = B7166 & B7165;
  assign new_n5184_ = ~new_n2005_ & ~new_n5183_;
  assign new_n5185_ = ~B7165 & ~new_n2003_;
  assign new_n5186_ = B7165 & new_n2003_;
  assign new_n5187_ = ~new_n5185_ & ~new_n5186_;
  assign new_n5188_ = new_n5184_ & ~new_n5187_;
  assign new_n5189_ = ~new_n3987_ & ~new_n5188_;
  assign new_n5190_ = B7199 & B7198;
  assign new_n5191_ = ~new_n2015_ & ~new_n5190_;
  assign new_n5192_ = ~B7198 & ~new_n2013_;
  assign new_n5193_ = B7198 & new_n2013_;
  assign new_n5194_ = ~new_n5192_ & ~new_n5193_;
  assign new_n5195_ = new_n5191_ & ~new_n5194_;
  assign new_n5196_ = ~new_n3994_ & ~new_n5195_;
  assign new_n5197_ = new_n5189_ & ~new_n5196_;
  assign new_n5198_ = ~new_n5189_ & new_n5196_;
  assign new_n5199_ = ~new_n5197_ & ~new_n5198_;
  assign new_n5200_ = B7232 & B7231;
  assign new_n5201_ = ~new_n2028_ & ~new_n5200_;
  assign new_n5202_ = ~B7231 & ~new_n2026_;
  assign new_n5203_ = B7231 & new_n2026_;
  assign new_n5204_ = ~new_n5202_ & ~new_n5203_;
  assign new_n5205_ = new_n5201_ & ~new_n5204_;
  assign new_n5206_ = ~new_n4004_ & ~new_n5205_;
  assign new_n5207_ = B7265 & B7264;
  assign new_n5208_ = ~new_n2038_ & ~new_n5207_;
  assign new_n5209_ = ~B7264 & ~new_n2036_;
  assign new_n5210_ = B7264 & new_n2036_;
  assign new_n5211_ = ~new_n5209_ & ~new_n5210_;
  assign new_n5212_ = new_n5208_ & ~new_n5211_;
  assign new_n5213_ = ~new_n4011_ & ~new_n5212_;
  assign new_n5214_ = new_n5199_ & new_n5213_;
  assign new_n5215_ = B7298 & B7297;
  assign new_n5216_ = ~new_n2049_ & ~new_n5215_;
  assign new_n5217_ = ~B7297 & ~new_n2047_;
  assign new_n5218_ = B7297 & new_n2047_;
  assign new_n5219_ = ~new_n5217_ & ~new_n5218_;
  assign new_n5220_ = new_n5216_ & ~new_n5219_;
  assign new_n5221_ = ~new_n4019_ & ~new_n5220_;
  assign new_n5222_ = new_n5213_ & new_n5221_;
  assign new_n5223_ = ~new_n5214_ & ~new_n5222_;
  assign new_n5224_ = ~new_n5206_ & new_n5223_;
  assign new_n5225_ = new_n5206_ & ~new_n5223_;
  assign new_n5226_ = ~new_n5224_ & ~new_n5225_;
  assign new_n5227_ = ~new_n5199_ & ~new_n5226_;
  assign new_n5228_ = B7331 & B7330;
  assign new_n5229_ = ~new_n2065_ & ~new_n5228_;
  assign new_n5230_ = ~B7330 & ~new_n2063_;
  assign new_n5231_ = B7330 & new_n2063_;
  assign new_n5232_ = ~new_n5230_ & ~new_n5231_;
  assign new_n5233_ = new_n5229_ & ~new_n5232_;
  assign new_n5234_ = ~new_n4032_ & ~new_n5233_;
  assign new_n5235_ = B7364 & B7363;
  assign new_n5236_ = ~new_n2075_ & ~new_n5235_;
  assign new_n5237_ = ~B7363 & ~new_n2073_;
  assign new_n5238_ = B7363 & new_n2073_;
  assign new_n5239_ = ~new_n5237_ & ~new_n5238_;
  assign new_n5240_ = new_n5236_ & ~new_n5239_;
  assign new_n5241_ = ~new_n4039_ & ~new_n5240_;
  assign new_n5242_ = new_n5234_ & ~new_n5241_;
  assign new_n5243_ = ~new_n5234_ & new_n5241_;
  assign new_n5244_ = ~new_n5242_ & ~new_n5243_;
  assign new_n5245_ = B7397 & B7396;
  assign new_n5246_ = ~new_n2088_ & ~new_n5245_;
  assign new_n5247_ = ~B7396 & ~new_n2086_;
  assign new_n5248_ = B7396 & new_n2086_;
  assign new_n5249_ = ~new_n5247_ & ~new_n5248_;
  assign new_n5250_ = new_n5246_ & ~new_n5249_;
  assign new_n5251_ = ~new_n4049_ & ~new_n5250_;
  assign new_n5252_ = B7430 & B7429;
  assign new_n5253_ = ~new_n2098_ & ~new_n5252_;
  assign new_n5254_ = ~B7429 & ~new_n2096_;
  assign new_n5255_ = B7429 & new_n2096_;
  assign new_n5256_ = ~new_n5254_ & ~new_n5255_;
  assign new_n5257_ = new_n5253_ & ~new_n5256_;
  assign new_n5258_ = ~new_n4056_ & ~new_n5257_;
  assign new_n5259_ = new_n5244_ & new_n5258_;
  assign new_n5260_ = B7463 & B7462;
  assign new_n5261_ = ~new_n2109_ & ~new_n5260_;
  assign new_n5262_ = ~B7462 & ~new_n2107_;
  assign new_n5263_ = B7462 & new_n2107_;
  assign new_n5264_ = ~new_n5262_ & ~new_n5263_;
  assign new_n5265_ = new_n5261_ & ~new_n5264_;
  assign new_n5266_ = ~new_n4064_ & ~new_n5265_;
  assign new_n5267_ = new_n5258_ & new_n5266_;
  assign new_n5268_ = ~new_n5259_ & ~new_n5267_;
  assign new_n5269_ = ~new_n5251_ & new_n5268_;
  assign new_n5270_ = new_n5251_ & ~new_n5268_;
  assign new_n5271_ = ~new_n5269_ & ~new_n5270_;
  assign new_n5272_ = ~new_n5244_ & ~new_n5271_;
  assign new_n5273_ = new_n5182_ & ~new_n5272_;
  assign new_n5274_ = B7496 & B7495;
  assign new_n5275_ = ~new_n2126_ & ~new_n5274_;
  assign new_n5276_ = ~B7495 & ~new_n2124_;
  assign new_n5277_ = B7495 & new_n2124_;
  assign new_n5278_ = ~new_n5276_ & ~new_n5277_;
  assign new_n5279_ = new_n5275_ & ~new_n5278_;
  assign new_n5280_ = ~new_n4078_ & ~new_n5279_;
  assign new_n5281_ = B7529 & B7528;
  assign new_n5282_ = ~new_n2136_ & ~new_n5281_;
  assign new_n5283_ = ~B7528 & ~new_n2134_;
  assign new_n5284_ = B7528 & new_n2134_;
  assign new_n5285_ = ~new_n5283_ & ~new_n5284_;
  assign new_n5286_ = new_n5282_ & ~new_n5285_;
  assign new_n5287_ = ~new_n4085_ & ~new_n5286_;
  assign new_n5288_ = new_n5280_ & ~new_n5287_;
  assign new_n5289_ = ~new_n5280_ & new_n5287_;
  assign new_n5290_ = ~new_n5288_ & ~new_n5289_;
  assign new_n5291_ = B7562 & B7561;
  assign new_n5292_ = ~new_n2149_ & ~new_n5291_;
  assign new_n5293_ = ~B7561 & ~new_n2147_;
  assign new_n5294_ = B7561 & new_n2147_;
  assign new_n5295_ = ~new_n5293_ & ~new_n5294_;
  assign new_n5296_ = new_n5292_ & ~new_n5295_;
  assign new_n5297_ = ~new_n4095_ & ~new_n5296_;
  assign new_n5298_ = B7595 & B7594;
  assign new_n5299_ = ~new_n2159_ & ~new_n5298_;
  assign new_n5300_ = ~B7594 & ~new_n2157_;
  assign new_n5301_ = B7594 & new_n2157_;
  assign new_n5302_ = ~new_n5300_ & ~new_n5301_;
  assign new_n5303_ = new_n5299_ & ~new_n5302_;
  assign new_n5304_ = ~new_n4102_ & ~new_n5303_;
  assign new_n5305_ = new_n5290_ & new_n5304_;
  assign new_n5306_ = B7628 & B7627;
  assign new_n5307_ = ~new_n2170_ & ~new_n5306_;
  assign new_n5308_ = ~B7627 & ~new_n2168_;
  assign new_n5309_ = B7627 & new_n2168_;
  assign new_n5310_ = ~new_n5308_ & ~new_n5309_;
  assign new_n5311_ = new_n5307_ & ~new_n5310_;
  assign new_n5312_ = ~new_n4110_ & ~new_n5311_;
  assign new_n5313_ = new_n5304_ & new_n5312_;
  assign new_n5314_ = ~new_n5305_ & ~new_n5313_;
  assign new_n5315_ = ~new_n5297_ & new_n5314_;
  assign new_n5316_ = new_n5297_ & ~new_n5314_;
  assign new_n5317_ = ~new_n5315_ & ~new_n5316_;
  assign new_n5318_ = ~new_n5290_ & ~new_n5317_;
  assign new_n5319_ = ~new_n5272_ & ~new_n5318_;
  assign new_n5320_ = ~new_n5273_ & ~new_n5319_;
  assign new_n5321_ = new_n5227_ & new_n5320_;
  assign new_n5322_ = ~new_n5227_ & ~new_n5320_;
  assign new_n5323_ = ~new_n5321_ & ~new_n5322_;
  assign new_n5324_ = ~new_n5182_ & ~new_n5323_;
  assign new_n5325_ = B7661 & B7660;
  assign new_n5326_ = ~new_n2192_ & ~new_n5325_;
  assign new_n5327_ = ~B7660 & ~new_n2190_;
  assign new_n5328_ = B7660 & new_n2190_;
  assign new_n5329_ = ~new_n5327_ & ~new_n5328_;
  assign new_n5330_ = new_n5326_ & ~new_n5329_;
  assign new_n5331_ = ~new_n4129_ & ~new_n5330_;
  assign new_n5332_ = B7694 & B7693;
  assign new_n5333_ = ~new_n2202_ & ~new_n5332_;
  assign new_n5334_ = ~B7693 & ~new_n2200_;
  assign new_n5335_ = B7693 & new_n2200_;
  assign new_n5336_ = ~new_n5334_ & ~new_n5335_;
  assign new_n5337_ = new_n5333_ & ~new_n5336_;
  assign new_n5338_ = ~new_n4136_ & ~new_n5337_;
  assign new_n5339_ = new_n5331_ & ~new_n5338_;
  assign new_n5340_ = ~new_n5331_ & new_n5338_;
  assign new_n5341_ = ~new_n5339_ & ~new_n5340_;
  assign new_n5342_ = B7727 & B7726;
  assign new_n5343_ = ~new_n2215_ & ~new_n5342_;
  assign new_n5344_ = ~B7726 & ~new_n2213_;
  assign new_n5345_ = B7726 & new_n2213_;
  assign new_n5346_ = ~new_n5344_ & ~new_n5345_;
  assign new_n5347_ = new_n5343_ & ~new_n5346_;
  assign new_n5348_ = ~new_n4146_ & ~new_n5347_;
  assign new_n5349_ = B7760 & B7759;
  assign new_n5350_ = ~new_n2225_ & ~new_n5349_;
  assign new_n5351_ = ~B7759 & ~new_n2223_;
  assign new_n5352_ = B7759 & new_n2223_;
  assign new_n5353_ = ~new_n5351_ & ~new_n5352_;
  assign new_n5354_ = new_n5350_ & ~new_n5353_;
  assign new_n5355_ = ~new_n4153_ & ~new_n5354_;
  assign new_n5356_ = new_n5341_ & new_n5355_;
  assign new_n5357_ = B7793 & B7792;
  assign new_n5358_ = ~new_n2236_ & ~new_n5357_;
  assign new_n5359_ = ~B7792 & ~new_n2234_;
  assign new_n5360_ = B7792 & new_n2234_;
  assign new_n5361_ = ~new_n5359_ & ~new_n5360_;
  assign new_n5362_ = new_n5358_ & ~new_n5361_;
  assign new_n5363_ = ~new_n4161_ & ~new_n5362_;
  assign new_n5364_ = new_n5355_ & new_n5363_;
  assign new_n5365_ = ~new_n5356_ & ~new_n5364_;
  assign new_n5366_ = ~new_n5348_ & new_n5365_;
  assign new_n5367_ = new_n5348_ & ~new_n5365_;
  assign new_n5368_ = ~new_n5366_ & ~new_n5367_;
  assign new_n5369_ = ~new_n5341_ & ~new_n5368_;
  assign new_n5370_ = B7826 & B7825;
  assign new_n5371_ = ~new_n2252_ & ~new_n5370_;
  assign new_n5372_ = ~B7825 & ~new_n2250_;
  assign new_n5373_ = B7825 & new_n2250_;
  assign new_n5374_ = ~new_n5372_ & ~new_n5373_;
  assign new_n5375_ = new_n5371_ & ~new_n5374_;
  assign new_n5376_ = ~new_n4174_ & ~new_n5375_;
  assign new_n5377_ = B7859 & B7858;
  assign new_n5378_ = ~new_n2262_ & ~new_n5377_;
  assign new_n5379_ = ~B7858 & ~new_n2260_;
  assign new_n5380_ = B7858 & new_n2260_;
  assign new_n5381_ = ~new_n5379_ & ~new_n5380_;
  assign new_n5382_ = new_n5378_ & ~new_n5381_;
  assign new_n5383_ = ~new_n4181_ & ~new_n5382_;
  assign new_n5384_ = new_n5376_ & ~new_n5383_;
  assign new_n5385_ = ~new_n5376_ & new_n5383_;
  assign new_n5386_ = ~new_n5384_ & ~new_n5385_;
  assign new_n5387_ = B7892 & B7891;
  assign new_n5388_ = ~new_n2275_ & ~new_n5387_;
  assign new_n5389_ = ~B7891 & ~new_n2273_;
  assign new_n5390_ = B7891 & new_n2273_;
  assign new_n5391_ = ~new_n5389_ & ~new_n5390_;
  assign new_n5392_ = new_n5388_ & ~new_n5391_;
  assign new_n5393_ = ~new_n4191_ & ~new_n5392_;
  assign new_n5394_ = B7925 & B7924;
  assign new_n5395_ = ~new_n2285_ & ~new_n5394_;
  assign new_n5396_ = ~B7924 & ~new_n2283_;
  assign new_n5397_ = B7924 & new_n2283_;
  assign new_n5398_ = ~new_n5396_ & ~new_n5397_;
  assign new_n5399_ = new_n5395_ & ~new_n5398_;
  assign new_n5400_ = ~new_n4198_ & ~new_n5399_;
  assign new_n5401_ = new_n5386_ & new_n5400_;
  assign new_n5402_ = B7958 & B7957;
  assign new_n5403_ = ~new_n2296_ & ~new_n5402_;
  assign new_n5404_ = ~B7957 & ~new_n2294_;
  assign new_n5405_ = B7957 & new_n2294_;
  assign new_n5406_ = ~new_n5404_ & ~new_n5405_;
  assign new_n5407_ = new_n5403_ & ~new_n5406_;
  assign new_n5408_ = ~new_n4206_ & ~new_n5407_;
  assign new_n5409_ = new_n5400_ & new_n5408_;
  assign new_n5410_ = ~new_n5401_ & ~new_n5409_;
  assign new_n5411_ = ~new_n5393_ & new_n5410_;
  assign new_n5412_ = new_n5393_ & ~new_n5410_;
  assign new_n5413_ = ~new_n5411_ & ~new_n5412_;
  assign new_n5414_ = ~new_n5386_ & ~new_n5413_;
  assign new_n5415_ = ~new_n5369_ & new_n5414_;
  assign new_n5416_ = new_n5369_ & ~new_n5414_;
  assign new_n5417_ = ~new_n5415_ & ~new_n5416_;
  assign new_n5418_ = B7991 & B7990;
  assign new_n5419_ = ~new_n2315_ & ~new_n5418_;
  assign new_n5420_ = ~B7990 & ~new_n2313_;
  assign new_n5421_ = B7990 & new_n2313_;
  assign new_n5422_ = ~new_n5420_ & ~new_n5421_;
  assign new_n5423_ = new_n5419_ & ~new_n5422_;
  assign new_n5424_ = ~new_n4222_ & ~new_n5423_;
  assign new_n5425_ = B8024 & B8023;
  assign new_n5426_ = ~new_n2325_ & ~new_n5425_;
  assign new_n5427_ = ~B8023 & ~new_n2323_;
  assign new_n5428_ = B8023 & new_n2323_;
  assign new_n5429_ = ~new_n5427_ & ~new_n5428_;
  assign new_n5430_ = new_n5426_ & ~new_n5429_;
  assign new_n5431_ = ~new_n4229_ & ~new_n5430_;
  assign new_n5432_ = new_n5424_ & ~new_n5431_;
  assign new_n5433_ = ~new_n5424_ & new_n5431_;
  assign new_n5434_ = ~new_n5432_ & ~new_n5433_;
  assign new_n5435_ = B8057 & B8056;
  assign new_n5436_ = ~new_n2338_ & ~new_n5435_;
  assign new_n5437_ = ~B8056 & ~new_n2336_;
  assign new_n5438_ = B8056 & new_n2336_;
  assign new_n5439_ = ~new_n5437_ & ~new_n5438_;
  assign new_n5440_ = new_n5436_ & ~new_n5439_;
  assign new_n5441_ = ~new_n4239_ & ~new_n5440_;
  assign new_n5442_ = B8090 & B8089;
  assign new_n5443_ = ~new_n2348_ & ~new_n5442_;
  assign new_n5444_ = ~B8089 & ~new_n2346_;
  assign new_n5445_ = B8089 & new_n2346_;
  assign new_n5446_ = ~new_n5444_ & ~new_n5445_;
  assign new_n5447_ = new_n5443_ & ~new_n5446_;
  assign new_n5448_ = ~new_n4246_ & ~new_n5447_;
  assign new_n5449_ = new_n5434_ & new_n5448_;
  assign new_n5450_ = B8123 & B8122;
  assign new_n5451_ = ~new_n2359_ & ~new_n5450_;
  assign new_n5452_ = ~B8122 & ~new_n2357_;
  assign new_n5453_ = B8122 & new_n2357_;
  assign new_n5454_ = ~new_n5452_ & ~new_n5453_;
  assign new_n5455_ = new_n5451_ & ~new_n5454_;
  assign new_n5456_ = ~new_n4254_ & ~new_n5455_;
  assign new_n5457_ = new_n5448_ & new_n5456_;
  assign new_n5458_ = ~new_n5449_ & ~new_n5457_;
  assign new_n5459_ = ~new_n5441_ & new_n5458_;
  assign new_n5460_ = new_n5441_ & ~new_n5458_;
  assign new_n5461_ = ~new_n5459_ & ~new_n5460_;
  assign new_n5462_ = ~new_n5434_ & ~new_n5461_;
  assign new_n5463_ = B8156 & B8155;
  assign new_n5464_ = ~new_n2375_ & ~new_n5463_;
  assign new_n5465_ = ~B8155 & ~new_n2373_;
  assign new_n5466_ = B8155 & new_n2373_;
  assign new_n5467_ = ~new_n5465_ & ~new_n5466_;
  assign new_n5468_ = new_n5464_ & ~new_n5467_;
  assign new_n5469_ = ~new_n4267_ & ~new_n5468_;
  assign new_n5470_ = B8189 & B8188;
  assign new_n5471_ = ~new_n2385_ & ~new_n5470_;
  assign new_n5472_ = ~B8188 & ~new_n2383_;
  assign new_n5473_ = B8188 & new_n2383_;
  assign new_n5474_ = ~new_n5472_ & ~new_n5473_;
  assign new_n5475_ = new_n5471_ & ~new_n5474_;
  assign new_n5476_ = ~new_n4274_ & ~new_n5475_;
  assign new_n5477_ = new_n5469_ & ~new_n5476_;
  assign new_n5478_ = ~new_n5469_ & new_n5476_;
  assign new_n5479_ = ~new_n5477_ & ~new_n5478_;
  assign new_n5480_ = B8222 & B8221;
  assign new_n5481_ = ~new_n2398_ & ~new_n5480_;
  assign new_n5482_ = ~B8221 & ~new_n2396_;
  assign new_n5483_ = B8221 & new_n2396_;
  assign new_n5484_ = ~new_n5482_ & ~new_n5483_;
  assign new_n5485_ = new_n5481_ & ~new_n5484_;
  assign new_n5486_ = ~new_n4284_ & ~new_n5485_;
  assign new_n5487_ = B8255 & B8254;
  assign new_n5488_ = ~new_n2408_ & ~new_n5487_;
  assign new_n5489_ = ~B8254 & ~new_n2406_;
  assign new_n5490_ = B8254 & new_n2406_;
  assign new_n5491_ = ~new_n5489_ & ~new_n5490_;
  assign new_n5492_ = new_n5488_ & ~new_n5491_;
  assign new_n5493_ = ~new_n4291_ & ~new_n5492_;
  assign new_n5494_ = new_n5479_ & new_n5493_;
  assign new_n5495_ = B8288 & B8287;
  assign new_n5496_ = ~new_n2419_ & ~new_n5495_;
  assign new_n5497_ = ~B8287 & ~new_n2417_;
  assign new_n5498_ = B8287 & new_n2417_;
  assign new_n5499_ = ~new_n5497_ & ~new_n5498_;
  assign new_n5500_ = new_n5496_ & ~new_n5499_;
  assign new_n5501_ = ~new_n4299_ & ~new_n5500_;
  assign new_n5502_ = new_n5493_ & new_n5501_;
  assign new_n5503_ = ~new_n5494_ & ~new_n5502_;
  assign new_n5504_ = ~new_n5486_ & new_n5503_;
  assign new_n5505_ = new_n5486_ & ~new_n5503_;
  assign new_n5506_ = ~new_n5504_ & ~new_n5505_;
  assign new_n5507_ = ~new_n5479_ & ~new_n5506_;
  assign new_n5508_ = new_n5417_ & ~new_n5507_;
  assign new_n5509_ = B8321 & B8320;
  assign new_n5510_ = ~new_n2436_ & ~new_n5509_;
  assign new_n5511_ = ~B8320 & ~new_n2434_;
  assign new_n5512_ = B8320 & new_n2434_;
  assign new_n5513_ = ~new_n5511_ & ~new_n5512_;
  assign new_n5514_ = new_n5510_ & ~new_n5513_;
  assign new_n5515_ = ~new_n4313_ & ~new_n5514_;
  assign new_n5516_ = B8354 & B8353;
  assign new_n5517_ = ~new_n2446_ & ~new_n5516_;
  assign new_n5518_ = ~B8353 & ~new_n2444_;
  assign new_n5519_ = B8353 & new_n2444_;
  assign new_n5520_ = ~new_n5518_ & ~new_n5519_;
  assign new_n5521_ = new_n5517_ & ~new_n5520_;
  assign new_n5522_ = ~new_n4320_ & ~new_n5521_;
  assign new_n5523_ = new_n5515_ & ~new_n5522_;
  assign new_n5524_ = ~new_n5515_ & new_n5522_;
  assign new_n5525_ = ~new_n5523_ & ~new_n5524_;
  assign new_n5526_ = B8387 & B8386;
  assign new_n5527_ = ~new_n2459_ & ~new_n5526_;
  assign new_n5528_ = ~B8386 & ~new_n2457_;
  assign new_n5529_ = B8386 & new_n2457_;
  assign new_n5530_ = ~new_n5528_ & ~new_n5529_;
  assign new_n5531_ = new_n5527_ & ~new_n5530_;
  assign new_n5532_ = ~new_n4330_ & ~new_n5531_;
  assign new_n5533_ = B8420 & B8419;
  assign new_n5534_ = ~new_n2469_ & ~new_n5533_;
  assign new_n5535_ = ~B8419 & ~new_n2467_;
  assign new_n5536_ = B8419 & new_n2467_;
  assign new_n5537_ = ~new_n5535_ & ~new_n5536_;
  assign new_n5538_ = new_n5534_ & ~new_n5537_;
  assign new_n5539_ = ~new_n4337_ & ~new_n5538_;
  assign new_n5540_ = new_n5525_ & new_n5539_;
  assign new_n5541_ = B8453 & B8452;
  assign new_n5542_ = ~new_n2480_ & ~new_n5541_;
  assign new_n5543_ = ~B8452 & ~new_n2478_;
  assign new_n5544_ = B8452 & new_n2478_;
  assign new_n5545_ = ~new_n5543_ & ~new_n5544_;
  assign new_n5546_ = new_n5542_ & ~new_n5545_;
  assign new_n5547_ = ~new_n4345_ & ~new_n5546_;
  assign new_n5548_ = new_n5539_ & new_n5547_;
  assign new_n5549_ = ~new_n5540_ & ~new_n5548_;
  assign new_n5550_ = ~new_n5532_ & new_n5549_;
  assign new_n5551_ = new_n5532_ & ~new_n5549_;
  assign new_n5552_ = ~new_n5550_ & ~new_n5551_;
  assign new_n5553_ = ~new_n5525_ & ~new_n5552_;
  assign new_n5554_ = ~new_n5507_ & ~new_n5553_;
  assign new_n5555_ = ~new_n5508_ & ~new_n5554_;
  assign new_n5556_ = new_n5462_ & new_n5555_;
  assign new_n5557_ = ~new_n5462_ & ~new_n5555_;
  assign new_n5558_ = ~new_n5556_ & ~new_n5557_;
  assign new_n5559_ = ~new_n5417_ & ~new_n5558_;
  assign new_n5560_ = new_n5089_ & ~new_n5559_;
  assign new_n5561_ = B8486 & B8485;
  assign new_n5562_ = ~new_n2503_ & ~new_n5561_;
  assign new_n5563_ = ~B8485 & ~new_n2501_;
  assign new_n5564_ = B8485 & new_n2501_;
  assign new_n5565_ = ~new_n5563_ & ~new_n5564_;
  assign new_n5566_ = new_n5562_ & ~new_n5565_;
  assign new_n5567_ = ~new_n4365_ & ~new_n5566_;
  assign new_n5568_ = B8519 & B8518;
  assign new_n5569_ = ~new_n2513_ & ~new_n5568_;
  assign new_n5570_ = ~B8518 & ~new_n2511_;
  assign new_n5571_ = B8518 & new_n2511_;
  assign new_n5572_ = ~new_n5570_ & ~new_n5571_;
  assign new_n5573_ = new_n5569_ & ~new_n5572_;
  assign new_n5574_ = ~new_n4372_ & ~new_n5573_;
  assign new_n5575_ = new_n5567_ & ~new_n5574_;
  assign new_n5576_ = ~new_n5567_ & new_n5574_;
  assign new_n5577_ = ~new_n5575_ & ~new_n5576_;
  assign new_n5578_ = B8552 & B8551;
  assign new_n5579_ = ~new_n2526_ & ~new_n5578_;
  assign new_n5580_ = ~B8551 & ~new_n2524_;
  assign new_n5581_ = B8551 & new_n2524_;
  assign new_n5582_ = ~new_n5580_ & ~new_n5581_;
  assign new_n5583_ = new_n5579_ & ~new_n5582_;
  assign new_n5584_ = ~new_n4382_ & ~new_n5583_;
  assign new_n5585_ = B8585 & B8584;
  assign new_n5586_ = ~new_n2536_ & ~new_n5585_;
  assign new_n5587_ = ~B8584 & ~new_n2534_;
  assign new_n5588_ = B8584 & new_n2534_;
  assign new_n5589_ = ~new_n5587_ & ~new_n5588_;
  assign new_n5590_ = new_n5586_ & ~new_n5589_;
  assign new_n5591_ = ~new_n4389_ & ~new_n5590_;
  assign new_n5592_ = new_n5577_ & new_n5591_;
  assign new_n5593_ = B8618 & B8617;
  assign new_n5594_ = ~new_n2547_ & ~new_n5593_;
  assign new_n5595_ = ~B8617 & ~new_n2545_;
  assign new_n5596_ = B8617 & new_n2545_;
  assign new_n5597_ = ~new_n5595_ & ~new_n5596_;
  assign new_n5598_ = new_n5594_ & ~new_n5597_;
  assign new_n5599_ = ~new_n4397_ & ~new_n5598_;
  assign new_n5600_ = new_n5591_ & new_n5599_;
  assign new_n5601_ = ~new_n5592_ & ~new_n5600_;
  assign new_n5602_ = ~new_n5584_ & new_n5601_;
  assign new_n5603_ = new_n5584_ & ~new_n5601_;
  assign new_n5604_ = ~new_n5602_ & ~new_n5603_;
  assign new_n5605_ = ~new_n5577_ & ~new_n5604_;
  assign new_n5606_ = B8651 & B8650;
  assign new_n5607_ = ~new_n2563_ & ~new_n5606_;
  assign new_n5608_ = ~B8650 & ~new_n2561_;
  assign new_n5609_ = B8650 & new_n2561_;
  assign new_n5610_ = ~new_n5608_ & ~new_n5609_;
  assign new_n5611_ = new_n5607_ & ~new_n5610_;
  assign new_n5612_ = ~new_n4410_ & ~new_n5611_;
  assign new_n5613_ = B8684 & B8683;
  assign new_n5614_ = ~new_n2573_ & ~new_n5613_;
  assign new_n5615_ = ~B8683 & ~new_n2571_;
  assign new_n5616_ = B8683 & new_n2571_;
  assign new_n5617_ = ~new_n5615_ & ~new_n5616_;
  assign new_n5618_ = new_n5614_ & ~new_n5617_;
  assign new_n5619_ = ~new_n4417_ & ~new_n5618_;
  assign new_n5620_ = new_n5612_ & ~new_n5619_;
  assign new_n5621_ = ~new_n5612_ & new_n5619_;
  assign new_n5622_ = ~new_n5620_ & ~new_n5621_;
  assign new_n5623_ = B8717 & B8716;
  assign new_n5624_ = ~new_n2586_ & ~new_n5623_;
  assign new_n5625_ = ~B8716 & ~new_n2584_;
  assign new_n5626_ = B8716 & new_n2584_;
  assign new_n5627_ = ~new_n5625_ & ~new_n5626_;
  assign new_n5628_ = new_n5624_ & ~new_n5627_;
  assign new_n5629_ = ~new_n4427_ & ~new_n5628_;
  assign new_n5630_ = B8750 & B8749;
  assign new_n5631_ = ~new_n2596_ & ~new_n5630_;
  assign new_n5632_ = ~B8749 & ~new_n2594_;
  assign new_n5633_ = B8749 & new_n2594_;
  assign new_n5634_ = ~new_n5632_ & ~new_n5633_;
  assign new_n5635_ = new_n5631_ & ~new_n5634_;
  assign new_n5636_ = ~new_n4434_ & ~new_n5635_;
  assign new_n5637_ = new_n5622_ & new_n5636_;
  assign new_n5638_ = B8783 & B8782;
  assign new_n5639_ = ~new_n2607_ & ~new_n5638_;
  assign new_n5640_ = ~B8782 & ~new_n2605_;
  assign new_n5641_ = B8782 & new_n2605_;
  assign new_n5642_ = ~new_n5640_ & ~new_n5641_;
  assign new_n5643_ = new_n5639_ & ~new_n5642_;
  assign new_n5644_ = ~new_n4442_ & ~new_n5643_;
  assign new_n5645_ = new_n5636_ & new_n5644_;
  assign new_n5646_ = ~new_n5637_ & ~new_n5645_;
  assign new_n5647_ = ~new_n5629_ & new_n5646_;
  assign new_n5648_ = new_n5629_ & ~new_n5646_;
  assign new_n5649_ = ~new_n5647_ & ~new_n5648_;
  assign new_n5650_ = ~new_n5622_ & ~new_n5649_;
  assign new_n5651_ = ~new_n5605_ & new_n5650_;
  assign new_n5652_ = new_n5605_ & ~new_n5650_;
  assign new_n5653_ = ~new_n5651_ & ~new_n5652_;
  assign new_n5654_ = B8816 & B8815;
  assign new_n5655_ = ~new_n2626_ & ~new_n5654_;
  assign new_n5656_ = ~B8815 & ~new_n2624_;
  assign new_n5657_ = B8815 & new_n2624_;
  assign new_n5658_ = ~new_n5656_ & ~new_n5657_;
  assign new_n5659_ = new_n5655_ & ~new_n5658_;
  assign new_n5660_ = ~new_n4458_ & ~new_n5659_;
  assign new_n5661_ = B8849 & B8848;
  assign new_n5662_ = ~new_n2636_ & ~new_n5661_;
  assign new_n5663_ = ~B8848 & ~new_n2634_;
  assign new_n5664_ = B8848 & new_n2634_;
  assign new_n5665_ = ~new_n5663_ & ~new_n5664_;
  assign new_n5666_ = new_n5662_ & ~new_n5665_;
  assign new_n5667_ = ~new_n4465_ & ~new_n5666_;
  assign new_n5668_ = new_n5660_ & ~new_n5667_;
  assign new_n5669_ = ~new_n5660_ & new_n5667_;
  assign new_n5670_ = ~new_n5668_ & ~new_n5669_;
  assign new_n5671_ = B8882 & B8881;
  assign new_n5672_ = ~new_n2649_ & ~new_n5671_;
  assign new_n5673_ = ~B8881 & ~new_n2647_;
  assign new_n5674_ = B8881 & new_n2647_;
  assign new_n5675_ = ~new_n5673_ & ~new_n5674_;
  assign new_n5676_ = new_n5672_ & ~new_n5675_;
  assign new_n5677_ = ~new_n4475_ & ~new_n5676_;
  assign new_n5678_ = B8915 & B8914;
  assign new_n5679_ = ~new_n2659_ & ~new_n5678_;
  assign new_n5680_ = ~B8914 & ~new_n2657_;
  assign new_n5681_ = B8914 & new_n2657_;
  assign new_n5682_ = ~new_n5680_ & ~new_n5681_;
  assign new_n5683_ = new_n5679_ & ~new_n5682_;
  assign new_n5684_ = ~new_n4482_ & ~new_n5683_;
  assign new_n5685_ = new_n5670_ & new_n5684_;
  assign new_n5686_ = B8948 & B8947;
  assign new_n5687_ = ~new_n2670_ & ~new_n5686_;
  assign new_n5688_ = ~B8947 & ~new_n2668_;
  assign new_n5689_ = B8947 & new_n2668_;
  assign new_n5690_ = ~new_n5688_ & ~new_n5689_;
  assign new_n5691_ = new_n5687_ & ~new_n5690_;
  assign new_n5692_ = ~new_n4490_ & ~new_n5691_;
  assign new_n5693_ = new_n5684_ & new_n5692_;
  assign new_n5694_ = ~new_n5685_ & ~new_n5693_;
  assign new_n5695_ = ~new_n5677_ & new_n5694_;
  assign new_n5696_ = new_n5677_ & ~new_n5694_;
  assign new_n5697_ = ~new_n5695_ & ~new_n5696_;
  assign new_n5698_ = ~new_n5670_ & ~new_n5697_;
  assign new_n5699_ = B8981 & B8980;
  assign new_n5700_ = ~new_n2686_ & ~new_n5699_;
  assign new_n5701_ = ~B8980 & ~new_n2684_;
  assign new_n5702_ = B8980 & new_n2684_;
  assign new_n5703_ = ~new_n5701_ & ~new_n5702_;
  assign new_n5704_ = new_n5700_ & ~new_n5703_;
  assign new_n5705_ = ~new_n4503_ & ~new_n5704_;
  assign new_n5706_ = B9014 & B9013;
  assign new_n5707_ = ~new_n2696_ & ~new_n5706_;
  assign new_n5708_ = ~B9013 & ~new_n2694_;
  assign new_n5709_ = B9013 & new_n2694_;
  assign new_n5710_ = ~new_n5708_ & ~new_n5709_;
  assign new_n5711_ = new_n5707_ & ~new_n5710_;
  assign new_n5712_ = ~new_n4510_ & ~new_n5711_;
  assign new_n5713_ = new_n5705_ & ~new_n5712_;
  assign new_n5714_ = ~new_n5705_ & new_n5712_;
  assign new_n5715_ = ~new_n5713_ & ~new_n5714_;
  assign new_n5716_ = B9047 & B9046;
  assign new_n5717_ = ~new_n2709_ & ~new_n5716_;
  assign new_n5718_ = ~B9046 & ~new_n2707_;
  assign new_n5719_ = B9046 & new_n2707_;
  assign new_n5720_ = ~new_n5718_ & ~new_n5719_;
  assign new_n5721_ = new_n5717_ & ~new_n5720_;
  assign new_n5722_ = ~new_n4520_ & ~new_n5721_;
  assign new_n5723_ = B9080 & B9079;
  assign new_n5724_ = ~new_n2719_ & ~new_n5723_;
  assign new_n5725_ = ~B9079 & ~new_n2717_;
  assign new_n5726_ = B9079 & new_n2717_;
  assign new_n5727_ = ~new_n5725_ & ~new_n5726_;
  assign new_n5728_ = new_n5724_ & ~new_n5727_;
  assign new_n5729_ = ~new_n4527_ & ~new_n5728_;
  assign new_n5730_ = new_n5715_ & new_n5729_;
  assign new_n5731_ = B9113 & B9112;
  assign new_n5732_ = ~new_n2730_ & ~new_n5731_;
  assign new_n5733_ = ~B9112 & ~new_n2728_;
  assign new_n5734_ = B9112 & new_n2728_;
  assign new_n5735_ = ~new_n5733_ & ~new_n5734_;
  assign new_n5736_ = new_n5732_ & ~new_n5735_;
  assign new_n5737_ = ~new_n4535_ & ~new_n5736_;
  assign new_n5738_ = new_n5729_ & new_n5737_;
  assign new_n5739_ = ~new_n5730_ & ~new_n5738_;
  assign new_n5740_ = ~new_n5722_ & new_n5739_;
  assign new_n5741_ = new_n5722_ & ~new_n5739_;
  assign new_n5742_ = ~new_n5740_ & ~new_n5741_;
  assign new_n5743_ = ~new_n5715_ & ~new_n5742_;
  assign new_n5744_ = new_n5653_ & ~new_n5743_;
  assign new_n5745_ = B9146 & B9145;
  assign new_n5746_ = ~new_n2747_ & ~new_n5745_;
  assign new_n5747_ = ~B9145 & ~new_n2745_;
  assign new_n5748_ = B9145 & new_n2745_;
  assign new_n5749_ = ~new_n5747_ & ~new_n5748_;
  assign new_n5750_ = new_n5746_ & ~new_n5749_;
  assign new_n5751_ = ~new_n4549_ & ~new_n5750_;
  assign new_n5752_ = B9179 & B9178;
  assign new_n5753_ = ~new_n2757_ & ~new_n5752_;
  assign new_n5754_ = ~B9178 & ~new_n2755_;
  assign new_n5755_ = B9178 & new_n2755_;
  assign new_n5756_ = ~new_n5754_ & ~new_n5755_;
  assign new_n5757_ = new_n5753_ & ~new_n5756_;
  assign new_n5758_ = ~new_n4556_ & ~new_n5757_;
  assign new_n5759_ = new_n5751_ & ~new_n5758_;
  assign new_n5760_ = ~new_n5751_ & new_n5758_;
  assign new_n5761_ = ~new_n5759_ & ~new_n5760_;
  assign new_n5762_ = B9212 & B9211;
  assign new_n5763_ = ~new_n2770_ & ~new_n5762_;
  assign new_n5764_ = ~B9211 & ~new_n2768_;
  assign new_n5765_ = B9211 & new_n2768_;
  assign new_n5766_ = ~new_n5764_ & ~new_n5765_;
  assign new_n5767_ = new_n5763_ & ~new_n5766_;
  assign new_n5768_ = ~new_n4566_ & ~new_n5767_;
  assign new_n5769_ = B9245 & B9244;
  assign new_n5770_ = ~new_n2780_ & ~new_n5769_;
  assign new_n5771_ = ~B9244 & ~new_n2778_;
  assign new_n5772_ = B9244 & new_n2778_;
  assign new_n5773_ = ~new_n5771_ & ~new_n5772_;
  assign new_n5774_ = new_n5770_ & ~new_n5773_;
  assign new_n5775_ = ~new_n4573_ & ~new_n5774_;
  assign new_n5776_ = new_n5761_ & new_n5775_;
  assign new_n5777_ = B9278 & B9277;
  assign new_n5778_ = ~new_n2791_ & ~new_n5777_;
  assign new_n5779_ = ~B9277 & ~new_n2789_;
  assign new_n5780_ = B9277 & new_n2789_;
  assign new_n5781_ = ~new_n5779_ & ~new_n5780_;
  assign new_n5782_ = new_n5778_ & ~new_n5781_;
  assign new_n5783_ = ~new_n4581_ & ~new_n5782_;
  assign new_n5784_ = new_n5775_ & new_n5783_;
  assign new_n5785_ = ~new_n5776_ & ~new_n5784_;
  assign new_n5786_ = ~new_n5768_ & new_n5785_;
  assign new_n5787_ = new_n5768_ & ~new_n5785_;
  assign new_n5788_ = ~new_n5786_ & ~new_n5787_;
  assign new_n5789_ = ~new_n5761_ & ~new_n5788_;
  assign new_n5790_ = ~new_n5743_ & ~new_n5789_;
  assign new_n5791_ = ~new_n5744_ & ~new_n5790_;
  assign new_n5792_ = new_n5698_ & new_n5791_;
  assign new_n5793_ = ~new_n5698_ & ~new_n5791_;
  assign new_n5794_ = ~new_n5792_ & ~new_n5793_;
  assign new_n5795_ = ~new_n5653_ & ~new_n5794_;
  assign new_n5796_ = ~new_n5559_ & ~new_n5795_;
  assign new_n5797_ = ~new_n5560_ & ~new_n5796_;
  assign new_n5798_ = new_n5324_ & new_n5797_;
  assign new_n5799_ = ~new_n5324_ & ~new_n5797_;
  assign new_n5800_ = ~new_n5798_ & ~new_n5799_;
  assign A6808 = ~new_n5089_ & ~new_n5800_;
  assign new_n5802_ = ~new_n5086_ & ~new_n5798_;
  assign A6807 = ~new_n5089_ & ~new_n5802_;
  assign new_n5804_ = new_n5086_ & new_n5324_;
  assign new_n5805_ = ~new_n5089_ & ~new_n5804_;
  assign new_n5806_ = new_n5089_ & ~new_n5805_;
  assign new_n5807_ = new_n5089_ & new_n5804_;
  assign new_n5808_ = new_n5806_ & ~new_n5807_;
  assign new_n5809_ = new_n5324_ & ~new_n5808_;
  assign A6806 = new_n5797_ | new_n5809_;
  assign new_n5811_ = new_n5559_ & new_n5795_;
  assign new_n5812_ = ~new_n5796_ & ~new_n5811_;
  assign new_n5813_ = ~new_n5089_ & ~new_n5559_;
  assign new_n5814_ = new_n5089_ & new_n5559_;
  assign new_n5815_ = ~new_n5813_ & ~new_n5814_;
  assign new_n5816_ = new_n5812_ & ~new_n5815_;
  assign A6805 = new_n5809_ | new_n5816_;
  assign new_n5818_ = new_n5324_ & ~new_n5816_;
  assign new_n5819_ = ~new_n5324_ & new_n5816_;
  assign new_n5820_ = ~new_n5818_ & ~new_n5819_;
  assign A6804 = ~new_n5089_ & ~new_n5820_;
  assign new_n5822_ = B5217 & ~new_n4629_;
  assign new_n5823_ = ~B5217 & new_n4629_;
  assign new_n5824_ = ~new_n5822_ & ~new_n5823_;
  assign new_n5825_ = ~new_n1267_ & ~new_n5824_;
  assign new_n5826_ = ~B5184 & ~new_n3421_;
  assign new_n5827_ = ~new_n4621_ & ~new_n5826_;
  assign new_n5828_ = ~new_n1256_ & ~new_n5827_;
  assign new_n5829_ = new_n5825_ & new_n5828_;
  assign new_n5830_ = ~new_n5825_ & ~new_n5828_;
  assign new_n5831_ = ~new_n5829_ & ~new_n5830_;
  assign new_n5832_ = B5316 & ~new_n4654_;
  assign new_n5833_ = ~B5316 & new_n4654_;
  assign new_n5834_ = ~new_n5832_ & ~new_n5833_;
  assign new_n5835_ = ~new_n1301_ & ~new_n5834_;
  assign new_n5836_ = B5283 & ~new_n4646_;
  assign new_n5837_ = ~B5283 & new_n4646_;
  assign new_n5838_ = ~new_n5836_ & ~new_n5837_;
  assign new_n5839_ = ~new_n1290_ & ~new_n5838_;
  assign new_n5840_ = ~new_n5835_ & new_n5839_;
  assign new_n5841_ = new_n5835_ & ~new_n5839_;
  assign new_n5842_ = ~new_n5840_ & ~new_n5841_;
  assign new_n5843_ = ~new_n5825_ & ~new_n5842_;
  assign new_n5844_ = new_n5825_ & new_n5842_;
  assign new_n5845_ = ~new_n5843_ & ~new_n5844_;
  assign new_n5846_ = new_n5831_ & ~new_n5845_;
  assign new_n5847_ = B5250 & ~new_n4639_;
  assign new_n5848_ = ~B5250 & new_n4639_;
  assign new_n5849_ = ~new_n5847_ & ~new_n5848_;
  assign new_n5850_ = ~new_n1280_ & ~new_n5849_;
  assign new_n5851_ = ~new_n5846_ & new_n5850_;
  assign new_n5852_ = new_n5846_ & ~new_n5850_;
  assign new_n5853_ = ~new_n5851_ & ~new_n5852_;
  assign new_n5854_ = ~new_n5842_ & ~new_n5853_;
  assign new_n5855_ = B5349 & ~new_n4667_;
  assign new_n5856_ = ~B5349 & new_n4667_;
  assign new_n5857_ = ~new_n5855_ & ~new_n5856_;
  assign new_n5858_ = ~new_n1317_ & ~new_n5857_;
  assign new_n5859_ = B5382 & ~new_n4674_;
  assign new_n5860_ = ~B5382 & new_n4674_;
  assign new_n5861_ = ~new_n5859_ & ~new_n5860_;
  assign new_n5862_ = ~new_n1327_ & ~new_n5861_;
  assign new_n5863_ = ~new_n5858_ & new_n5862_;
  assign new_n5864_ = new_n5858_ & ~new_n5862_;
  assign new_n5865_ = ~new_n5863_ & ~new_n5864_;
  assign new_n5866_ = B5415 & ~new_n4684_;
  assign new_n5867_ = ~B5415 & new_n4684_;
  assign new_n5868_ = ~new_n5866_ & ~new_n5867_;
  assign new_n5869_ = ~new_n1340_ & ~new_n5868_;
  assign new_n5870_ = B5448 & ~new_n4691_;
  assign new_n5871_ = ~B5448 & new_n4691_;
  assign new_n5872_ = ~new_n5870_ & ~new_n5871_;
  assign new_n5873_ = ~new_n1350_ & ~new_n5872_;
  assign new_n5874_ = new_n5865_ & ~new_n5873_;
  assign new_n5875_ = B5481 & ~new_n4699_;
  assign new_n5876_ = ~B5481 & new_n4699_;
  assign new_n5877_ = ~new_n5875_ & ~new_n5876_;
  assign new_n5878_ = ~new_n1361_ & ~new_n5877_;
  assign new_n5879_ = ~new_n5873_ & ~new_n5878_;
  assign new_n5880_ = ~new_n5874_ & ~new_n5879_;
  assign new_n5881_ = new_n5869_ & new_n5880_;
  assign new_n5882_ = ~new_n5869_ & ~new_n5880_;
  assign new_n5883_ = ~new_n5881_ & ~new_n5882_;
  assign new_n5884_ = ~new_n5865_ & ~new_n5883_;
  assign new_n5885_ = ~new_n5854_ & new_n5884_;
  assign new_n5886_ = new_n5854_ & ~new_n5884_;
  assign new_n5887_ = ~new_n5885_ & ~new_n5886_;
  assign new_n5888_ = B5514 & ~new_n4715_;
  assign new_n5889_ = ~B5514 & new_n4715_;
  assign new_n5890_ = ~new_n5888_ & ~new_n5889_;
  assign new_n5891_ = ~new_n1380_ & ~new_n5890_;
  assign new_n5892_ = B5547 & ~new_n4722_;
  assign new_n5893_ = ~B5547 & new_n4722_;
  assign new_n5894_ = ~new_n5892_ & ~new_n5893_;
  assign new_n5895_ = ~new_n1390_ & ~new_n5894_;
  assign new_n5896_ = ~new_n5891_ & new_n5895_;
  assign new_n5897_ = new_n5891_ & ~new_n5895_;
  assign new_n5898_ = ~new_n5896_ & ~new_n5897_;
  assign new_n5899_ = B5580 & ~new_n4732_;
  assign new_n5900_ = ~B5580 & new_n4732_;
  assign new_n5901_ = ~new_n5899_ & ~new_n5900_;
  assign new_n5902_ = ~new_n1403_ & ~new_n5901_;
  assign new_n5903_ = B5613 & ~new_n4739_;
  assign new_n5904_ = ~B5613 & new_n4739_;
  assign new_n5905_ = ~new_n5903_ & ~new_n5904_;
  assign new_n5906_ = ~new_n1413_ & ~new_n5905_;
  assign new_n5907_ = new_n5898_ & ~new_n5906_;
  assign new_n5908_ = B5646 & ~new_n4747_;
  assign new_n5909_ = ~B5646 & new_n4747_;
  assign new_n5910_ = ~new_n5908_ & ~new_n5909_;
  assign new_n5911_ = ~new_n1424_ & ~new_n5910_;
  assign new_n5912_ = ~new_n5906_ & ~new_n5911_;
  assign new_n5913_ = ~new_n5907_ & ~new_n5912_;
  assign new_n5914_ = new_n5902_ & new_n5913_;
  assign new_n5915_ = ~new_n5902_ & ~new_n5913_;
  assign new_n5916_ = ~new_n5914_ & ~new_n5915_;
  assign new_n5917_ = ~new_n5898_ & ~new_n5916_;
  assign new_n5918_ = B5679 & ~new_n4760_;
  assign new_n5919_ = ~B5679 & new_n4760_;
  assign new_n5920_ = ~new_n5918_ & ~new_n5919_;
  assign new_n5921_ = ~new_n1440_ & ~new_n5920_;
  assign new_n5922_ = B5712 & ~new_n4767_;
  assign new_n5923_ = ~B5712 & new_n4767_;
  assign new_n5924_ = ~new_n5922_ & ~new_n5923_;
  assign new_n5925_ = ~new_n1450_ & ~new_n5924_;
  assign new_n5926_ = ~new_n5921_ & new_n5925_;
  assign new_n5927_ = new_n5921_ & ~new_n5925_;
  assign new_n5928_ = ~new_n5926_ & ~new_n5927_;
  assign new_n5929_ = B5745 & ~new_n4777_;
  assign new_n5930_ = ~B5745 & new_n4777_;
  assign new_n5931_ = ~new_n5929_ & ~new_n5930_;
  assign new_n5932_ = ~new_n1463_ & ~new_n5931_;
  assign new_n5933_ = B5778 & ~new_n4784_;
  assign new_n5934_ = ~B5778 & new_n4784_;
  assign new_n5935_ = ~new_n5933_ & ~new_n5934_;
  assign new_n5936_ = ~new_n1473_ & ~new_n5935_;
  assign new_n5937_ = new_n5928_ & ~new_n5936_;
  assign new_n5938_ = B5811 & ~new_n4792_;
  assign new_n5939_ = ~B5811 & new_n4792_;
  assign new_n5940_ = ~new_n5938_ & ~new_n5939_;
  assign new_n5941_ = ~new_n1484_ & ~new_n5940_;
  assign new_n5942_ = ~new_n5936_ & ~new_n5941_;
  assign new_n5943_ = ~new_n5937_ & ~new_n5942_;
  assign new_n5944_ = new_n5932_ & new_n5943_;
  assign new_n5945_ = ~new_n5932_ & ~new_n5943_;
  assign new_n5946_ = ~new_n5944_ & ~new_n5945_;
  assign new_n5947_ = ~new_n5928_ & ~new_n5946_;
  assign new_n5948_ = new_n5887_ & ~new_n5947_;
  assign new_n5949_ = B5844 & ~new_n4806_;
  assign new_n5950_ = ~B5844 & new_n4806_;
  assign new_n5951_ = ~new_n5949_ & ~new_n5950_;
  assign new_n5952_ = ~new_n1501_ & ~new_n5951_;
  assign new_n5953_ = B5877 & ~new_n4813_;
  assign new_n5954_ = ~B5877 & new_n4813_;
  assign new_n5955_ = ~new_n5953_ & ~new_n5954_;
  assign new_n5956_ = ~new_n1511_ & ~new_n5955_;
  assign new_n5957_ = ~new_n5952_ & new_n5956_;
  assign new_n5958_ = new_n5952_ & ~new_n5956_;
  assign new_n5959_ = ~new_n5957_ & ~new_n5958_;
  assign new_n5960_ = B5910 & ~new_n4823_;
  assign new_n5961_ = ~B5910 & new_n4823_;
  assign new_n5962_ = ~new_n5960_ & ~new_n5961_;
  assign new_n5963_ = ~new_n1524_ & ~new_n5962_;
  assign new_n5964_ = B5943 & ~new_n4830_;
  assign new_n5965_ = ~B5943 & new_n4830_;
  assign new_n5966_ = ~new_n5964_ & ~new_n5965_;
  assign new_n5967_ = ~new_n1534_ & ~new_n5966_;
  assign new_n5968_ = new_n5959_ & ~new_n5967_;
  assign new_n5969_ = B5976 & ~new_n4838_;
  assign new_n5970_ = ~B5976 & new_n4838_;
  assign new_n5971_ = ~new_n5969_ & ~new_n5970_;
  assign new_n5972_ = ~new_n1545_ & ~new_n5971_;
  assign new_n5973_ = ~new_n5967_ & ~new_n5972_;
  assign new_n5974_ = ~new_n5968_ & ~new_n5973_;
  assign new_n5975_ = new_n5963_ & new_n5974_;
  assign new_n5976_ = ~new_n5963_ & ~new_n5974_;
  assign new_n5977_ = ~new_n5975_ & ~new_n5976_;
  assign new_n5978_ = ~new_n5959_ & ~new_n5977_;
  assign new_n5979_ = ~new_n5947_ & ~new_n5978_;
  assign new_n5980_ = ~new_n5948_ & ~new_n5979_;
  assign new_n5981_ = new_n5917_ & new_n5980_;
  assign new_n5982_ = ~new_n5917_ & ~new_n5980_;
  assign new_n5983_ = ~new_n5981_ & ~new_n5982_;
  assign new_n5984_ = ~new_n5887_ & ~new_n5983_;
  assign new_n5985_ = B6009 & ~new_n4857_;
  assign new_n5986_ = ~B6009 & new_n4857_;
  assign new_n5987_ = ~new_n5985_ & ~new_n5986_;
  assign new_n5988_ = ~new_n1567_ & ~new_n5987_;
  assign new_n5989_ = B6042 & ~new_n4864_;
  assign new_n5990_ = ~B6042 & new_n4864_;
  assign new_n5991_ = ~new_n5989_ & ~new_n5990_;
  assign new_n5992_ = ~new_n1577_ & ~new_n5991_;
  assign new_n5993_ = ~new_n5988_ & new_n5992_;
  assign new_n5994_ = new_n5988_ & ~new_n5992_;
  assign new_n5995_ = ~new_n5993_ & ~new_n5994_;
  assign new_n5996_ = B6075 & ~new_n4874_;
  assign new_n5997_ = ~B6075 & new_n4874_;
  assign new_n5998_ = ~new_n5996_ & ~new_n5997_;
  assign new_n5999_ = ~new_n1590_ & ~new_n5998_;
  assign new_n6000_ = B6108 & ~new_n4881_;
  assign new_n6001_ = ~B6108 & new_n4881_;
  assign new_n6002_ = ~new_n6000_ & ~new_n6001_;
  assign new_n6003_ = ~new_n1600_ & ~new_n6002_;
  assign new_n6004_ = new_n5995_ & ~new_n6003_;
  assign new_n6005_ = B6141 & ~new_n4889_;
  assign new_n6006_ = ~B6141 & new_n4889_;
  assign new_n6007_ = ~new_n6005_ & ~new_n6006_;
  assign new_n6008_ = ~new_n1611_ & ~new_n6007_;
  assign new_n6009_ = ~new_n6003_ & ~new_n6008_;
  assign new_n6010_ = ~new_n6004_ & ~new_n6009_;
  assign new_n6011_ = new_n5999_ & new_n6010_;
  assign new_n6012_ = ~new_n5999_ & ~new_n6010_;
  assign new_n6013_ = ~new_n6011_ & ~new_n6012_;
  assign new_n6014_ = ~new_n5995_ & ~new_n6013_;
  assign new_n6015_ = B6174 & ~new_n4902_;
  assign new_n6016_ = ~B6174 & new_n4902_;
  assign new_n6017_ = ~new_n6015_ & ~new_n6016_;
  assign new_n6018_ = ~new_n1627_ & ~new_n6017_;
  assign new_n6019_ = B6207 & ~new_n4909_;
  assign new_n6020_ = ~B6207 & new_n4909_;
  assign new_n6021_ = ~new_n6019_ & ~new_n6020_;
  assign new_n6022_ = ~new_n1637_ & ~new_n6021_;
  assign new_n6023_ = ~new_n6018_ & new_n6022_;
  assign new_n6024_ = new_n6018_ & ~new_n6022_;
  assign new_n6025_ = ~new_n6023_ & ~new_n6024_;
  assign new_n6026_ = B6240 & ~new_n4919_;
  assign new_n6027_ = ~B6240 & new_n4919_;
  assign new_n6028_ = ~new_n6026_ & ~new_n6027_;
  assign new_n6029_ = ~new_n1650_ & ~new_n6028_;
  assign new_n6030_ = B6273 & ~new_n4926_;
  assign new_n6031_ = ~B6273 & new_n4926_;
  assign new_n6032_ = ~new_n6030_ & ~new_n6031_;
  assign new_n6033_ = ~new_n1660_ & ~new_n6032_;
  assign new_n6034_ = new_n6025_ & ~new_n6033_;
  assign new_n6035_ = B6306 & ~new_n4934_;
  assign new_n6036_ = ~B6306 & new_n4934_;
  assign new_n6037_ = ~new_n6035_ & ~new_n6036_;
  assign new_n6038_ = ~new_n1671_ & ~new_n6037_;
  assign new_n6039_ = ~new_n6033_ & ~new_n6038_;
  assign new_n6040_ = ~new_n6034_ & ~new_n6039_;
  assign new_n6041_ = new_n6029_ & new_n6040_;
  assign new_n6042_ = ~new_n6029_ & ~new_n6040_;
  assign new_n6043_ = ~new_n6041_ & ~new_n6042_;
  assign new_n6044_ = ~new_n6025_ & ~new_n6043_;
  assign new_n6045_ = ~new_n6014_ & new_n6044_;
  assign new_n6046_ = new_n6014_ & ~new_n6044_;
  assign new_n6047_ = ~new_n6045_ & ~new_n6046_;
  assign new_n6048_ = B6339 & ~new_n4950_;
  assign new_n6049_ = ~B6339 & new_n4950_;
  assign new_n6050_ = ~new_n6048_ & ~new_n6049_;
  assign new_n6051_ = ~new_n1690_ & ~new_n6050_;
  assign new_n6052_ = B6372 & ~new_n4957_;
  assign new_n6053_ = ~B6372 & new_n4957_;
  assign new_n6054_ = ~new_n6052_ & ~new_n6053_;
  assign new_n6055_ = ~new_n1700_ & ~new_n6054_;
  assign new_n6056_ = ~new_n6051_ & new_n6055_;
  assign new_n6057_ = new_n6051_ & ~new_n6055_;
  assign new_n6058_ = ~new_n6056_ & ~new_n6057_;
  assign new_n6059_ = B6405 & ~new_n4967_;
  assign new_n6060_ = ~B6405 & new_n4967_;
  assign new_n6061_ = ~new_n6059_ & ~new_n6060_;
  assign new_n6062_ = ~new_n1713_ & ~new_n6061_;
  assign new_n6063_ = B6438 & ~new_n4974_;
  assign new_n6064_ = ~B6438 & new_n4974_;
  assign new_n6065_ = ~new_n6063_ & ~new_n6064_;
  assign new_n6066_ = ~new_n1723_ & ~new_n6065_;
  assign new_n6067_ = new_n6058_ & ~new_n6066_;
  assign new_n6068_ = B6471 & ~new_n4982_;
  assign new_n6069_ = ~B6471 & new_n4982_;
  assign new_n6070_ = ~new_n6068_ & ~new_n6069_;
  assign new_n6071_ = ~new_n1734_ & ~new_n6070_;
  assign new_n6072_ = ~new_n6066_ & ~new_n6071_;
  assign new_n6073_ = ~new_n6067_ & ~new_n6072_;
  assign new_n6074_ = new_n6062_ & new_n6073_;
  assign new_n6075_ = ~new_n6062_ & ~new_n6073_;
  assign new_n6076_ = ~new_n6074_ & ~new_n6075_;
  assign new_n6077_ = ~new_n6058_ & ~new_n6076_;
  assign new_n6078_ = B6504 & ~new_n4995_;
  assign new_n6079_ = ~B6504 & new_n4995_;
  assign new_n6080_ = ~new_n6078_ & ~new_n6079_;
  assign new_n6081_ = ~new_n1750_ & ~new_n6080_;
  assign new_n6082_ = B6537 & ~new_n5002_;
  assign new_n6083_ = ~B6537 & new_n5002_;
  assign new_n6084_ = ~new_n6082_ & ~new_n6083_;
  assign new_n6085_ = ~new_n1760_ & ~new_n6084_;
  assign new_n6086_ = ~new_n6081_ & new_n6085_;
  assign new_n6087_ = new_n6081_ & ~new_n6085_;
  assign new_n6088_ = ~new_n6086_ & ~new_n6087_;
  assign new_n6089_ = B6570 & ~new_n5012_;
  assign new_n6090_ = ~B6570 & new_n5012_;
  assign new_n6091_ = ~new_n6089_ & ~new_n6090_;
  assign new_n6092_ = ~new_n1773_ & ~new_n6091_;
  assign new_n6093_ = B6603 & ~new_n5019_;
  assign new_n6094_ = ~B6603 & new_n5019_;
  assign new_n6095_ = ~new_n6093_ & ~new_n6094_;
  assign new_n6096_ = ~new_n1783_ & ~new_n6095_;
  assign new_n6097_ = new_n6088_ & ~new_n6096_;
  assign new_n6098_ = B6636 & ~new_n5027_;
  assign new_n6099_ = ~B6636 & new_n5027_;
  assign new_n6100_ = ~new_n6098_ & ~new_n6099_;
  assign new_n6101_ = ~new_n1794_ & ~new_n6100_;
  assign new_n6102_ = ~new_n6096_ & ~new_n6101_;
  assign new_n6103_ = ~new_n6097_ & ~new_n6102_;
  assign new_n6104_ = new_n6092_ & new_n6103_;
  assign new_n6105_ = ~new_n6092_ & ~new_n6103_;
  assign new_n6106_ = ~new_n6104_ & ~new_n6105_;
  assign new_n6107_ = ~new_n6088_ & ~new_n6106_;
  assign new_n6108_ = new_n6047_ & ~new_n6107_;
  assign new_n6109_ = B6669 & ~new_n5041_;
  assign new_n6110_ = ~B6669 & new_n5041_;
  assign new_n6111_ = ~new_n6109_ & ~new_n6110_;
  assign new_n6112_ = ~new_n1811_ & ~new_n6111_;
  assign new_n6113_ = B6702 & ~new_n5048_;
  assign new_n6114_ = ~B6702 & new_n5048_;
  assign new_n6115_ = ~new_n6113_ & ~new_n6114_;
  assign new_n6116_ = ~new_n1821_ & ~new_n6115_;
  assign new_n6117_ = ~new_n6112_ & new_n6116_;
  assign new_n6118_ = new_n6112_ & ~new_n6116_;
  assign new_n6119_ = ~new_n6117_ & ~new_n6118_;
  assign new_n6120_ = B6735 & ~new_n5058_;
  assign new_n6121_ = ~B6735 & new_n5058_;
  assign new_n6122_ = ~new_n6120_ & ~new_n6121_;
  assign new_n6123_ = ~new_n1834_ & ~new_n6122_;
  assign new_n6124_ = B6768 & ~new_n5065_;
  assign new_n6125_ = ~B6768 & new_n5065_;
  assign new_n6126_ = ~new_n6124_ & ~new_n6125_;
  assign new_n6127_ = ~new_n1844_ & ~new_n6126_;
  assign new_n6128_ = new_n6119_ & ~new_n6127_;
  assign new_n6129_ = B6801 & ~new_n5073_;
  assign new_n6130_ = ~B6801 & new_n5073_;
  assign new_n6131_ = ~new_n6129_ & ~new_n6130_;
  assign new_n6132_ = ~new_n1855_ & ~new_n6131_;
  assign new_n6133_ = ~new_n6127_ & ~new_n6132_;
  assign new_n6134_ = ~new_n6128_ & ~new_n6133_;
  assign new_n6135_ = new_n6123_ & new_n6134_;
  assign new_n6136_ = ~new_n6123_ & ~new_n6134_;
  assign new_n6137_ = ~new_n6135_ & ~new_n6136_;
  assign new_n6138_ = ~new_n6119_ & ~new_n6137_;
  assign new_n6139_ = ~new_n6107_ & ~new_n6138_;
  assign new_n6140_ = ~new_n6108_ & ~new_n6139_;
  assign new_n6141_ = new_n6077_ & new_n6140_;
  assign new_n6142_ = ~new_n6077_ & ~new_n6140_;
  assign new_n6143_ = ~new_n6141_ & ~new_n6142_;
  assign new_n6144_ = ~new_n6047_ & ~new_n6143_;
  assign new_n6145_ = ~new_n5984_ & new_n6144_;
  assign new_n6146_ = new_n5984_ & ~new_n6144_;
  assign new_n6147_ = ~new_n6145_ & ~new_n6146_;
  assign new_n6148_ = B6834 & ~new_n5095_;
  assign new_n6149_ = ~B6834 & new_n5095_;
  assign new_n6150_ = ~new_n6148_ & ~new_n6149_;
  assign new_n6151_ = ~new_n1880_ & ~new_n6150_;
  assign new_n6152_ = B6867 & ~new_n5102_;
  assign new_n6153_ = ~B6867 & new_n5102_;
  assign new_n6154_ = ~new_n6152_ & ~new_n6153_;
  assign new_n6155_ = ~new_n1890_ & ~new_n6154_;
  assign new_n6156_ = ~new_n6151_ & new_n6155_;
  assign new_n6157_ = new_n6151_ & ~new_n6155_;
  assign new_n6158_ = ~new_n6156_ & ~new_n6157_;
  assign new_n6159_ = B6900 & ~new_n5112_;
  assign new_n6160_ = ~B6900 & new_n5112_;
  assign new_n6161_ = ~new_n6159_ & ~new_n6160_;
  assign new_n6162_ = ~new_n1903_ & ~new_n6161_;
  assign new_n6163_ = B6933 & ~new_n5119_;
  assign new_n6164_ = ~B6933 & new_n5119_;
  assign new_n6165_ = ~new_n6163_ & ~new_n6164_;
  assign new_n6166_ = ~new_n1913_ & ~new_n6165_;
  assign new_n6167_ = new_n6158_ & ~new_n6166_;
  assign new_n6168_ = B6966 & ~new_n5127_;
  assign new_n6169_ = ~B6966 & new_n5127_;
  assign new_n6170_ = ~new_n6168_ & ~new_n6169_;
  assign new_n6171_ = ~new_n1924_ & ~new_n6170_;
  assign new_n6172_ = ~new_n6166_ & ~new_n6171_;
  assign new_n6173_ = ~new_n6167_ & ~new_n6172_;
  assign new_n6174_ = new_n6162_ & new_n6173_;
  assign new_n6175_ = ~new_n6162_ & ~new_n6173_;
  assign new_n6176_ = ~new_n6174_ & ~new_n6175_;
  assign new_n6177_ = ~new_n6158_ & ~new_n6176_;
  assign new_n6178_ = B6999 & ~new_n5140_;
  assign new_n6179_ = ~B6999 & new_n5140_;
  assign new_n6180_ = ~new_n6178_ & ~new_n6179_;
  assign new_n6181_ = ~new_n1940_ & ~new_n6180_;
  assign new_n6182_ = B7032 & ~new_n5147_;
  assign new_n6183_ = ~B7032 & new_n5147_;
  assign new_n6184_ = ~new_n6182_ & ~new_n6183_;
  assign new_n6185_ = ~new_n1950_ & ~new_n6184_;
  assign new_n6186_ = ~new_n6181_ & new_n6185_;
  assign new_n6187_ = new_n6181_ & ~new_n6185_;
  assign new_n6188_ = ~new_n6186_ & ~new_n6187_;
  assign new_n6189_ = B7065 & ~new_n5157_;
  assign new_n6190_ = ~B7065 & new_n5157_;
  assign new_n6191_ = ~new_n6189_ & ~new_n6190_;
  assign new_n6192_ = ~new_n1963_ & ~new_n6191_;
  assign new_n6193_ = B7098 & ~new_n5164_;
  assign new_n6194_ = ~B7098 & new_n5164_;
  assign new_n6195_ = ~new_n6193_ & ~new_n6194_;
  assign new_n6196_ = ~new_n1973_ & ~new_n6195_;
  assign new_n6197_ = new_n6188_ & ~new_n6196_;
  assign new_n6198_ = B7131 & ~new_n5172_;
  assign new_n6199_ = ~B7131 & new_n5172_;
  assign new_n6200_ = ~new_n6198_ & ~new_n6199_;
  assign new_n6201_ = ~new_n1984_ & ~new_n6200_;
  assign new_n6202_ = ~new_n6196_ & ~new_n6201_;
  assign new_n6203_ = ~new_n6197_ & ~new_n6202_;
  assign new_n6204_ = new_n6192_ & new_n6203_;
  assign new_n6205_ = ~new_n6192_ & ~new_n6203_;
  assign new_n6206_ = ~new_n6204_ & ~new_n6205_;
  assign new_n6207_ = ~new_n6188_ & ~new_n6206_;
  assign new_n6208_ = ~new_n6177_ & new_n6207_;
  assign new_n6209_ = new_n6177_ & ~new_n6207_;
  assign new_n6210_ = ~new_n6208_ & ~new_n6209_;
  assign new_n6211_ = B7164 & ~new_n5188_;
  assign new_n6212_ = ~B7164 & new_n5188_;
  assign new_n6213_ = ~new_n6211_ & ~new_n6212_;
  assign new_n6214_ = ~new_n2003_ & ~new_n6213_;
  assign new_n6215_ = B7197 & ~new_n5195_;
  assign new_n6216_ = ~B7197 & new_n5195_;
  assign new_n6217_ = ~new_n6215_ & ~new_n6216_;
  assign new_n6218_ = ~new_n2013_ & ~new_n6217_;
  assign new_n6219_ = ~new_n6214_ & new_n6218_;
  assign new_n6220_ = new_n6214_ & ~new_n6218_;
  assign new_n6221_ = ~new_n6219_ & ~new_n6220_;
  assign new_n6222_ = B7230 & ~new_n5205_;
  assign new_n6223_ = ~B7230 & new_n5205_;
  assign new_n6224_ = ~new_n6222_ & ~new_n6223_;
  assign new_n6225_ = ~new_n2026_ & ~new_n6224_;
  assign new_n6226_ = B7263 & ~new_n5212_;
  assign new_n6227_ = ~B7263 & new_n5212_;
  assign new_n6228_ = ~new_n6226_ & ~new_n6227_;
  assign new_n6229_ = ~new_n2036_ & ~new_n6228_;
  assign new_n6230_ = new_n6221_ & ~new_n6229_;
  assign new_n6231_ = B7296 & ~new_n5220_;
  assign new_n6232_ = ~B7296 & new_n5220_;
  assign new_n6233_ = ~new_n6231_ & ~new_n6232_;
  assign new_n6234_ = ~new_n2047_ & ~new_n6233_;
  assign new_n6235_ = ~new_n6229_ & ~new_n6234_;
  assign new_n6236_ = ~new_n6230_ & ~new_n6235_;
  assign new_n6237_ = new_n6225_ & new_n6236_;
  assign new_n6238_ = ~new_n6225_ & ~new_n6236_;
  assign new_n6239_ = ~new_n6237_ & ~new_n6238_;
  assign new_n6240_ = ~new_n6221_ & ~new_n6239_;
  assign new_n6241_ = B7329 & ~new_n5233_;
  assign new_n6242_ = ~B7329 & new_n5233_;
  assign new_n6243_ = ~new_n6241_ & ~new_n6242_;
  assign new_n6244_ = ~new_n2063_ & ~new_n6243_;
  assign new_n6245_ = B7362 & ~new_n5240_;
  assign new_n6246_ = ~B7362 & new_n5240_;
  assign new_n6247_ = ~new_n6245_ & ~new_n6246_;
  assign new_n6248_ = ~new_n2073_ & ~new_n6247_;
  assign new_n6249_ = ~new_n6244_ & new_n6248_;
  assign new_n6250_ = new_n6244_ & ~new_n6248_;
  assign new_n6251_ = ~new_n6249_ & ~new_n6250_;
  assign new_n6252_ = B7395 & ~new_n5250_;
  assign new_n6253_ = ~B7395 & new_n5250_;
  assign new_n6254_ = ~new_n6252_ & ~new_n6253_;
  assign new_n6255_ = ~new_n2086_ & ~new_n6254_;
  assign new_n6256_ = B7428 & ~new_n5257_;
  assign new_n6257_ = ~B7428 & new_n5257_;
  assign new_n6258_ = ~new_n6256_ & ~new_n6257_;
  assign new_n6259_ = ~new_n2096_ & ~new_n6258_;
  assign new_n6260_ = new_n6251_ & ~new_n6259_;
  assign new_n6261_ = B7461 & ~new_n5265_;
  assign new_n6262_ = ~B7461 & new_n5265_;
  assign new_n6263_ = ~new_n6261_ & ~new_n6262_;
  assign new_n6264_ = ~new_n2107_ & ~new_n6263_;
  assign new_n6265_ = ~new_n6259_ & ~new_n6264_;
  assign new_n6266_ = ~new_n6260_ & ~new_n6265_;
  assign new_n6267_ = new_n6255_ & new_n6266_;
  assign new_n6268_ = ~new_n6255_ & ~new_n6266_;
  assign new_n6269_ = ~new_n6267_ & ~new_n6268_;
  assign new_n6270_ = ~new_n6251_ & ~new_n6269_;
  assign new_n6271_ = new_n6210_ & ~new_n6270_;
  assign new_n6272_ = B7494 & ~new_n5279_;
  assign new_n6273_ = ~B7494 & new_n5279_;
  assign new_n6274_ = ~new_n6272_ & ~new_n6273_;
  assign new_n6275_ = ~new_n2124_ & ~new_n6274_;
  assign new_n6276_ = B7527 & ~new_n5286_;
  assign new_n6277_ = ~B7527 & new_n5286_;
  assign new_n6278_ = ~new_n6276_ & ~new_n6277_;
  assign new_n6279_ = ~new_n2134_ & ~new_n6278_;
  assign new_n6280_ = ~new_n6275_ & new_n6279_;
  assign new_n6281_ = new_n6275_ & ~new_n6279_;
  assign new_n6282_ = ~new_n6280_ & ~new_n6281_;
  assign new_n6283_ = B7560 & ~new_n5296_;
  assign new_n6284_ = ~B7560 & new_n5296_;
  assign new_n6285_ = ~new_n6283_ & ~new_n6284_;
  assign new_n6286_ = ~new_n2147_ & ~new_n6285_;
  assign new_n6287_ = B7593 & ~new_n5303_;
  assign new_n6288_ = ~B7593 & new_n5303_;
  assign new_n6289_ = ~new_n6287_ & ~new_n6288_;
  assign new_n6290_ = ~new_n2157_ & ~new_n6289_;
  assign new_n6291_ = new_n6282_ & ~new_n6290_;
  assign new_n6292_ = B7626 & ~new_n5311_;
  assign new_n6293_ = ~B7626 & new_n5311_;
  assign new_n6294_ = ~new_n6292_ & ~new_n6293_;
  assign new_n6295_ = ~new_n2168_ & ~new_n6294_;
  assign new_n6296_ = ~new_n6290_ & ~new_n6295_;
  assign new_n6297_ = ~new_n6291_ & ~new_n6296_;
  assign new_n6298_ = new_n6286_ & new_n6297_;
  assign new_n6299_ = ~new_n6286_ & ~new_n6297_;
  assign new_n6300_ = ~new_n6298_ & ~new_n6299_;
  assign new_n6301_ = ~new_n6282_ & ~new_n6300_;
  assign new_n6302_ = ~new_n6270_ & ~new_n6301_;
  assign new_n6303_ = ~new_n6271_ & ~new_n6302_;
  assign new_n6304_ = new_n6240_ & new_n6303_;
  assign new_n6305_ = ~new_n6240_ & ~new_n6303_;
  assign new_n6306_ = ~new_n6304_ & ~new_n6305_;
  assign new_n6307_ = ~new_n6210_ & ~new_n6306_;
  assign new_n6308_ = B7659 & ~new_n5330_;
  assign new_n6309_ = ~B7659 & new_n5330_;
  assign new_n6310_ = ~new_n6308_ & ~new_n6309_;
  assign new_n6311_ = ~new_n2190_ & ~new_n6310_;
  assign new_n6312_ = B7692 & ~new_n5337_;
  assign new_n6313_ = ~B7692 & new_n5337_;
  assign new_n6314_ = ~new_n6312_ & ~new_n6313_;
  assign new_n6315_ = ~new_n2200_ & ~new_n6314_;
  assign new_n6316_ = ~new_n6311_ & new_n6315_;
  assign new_n6317_ = new_n6311_ & ~new_n6315_;
  assign new_n6318_ = ~new_n6316_ & ~new_n6317_;
  assign new_n6319_ = B7725 & ~new_n5347_;
  assign new_n6320_ = ~B7725 & new_n5347_;
  assign new_n6321_ = ~new_n6319_ & ~new_n6320_;
  assign new_n6322_ = ~new_n2213_ & ~new_n6321_;
  assign new_n6323_ = B7758 & ~new_n5354_;
  assign new_n6324_ = ~B7758 & new_n5354_;
  assign new_n6325_ = ~new_n6323_ & ~new_n6324_;
  assign new_n6326_ = ~new_n2223_ & ~new_n6325_;
  assign new_n6327_ = new_n6318_ & ~new_n6326_;
  assign new_n6328_ = B7791 & ~new_n5362_;
  assign new_n6329_ = ~B7791 & new_n5362_;
  assign new_n6330_ = ~new_n6328_ & ~new_n6329_;
  assign new_n6331_ = ~new_n2234_ & ~new_n6330_;
  assign new_n6332_ = ~new_n6326_ & ~new_n6331_;
  assign new_n6333_ = ~new_n6327_ & ~new_n6332_;
  assign new_n6334_ = new_n6322_ & new_n6333_;
  assign new_n6335_ = ~new_n6322_ & ~new_n6333_;
  assign new_n6336_ = ~new_n6334_ & ~new_n6335_;
  assign new_n6337_ = ~new_n6318_ & ~new_n6336_;
  assign new_n6338_ = B7824 & ~new_n5375_;
  assign new_n6339_ = ~B7824 & new_n5375_;
  assign new_n6340_ = ~new_n6338_ & ~new_n6339_;
  assign new_n6341_ = ~new_n2250_ & ~new_n6340_;
  assign new_n6342_ = B7857 & ~new_n5382_;
  assign new_n6343_ = ~B7857 & new_n5382_;
  assign new_n6344_ = ~new_n6342_ & ~new_n6343_;
  assign new_n6345_ = ~new_n2260_ & ~new_n6344_;
  assign new_n6346_ = ~new_n6341_ & new_n6345_;
  assign new_n6347_ = new_n6341_ & ~new_n6345_;
  assign new_n6348_ = ~new_n6346_ & ~new_n6347_;
  assign new_n6349_ = B7890 & ~new_n5392_;
  assign new_n6350_ = ~B7890 & new_n5392_;
  assign new_n6351_ = ~new_n6349_ & ~new_n6350_;
  assign new_n6352_ = ~new_n2273_ & ~new_n6351_;
  assign new_n6353_ = B7923 & ~new_n5399_;
  assign new_n6354_ = ~B7923 & new_n5399_;
  assign new_n6355_ = ~new_n6353_ & ~new_n6354_;
  assign new_n6356_ = ~new_n2283_ & ~new_n6355_;
  assign new_n6357_ = new_n6348_ & ~new_n6356_;
  assign new_n6358_ = B7956 & ~new_n5407_;
  assign new_n6359_ = ~B7956 & new_n5407_;
  assign new_n6360_ = ~new_n6358_ & ~new_n6359_;
  assign new_n6361_ = ~new_n2294_ & ~new_n6360_;
  assign new_n6362_ = ~new_n6356_ & ~new_n6361_;
  assign new_n6363_ = ~new_n6357_ & ~new_n6362_;
  assign new_n6364_ = new_n6352_ & new_n6363_;
  assign new_n6365_ = ~new_n6352_ & ~new_n6363_;
  assign new_n6366_ = ~new_n6364_ & ~new_n6365_;
  assign new_n6367_ = ~new_n6348_ & ~new_n6366_;
  assign new_n6368_ = ~new_n6337_ & new_n6367_;
  assign new_n6369_ = new_n6337_ & ~new_n6367_;
  assign new_n6370_ = ~new_n6368_ & ~new_n6369_;
  assign new_n6371_ = B7989 & ~new_n5423_;
  assign new_n6372_ = ~B7989 & new_n5423_;
  assign new_n6373_ = ~new_n6371_ & ~new_n6372_;
  assign new_n6374_ = ~new_n2313_ & ~new_n6373_;
  assign new_n6375_ = B8022 & ~new_n5430_;
  assign new_n6376_ = ~B8022 & new_n5430_;
  assign new_n6377_ = ~new_n6375_ & ~new_n6376_;
  assign new_n6378_ = ~new_n2323_ & ~new_n6377_;
  assign new_n6379_ = ~new_n6374_ & new_n6378_;
  assign new_n6380_ = new_n6374_ & ~new_n6378_;
  assign new_n6381_ = ~new_n6379_ & ~new_n6380_;
  assign new_n6382_ = B8055 & ~new_n5440_;
  assign new_n6383_ = ~B8055 & new_n5440_;
  assign new_n6384_ = ~new_n6382_ & ~new_n6383_;
  assign new_n6385_ = ~new_n2336_ & ~new_n6384_;
  assign new_n6386_ = B8088 & ~new_n5447_;
  assign new_n6387_ = ~B8088 & new_n5447_;
  assign new_n6388_ = ~new_n6386_ & ~new_n6387_;
  assign new_n6389_ = ~new_n2346_ & ~new_n6388_;
  assign new_n6390_ = new_n6381_ & ~new_n6389_;
  assign new_n6391_ = B8121 & ~new_n5455_;
  assign new_n6392_ = ~B8121 & new_n5455_;
  assign new_n6393_ = ~new_n6391_ & ~new_n6392_;
  assign new_n6394_ = ~new_n2357_ & ~new_n6393_;
  assign new_n6395_ = ~new_n6389_ & ~new_n6394_;
  assign new_n6396_ = ~new_n6390_ & ~new_n6395_;
  assign new_n6397_ = new_n6385_ & new_n6396_;
  assign new_n6398_ = ~new_n6385_ & ~new_n6396_;
  assign new_n6399_ = ~new_n6397_ & ~new_n6398_;
  assign new_n6400_ = ~new_n6381_ & ~new_n6399_;
  assign new_n6401_ = B8154 & ~new_n5468_;
  assign new_n6402_ = ~B8154 & new_n5468_;
  assign new_n6403_ = ~new_n6401_ & ~new_n6402_;
  assign new_n6404_ = ~new_n2373_ & ~new_n6403_;
  assign new_n6405_ = B8187 & ~new_n5475_;
  assign new_n6406_ = ~B8187 & new_n5475_;
  assign new_n6407_ = ~new_n6405_ & ~new_n6406_;
  assign new_n6408_ = ~new_n2383_ & ~new_n6407_;
  assign new_n6409_ = ~new_n6404_ & new_n6408_;
  assign new_n6410_ = new_n6404_ & ~new_n6408_;
  assign new_n6411_ = ~new_n6409_ & ~new_n6410_;
  assign new_n6412_ = B8220 & ~new_n5485_;
  assign new_n6413_ = ~B8220 & new_n5485_;
  assign new_n6414_ = ~new_n6412_ & ~new_n6413_;
  assign new_n6415_ = ~new_n2396_ & ~new_n6414_;
  assign new_n6416_ = B8253 & ~new_n5492_;
  assign new_n6417_ = ~B8253 & new_n5492_;
  assign new_n6418_ = ~new_n6416_ & ~new_n6417_;
  assign new_n6419_ = ~new_n2406_ & ~new_n6418_;
  assign new_n6420_ = new_n6411_ & ~new_n6419_;
  assign new_n6421_ = B8286 & ~new_n5500_;
  assign new_n6422_ = ~B8286 & new_n5500_;
  assign new_n6423_ = ~new_n6421_ & ~new_n6422_;
  assign new_n6424_ = ~new_n2417_ & ~new_n6423_;
  assign new_n6425_ = ~new_n6419_ & ~new_n6424_;
  assign new_n6426_ = ~new_n6420_ & ~new_n6425_;
  assign new_n6427_ = new_n6415_ & new_n6426_;
  assign new_n6428_ = ~new_n6415_ & ~new_n6426_;
  assign new_n6429_ = ~new_n6427_ & ~new_n6428_;
  assign new_n6430_ = ~new_n6411_ & ~new_n6429_;
  assign new_n6431_ = new_n6370_ & ~new_n6430_;
  assign new_n6432_ = B8319 & ~new_n5514_;
  assign new_n6433_ = ~B8319 & new_n5514_;
  assign new_n6434_ = ~new_n6432_ & ~new_n6433_;
  assign new_n6435_ = ~new_n2434_ & ~new_n6434_;
  assign new_n6436_ = B8352 & ~new_n5521_;
  assign new_n6437_ = ~B8352 & new_n5521_;
  assign new_n6438_ = ~new_n6436_ & ~new_n6437_;
  assign new_n6439_ = ~new_n2444_ & ~new_n6438_;
  assign new_n6440_ = ~new_n6435_ & new_n6439_;
  assign new_n6441_ = new_n6435_ & ~new_n6439_;
  assign new_n6442_ = ~new_n6440_ & ~new_n6441_;
  assign new_n6443_ = B8385 & ~new_n5531_;
  assign new_n6444_ = ~B8385 & new_n5531_;
  assign new_n6445_ = ~new_n6443_ & ~new_n6444_;
  assign new_n6446_ = ~new_n2457_ & ~new_n6445_;
  assign new_n6447_ = B8418 & ~new_n5538_;
  assign new_n6448_ = ~B8418 & new_n5538_;
  assign new_n6449_ = ~new_n6447_ & ~new_n6448_;
  assign new_n6450_ = ~new_n2467_ & ~new_n6449_;
  assign new_n6451_ = new_n6442_ & ~new_n6450_;
  assign new_n6452_ = B8451 & ~new_n5546_;
  assign new_n6453_ = ~B8451 & new_n5546_;
  assign new_n6454_ = ~new_n6452_ & ~new_n6453_;
  assign new_n6455_ = ~new_n2478_ & ~new_n6454_;
  assign new_n6456_ = ~new_n6450_ & ~new_n6455_;
  assign new_n6457_ = ~new_n6451_ & ~new_n6456_;
  assign new_n6458_ = new_n6446_ & new_n6457_;
  assign new_n6459_ = ~new_n6446_ & ~new_n6457_;
  assign new_n6460_ = ~new_n6458_ & ~new_n6459_;
  assign new_n6461_ = ~new_n6442_ & ~new_n6460_;
  assign new_n6462_ = ~new_n6430_ & ~new_n6461_;
  assign new_n6463_ = ~new_n6431_ & ~new_n6462_;
  assign new_n6464_ = new_n6400_ & new_n6463_;
  assign new_n6465_ = ~new_n6400_ & ~new_n6463_;
  assign new_n6466_ = ~new_n6464_ & ~new_n6465_;
  assign new_n6467_ = ~new_n6370_ & ~new_n6466_;
  assign new_n6468_ = new_n6147_ & ~new_n6467_;
  assign new_n6469_ = B8484 & ~new_n5566_;
  assign new_n6470_ = ~B8484 & new_n5566_;
  assign new_n6471_ = ~new_n6469_ & ~new_n6470_;
  assign new_n6472_ = ~new_n2501_ & ~new_n6471_;
  assign new_n6473_ = B8517 & ~new_n5573_;
  assign new_n6474_ = ~B8517 & new_n5573_;
  assign new_n6475_ = ~new_n6473_ & ~new_n6474_;
  assign new_n6476_ = ~new_n2511_ & ~new_n6475_;
  assign new_n6477_ = ~new_n6472_ & new_n6476_;
  assign new_n6478_ = new_n6472_ & ~new_n6476_;
  assign new_n6479_ = ~new_n6477_ & ~new_n6478_;
  assign new_n6480_ = B8550 & ~new_n5583_;
  assign new_n6481_ = ~B8550 & new_n5583_;
  assign new_n6482_ = ~new_n6480_ & ~new_n6481_;
  assign new_n6483_ = ~new_n2524_ & ~new_n6482_;
  assign new_n6484_ = B8583 & ~new_n5590_;
  assign new_n6485_ = ~B8583 & new_n5590_;
  assign new_n6486_ = ~new_n6484_ & ~new_n6485_;
  assign new_n6487_ = ~new_n2534_ & ~new_n6486_;
  assign new_n6488_ = new_n6479_ & ~new_n6487_;
  assign new_n6489_ = B8616 & ~new_n5598_;
  assign new_n6490_ = ~B8616 & new_n5598_;
  assign new_n6491_ = ~new_n6489_ & ~new_n6490_;
  assign new_n6492_ = ~new_n2545_ & ~new_n6491_;
  assign new_n6493_ = ~new_n6487_ & ~new_n6492_;
  assign new_n6494_ = ~new_n6488_ & ~new_n6493_;
  assign new_n6495_ = new_n6483_ & new_n6494_;
  assign new_n6496_ = ~new_n6483_ & ~new_n6494_;
  assign new_n6497_ = ~new_n6495_ & ~new_n6496_;
  assign new_n6498_ = ~new_n6479_ & ~new_n6497_;
  assign new_n6499_ = B8649 & ~new_n5611_;
  assign new_n6500_ = ~B8649 & new_n5611_;
  assign new_n6501_ = ~new_n6499_ & ~new_n6500_;
  assign new_n6502_ = ~new_n2561_ & ~new_n6501_;
  assign new_n6503_ = B8682 & ~new_n5618_;
  assign new_n6504_ = ~B8682 & new_n5618_;
  assign new_n6505_ = ~new_n6503_ & ~new_n6504_;
  assign new_n6506_ = ~new_n2571_ & ~new_n6505_;
  assign new_n6507_ = ~new_n6502_ & new_n6506_;
  assign new_n6508_ = new_n6502_ & ~new_n6506_;
  assign new_n6509_ = ~new_n6507_ & ~new_n6508_;
  assign new_n6510_ = B8715 & ~new_n5628_;
  assign new_n6511_ = ~B8715 & new_n5628_;
  assign new_n6512_ = ~new_n6510_ & ~new_n6511_;
  assign new_n6513_ = ~new_n2584_ & ~new_n6512_;
  assign new_n6514_ = B8748 & ~new_n5635_;
  assign new_n6515_ = ~B8748 & new_n5635_;
  assign new_n6516_ = ~new_n6514_ & ~new_n6515_;
  assign new_n6517_ = ~new_n2594_ & ~new_n6516_;
  assign new_n6518_ = new_n6509_ & ~new_n6517_;
  assign new_n6519_ = B8781 & ~new_n5643_;
  assign new_n6520_ = ~B8781 & new_n5643_;
  assign new_n6521_ = ~new_n6519_ & ~new_n6520_;
  assign new_n6522_ = ~new_n2605_ & ~new_n6521_;
  assign new_n6523_ = ~new_n6517_ & ~new_n6522_;
  assign new_n6524_ = ~new_n6518_ & ~new_n6523_;
  assign new_n6525_ = new_n6513_ & new_n6524_;
  assign new_n6526_ = ~new_n6513_ & ~new_n6524_;
  assign new_n6527_ = ~new_n6525_ & ~new_n6526_;
  assign new_n6528_ = ~new_n6509_ & ~new_n6527_;
  assign new_n6529_ = ~new_n6498_ & new_n6528_;
  assign new_n6530_ = new_n6498_ & ~new_n6528_;
  assign new_n6531_ = ~new_n6529_ & ~new_n6530_;
  assign new_n6532_ = B8814 & ~new_n5659_;
  assign new_n6533_ = ~B8814 & new_n5659_;
  assign new_n6534_ = ~new_n6532_ & ~new_n6533_;
  assign new_n6535_ = ~new_n2624_ & ~new_n6534_;
  assign new_n6536_ = B8847 & ~new_n5666_;
  assign new_n6537_ = ~B8847 & new_n5666_;
  assign new_n6538_ = ~new_n6536_ & ~new_n6537_;
  assign new_n6539_ = ~new_n2634_ & ~new_n6538_;
  assign new_n6540_ = ~new_n6535_ & new_n6539_;
  assign new_n6541_ = new_n6535_ & ~new_n6539_;
  assign new_n6542_ = ~new_n6540_ & ~new_n6541_;
  assign new_n6543_ = B8880 & ~new_n5676_;
  assign new_n6544_ = ~B8880 & new_n5676_;
  assign new_n6545_ = ~new_n6543_ & ~new_n6544_;
  assign new_n6546_ = ~new_n2647_ & ~new_n6545_;
  assign new_n6547_ = B8913 & ~new_n5683_;
  assign new_n6548_ = ~B8913 & new_n5683_;
  assign new_n6549_ = ~new_n6547_ & ~new_n6548_;
  assign new_n6550_ = ~new_n2657_ & ~new_n6549_;
  assign new_n6551_ = new_n6542_ & ~new_n6550_;
  assign new_n6552_ = B8946 & ~new_n5691_;
  assign new_n6553_ = ~B8946 & new_n5691_;
  assign new_n6554_ = ~new_n6552_ & ~new_n6553_;
  assign new_n6555_ = ~new_n2668_ & ~new_n6554_;
  assign new_n6556_ = ~new_n6550_ & ~new_n6555_;
  assign new_n6557_ = ~new_n6551_ & ~new_n6556_;
  assign new_n6558_ = new_n6546_ & new_n6557_;
  assign new_n6559_ = ~new_n6546_ & ~new_n6557_;
  assign new_n6560_ = ~new_n6558_ & ~new_n6559_;
  assign new_n6561_ = ~new_n6542_ & ~new_n6560_;
  assign new_n6562_ = B8979 & ~new_n5704_;
  assign new_n6563_ = ~B8979 & new_n5704_;
  assign new_n6564_ = ~new_n6562_ & ~new_n6563_;
  assign new_n6565_ = ~new_n2684_ & ~new_n6564_;
  assign new_n6566_ = B9012 & ~new_n5711_;
  assign new_n6567_ = ~B9012 & new_n5711_;
  assign new_n6568_ = ~new_n6566_ & ~new_n6567_;
  assign new_n6569_ = ~new_n2694_ & ~new_n6568_;
  assign new_n6570_ = ~new_n6565_ & new_n6569_;
  assign new_n6571_ = new_n6565_ & ~new_n6569_;
  assign new_n6572_ = ~new_n6570_ & ~new_n6571_;
  assign new_n6573_ = B9045 & ~new_n5721_;
  assign new_n6574_ = ~B9045 & new_n5721_;
  assign new_n6575_ = ~new_n6573_ & ~new_n6574_;
  assign new_n6576_ = ~new_n2707_ & ~new_n6575_;
  assign new_n6577_ = B9078 & ~new_n5728_;
  assign new_n6578_ = ~B9078 & new_n5728_;
  assign new_n6579_ = ~new_n6577_ & ~new_n6578_;
  assign new_n6580_ = ~new_n2717_ & ~new_n6579_;
  assign new_n6581_ = new_n6572_ & ~new_n6580_;
  assign new_n6582_ = B9111 & ~new_n5736_;
  assign new_n6583_ = ~B9111 & new_n5736_;
  assign new_n6584_ = ~new_n6582_ & ~new_n6583_;
  assign new_n6585_ = ~new_n2728_ & ~new_n6584_;
  assign new_n6586_ = ~new_n6580_ & ~new_n6585_;
  assign new_n6587_ = ~new_n6581_ & ~new_n6586_;
  assign new_n6588_ = new_n6576_ & new_n6587_;
  assign new_n6589_ = ~new_n6576_ & ~new_n6587_;
  assign new_n6590_ = ~new_n6588_ & ~new_n6589_;
  assign new_n6591_ = ~new_n6572_ & ~new_n6590_;
  assign new_n6592_ = new_n6531_ & ~new_n6591_;
  assign new_n6593_ = B9144 & ~new_n5750_;
  assign new_n6594_ = ~B9144 & new_n5750_;
  assign new_n6595_ = ~new_n6593_ & ~new_n6594_;
  assign new_n6596_ = ~new_n2745_ & ~new_n6595_;
  assign new_n6597_ = B9177 & ~new_n5757_;
  assign new_n6598_ = ~B9177 & new_n5757_;
  assign new_n6599_ = ~new_n6597_ & ~new_n6598_;
  assign new_n6600_ = ~new_n2755_ & ~new_n6599_;
  assign new_n6601_ = ~new_n6596_ & new_n6600_;
  assign new_n6602_ = new_n6596_ & ~new_n6600_;
  assign new_n6603_ = ~new_n6601_ & ~new_n6602_;
  assign new_n6604_ = B9210 & ~new_n5767_;
  assign new_n6605_ = ~B9210 & new_n5767_;
  assign new_n6606_ = ~new_n6604_ & ~new_n6605_;
  assign new_n6607_ = ~new_n2768_ & ~new_n6606_;
  assign new_n6608_ = B9243 & ~new_n5774_;
  assign new_n6609_ = ~B9243 & new_n5774_;
  assign new_n6610_ = ~new_n6608_ & ~new_n6609_;
  assign new_n6611_ = ~new_n2778_ & ~new_n6610_;
  assign new_n6612_ = new_n6603_ & ~new_n6611_;
  assign new_n6613_ = B9276 & ~new_n5782_;
  assign new_n6614_ = ~B9276 & new_n5782_;
  assign new_n6615_ = ~new_n6613_ & ~new_n6614_;
  assign new_n6616_ = ~new_n2789_ & ~new_n6615_;
  assign new_n6617_ = ~new_n6611_ & ~new_n6616_;
  assign new_n6618_ = ~new_n6612_ & ~new_n6617_;
  assign new_n6619_ = new_n6607_ & new_n6618_;
  assign new_n6620_ = ~new_n6607_ & ~new_n6618_;
  assign new_n6621_ = ~new_n6619_ & ~new_n6620_;
  assign new_n6622_ = ~new_n6603_ & ~new_n6621_;
  assign new_n6623_ = ~new_n6591_ & ~new_n6622_;
  assign new_n6624_ = ~new_n6592_ & ~new_n6623_;
  assign new_n6625_ = new_n6561_ & new_n6624_;
  assign new_n6626_ = ~new_n6561_ & ~new_n6624_;
  assign new_n6627_ = ~new_n6625_ & ~new_n6626_;
  assign new_n6628_ = ~new_n6531_ & ~new_n6627_;
  assign new_n6629_ = ~new_n6467_ & ~new_n6628_;
  assign new_n6630_ = ~new_n6468_ & ~new_n6629_;
  assign new_n6631_ = new_n6307_ & new_n6630_;
  assign new_n6632_ = ~new_n6307_ & ~new_n6630_;
  assign new_n6633_ = ~new_n6631_ & ~new_n6632_;
  assign A6775 = ~new_n6147_ & ~new_n6633_;
  assign new_n6635_ = ~new_n6144_ & ~new_n6631_;
  assign A6774 = ~new_n6147_ & ~new_n6635_;
  assign new_n6637_ = new_n6144_ & new_n6307_;
  assign new_n6638_ = ~new_n6147_ & ~new_n6637_;
  assign new_n6639_ = new_n6147_ & ~new_n6638_;
  assign new_n6640_ = new_n6147_ & new_n6637_;
  assign new_n6641_ = new_n6639_ & ~new_n6640_;
  assign new_n6642_ = new_n6307_ & ~new_n6641_;
  assign A6773 = new_n6630_ | new_n6642_;
  assign new_n6644_ = new_n6467_ & new_n6628_;
  assign new_n6645_ = ~new_n6629_ & ~new_n6644_;
  assign new_n6646_ = ~new_n6147_ & ~new_n6467_;
  assign new_n6647_ = new_n6147_ & new_n6467_;
  assign new_n6648_ = ~new_n6646_ & ~new_n6647_;
  assign new_n6649_ = new_n6645_ & ~new_n6648_;
  assign A6772 = new_n6642_ | new_n6649_;
  assign new_n6651_ = new_n6307_ & ~new_n6649_;
  assign new_n6652_ = ~new_n6307_ & new_n6649_;
  assign new_n6653_ = ~new_n6651_ & ~new_n6652_;
  assign A6771 = ~new_n6147_ & ~new_n6653_;
  assign new_n6655_ = ~new_n1274_ & ~new_n1311_;
  assign new_n6656_ = ~new_n1277_ & ~new_n6655_;
  assign new_n6657_ = ~new_n1334_ & ~new_n1371_;
  assign new_n6658_ = ~new_n1337_ & ~new_n6657_;
  assign new_n6659_ = ~new_n6656_ & new_n6658_;
  assign new_n6660_ = new_n6656_ & ~new_n6658_;
  assign new_n6661_ = ~new_n6659_ & ~new_n6660_;
  assign new_n6662_ = ~new_n1397_ & ~new_n1434_;
  assign new_n6663_ = ~new_n1400_ & ~new_n6662_;
  assign new_n6664_ = ~new_n1457_ & ~new_n1494_;
  assign new_n6665_ = ~new_n1460_ & ~new_n6664_;
  assign new_n6666_ = new_n6661_ & ~new_n6665_;
  assign new_n6667_ = ~new_n1518_ & ~new_n1555_;
  assign new_n6668_ = ~new_n1521_ & ~new_n6667_;
  assign new_n6669_ = ~new_n6665_ & ~new_n6668_;
  assign new_n6670_ = ~new_n6666_ & ~new_n6669_;
  assign new_n6671_ = new_n6663_ & new_n6670_;
  assign new_n6672_ = ~new_n6663_ & ~new_n6670_;
  assign new_n6673_ = ~new_n6671_ & ~new_n6672_;
  assign new_n6674_ = ~new_n6661_ & ~new_n6673_;
  assign new_n6675_ = ~new_n1584_ & ~new_n1621_;
  assign new_n6676_ = ~new_n1587_ & ~new_n6675_;
  assign new_n6677_ = ~new_n1644_ & ~new_n1681_;
  assign new_n6678_ = ~new_n1647_ & ~new_n6677_;
  assign new_n6679_ = ~new_n6676_ & new_n6678_;
  assign new_n6680_ = new_n6676_ & ~new_n6678_;
  assign new_n6681_ = ~new_n6679_ & ~new_n6680_;
  assign new_n6682_ = ~new_n1707_ & ~new_n1744_;
  assign new_n6683_ = ~new_n1710_ & ~new_n6682_;
  assign new_n6684_ = ~new_n1767_ & ~new_n1804_;
  assign new_n6685_ = ~new_n1770_ & ~new_n6684_;
  assign new_n6686_ = new_n6681_ & ~new_n6685_;
  assign new_n6687_ = ~new_n1828_ & ~new_n1865_;
  assign new_n6688_ = ~new_n1831_ & ~new_n6687_;
  assign new_n6689_ = ~new_n6685_ & ~new_n6688_;
  assign new_n6690_ = ~new_n6686_ & ~new_n6689_;
  assign new_n6691_ = new_n6683_ & new_n6690_;
  assign new_n6692_ = ~new_n6683_ & ~new_n6690_;
  assign new_n6693_ = ~new_n6691_ & ~new_n6692_;
  assign new_n6694_ = ~new_n6681_ & ~new_n6693_;
  assign new_n6695_ = ~new_n6674_ & new_n6694_;
  assign new_n6696_ = new_n6674_ & ~new_n6694_;
  assign new_n6697_ = ~new_n6695_ & ~new_n6696_;
  assign new_n6698_ = ~new_n1897_ & ~new_n1934_;
  assign new_n6699_ = ~new_n1900_ & ~new_n6698_;
  assign new_n6700_ = ~new_n1957_ & ~new_n1994_;
  assign new_n6701_ = ~new_n1960_ & ~new_n6700_;
  assign new_n6702_ = ~new_n6699_ & new_n6701_;
  assign new_n6703_ = new_n6699_ & ~new_n6701_;
  assign new_n6704_ = ~new_n6702_ & ~new_n6703_;
  assign new_n6705_ = ~new_n2020_ & ~new_n2057_;
  assign new_n6706_ = ~new_n2023_ & ~new_n6705_;
  assign new_n6707_ = ~new_n2080_ & ~new_n2117_;
  assign new_n6708_ = ~new_n2083_ & ~new_n6707_;
  assign new_n6709_ = new_n6704_ & ~new_n6708_;
  assign new_n6710_ = ~new_n2141_ & ~new_n2178_;
  assign new_n6711_ = ~new_n2144_ & ~new_n6710_;
  assign new_n6712_ = ~new_n6708_ & ~new_n6711_;
  assign new_n6713_ = ~new_n6709_ & ~new_n6712_;
  assign new_n6714_ = new_n6706_ & new_n6713_;
  assign new_n6715_ = ~new_n6706_ & ~new_n6713_;
  assign new_n6716_ = ~new_n6714_ & ~new_n6715_;
  assign new_n6717_ = ~new_n6704_ & ~new_n6716_;
  assign new_n6718_ = ~new_n2207_ & ~new_n2244_;
  assign new_n6719_ = ~new_n2210_ & ~new_n6718_;
  assign new_n6720_ = ~new_n2267_ & ~new_n2304_;
  assign new_n6721_ = ~new_n2270_ & ~new_n6720_;
  assign new_n6722_ = ~new_n6719_ & new_n6721_;
  assign new_n6723_ = new_n6719_ & ~new_n6721_;
  assign new_n6724_ = ~new_n6722_ & ~new_n6723_;
  assign new_n6725_ = ~new_n2330_ & ~new_n2367_;
  assign new_n6726_ = ~new_n2333_ & ~new_n6725_;
  assign new_n6727_ = ~new_n2390_ & ~new_n2427_;
  assign new_n6728_ = ~new_n2393_ & ~new_n6727_;
  assign new_n6729_ = new_n6724_ & ~new_n6728_;
  assign new_n6730_ = ~new_n2451_ & ~new_n2488_;
  assign new_n6731_ = ~new_n2454_ & ~new_n6730_;
  assign new_n6732_ = ~new_n6728_ & ~new_n6731_;
  assign new_n6733_ = ~new_n6729_ & ~new_n6732_;
  assign new_n6734_ = new_n6726_ & new_n6733_;
  assign new_n6735_ = ~new_n6726_ & ~new_n6733_;
  assign new_n6736_ = ~new_n6734_ & ~new_n6735_;
  assign new_n6737_ = ~new_n6724_ & ~new_n6736_;
  assign new_n6738_ = new_n6697_ & ~new_n6737_;
  assign new_n6739_ = ~new_n2518_ & ~new_n2555_;
  assign new_n6740_ = ~new_n2521_ & ~new_n6739_;
  assign new_n6741_ = ~new_n2578_ & ~new_n2615_;
  assign new_n6742_ = ~new_n2581_ & ~new_n6741_;
  assign new_n6743_ = ~new_n6740_ & new_n6742_;
  assign new_n6744_ = new_n6740_ & ~new_n6742_;
  assign new_n6745_ = ~new_n6743_ & ~new_n6744_;
  assign new_n6746_ = ~new_n2641_ & ~new_n2678_;
  assign new_n6747_ = ~new_n2644_ & ~new_n6746_;
  assign new_n6748_ = ~new_n2701_ & ~new_n2738_;
  assign new_n6749_ = ~new_n2704_ & ~new_n6748_;
  assign new_n6750_ = new_n6745_ & ~new_n6749_;
  assign new_n6751_ = ~new_n2762_ & ~new_n2799_;
  assign new_n6752_ = ~new_n2765_ & ~new_n6751_;
  assign new_n6753_ = ~new_n6749_ & ~new_n6752_;
  assign new_n6754_ = ~new_n6750_ & ~new_n6753_;
  assign new_n6755_ = new_n6747_ & new_n6754_;
  assign new_n6756_ = ~new_n6747_ & ~new_n6754_;
  assign new_n6757_ = ~new_n6755_ & ~new_n6756_;
  assign new_n6758_ = ~new_n6745_ & ~new_n6757_;
  assign new_n6759_ = ~new_n6737_ & ~new_n6758_;
  assign new_n6760_ = ~new_n6738_ & ~new_n6759_;
  assign new_n6761_ = new_n6717_ & new_n6760_;
  assign new_n6762_ = ~new_n6717_ & ~new_n6760_;
  assign new_n6763_ = ~new_n6761_ & ~new_n6762_;
  assign A6742 = ~new_n6697_ & ~new_n6763_;
  assign new_n6765_ = ~new_n6694_ & ~new_n6761_;
  assign A6741 = ~new_n6697_ & ~new_n6765_;
  assign new_n6767_ = new_n6694_ & new_n6717_;
  assign new_n6768_ = ~new_n6697_ & ~new_n6767_;
  assign new_n6769_ = new_n6697_ & ~new_n6768_;
  assign new_n6770_ = new_n6697_ & new_n6767_;
  assign new_n6771_ = new_n6769_ & ~new_n6770_;
  assign new_n6772_ = new_n6717_ & ~new_n6771_;
  assign A6740 = new_n6760_ | new_n6772_;
  assign new_n6774_ = new_n6737_ & new_n6758_;
  assign new_n6775_ = ~new_n6759_ & ~new_n6774_;
  assign new_n6776_ = ~new_n6697_ & ~new_n6737_;
  assign new_n6777_ = new_n6697_ & new_n6737_;
  assign new_n6778_ = ~new_n6776_ & ~new_n6777_;
  assign new_n6779_ = new_n6775_ & ~new_n6778_;
  assign A6739 = new_n6772_ | new_n6779_;
  assign new_n6781_ = new_n6717_ & ~new_n6779_;
  assign new_n6782_ = ~new_n6717_ & new_n6779_;
  assign new_n6783_ = ~new_n6781_ & ~new_n6782_;
  assign A6738 = ~new_n6697_ & ~new_n6783_;
  assign new_n6785_ = ~new_n2843_ & ~new_n2856_;
  assign new_n6786_ = ~new_n2846_ & ~new_n6785_;
  assign new_n6787_ = ~new_n2863_ & ~new_n2876_;
  assign new_n6788_ = ~new_n2866_ & ~new_n6787_;
  assign new_n6789_ = ~new_n6786_ & new_n6788_;
  assign new_n6790_ = new_n6786_ & ~new_n6788_;
  assign new_n6791_ = ~new_n6789_ & ~new_n6790_;
  assign new_n6792_ = ~new_n2886_ & ~new_n2899_;
  assign new_n6793_ = ~new_n2889_ & ~new_n6792_;
  assign new_n6794_ = ~new_n2906_ & ~new_n2919_;
  assign new_n6795_ = ~new_n2909_ & ~new_n6794_;
  assign new_n6796_ = new_n6791_ & ~new_n6795_;
  assign new_n6797_ = ~new_n2927_ & ~new_n2940_;
  assign new_n6798_ = ~new_n2930_ & ~new_n6797_;
  assign new_n6799_ = ~new_n6795_ & ~new_n6798_;
  assign new_n6800_ = ~new_n6796_ & ~new_n6799_;
  assign new_n6801_ = new_n6793_ & new_n6800_;
  assign new_n6802_ = ~new_n6793_ & ~new_n6800_;
  assign new_n6803_ = ~new_n6801_ & ~new_n6802_;
  assign new_n6804_ = ~new_n6791_ & ~new_n6803_;
  assign new_n6805_ = ~new_n2953_ & ~new_n2966_;
  assign new_n6806_ = ~new_n2956_ & ~new_n6805_;
  assign new_n6807_ = ~new_n2973_ & ~new_n2986_;
  assign new_n6808_ = ~new_n2976_ & ~new_n6807_;
  assign new_n6809_ = ~new_n6806_ & new_n6808_;
  assign new_n6810_ = new_n6806_ & ~new_n6808_;
  assign new_n6811_ = ~new_n6809_ & ~new_n6810_;
  assign new_n6812_ = ~new_n2996_ & ~new_n3009_;
  assign new_n6813_ = ~new_n2999_ & ~new_n6812_;
  assign new_n6814_ = ~new_n3016_ & ~new_n3029_;
  assign new_n6815_ = ~new_n3019_ & ~new_n6814_;
  assign new_n6816_ = new_n6811_ & ~new_n6815_;
  assign new_n6817_ = ~new_n3037_ & ~new_n3050_;
  assign new_n6818_ = ~new_n3040_ & ~new_n6817_;
  assign new_n6819_ = ~new_n6815_ & ~new_n6818_;
  assign new_n6820_ = ~new_n6816_ & ~new_n6819_;
  assign new_n6821_ = new_n6813_ & new_n6820_;
  assign new_n6822_ = ~new_n6813_ & ~new_n6820_;
  assign new_n6823_ = ~new_n6821_ & ~new_n6822_;
  assign new_n6824_ = ~new_n6811_ & ~new_n6823_;
  assign new_n6825_ = ~new_n6804_ & new_n6824_;
  assign new_n6826_ = new_n6804_ & ~new_n6824_;
  assign new_n6827_ = ~new_n6825_ & ~new_n6826_;
  assign new_n6828_ = ~new_n3066_ & ~new_n3079_;
  assign new_n6829_ = ~new_n3069_ & ~new_n6828_;
  assign new_n6830_ = ~new_n3086_ & ~new_n3099_;
  assign new_n6831_ = ~new_n3089_ & ~new_n6830_;
  assign new_n6832_ = ~new_n6829_ & new_n6831_;
  assign new_n6833_ = new_n6829_ & ~new_n6831_;
  assign new_n6834_ = ~new_n6832_ & ~new_n6833_;
  assign new_n6835_ = ~new_n3109_ & ~new_n3122_;
  assign new_n6836_ = ~new_n3112_ & ~new_n6835_;
  assign new_n6837_ = ~new_n3129_ & ~new_n3142_;
  assign new_n6838_ = ~new_n3132_ & ~new_n6837_;
  assign new_n6839_ = new_n6834_ & ~new_n6838_;
  assign new_n6840_ = ~new_n3150_ & ~new_n3163_;
  assign new_n6841_ = ~new_n3153_ & ~new_n6840_;
  assign new_n6842_ = ~new_n6838_ & ~new_n6841_;
  assign new_n6843_ = ~new_n6839_ & ~new_n6842_;
  assign new_n6844_ = new_n6836_ & new_n6843_;
  assign new_n6845_ = ~new_n6836_ & ~new_n6843_;
  assign new_n6846_ = ~new_n6844_ & ~new_n6845_;
  assign new_n6847_ = ~new_n6834_ & ~new_n6846_;
  assign new_n6848_ = ~new_n3176_ & ~new_n3189_;
  assign new_n6849_ = ~new_n3179_ & ~new_n6848_;
  assign new_n6850_ = ~new_n3196_ & ~new_n3209_;
  assign new_n6851_ = ~new_n3199_ & ~new_n6850_;
  assign new_n6852_ = ~new_n6849_ & new_n6851_;
  assign new_n6853_ = new_n6849_ & ~new_n6851_;
  assign new_n6854_ = ~new_n6852_ & ~new_n6853_;
  assign new_n6855_ = ~new_n3219_ & ~new_n3232_;
  assign new_n6856_ = ~new_n3222_ & ~new_n6855_;
  assign new_n6857_ = ~new_n3239_ & ~new_n3252_;
  assign new_n6858_ = ~new_n3242_ & ~new_n6857_;
  assign new_n6859_ = new_n6854_ & ~new_n6858_;
  assign new_n6860_ = ~new_n3260_ & ~new_n3273_;
  assign new_n6861_ = ~new_n3263_ & ~new_n6860_;
  assign new_n6862_ = ~new_n6858_ & ~new_n6861_;
  assign new_n6863_ = ~new_n6859_ & ~new_n6862_;
  assign new_n6864_ = new_n6856_ & new_n6863_;
  assign new_n6865_ = ~new_n6856_ & ~new_n6863_;
  assign new_n6866_ = ~new_n6864_ & ~new_n6865_;
  assign new_n6867_ = ~new_n6854_ & ~new_n6866_;
  assign new_n6868_ = new_n6827_ & ~new_n6867_;
  assign new_n6869_ = ~new_n3287_ & ~new_n3300_;
  assign new_n6870_ = ~new_n3290_ & ~new_n6869_;
  assign new_n6871_ = ~new_n3307_ & ~new_n3320_;
  assign new_n6872_ = ~new_n3310_ & ~new_n6871_;
  assign new_n6873_ = ~new_n6870_ & new_n6872_;
  assign new_n6874_ = new_n6870_ & ~new_n6872_;
  assign new_n6875_ = ~new_n6873_ & ~new_n6874_;
  assign new_n6876_ = ~new_n3330_ & ~new_n3343_;
  assign new_n6877_ = ~new_n3333_ & ~new_n6876_;
  assign new_n6878_ = ~new_n3350_ & ~new_n3363_;
  assign new_n6879_ = ~new_n3353_ & ~new_n6878_;
  assign new_n6880_ = new_n6875_ & ~new_n6879_;
  assign new_n6881_ = ~new_n3371_ & ~new_n3384_;
  assign new_n6882_ = ~new_n3374_ & ~new_n6881_;
  assign new_n6883_ = ~new_n6879_ & ~new_n6882_;
  assign new_n6884_ = ~new_n6880_ & ~new_n6883_;
  assign new_n6885_ = new_n6877_ & new_n6884_;
  assign new_n6886_ = ~new_n6877_ & ~new_n6884_;
  assign new_n6887_ = ~new_n6885_ & ~new_n6886_;
  assign new_n6888_ = ~new_n6875_ & ~new_n6887_;
  assign new_n6889_ = ~new_n6867_ & ~new_n6888_;
  assign new_n6890_ = ~new_n6868_ & ~new_n6889_;
  assign new_n6891_ = new_n6847_ & new_n6890_;
  assign new_n6892_ = ~new_n6847_ & ~new_n6890_;
  assign new_n6893_ = ~new_n6891_ & ~new_n6892_;
  assign A6709 = ~new_n6827_ & ~new_n6893_;
  assign new_n6895_ = ~new_n6824_ & ~new_n6891_;
  assign A6708 = ~new_n6827_ & ~new_n6895_;
  assign new_n6897_ = new_n6824_ & new_n6847_;
  assign new_n6898_ = ~new_n6827_ & ~new_n6897_;
  assign new_n6899_ = new_n6827_ & ~new_n6898_;
  assign new_n6900_ = new_n6827_ & new_n6897_;
  assign new_n6901_ = new_n6899_ & ~new_n6900_;
  assign new_n6902_ = new_n6847_ & ~new_n6901_;
  assign A6707 = new_n6890_ | new_n6902_;
  assign new_n6904_ = new_n6867_ & new_n6888_;
  assign new_n6905_ = ~new_n6889_ & ~new_n6904_;
  assign new_n6906_ = ~new_n6827_ & ~new_n6867_;
  assign new_n6907_ = new_n6827_ & new_n6867_;
  assign new_n6908_ = ~new_n6906_ & ~new_n6907_;
  assign new_n6909_ = new_n6905_ & ~new_n6908_;
  assign A6706 = new_n6902_ | new_n6909_;
  assign new_n6911_ = new_n6847_ & ~new_n6909_;
  assign new_n6912_ = ~new_n6847_ & new_n6909_;
  assign new_n6913_ = ~new_n6911_ & ~new_n6912_;
  assign A6705 = ~new_n6827_ & ~new_n6913_;
  assign new_n6915_ = new_n3429_ & ~new_n3457_;
  assign new_n6916_ = ~new_n3432_ & ~new_n6915_;
  assign new_n6917_ = new_n3474_ & ~new_n3502_;
  assign new_n6918_ = ~new_n3477_ & ~new_n6917_;
  assign new_n6919_ = ~new_n6916_ & new_n6918_;
  assign new_n6920_ = new_n6916_ & ~new_n6918_;
  assign new_n6921_ = ~new_n6919_ & ~new_n6920_;
  assign new_n6922_ = new_n3522_ & ~new_n3550_;
  assign new_n6923_ = ~new_n3525_ & ~new_n6922_;
  assign new_n6924_ = new_n3567_ & ~new_n3595_;
  assign new_n6925_ = ~new_n3570_ & ~new_n6924_;
  assign new_n6926_ = new_n6921_ & ~new_n6925_;
  assign new_n6927_ = new_n3613_ & ~new_n3641_;
  assign new_n6928_ = ~new_n3616_ & ~new_n6927_;
  assign new_n6929_ = ~new_n6925_ & ~new_n6928_;
  assign new_n6930_ = ~new_n6926_ & ~new_n6929_;
  assign new_n6931_ = new_n6923_ & new_n6930_;
  assign new_n6932_ = ~new_n6923_ & ~new_n6930_;
  assign new_n6933_ = ~new_n6931_ & ~new_n6932_;
  assign new_n6934_ = ~new_n6921_ & ~new_n6933_;
  assign new_n6935_ = new_n3664_ & ~new_n3692_;
  assign new_n6936_ = ~new_n3667_ & ~new_n6935_;
  assign new_n6937_ = new_n3709_ & ~new_n3737_;
  assign new_n6938_ = ~new_n3712_ & ~new_n6937_;
  assign new_n6939_ = ~new_n6936_ & new_n6938_;
  assign new_n6940_ = new_n6936_ & ~new_n6938_;
  assign new_n6941_ = ~new_n6939_ & ~new_n6940_;
  assign new_n6942_ = new_n3757_ & ~new_n3785_;
  assign new_n6943_ = ~new_n3760_ & ~new_n6942_;
  assign new_n6944_ = new_n3802_ & ~new_n3830_;
  assign new_n6945_ = ~new_n3805_ & ~new_n6944_;
  assign new_n6946_ = new_n6941_ & ~new_n6945_;
  assign new_n6947_ = new_n3848_ & ~new_n3876_;
  assign new_n6948_ = ~new_n3851_ & ~new_n6947_;
  assign new_n6949_ = ~new_n6945_ & ~new_n6948_;
  assign new_n6950_ = ~new_n6946_ & ~new_n6949_;
  assign new_n6951_ = new_n6943_ & new_n6950_;
  assign new_n6952_ = ~new_n6943_ & ~new_n6950_;
  assign new_n6953_ = ~new_n6951_ & ~new_n6952_;
  assign new_n6954_ = ~new_n6941_ & ~new_n6953_;
  assign new_n6955_ = ~new_n6934_ & new_n6954_;
  assign new_n6956_ = new_n6934_ & ~new_n6954_;
  assign new_n6957_ = ~new_n6955_ & ~new_n6956_;
  assign new_n6958_ = new_n3902_ & ~new_n3930_;
  assign new_n6959_ = ~new_n3905_ & ~new_n6958_;
  assign new_n6960_ = new_n3947_ & ~new_n3975_;
  assign new_n6961_ = ~new_n3950_ & ~new_n6960_;
  assign new_n6962_ = ~new_n6959_ & new_n6961_;
  assign new_n6963_ = new_n6959_ & ~new_n6961_;
  assign new_n6964_ = ~new_n6962_ & ~new_n6963_;
  assign new_n6965_ = new_n3995_ & ~new_n4023_;
  assign new_n6966_ = ~new_n3998_ & ~new_n6965_;
  assign new_n6967_ = new_n4040_ & ~new_n4068_;
  assign new_n6968_ = ~new_n4043_ & ~new_n6967_;
  assign new_n6969_ = new_n6964_ & ~new_n6968_;
  assign new_n6970_ = new_n4086_ & ~new_n4114_;
  assign new_n6971_ = ~new_n4089_ & ~new_n6970_;
  assign new_n6972_ = ~new_n6968_ & ~new_n6971_;
  assign new_n6973_ = ~new_n6969_ & ~new_n6972_;
  assign new_n6974_ = new_n6966_ & new_n6973_;
  assign new_n6975_ = ~new_n6966_ & ~new_n6973_;
  assign new_n6976_ = ~new_n6974_ & ~new_n6975_;
  assign new_n6977_ = ~new_n6964_ & ~new_n6976_;
  assign new_n6978_ = new_n4137_ & ~new_n4165_;
  assign new_n6979_ = ~new_n4140_ & ~new_n6978_;
  assign new_n6980_ = new_n4182_ & ~new_n4210_;
  assign new_n6981_ = ~new_n4185_ & ~new_n6980_;
  assign new_n6982_ = ~new_n6979_ & new_n6981_;
  assign new_n6983_ = new_n6979_ & ~new_n6981_;
  assign new_n6984_ = ~new_n6982_ & ~new_n6983_;
  assign new_n6985_ = new_n4230_ & ~new_n4258_;
  assign new_n6986_ = ~new_n4233_ & ~new_n6985_;
  assign new_n6987_ = new_n4275_ & ~new_n4303_;
  assign new_n6988_ = ~new_n4278_ & ~new_n6987_;
  assign new_n6989_ = new_n6984_ & ~new_n6988_;
  assign new_n6990_ = new_n4321_ & ~new_n4349_;
  assign new_n6991_ = ~new_n4324_ & ~new_n6990_;
  assign new_n6992_ = ~new_n6988_ & ~new_n6991_;
  assign new_n6993_ = ~new_n6989_ & ~new_n6992_;
  assign new_n6994_ = new_n6986_ & new_n6993_;
  assign new_n6995_ = ~new_n6986_ & ~new_n6993_;
  assign new_n6996_ = ~new_n6994_ & ~new_n6995_;
  assign new_n6997_ = ~new_n6984_ & ~new_n6996_;
  assign new_n6998_ = new_n6957_ & ~new_n6997_;
  assign new_n6999_ = new_n4373_ & ~new_n4401_;
  assign new_n7000_ = ~new_n4376_ & ~new_n6999_;
  assign new_n7001_ = new_n4418_ & ~new_n4446_;
  assign new_n7002_ = ~new_n4421_ & ~new_n7001_;
  assign new_n7003_ = ~new_n7000_ & new_n7002_;
  assign new_n7004_ = new_n7000_ & ~new_n7002_;
  assign new_n7005_ = ~new_n7003_ & ~new_n7004_;
  assign new_n7006_ = new_n4466_ & ~new_n4494_;
  assign new_n7007_ = ~new_n4469_ & ~new_n7006_;
  assign new_n7008_ = new_n4511_ & ~new_n4539_;
  assign new_n7009_ = ~new_n4514_ & ~new_n7008_;
  assign new_n7010_ = new_n7005_ & ~new_n7009_;
  assign new_n7011_ = new_n4557_ & ~new_n4585_;
  assign new_n7012_ = ~new_n4560_ & ~new_n7011_;
  assign new_n7013_ = ~new_n7009_ & ~new_n7012_;
  assign new_n7014_ = ~new_n7010_ & ~new_n7013_;
  assign new_n7015_ = new_n7007_ & new_n7014_;
  assign new_n7016_ = ~new_n7007_ & ~new_n7014_;
  assign new_n7017_ = ~new_n7015_ & ~new_n7016_;
  assign new_n7018_ = ~new_n7005_ & ~new_n7017_;
  assign new_n7019_ = ~new_n6997_ & ~new_n7018_;
  assign new_n7020_ = ~new_n6998_ & ~new_n7019_;
  assign new_n7021_ = new_n6977_ & new_n7020_;
  assign new_n7022_ = ~new_n6977_ & ~new_n7020_;
  assign new_n7023_ = ~new_n7021_ & ~new_n7022_;
  assign A6676 = ~new_n6957_ & ~new_n7023_;
  assign new_n7025_ = ~new_n6954_ & ~new_n7021_;
  assign A6675 = ~new_n6957_ & ~new_n7025_;
  assign new_n7027_ = new_n6954_ & new_n6977_;
  assign new_n7028_ = ~new_n6957_ & ~new_n7027_;
  assign new_n7029_ = new_n6957_ & ~new_n7028_;
  assign new_n7030_ = new_n6957_ & new_n7027_;
  assign new_n7031_ = new_n7029_ & ~new_n7030_;
  assign new_n7032_ = new_n6977_ & ~new_n7031_;
  assign A6674 = new_n7020_ | new_n7032_;
  assign new_n7034_ = new_n6997_ & new_n7018_;
  assign new_n7035_ = ~new_n7019_ & ~new_n7034_;
  assign new_n7036_ = ~new_n6957_ & ~new_n6997_;
  assign new_n7037_ = new_n6957_ & new_n6997_;
  assign new_n7038_ = ~new_n7036_ & ~new_n7037_;
  assign new_n7039_ = new_n7035_ & ~new_n7038_;
  assign A6673 = new_n7032_ | new_n7039_;
  assign new_n7041_ = new_n6977_ & ~new_n7039_;
  assign new_n7042_ = ~new_n6977_ & new_n7039_;
  assign new_n7043_ = ~new_n7041_ & ~new_n7042_;
  assign A6672 = ~new_n6957_ & ~new_n7043_;
  assign new_n7045_ = new_n4630_ & ~new_n4658_;
  assign new_n7046_ = ~new_n4633_ & ~new_n7045_;
  assign new_n7047_ = new_n4675_ & ~new_n4703_;
  assign new_n7048_ = ~new_n4678_ & ~new_n7047_;
  assign new_n7049_ = ~new_n7046_ & new_n7048_;
  assign new_n7050_ = new_n7046_ & ~new_n7048_;
  assign new_n7051_ = ~new_n7049_ & ~new_n7050_;
  assign new_n7052_ = new_n4723_ & ~new_n4751_;
  assign new_n7053_ = ~new_n4726_ & ~new_n7052_;
  assign new_n7054_ = new_n4768_ & ~new_n4796_;
  assign new_n7055_ = ~new_n4771_ & ~new_n7054_;
  assign new_n7056_ = new_n7051_ & ~new_n7055_;
  assign new_n7057_ = new_n4814_ & ~new_n4842_;
  assign new_n7058_ = ~new_n4817_ & ~new_n7057_;
  assign new_n7059_ = ~new_n7055_ & ~new_n7058_;
  assign new_n7060_ = ~new_n7056_ & ~new_n7059_;
  assign new_n7061_ = new_n7053_ & new_n7060_;
  assign new_n7062_ = ~new_n7053_ & ~new_n7060_;
  assign new_n7063_ = ~new_n7061_ & ~new_n7062_;
  assign new_n7064_ = ~new_n7051_ & ~new_n7063_;
  assign new_n7065_ = new_n4865_ & ~new_n4893_;
  assign new_n7066_ = ~new_n4868_ & ~new_n7065_;
  assign new_n7067_ = new_n4910_ & ~new_n4938_;
  assign new_n7068_ = ~new_n4913_ & ~new_n7067_;
  assign new_n7069_ = ~new_n7066_ & new_n7068_;
  assign new_n7070_ = new_n7066_ & ~new_n7068_;
  assign new_n7071_ = ~new_n7069_ & ~new_n7070_;
  assign new_n7072_ = new_n4958_ & ~new_n4986_;
  assign new_n7073_ = ~new_n4961_ & ~new_n7072_;
  assign new_n7074_ = new_n5003_ & ~new_n5031_;
  assign new_n7075_ = ~new_n5006_ & ~new_n7074_;
  assign new_n7076_ = new_n7071_ & ~new_n7075_;
  assign new_n7077_ = new_n5049_ & ~new_n5077_;
  assign new_n7078_ = ~new_n5052_ & ~new_n7077_;
  assign new_n7079_ = ~new_n7075_ & ~new_n7078_;
  assign new_n7080_ = ~new_n7076_ & ~new_n7079_;
  assign new_n7081_ = new_n7073_ & new_n7080_;
  assign new_n7082_ = ~new_n7073_ & ~new_n7080_;
  assign new_n7083_ = ~new_n7081_ & ~new_n7082_;
  assign new_n7084_ = ~new_n7071_ & ~new_n7083_;
  assign new_n7085_ = ~new_n7064_ & new_n7084_;
  assign new_n7086_ = new_n7064_ & ~new_n7084_;
  assign new_n7087_ = ~new_n7085_ & ~new_n7086_;
  assign new_n7088_ = new_n5103_ & ~new_n5131_;
  assign new_n7089_ = ~new_n5106_ & ~new_n7088_;
  assign new_n7090_ = new_n5148_ & ~new_n5176_;
  assign new_n7091_ = ~new_n5151_ & ~new_n7090_;
  assign new_n7092_ = ~new_n7089_ & new_n7091_;
  assign new_n7093_ = new_n7089_ & ~new_n7091_;
  assign new_n7094_ = ~new_n7092_ & ~new_n7093_;
  assign new_n7095_ = new_n5196_ & ~new_n5224_;
  assign new_n7096_ = ~new_n5199_ & ~new_n7095_;
  assign new_n7097_ = new_n5241_ & ~new_n5269_;
  assign new_n7098_ = ~new_n5244_ & ~new_n7097_;
  assign new_n7099_ = new_n7094_ & ~new_n7098_;
  assign new_n7100_ = new_n5287_ & ~new_n5315_;
  assign new_n7101_ = ~new_n5290_ & ~new_n7100_;
  assign new_n7102_ = ~new_n7098_ & ~new_n7101_;
  assign new_n7103_ = ~new_n7099_ & ~new_n7102_;
  assign new_n7104_ = new_n7096_ & new_n7103_;
  assign new_n7105_ = ~new_n7096_ & ~new_n7103_;
  assign new_n7106_ = ~new_n7104_ & ~new_n7105_;
  assign new_n7107_ = ~new_n7094_ & ~new_n7106_;
  assign new_n7108_ = new_n5338_ & ~new_n5366_;
  assign new_n7109_ = ~new_n5341_ & ~new_n7108_;
  assign new_n7110_ = new_n5383_ & ~new_n5411_;
  assign new_n7111_ = ~new_n5386_ & ~new_n7110_;
  assign new_n7112_ = ~new_n7109_ & new_n7111_;
  assign new_n7113_ = new_n7109_ & ~new_n7111_;
  assign new_n7114_ = ~new_n7112_ & ~new_n7113_;
  assign new_n7115_ = new_n5431_ & ~new_n5459_;
  assign new_n7116_ = ~new_n5434_ & ~new_n7115_;
  assign new_n7117_ = new_n5476_ & ~new_n5504_;
  assign new_n7118_ = ~new_n5479_ & ~new_n7117_;
  assign new_n7119_ = new_n7114_ & ~new_n7118_;
  assign new_n7120_ = new_n5522_ & ~new_n5550_;
  assign new_n7121_ = ~new_n5525_ & ~new_n7120_;
  assign new_n7122_ = ~new_n7118_ & ~new_n7121_;
  assign new_n7123_ = ~new_n7119_ & ~new_n7122_;
  assign new_n7124_ = new_n7116_ & new_n7123_;
  assign new_n7125_ = ~new_n7116_ & ~new_n7123_;
  assign new_n7126_ = ~new_n7124_ & ~new_n7125_;
  assign new_n7127_ = ~new_n7114_ & ~new_n7126_;
  assign new_n7128_ = new_n7087_ & ~new_n7127_;
  assign new_n7129_ = new_n5574_ & ~new_n5602_;
  assign new_n7130_ = ~new_n5577_ & ~new_n7129_;
  assign new_n7131_ = new_n5619_ & ~new_n5647_;
  assign new_n7132_ = ~new_n5622_ & ~new_n7131_;
  assign new_n7133_ = ~new_n7130_ & new_n7132_;
  assign new_n7134_ = new_n7130_ & ~new_n7132_;
  assign new_n7135_ = ~new_n7133_ & ~new_n7134_;
  assign new_n7136_ = new_n5667_ & ~new_n5695_;
  assign new_n7137_ = ~new_n5670_ & ~new_n7136_;
  assign new_n7138_ = new_n5712_ & ~new_n5740_;
  assign new_n7139_ = ~new_n5715_ & ~new_n7138_;
  assign new_n7140_ = new_n7135_ & ~new_n7139_;
  assign new_n7141_ = new_n5758_ & ~new_n5786_;
  assign new_n7142_ = ~new_n5761_ & ~new_n7141_;
  assign new_n7143_ = ~new_n7139_ & ~new_n7142_;
  assign new_n7144_ = ~new_n7140_ & ~new_n7143_;
  assign new_n7145_ = new_n7137_ & new_n7144_;
  assign new_n7146_ = ~new_n7137_ & ~new_n7144_;
  assign new_n7147_ = ~new_n7145_ & ~new_n7146_;
  assign new_n7148_ = ~new_n7135_ & ~new_n7147_;
  assign new_n7149_ = ~new_n7127_ & ~new_n7148_;
  assign new_n7150_ = ~new_n7128_ & ~new_n7149_;
  assign new_n7151_ = new_n7107_ & new_n7150_;
  assign new_n7152_ = ~new_n7107_ & ~new_n7150_;
  assign new_n7153_ = ~new_n7151_ & ~new_n7152_;
  assign A6643 = ~new_n7087_ & ~new_n7153_;
  assign new_n7155_ = ~new_n7084_ & ~new_n7151_;
  assign A6642 = ~new_n7087_ & ~new_n7155_;
  assign new_n7157_ = new_n7084_ & new_n7107_;
  assign new_n7158_ = ~new_n7087_ & ~new_n7157_;
  assign new_n7159_ = new_n7087_ & ~new_n7158_;
  assign new_n7160_ = new_n7087_ & new_n7157_;
  assign new_n7161_ = new_n7159_ & ~new_n7160_;
  assign new_n7162_ = new_n7107_ & ~new_n7161_;
  assign A6641 = new_n7150_ | new_n7162_;
  assign new_n7164_ = new_n7127_ & new_n7148_;
  assign new_n7165_ = ~new_n7149_ & ~new_n7164_;
  assign new_n7166_ = ~new_n7087_ & ~new_n7127_;
  assign new_n7167_ = new_n7087_ & new_n7127_;
  assign new_n7168_ = ~new_n7166_ & ~new_n7167_;
  assign new_n7169_ = new_n7165_ & ~new_n7168_;
  assign A6640 = new_n7162_ | new_n7169_;
  assign new_n7171_ = new_n7107_ & ~new_n7169_;
  assign new_n7172_ = ~new_n7107_ & new_n7169_;
  assign new_n7173_ = ~new_n7171_ & ~new_n7172_;
  assign A6639 = ~new_n7087_ & ~new_n7173_;
  assign new_n7175_ = new_n5839_ & new_n5850_;
  assign new_n7176_ = ~new_n5842_ & ~new_n7175_;
  assign new_n7177_ = new_n5842_ & ~new_n7176_;
  assign new_n7178_ = new_n5842_ & new_n7175_;
  assign new_n7179_ = new_n7177_ & ~new_n7178_;
  assign new_n7180_ = new_n5850_ & ~new_n7179_;
  assign new_n7181_ = ~new_n5846_ & ~new_n7180_;
  assign new_n7182_ = ~new_n5862_ & ~new_n5881_;
  assign new_n7183_ = ~new_n5865_ & ~new_n7182_;
  assign new_n7184_ = new_n7181_ & new_n7183_;
  assign new_n7185_ = ~new_n7181_ & ~new_n7183_;
  assign new_n7186_ = ~new_n7184_ & ~new_n7185_;
  assign new_n7187_ = ~new_n5895_ & ~new_n5914_;
  assign new_n7188_ = ~new_n5898_ & ~new_n7187_;
  assign new_n7189_ = ~new_n5925_ & ~new_n5944_;
  assign new_n7190_ = ~new_n5928_ & ~new_n7189_;
  assign new_n7191_ = new_n7186_ & ~new_n7190_;
  assign new_n7192_ = ~new_n5956_ & ~new_n5975_;
  assign new_n7193_ = ~new_n5959_ & ~new_n7192_;
  assign new_n7194_ = ~new_n7190_ & ~new_n7193_;
  assign new_n7195_ = ~new_n7191_ & ~new_n7194_;
  assign new_n7196_ = new_n7188_ & new_n7195_;
  assign new_n7197_ = ~new_n7188_ & ~new_n7195_;
  assign new_n7198_ = ~new_n7196_ & ~new_n7197_;
  assign new_n7199_ = ~new_n7186_ & ~new_n7198_;
  assign new_n7200_ = ~new_n5992_ & ~new_n6011_;
  assign new_n7201_ = ~new_n5995_ & ~new_n7200_;
  assign new_n7202_ = ~new_n6022_ & ~new_n6041_;
  assign new_n7203_ = ~new_n6025_ & ~new_n7202_;
  assign new_n7204_ = ~new_n7201_ & new_n7203_;
  assign new_n7205_ = new_n7201_ & ~new_n7203_;
  assign new_n7206_ = ~new_n7204_ & ~new_n7205_;
  assign new_n7207_ = ~new_n6055_ & ~new_n6074_;
  assign new_n7208_ = ~new_n6058_ & ~new_n7207_;
  assign new_n7209_ = ~new_n6085_ & ~new_n6104_;
  assign new_n7210_ = ~new_n6088_ & ~new_n7209_;
  assign new_n7211_ = new_n7206_ & ~new_n7210_;
  assign new_n7212_ = ~new_n6116_ & ~new_n6135_;
  assign new_n7213_ = ~new_n6119_ & ~new_n7212_;
  assign new_n7214_ = ~new_n7210_ & ~new_n7213_;
  assign new_n7215_ = ~new_n7211_ & ~new_n7214_;
  assign new_n7216_ = new_n7208_ & new_n7215_;
  assign new_n7217_ = ~new_n7208_ & ~new_n7215_;
  assign new_n7218_ = ~new_n7216_ & ~new_n7217_;
  assign new_n7219_ = ~new_n7206_ & ~new_n7218_;
  assign new_n7220_ = ~new_n7199_ & new_n7219_;
  assign new_n7221_ = new_n7199_ & ~new_n7219_;
  assign new_n7222_ = ~new_n7220_ & ~new_n7221_;
  assign new_n7223_ = ~new_n6155_ & ~new_n6174_;
  assign new_n7224_ = ~new_n6158_ & ~new_n7223_;
  assign new_n7225_ = ~new_n6185_ & ~new_n6204_;
  assign new_n7226_ = ~new_n6188_ & ~new_n7225_;
  assign new_n7227_ = ~new_n7224_ & new_n7226_;
  assign new_n7228_ = new_n7224_ & ~new_n7226_;
  assign new_n7229_ = ~new_n7227_ & ~new_n7228_;
  assign new_n7230_ = ~new_n6218_ & ~new_n6237_;
  assign new_n7231_ = ~new_n6221_ & ~new_n7230_;
  assign new_n7232_ = ~new_n6248_ & ~new_n6267_;
  assign new_n7233_ = ~new_n6251_ & ~new_n7232_;
  assign new_n7234_ = new_n7229_ & ~new_n7233_;
  assign new_n7235_ = ~new_n6279_ & ~new_n6298_;
  assign new_n7236_ = ~new_n6282_ & ~new_n7235_;
  assign new_n7237_ = ~new_n7233_ & ~new_n7236_;
  assign new_n7238_ = ~new_n7234_ & ~new_n7237_;
  assign new_n7239_ = new_n7231_ & new_n7238_;
  assign new_n7240_ = ~new_n7231_ & ~new_n7238_;
  assign new_n7241_ = ~new_n7239_ & ~new_n7240_;
  assign new_n7242_ = ~new_n7229_ & ~new_n7241_;
  assign new_n7243_ = ~new_n6315_ & ~new_n6334_;
  assign new_n7244_ = ~new_n6318_ & ~new_n7243_;
  assign new_n7245_ = ~new_n6345_ & ~new_n6364_;
  assign new_n7246_ = ~new_n6348_ & ~new_n7245_;
  assign new_n7247_ = ~new_n7244_ & new_n7246_;
  assign new_n7248_ = new_n7244_ & ~new_n7246_;
  assign new_n7249_ = ~new_n7247_ & ~new_n7248_;
  assign new_n7250_ = ~new_n6378_ & ~new_n6397_;
  assign new_n7251_ = ~new_n6381_ & ~new_n7250_;
  assign new_n7252_ = ~new_n6408_ & ~new_n6427_;
  assign new_n7253_ = ~new_n6411_ & ~new_n7252_;
  assign new_n7254_ = new_n7249_ & ~new_n7253_;
  assign new_n7255_ = ~new_n6439_ & ~new_n6458_;
  assign new_n7256_ = ~new_n6442_ & ~new_n7255_;
  assign new_n7257_ = ~new_n7253_ & ~new_n7256_;
  assign new_n7258_ = ~new_n7254_ & ~new_n7257_;
  assign new_n7259_ = new_n7251_ & new_n7258_;
  assign new_n7260_ = ~new_n7251_ & ~new_n7258_;
  assign new_n7261_ = ~new_n7259_ & ~new_n7260_;
  assign new_n7262_ = ~new_n7249_ & ~new_n7261_;
  assign new_n7263_ = new_n7222_ & ~new_n7262_;
  assign new_n7264_ = ~new_n6476_ & ~new_n6495_;
  assign new_n7265_ = ~new_n6479_ & ~new_n7264_;
  assign new_n7266_ = ~new_n6506_ & ~new_n6525_;
  assign new_n7267_ = ~new_n6509_ & ~new_n7266_;
  assign new_n7268_ = ~new_n7265_ & new_n7267_;
  assign new_n7269_ = new_n7265_ & ~new_n7267_;
  assign new_n7270_ = ~new_n7268_ & ~new_n7269_;
  assign new_n7271_ = ~new_n6539_ & ~new_n6558_;
  assign new_n7272_ = ~new_n6542_ & ~new_n7271_;
  assign new_n7273_ = ~new_n6569_ & ~new_n6588_;
  assign new_n7274_ = ~new_n6572_ & ~new_n7273_;
  assign new_n7275_ = new_n7270_ & ~new_n7274_;
  assign new_n7276_ = ~new_n6600_ & ~new_n6619_;
  assign new_n7277_ = ~new_n6603_ & ~new_n7276_;
  assign new_n7278_ = ~new_n7274_ & ~new_n7277_;
  assign new_n7279_ = ~new_n7275_ & ~new_n7278_;
  assign new_n7280_ = new_n7272_ & new_n7279_;
  assign new_n7281_ = ~new_n7272_ & ~new_n7279_;
  assign new_n7282_ = ~new_n7280_ & ~new_n7281_;
  assign new_n7283_ = ~new_n7270_ & ~new_n7282_;
  assign new_n7284_ = ~new_n7262_ & ~new_n7283_;
  assign new_n7285_ = ~new_n7263_ & ~new_n7284_;
  assign new_n7286_ = new_n7242_ & new_n7285_;
  assign new_n7287_ = ~new_n7242_ & ~new_n7285_;
  assign new_n7288_ = ~new_n7286_ & ~new_n7287_;
  assign A6610 = ~new_n7222_ & ~new_n7288_;
  assign new_n7290_ = ~new_n7219_ & ~new_n7286_;
  assign A6609 = ~new_n7222_ & ~new_n7290_;
  assign new_n7292_ = new_n7219_ & new_n7242_;
  assign new_n7293_ = ~new_n7222_ & ~new_n7292_;
  assign new_n7294_ = new_n7222_ & ~new_n7293_;
  assign new_n7295_ = new_n7222_ & new_n7292_;
  assign new_n7296_ = new_n7294_ & ~new_n7295_;
  assign new_n7297_ = new_n7242_ & ~new_n7296_;
  assign A6608 = new_n7285_ | new_n7297_;
  assign new_n7299_ = new_n7262_ & new_n7283_;
  assign new_n7300_ = ~new_n7284_ & ~new_n7299_;
  assign new_n7301_ = ~new_n7222_ & ~new_n7262_;
  assign new_n7302_ = new_n7222_ & new_n7262_;
  assign new_n7303_ = ~new_n7301_ & ~new_n7302_;
  assign new_n7304_ = new_n7300_ & ~new_n7303_;
  assign A6607 = new_n7297_ | new_n7304_;
  assign new_n7306_ = new_n7242_ & ~new_n7304_;
  assign new_n7307_ = ~new_n7242_ & new_n7304_;
  assign new_n7308_ = ~new_n7306_ & ~new_n7307_;
  assign A6606 = ~new_n7222_ & ~new_n7308_;
  assign new_n7310_ = new_n1274_ & new_n1287_;
  assign new_n7311_ = ~new_n1277_ & ~new_n7310_;
  assign new_n7312_ = new_n1277_ & ~new_n7311_;
  assign new_n7313_ = new_n1277_ & new_n7310_;
  assign new_n7314_ = new_n7312_ & ~new_n7313_;
  assign new_n7315_ = new_n1287_ & ~new_n7314_;
  assign new_n7316_ = ~new_n1310_ & ~new_n7315_;
  assign new_n7317_ = new_n1334_ & new_n1347_;
  assign new_n7318_ = ~new_n1337_ & ~new_n7317_;
  assign new_n7319_ = new_n1337_ & ~new_n7318_;
  assign new_n7320_ = new_n1337_ & new_n7317_;
  assign new_n7321_ = new_n7319_ & ~new_n7320_;
  assign new_n7322_ = new_n1347_ & ~new_n7321_;
  assign new_n7323_ = ~new_n1370_ & ~new_n7322_;
  assign new_n7324_ = new_n7316_ & ~new_n7323_;
  assign new_n7325_ = ~new_n7316_ & new_n7323_;
  assign new_n7326_ = ~new_n7324_ & ~new_n7325_;
  assign new_n7327_ = new_n1397_ & new_n1410_;
  assign new_n7328_ = ~new_n1400_ & ~new_n7327_;
  assign new_n7329_ = new_n1400_ & ~new_n7328_;
  assign new_n7330_ = new_n1400_ & new_n7327_;
  assign new_n7331_ = new_n7329_ & ~new_n7330_;
  assign new_n7332_ = new_n1410_ & ~new_n7331_;
  assign new_n7333_ = ~new_n1433_ & ~new_n7332_;
  assign new_n7334_ = new_n1457_ & new_n1470_;
  assign new_n7335_ = ~new_n1460_ & ~new_n7334_;
  assign new_n7336_ = new_n1460_ & ~new_n7335_;
  assign new_n7337_ = new_n1460_ & new_n7334_;
  assign new_n7338_ = new_n7336_ & ~new_n7337_;
  assign new_n7339_ = new_n1470_ & ~new_n7338_;
  assign new_n7340_ = ~new_n1493_ & ~new_n7339_;
  assign new_n7341_ = new_n7326_ & new_n7340_;
  assign new_n7342_ = new_n1518_ & new_n1531_;
  assign new_n7343_ = ~new_n1521_ & ~new_n7342_;
  assign new_n7344_ = new_n1521_ & ~new_n7343_;
  assign new_n7345_ = new_n1521_ & new_n7342_;
  assign new_n7346_ = new_n7344_ & ~new_n7345_;
  assign new_n7347_ = new_n1531_ & ~new_n7346_;
  assign new_n7348_ = ~new_n1554_ & ~new_n7347_;
  assign new_n7349_ = new_n7340_ & new_n7348_;
  assign new_n7350_ = ~new_n7341_ & ~new_n7349_;
  assign new_n7351_ = ~new_n7333_ & new_n7350_;
  assign new_n7352_ = new_n7333_ & ~new_n7350_;
  assign new_n7353_ = ~new_n7351_ & ~new_n7352_;
  assign new_n7354_ = ~new_n7326_ & ~new_n7353_;
  assign new_n7355_ = new_n1584_ & new_n1597_;
  assign new_n7356_ = ~new_n1587_ & ~new_n7355_;
  assign new_n7357_ = new_n1587_ & ~new_n7356_;
  assign new_n7358_ = new_n1587_ & new_n7355_;
  assign new_n7359_ = new_n7357_ & ~new_n7358_;
  assign new_n7360_ = new_n1597_ & ~new_n7359_;
  assign new_n7361_ = ~new_n1620_ & ~new_n7360_;
  assign new_n7362_ = new_n1644_ & new_n1657_;
  assign new_n7363_ = ~new_n1647_ & ~new_n7362_;
  assign new_n7364_ = new_n1647_ & ~new_n7363_;
  assign new_n7365_ = new_n1647_ & new_n7362_;
  assign new_n7366_ = new_n7364_ & ~new_n7365_;
  assign new_n7367_ = new_n1657_ & ~new_n7366_;
  assign new_n7368_ = ~new_n1680_ & ~new_n7367_;
  assign new_n7369_ = new_n7361_ & ~new_n7368_;
  assign new_n7370_ = ~new_n7361_ & new_n7368_;
  assign new_n7371_ = ~new_n7369_ & ~new_n7370_;
  assign new_n7372_ = new_n1707_ & new_n1720_;
  assign new_n7373_ = ~new_n1710_ & ~new_n7372_;
  assign new_n7374_ = new_n1710_ & ~new_n7373_;
  assign new_n7375_ = new_n1710_ & new_n7372_;
  assign new_n7376_ = new_n7374_ & ~new_n7375_;
  assign new_n7377_ = new_n1720_ & ~new_n7376_;
  assign new_n7378_ = ~new_n1743_ & ~new_n7377_;
  assign new_n7379_ = new_n1767_ & new_n1780_;
  assign new_n7380_ = ~new_n1770_ & ~new_n7379_;
  assign new_n7381_ = new_n1770_ & ~new_n7380_;
  assign new_n7382_ = new_n1770_ & new_n7379_;
  assign new_n7383_ = new_n7381_ & ~new_n7382_;
  assign new_n7384_ = new_n1780_ & ~new_n7383_;
  assign new_n7385_ = ~new_n1803_ & ~new_n7384_;
  assign new_n7386_ = new_n7371_ & new_n7385_;
  assign new_n7387_ = new_n1828_ & new_n1841_;
  assign new_n7388_ = ~new_n1831_ & ~new_n7387_;
  assign new_n7389_ = new_n1831_ & ~new_n7388_;
  assign new_n7390_ = new_n1831_ & new_n7387_;
  assign new_n7391_ = new_n7389_ & ~new_n7390_;
  assign new_n7392_ = new_n1841_ & ~new_n7391_;
  assign new_n7393_ = ~new_n1864_ & ~new_n7392_;
  assign new_n7394_ = new_n7385_ & new_n7393_;
  assign new_n7395_ = ~new_n7386_ & ~new_n7394_;
  assign new_n7396_ = ~new_n7378_ & new_n7395_;
  assign new_n7397_ = new_n7378_ & ~new_n7395_;
  assign new_n7398_ = ~new_n7396_ & ~new_n7397_;
  assign new_n7399_ = ~new_n7371_ & ~new_n7398_;
  assign new_n7400_ = ~new_n7354_ & new_n7399_;
  assign new_n7401_ = new_n7354_ & ~new_n7399_;
  assign new_n7402_ = ~new_n7400_ & ~new_n7401_;
  assign new_n7403_ = new_n1897_ & new_n1910_;
  assign new_n7404_ = ~new_n1900_ & ~new_n7403_;
  assign new_n7405_ = new_n1900_ & ~new_n7404_;
  assign new_n7406_ = new_n1900_ & new_n7403_;
  assign new_n7407_ = new_n7405_ & ~new_n7406_;
  assign new_n7408_ = new_n1910_ & ~new_n7407_;
  assign new_n7409_ = ~new_n1933_ & ~new_n7408_;
  assign new_n7410_ = new_n1957_ & new_n1970_;
  assign new_n7411_ = ~new_n1960_ & ~new_n7410_;
  assign new_n7412_ = new_n1960_ & ~new_n7411_;
  assign new_n7413_ = new_n1960_ & new_n7410_;
  assign new_n7414_ = new_n7412_ & ~new_n7413_;
  assign new_n7415_ = new_n1970_ & ~new_n7414_;
  assign new_n7416_ = ~new_n1993_ & ~new_n7415_;
  assign new_n7417_ = new_n7409_ & ~new_n7416_;
  assign new_n7418_ = ~new_n7409_ & new_n7416_;
  assign new_n7419_ = ~new_n7417_ & ~new_n7418_;
  assign new_n7420_ = new_n2020_ & new_n2033_;
  assign new_n7421_ = ~new_n2023_ & ~new_n7420_;
  assign new_n7422_ = new_n2023_ & ~new_n7421_;
  assign new_n7423_ = new_n2023_ & new_n7420_;
  assign new_n7424_ = new_n7422_ & ~new_n7423_;
  assign new_n7425_ = new_n2033_ & ~new_n7424_;
  assign new_n7426_ = ~new_n2056_ & ~new_n7425_;
  assign new_n7427_ = new_n2080_ & new_n2093_;
  assign new_n7428_ = ~new_n2083_ & ~new_n7427_;
  assign new_n7429_ = new_n2083_ & ~new_n7428_;
  assign new_n7430_ = new_n2083_ & new_n7427_;
  assign new_n7431_ = new_n7429_ & ~new_n7430_;
  assign new_n7432_ = new_n2093_ & ~new_n7431_;
  assign new_n7433_ = ~new_n2116_ & ~new_n7432_;
  assign new_n7434_ = new_n7419_ & new_n7433_;
  assign new_n7435_ = new_n2141_ & new_n2154_;
  assign new_n7436_ = ~new_n2144_ & ~new_n7435_;
  assign new_n7437_ = new_n2144_ & ~new_n7436_;
  assign new_n7438_ = new_n2144_ & new_n7435_;
  assign new_n7439_ = new_n7437_ & ~new_n7438_;
  assign new_n7440_ = new_n2154_ & ~new_n7439_;
  assign new_n7441_ = ~new_n2177_ & ~new_n7440_;
  assign new_n7442_ = new_n7433_ & new_n7441_;
  assign new_n7443_ = ~new_n7434_ & ~new_n7442_;
  assign new_n7444_ = ~new_n7426_ & new_n7443_;
  assign new_n7445_ = new_n7426_ & ~new_n7443_;
  assign new_n7446_ = ~new_n7444_ & ~new_n7445_;
  assign new_n7447_ = ~new_n7419_ & ~new_n7446_;
  assign new_n7448_ = new_n2207_ & new_n2220_;
  assign new_n7449_ = ~new_n2210_ & ~new_n7448_;
  assign new_n7450_ = new_n2210_ & ~new_n7449_;
  assign new_n7451_ = new_n2210_ & new_n7448_;
  assign new_n7452_ = new_n7450_ & ~new_n7451_;
  assign new_n7453_ = new_n2220_ & ~new_n7452_;
  assign new_n7454_ = ~new_n2243_ & ~new_n7453_;
  assign new_n7455_ = new_n2267_ & new_n2280_;
  assign new_n7456_ = ~new_n2270_ & ~new_n7455_;
  assign new_n7457_ = new_n2270_ & ~new_n7456_;
  assign new_n7458_ = new_n2270_ & new_n7455_;
  assign new_n7459_ = new_n7457_ & ~new_n7458_;
  assign new_n7460_ = new_n2280_ & ~new_n7459_;
  assign new_n7461_ = ~new_n2303_ & ~new_n7460_;
  assign new_n7462_ = new_n7454_ & ~new_n7461_;
  assign new_n7463_ = ~new_n7454_ & new_n7461_;
  assign new_n7464_ = ~new_n7462_ & ~new_n7463_;
  assign new_n7465_ = new_n2330_ & new_n2343_;
  assign new_n7466_ = ~new_n2333_ & ~new_n7465_;
  assign new_n7467_ = new_n2333_ & ~new_n7466_;
  assign new_n7468_ = new_n2333_ & new_n7465_;
  assign new_n7469_ = new_n7467_ & ~new_n7468_;
  assign new_n7470_ = new_n2343_ & ~new_n7469_;
  assign new_n7471_ = ~new_n2366_ & ~new_n7470_;
  assign new_n7472_ = new_n2390_ & new_n2403_;
  assign new_n7473_ = ~new_n2393_ & ~new_n7472_;
  assign new_n7474_ = new_n2393_ & ~new_n7473_;
  assign new_n7475_ = new_n2393_ & new_n7472_;
  assign new_n7476_ = new_n7474_ & ~new_n7475_;
  assign new_n7477_ = new_n2403_ & ~new_n7476_;
  assign new_n7478_ = ~new_n2426_ & ~new_n7477_;
  assign new_n7479_ = new_n7464_ & new_n7478_;
  assign new_n7480_ = new_n2451_ & new_n2464_;
  assign new_n7481_ = ~new_n2454_ & ~new_n7480_;
  assign new_n7482_ = new_n2454_ & ~new_n7481_;
  assign new_n7483_ = new_n2454_ & new_n7480_;
  assign new_n7484_ = new_n7482_ & ~new_n7483_;
  assign new_n7485_ = new_n2464_ & ~new_n7484_;
  assign new_n7486_ = ~new_n2487_ & ~new_n7485_;
  assign new_n7487_ = new_n7478_ & new_n7486_;
  assign new_n7488_ = ~new_n7479_ & ~new_n7487_;
  assign new_n7489_ = ~new_n7471_ & new_n7488_;
  assign new_n7490_ = new_n7471_ & ~new_n7488_;
  assign new_n7491_ = ~new_n7489_ & ~new_n7490_;
  assign new_n7492_ = ~new_n7464_ & ~new_n7491_;
  assign new_n7493_ = new_n7402_ & ~new_n7492_;
  assign new_n7494_ = new_n2518_ & new_n2531_;
  assign new_n7495_ = ~new_n2521_ & ~new_n7494_;
  assign new_n7496_ = new_n2521_ & ~new_n7495_;
  assign new_n7497_ = new_n2521_ & new_n7494_;
  assign new_n7498_ = new_n7496_ & ~new_n7497_;
  assign new_n7499_ = new_n2531_ & ~new_n7498_;
  assign new_n7500_ = ~new_n2554_ & ~new_n7499_;
  assign new_n7501_ = new_n2578_ & new_n2591_;
  assign new_n7502_ = ~new_n2581_ & ~new_n7501_;
  assign new_n7503_ = new_n2581_ & ~new_n7502_;
  assign new_n7504_ = new_n2581_ & new_n7501_;
  assign new_n7505_ = new_n7503_ & ~new_n7504_;
  assign new_n7506_ = new_n2591_ & ~new_n7505_;
  assign new_n7507_ = ~new_n2614_ & ~new_n7506_;
  assign new_n7508_ = new_n7500_ & ~new_n7507_;
  assign new_n7509_ = ~new_n7500_ & new_n7507_;
  assign new_n7510_ = ~new_n7508_ & ~new_n7509_;
  assign new_n7511_ = new_n2641_ & new_n2654_;
  assign new_n7512_ = ~new_n2644_ & ~new_n7511_;
  assign new_n7513_ = new_n2644_ & ~new_n7512_;
  assign new_n7514_ = new_n2644_ & new_n7511_;
  assign new_n7515_ = new_n7513_ & ~new_n7514_;
  assign new_n7516_ = new_n2654_ & ~new_n7515_;
  assign new_n7517_ = ~new_n2677_ & ~new_n7516_;
  assign new_n7518_ = new_n2701_ & new_n2714_;
  assign new_n7519_ = ~new_n2704_ & ~new_n7518_;
  assign new_n7520_ = new_n2704_ & ~new_n7519_;
  assign new_n7521_ = new_n2704_ & new_n7518_;
  assign new_n7522_ = new_n7520_ & ~new_n7521_;
  assign new_n7523_ = new_n2714_ & ~new_n7522_;
  assign new_n7524_ = ~new_n2737_ & ~new_n7523_;
  assign new_n7525_ = new_n7510_ & new_n7524_;
  assign new_n7526_ = new_n2762_ & new_n2775_;
  assign new_n7527_ = ~new_n2765_ & ~new_n7526_;
  assign new_n7528_ = new_n2765_ & ~new_n7527_;
  assign new_n7529_ = new_n2765_ & new_n7526_;
  assign new_n7530_ = new_n7528_ & ~new_n7529_;
  assign new_n7531_ = new_n2775_ & ~new_n7530_;
  assign new_n7532_ = ~new_n2798_ & ~new_n7531_;
  assign new_n7533_ = new_n7524_ & new_n7532_;
  assign new_n7534_ = ~new_n7525_ & ~new_n7533_;
  assign new_n7535_ = ~new_n7517_ & new_n7534_;
  assign new_n7536_ = new_n7517_ & ~new_n7534_;
  assign new_n7537_ = ~new_n7535_ & ~new_n7536_;
  assign new_n7538_ = ~new_n7510_ & ~new_n7537_;
  assign new_n7539_ = ~new_n7492_ & ~new_n7538_;
  assign new_n7540_ = ~new_n7493_ & ~new_n7539_;
  assign new_n7541_ = new_n7447_ & new_n7540_;
  assign new_n7542_ = ~new_n7447_ & ~new_n7540_;
  assign new_n7543_ = ~new_n7541_ & ~new_n7542_;
  assign A6577 = ~new_n7402_ & ~new_n7543_;
  assign new_n7545_ = ~new_n7399_ & ~new_n7541_;
  assign A6576 = ~new_n7402_ & ~new_n7545_;
  assign new_n7547_ = new_n7399_ & new_n7447_;
  assign new_n7548_ = ~new_n7402_ & ~new_n7547_;
  assign new_n7549_ = new_n7402_ & ~new_n7548_;
  assign new_n7550_ = new_n7402_ & new_n7547_;
  assign new_n7551_ = new_n7549_ & ~new_n7550_;
  assign new_n7552_ = new_n7447_ & ~new_n7551_;
  assign A6575 = new_n7540_ | new_n7552_;
  assign new_n7554_ = new_n7492_ & new_n7538_;
  assign new_n7555_ = ~new_n7539_ & ~new_n7554_;
  assign new_n7556_ = ~new_n7402_ & ~new_n7492_;
  assign new_n7557_ = new_n7402_ & new_n7492_;
  assign new_n7558_ = ~new_n7556_ & ~new_n7557_;
  assign new_n7559_ = new_n7555_ & ~new_n7558_;
  assign A6574 = new_n7552_ | new_n7559_;
  assign new_n7561_ = new_n7447_ & ~new_n7559_;
  assign new_n7562_ = ~new_n7447_ & new_n7559_;
  assign new_n7563_ = ~new_n7561_ & ~new_n7562_;
  assign A6573 = ~new_n7402_ & ~new_n7563_;
  assign new_n7565_ = new_n2843_ & new_n2848_;
  assign new_n7566_ = ~new_n2846_ & ~new_n7565_;
  assign new_n7567_ = new_n2846_ & ~new_n7566_;
  assign new_n7568_ = new_n2846_ & new_n7565_;
  assign new_n7569_ = new_n7567_ & ~new_n7568_;
  assign new_n7570_ = new_n2848_ & ~new_n7569_;
  assign new_n7571_ = ~new_n2855_ & ~new_n7570_;
  assign new_n7572_ = new_n2863_ & new_n2868_;
  assign new_n7573_ = ~new_n2866_ & ~new_n7572_;
  assign new_n7574_ = new_n2866_ & ~new_n7573_;
  assign new_n7575_ = new_n2866_ & new_n7572_;
  assign new_n7576_ = new_n7574_ & ~new_n7575_;
  assign new_n7577_ = new_n2868_ & ~new_n7576_;
  assign new_n7578_ = ~new_n2875_ & ~new_n7577_;
  assign new_n7579_ = new_n7571_ & ~new_n7578_;
  assign new_n7580_ = ~new_n7571_ & new_n7578_;
  assign new_n7581_ = ~new_n7579_ & ~new_n7580_;
  assign new_n7582_ = new_n2886_ & new_n2891_;
  assign new_n7583_ = ~new_n2889_ & ~new_n7582_;
  assign new_n7584_ = new_n2889_ & ~new_n7583_;
  assign new_n7585_ = new_n2889_ & new_n7582_;
  assign new_n7586_ = new_n7584_ & ~new_n7585_;
  assign new_n7587_ = new_n2891_ & ~new_n7586_;
  assign new_n7588_ = ~new_n2898_ & ~new_n7587_;
  assign new_n7589_ = new_n2906_ & new_n2911_;
  assign new_n7590_ = ~new_n2909_ & ~new_n7589_;
  assign new_n7591_ = new_n2909_ & ~new_n7590_;
  assign new_n7592_ = new_n2909_ & new_n7589_;
  assign new_n7593_ = new_n7591_ & ~new_n7592_;
  assign new_n7594_ = new_n2911_ & ~new_n7593_;
  assign new_n7595_ = ~new_n2918_ & ~new_n7594_;
  assign new_n7596_ = new_n7581_ & new_n7595_;
  assign new_n7597_ = new_n2927_ & new_n2932_;
  assign new_n7598_ = ~new_n2930_ & ~new_n7597_;
  assign new_n7599_ = new_n2930_ & ~new_n7598_;
  assign new_n7600_ = new_n2930_ & new_n7597_;
  assign new_n7601_ = new_n7599_ & ~new_n7600_;
  assign new_n7602_ = new_n2932_ & ~new_n7601_;
  assign new_n7603_ = ~new_n2939_ & ~new_n7602_;
  assign new_n7604_ = new_n7595_ & new_n7603_;
  assign new_n7605_ = ~new_n7596_ & ~new_n7604_;
  assign new_n7606_ = ~new_n7588_ & new_n7605_;
  assign new_n7607_ = new_n7588_ & ~new_n7605_;
  assign new_n7608_ = ~new_n7606_ & ~new_n7607_;
  assign new_n7609_ = ~new_n7581_ & ~new_n7608_;
  assign new_n7610_ = new_n2953_ & new_n2958_;
  assign new_n7611_ = ~new_n2956_ & ~new_n7610_;
  assign new_n7612_ = new_n2956_ & ~new_n7611_;
  assign new_n7613_ = new_n2956_ & new_n7610_;
  assign new_n7614_ = new_n7612_ & ~new_n7613_;
  assign new_n7615_ = new_n2958_ & ~new_n7614_;
  assign new_n7616_ = ~new_n2965_ & ~new_n7615_;
  assign new_n7617_ = new_n2973_ & new_n2978_;
  assign new_n7618_ = ~new_n2976_ & ~new_n7617_;
  assign new_n7619_ = new_n2976_ & ~new_n7618_;
  assign new_n7620_ = new_n2976_ & new_n7617_;
  assign new_n7621_ = new_n7619_ & ~new_n7620_;
  assign new_n7622_ = new_n2978_ & ~new_n7621_;
  assign new_n7623_ = ~new_n2985_ & ~new_n7622_;
  assign new_n7624_ = new_n7616_ & ~new_n7623_;
  assign new_n7625_ = ~new_n7616_ & new_n7623_;
  assign new_n7626_ = ~new_n7624_ & ~new_n7625_;
  assign new_n7627_ = new_n2996_ & new_n3001_;
  assign new_n7628_ = ~new_n2999_ & ~new_n7627_;
  assign new_n7629_ = new_n2999_ & ~new_n7628_;
  assign new_n7630_ = new_n2999_ & new_n7627_;
  assign new_n7631_ = new_n7629_ & ~new_n7630_;
  assign new_n7632_ = new_n3001_ & ~new_n7631_;
  assign new_n7633_ = ~new_n3008_ & ~new_n7632_;
  assign new_n7634_ = new_n3016_ & new_n3021_;
  assign new_n7635_ = ~new_n3019_ & ~new_n7634_;
  assign new_n7636_ = new_n3019_ & ~new_n7635_;
  assign new_n7637_ = new_n3019_ & new_n7634_;
  assign new_n7638_ = new_n7636_ & ~new_n7637_;
  assign new_n7639_ = new_n3021_ & ~new_n7638_;
  assign new_n7640_ = ~new_n3028_ & ~new_n7639_;
  assign new_n7641_ = new_n7626_ & new_n7640_;
  assign new_n7642_ = new_n3037_ & new_n3042_;
  assign new_n7643_ = ~new_n3040_ & ~new_n7642_;
  assign new_n7644_ = new_n3040_ & ~new_n7643_;
  assign new_n7645_ = new_n3040_ & new_n7642_;
  assign new_n7646_ = new_n7644_ & ~new_n7645_;
  assign new_n7647_ = new_n3042_ & ~new_n7646_;
  assign new_n7648_ = ~new_n3049_ & ~new_n7647_;
  assign new_n7649_ = new_n7640_ & new_n7648_;
  assign new_n7650_ = ~new_n7641_ & ~new_n7649_;
  assign new_n7651_ = ~new_n7633_ & new_n7650_;
  assign new_n7652_ = new_n7633_ & ~new_n7650_;
  assign new_n7653_ = ~new_n7651_ & ~new_n7652_;
  assign new_n7654_ = ~new_n7626_ & ~new_n7653_;
  assign new_n7655_ = ~new_n7609_ & new_n7654_;
  assign new_n7656_ = new_n7609_ & ~new_n7654_;
  assign new_n7657_ = ~new_n7655_ & ~new_n7656_;
  assign new_n7658_ = new_n3066_ & new_n3071_;
  assign new_n7659_ = ~new_n3069_ & ~new_n7658_;
  assign new_n7660_ = new_n3069_ & ~new_n7659_;
  assign new_n7661_ = new_n3069_ & new_n7658_;
  assign new_n7662_ = new_n7660_ & ~new_n7661_;
  assign new_n7663_ = new_n3071_ & ~new_n7662_;
  assign new_n7664_ = ~new_n3078_ & ~new_n7663_;
  assign new_n7665_ = new_n3086_ & new_n3091_;
  assign new_n7666_ = ~new_n3089_ & ~new_n7665_;
  assign new_n7667_ = new_n3089_ & ~new_n7666_;
  assign new_n7668_ = new_n3089_ & new_n7665_;
  assign new_n7669_ = new_n7667_ & ~new_n7668_;
  assign new_n7670_ = new_n3091_ & ~new_n7669_;
  assign new_n7671_ = ~new_n3098_ & ~new_n7670_;
  assign new_n7672_ = new_n7664_ & ~new_n7671_;
  assign new_n7673_ = ~new_n7664_ & new_n7671_;
  assign new_n7674_ = ~new_n7672_ & ~new_n7673_;
  assign new_n7675_ = new_n3109_ & new_n3114_;
  assign new_n7676_ = ~new_n3112_ & ~new_n7675_;
  assign new_n7677_ = new_n3112_ & ~new_n7676_;
  assign new_n7678_ = new_n3112_ & new_n7675_;
  assign new_n7679_ = new_n7677_ & ~new_n7678_;
  assign new_n7680_ = new_n3114_ & ~new_n7679_;
  assign new_n7681_ = ~new_n3121_ & ~new_n7680_;
  assign new_n7682_ = new_n3129_ & new_n3134_;
  assign new_n7683_ = ~new_n3132_ & ~new_n7682_;
  assign new_n7684_ = new_n3132_ & ~new_n7683_;
  assign new_n7685_ = new_n3132_ & new_n7682_;
  assign new_n7686_ = new_n7684_ & ~new_n7685_;
  assign new_n7687_ = new_n3134_ & ~new_n7686_;
  assign new_n7688_ = ~new_n3141_ & ~new_n7687_;
  assign new_n7689_ = new_n7674_ & new_n7688_;
  assign new_n7690_ = new_n3150_ & new_n3155_;
  assign new_n7691_ = ~new_n3153_ & ~new_n7690_;
  assign new_n7692_ = new_n3153_ & ~new_n7691_;
  assign new_n7693_ = new_n3153_ & new_n7690_;
  assign new_n7694_ = new_n7692_ & ~new_n7693_;
  assign new_n7695_ = new_n3155_ & ~new_n7694_;
  assign new_n7696_ = ~new_n3162_ & ~new_n7695_;
  assign new_n7697_ = new_n7688_ & new_n7696_;
  assign new_n7698_ = ~new_n7689_ & ~new_n7697_;
  assign new_n7699_ = ~new_n7681_ & new_n7698_;
  assign new_n7700_ = new_n7681_ & ~new_n7698_;
  assign new_n7701_ = ~new_n7699_ & ~new_n7700_;
  assign new_n7702_ = ~new_n7674_ & ~new_n7701_;
  assign new_n7703_ = new_n3176_ & new_n3181_;
  assign new_n7704_ = ~new_n3179_ & ~new_n7703_;
  assign new_n7705_ = new_n3179_ & ~new_n7704_;
  assign new_n7706_ = new_n3179_ & new_n7703_;
  assign new_n7707_ = new_n7705_ & ~new_n7706_;
  assign new_n7708_ = new_n3181_ & ~new_n7707_;
  assign new_n7709_ = ~new_n3188_ & ~new_n7708_;
  assign new_n7710_ = new_n3196_ & new_n3201_;
  assign new_n7711_ = ~new_n3199_ & ~new_n7710_;
  assign new_n7712_ = new_n3199_ & ~new_n7711_;
  assign new_n7713_ = new_n3199_ & new_n7710_;
  assign new_n7714_ = new_n7712_ & ~new_n7713_;
  assign new_n7715_ = new_n3201_ & ~new_n7714_;
  assign new_n7716_ = ~new_n3208_ & ~new_n7715_;
  assign new_n7717_ = new_n7709_ & ~new_n7716_;
  assign new_n7718_ = ~new_n7709_ & new_n7716_;
  assign new_n7719_ = ~new_n7717_ & ~new_n7718_;
  assign new_n7720_ = new_n3219_ & new_n3224_;
  assign new_n7721_ = ~new_n3222_ & ~new_n7720_;
  assign new_n7722_ = new_n3222_ & ~new_n7721_;
  assign new_n7723_ = new_n3222_ & new_n7720_;
  assign new_n7724_ = new_n7722_ & ~new_n7723_;
  assign new_n7725_ = new_n3224_ & ~new_n7724_;
  assign new_n7726_ = ~new_n3231_ & ~new_n7725_;
  assign new_n7727_ = new_n3239_ & new_n3244_;
  assign new_n7728_ = ~new_n3242_ & ~new_n7727_;
  assign new_n7729_ = new_n3242_ & ~new_n7728_;
  assign new_n7730_ = new_n3242_ & new_n7727_;
  assign new_n7731_ = new_n7729_ & ~new_n7730_;
  assign new_n7732_ = new_n3244_ & ~new_n7731_;
  assign new_n7733_ = ~new_n3251_ & ~new_n7732_;
  assign new_n7734_ = new_n7719_ & new_n7733_;
  assign new_n7735_ = new_n3260_ & new_n3265_;
  assign new_n7736_ = ~new_n3263_ & ~new_n7735_;
  assign new_n7737_ = new_n3263_ & ~new_n7736_;
  assign new_n7738_ = new_n3263_ & new_n7735_;
  assign new_n7739_ = new_n7737_ & ~new_n7738_;
  assign new_n7740_ = new_n3265_ & ~new_n7739_;
  assign new_n7741_ = ~new_n3272_ & ~new_n7740_;
  assign new_n7742_ = new_n7733_ & new_n7741_;
  assign new_n7743_ = ~new_n7734_ & ~new_n7742_;
  assign new_n7744_ = ~new_n7726_ & new_n7743_;
  assign new_n7745_ = new_n7726_ & ~new_n7743_;
  assign new_n7746_ = ~new_n7744_ & ~new_n7745_;
  assign new_n7747_ = ~new_n7719_ & ~new_n7746_;
  assign new_n7748_ = new_n7657_ & ~new_n7747_;
  assign new_n7749_ = new_n3287_ & new_n3292_;
  assign new_n7750_ = ~new_n3290_ & ~new_n7749_;
  assign new_n7751_ = new_n3290_ & ~new_n7750_;
  assign new_n7752_ = new_n3290_ & new_n7749_;
  assign new_n7753_ = new_n7751_ & ~new_n7752_;
  assign new_n7754_ = new_n3292_ & ~new_n7753_;
  assign new_n7755_ = ~new_n3299_ & ~new_n7754_;
  assign new_n7756_ = new_n3307_ & new_n3312_;
  assign new_n7757_ = ~new_n3310_ & ~new_n7756_;
  assign new_n7758_ = new_n3310_ & ~new_n7757_;
  assign new_n7759_ = new_n3310_ & new_n7756_;
  assign new_n7760_ = new_n7758_ & ~new_n7759_;
  assign new_n7761_ = new_n3312_ & ~new_n7760_;
  assign new_n7762_ = ~new_n3319_ & ~new_n7761_;
  assign new_n7763_ = new_n7755_ & ~new_n7762_;
  assign new_n7764_ = ~new_n7755_ & new_n7762_;
  assign new_n7765_ = ~new_n7763_ & ~new_n7764_;
  assign new_n7766_ = new_n3330_ & new_n3335_;
  assign new_n7767_ = ~new_n3333_ & ~new_n7766_;
  assign new_n7768_ = new_n3333_ & ~new_n7767_;
  assign new_n7769_ = new_n3333_ & new_n7766_;
  assign new_n7770_ = new_n7768_ & ~new_n7769_;
  assign new_n7771_ = new_n3335_ & ~new_n7770_;
  assign new_n7772_ = ~new_n3342_ & ~new_n7771_;
  assign new_n7773_ = new_n3350_ & new_n3355_;
  assign new_n7774_ = ~new_n3353_ & ~new_n7773_;
  assign new_n7775_ = new_n3353_ & ~new_n7774_;
  assign new_n7776_ = new_n3353_ & new_n7773_;
  assign new_n7777_ = new_n7775_ & ~new_n7776_;
  assign new_n7778_ = new_n3355_ & ~new_n7777_;
  assign new_n7779_ = ~new_n3362_ & ~new_n7778_;
  assign new_n7780_ = new_n7765_ & new_n7779_;
  assign new_n7781_ = new_n3371_ & new_n3376_;
  assign new_n7782_ = ~new_n3374_ & ~new_n7781_;
  assign new_n7783_ = new_n3374_ & ~new_n7782_;
  assign new_n7784_ = new_n3374_ & new_n7781_;
  assign new_n7785_ = new_n7783_ & ~new_n7784_;
  assign new_n7786_ = new_n3376_ & ~new_n7785_;
  assign new_n7787_ = ~new_n3383_ & ~new_n7786_;
  assign new_n7788_ = new_n7779_ & new_n7787_;
  assign new_n7789_ = ~new_n7780_ & ~new_n7788_;
  assign new_n7790_ = ~new_n7772_ & new_n7789_;
  assign new_n7791_ = new_n7772_ & ~new_n7789_;
  assign new_n7792_ = ~new_n7790_ & ~new_n7791_;
  assign new_n7793_ = ~new_n7765_ & ~new_n7792_;
  assign new_n7794_ = ~new_n7747_ & ~new_n7793_;
  assign new_n7795_ = ~new_n7748_ & ~new_n7794_;
  assign new_n7796_ = new_n7702_ & new_n7795_;
  assign new_n7797_ = ~new_n7702_ & ~new_n7795_;
  assign new_n7798_ = ~new_n7796_ & ~new_n7797_;
  assign A6544 = ~new_n7657_ & ~new_n7798_;
  assign new_n7800_ = ~new_n7654_ & ~new_n7796_;
  assign A6543 = ~new_n7657_ & ~new_n7800_;
  assign new_n7802_ = new_n7654_ & new_n7702_;
  assign new_n7803_ = ~new_n7657_ & ~new_n7802_;
  assign new_n7804_ = new_n7657_ & ~new_n7803_;
  assign new_n7805_ = new_n7657_ & new_n7802_;
  assign new_n7806_ = new_n7804_ & ~new_n7805_;
  assign new_n7807_ = new_n7702_ & ~new_n7806_;
  assign A6542 = new_n7795_ | new_n7807_;
  assign new_n7809_ = new_n7747_ & new_n7793_;
  assign new_n7810_ = ~new_n7794_ & ~new_n7809_;
  assign new_n7811_ = ~new_n7657_ & ~new_n7747_;
  assign new_n7812_ = new_n7657_ & new_n7747_;
  assign new_n7813_ = ~new_n7811_ & ~new_n7812_;
  assign new_n7814_ = new_n7810_ & ~new_n7813_;
  assign A6541 = new_n7807_ | new_n7814_;
  assign new_n7816_ = new_n7702_ & ~new_n7814_;
  assign new_n7817_ = ~new_n7702_ & new_n7814_;
  assign new_n7818_ = ~new_n7816_ & ~new_n7817_;
  assign A6540 = ~new_n7657_ & ~new_n7818_;
  assign new_n7820_ = ~new_n3429_ & ~new_n3439_;
  assign new_n7821_ = ~new_n3432_ & ~new_n7820_;
  assign new_n7822_ = new_n3432_ & ~new_n7821_;
  assign new_n7823_ = new_n3432_ & new_n7820_;
  assign new_n7824_ = new_n7822_ & ~new_n7823_;
  assign new_n7825_ = ~new_n3439_ & ~new_n7824_;
  assign new_n7826_ = ~new_n3456_ & ~new_n7825_;
  assign new_n7827_ = ~new_n3474_ & ~new_n3484_;
  assign new_n7828_ = ~new_n3477_ & ~new_n7827_;
  assign new_n7829_ = new_n3477_ & ~new_n7828_;
  assign new_n7830_ = new_n3477_ & new_n7827_;
  assign new_n7831_ = new_n7829_ & ~new_n7830_;
  assign new_n7832_ = ~new_n3484_ & ~new_n7831_;
  assign new_n7833_ = ~new_n3501_ & ~new_n7832_;
  assign new_n7834_ = new_n7826_ & ~new_n7833_;
  assign new_n7835_ = ~new_n7826_ & new_n7833_;
  assign new_n7836_ = ~new_n7834_ & ~new_n7835_;
  assign new_n7837_ = ~new_n3522_ & ~new_n3532_;
  assign new_n7838_ = ~new_n3525_ & ~new_n7837_;
  assign new_n7839_ = new_n3525_ & ~new_n7838_;
  assign new_n7840_ = new_n3525_ & new_n7837_;
  assign new_n7841_ = new_n7839_ & ~new_n7840_;
  assign new_n7842_ = ~new_n3532_ & ~new_n7841_;
  assign new_n7843_ = ~new_n3549_ & ~new_n7842_;
  assign new_n7844_ = ~new_n3567_ & ~new_n3577_;
  assign new_n7845_ = ~new_n3570_ & ~new_n7844_;
  assign new_n7846_ = new_n3570_ & ~new_n7845_;
  assign new_n7847_ = new_n3570_ & new_n7844_;
  assign new_n7848_ = new_n7846_ & ~new_n7847_;
  assign new_n7849_ = ~new_n3577_ & ~new_n7848_;
  assign new_n7850_ = ~new_n3594_ & ~new_n7849_;
  assign new_n7851_ = new_n7836_ & new_n7850_;
  assign new_n7852_ = ~new_n3613_ & ~new_n3623_;
  assign new_n7853_ = ~new_n3616_ & ~new_n7852_;
  assign new_n7854_ = new_n3616_ & ~new_n7853_;
  assign new_n7855_ = new_n3616_ & new_n7852_;
  assign new_n7856_ = new_n7854_ & ~new_n7855_;
  assign new_n7857_ = ~new_n3623_ & ~new_n7856_;
  assign new_n7858_ = ~new_n3640_ & ~new_n7857_;
  assign new_n7859_ = new_n7850_ & new_n7858_;
  assign new_n7860_ = ~new_n7851_ & ~new_n7859_;
  assign new_n7861_ = ~new_n7843_ & new_n7860_;
  assign new_n7862_ = new_n7843_ & ~new_n7860_;
  assign new_n7863_ = ~new_n7861_ & ~new_n7862_;
  assign new_n7864_ = ~new_n7836_ & ~new_n7863_;
  assign new_n7865_ = ~new_n3664_ & ~new_n3674_;
  assign new_n7866_ = ~new_n3667_ & ~new_n7865_;
  assign new_n7867_ = new_n3667_ & ~new_n7866_;
  assign new_n7868_ = new_n3667_ & new_n7865_;
  assign new_n7869_ = new_n7867_ & ~new_n7868_;
  assign new_n7870_ = ~new_n3674_ & ~new_n7869_;
  assign new_n7871_ = ~new_n3691_ & ~new_n7870_;
  assign new_n7872_ = ~new_n3709_ & ~new_n3719_;
  assign new_n7873_ = ~new_n3712_ & ~new_n7872_;
  assign new_n7874_ = new_n3712_ & ~new_n7873_;
  assign new_n7875_ = new_n3712_ & new_n7872_;
  assign new_n7876_ = new_n7874_ & ~new_n7875_;
  assign new_n7877_ = ~new_n3719_ & ~new_n7876_;
  assign new_n7878_ = ~new_n3736_ & ~new_n7877_;
  assign new_n7879_ = new_n7871_ & ~new_n7878_;
  assign new_n7880_ = ~new_n7871_ & new_n7878_;
  assign new_n7881_ = ~new_n7879_ & ~new_n7880_;
  assign new_n7882_ = ~new_n3757_ & ~new_n3767_;
  assign new_n7883_ = ~new_n3760_ & ~new_n7882_;
  assign new_n7884_ = new_n3760_ & ~new_n7883_;
  assign new_n7885_ = new_n3760_ & new_n7882_;
  assign new_n7886_ = new_n7884_ & ~new_n7885_;
  assign new_n7887_ = ~new_n3767_ & ~new_n7886_;
  assign new_n7888_ = ~new_n3784_ & ~new_n7887_;
  assign new_n7889_ = ~new_n3802_ & ~new_n3812_;
  assign new_n7890_ = ~new_n3805_ & ~new_n7889_;
  assign new_n7891_ = new_n3805_ & ~new_n7890_;
  assign new_n7892_ = new_n3805_ & new_n7889_;
  assign new_n7893_ = new_n7891_ & ~new_n7892_;
  assign new_n7894_ = ~new_n3812_ & ~new_n7893_;
  assign new_n7895_ = ~new_n3829_ & ~new_n7894_;
  assign new_n7896_ = new_n7881_ & new_n7895_;
  assign new_n7897_ = ~new_n3848_ & ~new_n3858_;
  assign new_n7898_ = ~new_n3851_ & ~new_n7897_;
  assign new_n7899_ = new_n3851_ & ~new_n7898_;
  assign new_n7900_ = new_n3851_ & new_n7897_;
  assign new_n7901_ = new_n7899_ & ~new_n7900_;
  assign new_n7902_ = ~new_n3858_ & ~new_n7901_;
  assign new_n7903_ = ~new_n3875_ & ~new_n7902_;
  assign new_n7904_ = new_n7895_ & new_n7903_;
  assign new_n7905_ = ~new_n7896_ & ~new_n7904_;
  assign new_n7906_ = ~new_n7888_ & new_n7905_;
  assign new_n7907_ = new_n7888_ & ~new_n7905_;
  assign new_n7908_ = ~new_n7906_ & ~new_n7907_;
  assign new_n7909_ = ~new_n7881_ & ~new_n7908_;
  assign new_n7910_ = ~new_n7864_ & new_n7909_;
  assign new_n7911_ = new_n7864_ & ~new_n7909_;
  assign new_n7912_ = ~new_n7910_ & ~new_n7911_;
  assign new_n7913_ = ~new_n3902_ & ~new_n3912_;
  assign new_n7914_ = ~new_n3905_ & ~new_n7913_;
  assign new_n7915_ = new_n3905_ & ~new_n7914_;
  assign new_n7916_ = new_n3905_ & new_n7913_;
  assign new_n7917_ = new_n7915_ & ~new_n7916_;
  assign new_n7918_ = ~new_n3912_ & ~new_n7917_;
  assign new_n7919_ = ~new_n3929_ & ~new_n7918_;
  assign new_n7920_ = ~new_n3947_ & ~new_n3957_;
  assign new_n7921_ = ~new_n3950_ & ~new_n7920_;
  assign new_n7922_ = new_n3950_ & ~new_n7921_;
  assign new_n7923_ = new_n3950_ & new_n7920_;
  assign new_n7924_ = new_n7922_ & ~new_n7923_;
  assign new_n7925_ = ~new_n3957_ & ~new_n7924_;
  assign new_n7926_ = ~new_n3974_ & ~new_n7925_;
  assign new_n7927_ = new_n7919_ & ~new_n7926_;
  assign new_n7928_ = ~new_n7919_ & new_n7926_;
  assign new_n7929_ = ~new_n7927_ & ~new_n7928_;
  assign new_n7930_ = ~new_n3995_ & ~new_n4005_;
  assign new_n7931_ = ~new_n3998_ & ~new_n7930_;
  assign new_n7932_ = new_n3998_ & ~new_n7931_;
  assign new_n7933_ = new_n3998_ & new_n7930_;
  assign new_n7934_ = new_n7932_ & ~new_n7933_;
  assign new_n7935_ = ~new_n4005_ & ~new_n7934_;
  assign new_n7936_ = ~new_n4022_ & ~new_n7935_;
  assign new_n7937_ = ~new_n4040_ & ~new_n4050_;
  assign new_n7938_ = ~new_n4043_ & ~new_n7937_;
  assign new_n7939_ = new_n4043_ & ~new_n7938_;
  assign new_n7940_ = new_n4043_ & new_n7937_;
  assign new_n7941_ = new_n7939_ & ~new_n7940_;
  assign new_n7942_ = ~new_n4050_ & ~new_n7941_;
  assign new_n7943_ = ~new_n4067_ & ~new_n7942_;
  assign new_n7944_ = new_n7929_ & new_n7943_;
  assign new_n7945_ = ~new_n4086_ & ~new_n4096_;
  assign new_n7946_ = ~new_n4089_ & ~new_n7945_;
  assign new_n7947_ = new_n4089_ & ~new_n7946_;
  assign new_n7948_ = new_n4089_ & new_n7945_;
  assign new_n7949_ = new_n7947_ & ~new_n7948_;
  assign new_n7950_ = ~new_n4096_ & ~new_n7949_;
  assign new_n7951_ = ~new_n4113_ & ~new_n7950_;
  assign new_n7952_ = new_n7943_ & new_n7951_;
  assign new_n7953_ = ~new_n7944_ & ~new_n7952_;
  assign new_n7954_ = ~new_n7936_ & new_n7953_;
  assign new_n7955_ = new_n7936_ & ~new_n7953_;
  assign new_n7956_ = ~new_n7954_ & ~new_n7955_;
  assign new_n7957_ = ~new_n7929_ & ~new_n7956_;
  assign new_n7958_ = ~new_n4137_ & ~new_n4147_;
  assign new_n7959_ = ~new_n4140_ & ~new_n7958_;
  assign new_n7960_ = new_n4140_ & ~new_n7959_;
  assign new_n7961_ = new_n4140_ & new_n7958_;
  assign new_n7962_ = new_n7960_ & ~new_n7961_;
  assign new_n7963_ = ~new_n4147_ & ~new_n7962_;
  assign new_n7964_ = ~new_n4164_ & ~new_n7963_;
  assign new_n7965_ = ~new_n4182_ & ~new_n4192_;
  assign new_n7966_ = ~new_n4185_ & ~new_n7965_;
  assign new_n7967_ = new_n4185_ & ~new_n7966_;
  assign new_n7968_ = new_n4185_ & new_n7965_;
  assign new_n7969_ = new_n7967_ & ~new_n7968_;
  assign new_n7970_ = ~new_n4192_ & ~new_n7969_;
  assign new_n7971_ = ~new_n4209_ & ~new_n7970_;
  assign new_n7972_ = new_n7964_ & ~new_n7971_;
  assign new_n7973_ = ~new_n7964_ & new_n7971_;
  assign new_n7974_ = ~new_n7972_ & ~new_n7973_;
  assign new_n7975_ = ~new_n4230_ & ~new_n4240_;
  assign new_n7976_ = ~new_n4233_ & ~new_n7975_;
  assign new_n7977_ = new_n4233_ & ~new_n7976_;
  assign new_n7978_ = new_n4233_ & new_n7975_;
  assign new_n7979_ = new_n7977_ & ~new_n7978_;
  assign new_n7980_ = ~new_n4240_ & ~new_n7979_;
  assign new_n7981_ = ~new_n4257_ & ~new_n7980_;
  assign new_n7982_ = ~new_n4275_ & ~new_n4285_;
  assign new_n7983_ = ~new_n4278_ & ~new_n7982_;
  assign new_n7984_ = new_n4278_ & ~new_n7983_;
  assign new_n7985_ = new_n4278_ & new_n7982_;
  assign new_n7986_ = new_n7984_ & ~new_n7985_;
  assign new_n7987_ = ~new_n4285_ & ~new_n7986_;
  assign new_n7988_ = ~new_n4302_ & ~new_n7987_;
  assign new_n7989_ = new_n7974_ & new_n7988_;
  assign new_n7990_ = ~new_n4321_ & ~new_n4331_;
  assign new_n7991_ = ~new_n4324_ & ~new_n7990_;
  assign new_n7992_ = new_n4324_ & ~new_n7991_;
  assign new_n7993_ = new_n4324_ & new_n7990_;
  assign new_n7994_ = new_n7992_ & ~new_n7993_;
  assign new_n7995_ = ~new_n4331_ & ~new_n7994_;
  assign new_n7996_ = ~new_n4348_ & ~new_n7995_;
  assign new_n7997_ = new_n7988_ & new_n7996_;
  assign new_n7998_ = ~new_n7989_ & ~new_n7997_;
  assign new_n7999_ = ~new_n7981_ & new_n7998_;
  assign new_n8000_ = new_n7981_ & ~new_n7998_;
  assign new_n8001_ = ~new_n7999_ & ~new_n8000_;
  assign new_n8002_ = ~new_n7974_ & ~new_n8001_;
  assign new_n8003_ = new_n7912_ & ~new_n8002_;
  assign new_n8004_ = ~new_n4373_ & ~new_n4383_;
  assign new_n8005_ = ~new_n4376_ & ~new_n8004_;
  assign new_n8006_ = new_n4376_ & ~new_n8005_;
  assign new_n8007_ = new_n4376_ & new_n8004_;
  assign new_n8008_ = new_n8006_ & ~new_n8007_;
  assign new_n8009_ = ~new_n4383_ & ~new_n8008_;
  assign new_n8010_ = ~new_n4400_ & ~new_n8009_;
  assign new_n8011_ = ~new_n4418_ & ~new_n4428_;
  assign new_n8012_ = ~new_n4421_ & ~new_n8011_;
  assign new_n8013_ = new_n4421_ & ~new_n8012_;
  assign new_n8014_ = new_n4421_ & new_n8011_;
  assign new_n8015_ = new_n8013_ & ~new_n8014_;
  assign new_n8016_ = ~new_n4428_ & ~new_n8015_;
  assign new_n8017_ = ~new_n4445_ & ~new_n8016_;
  assign new_n8018_ = new_n8010_ & ~new_n8017_;
  assign new_n8019_ = ~new_n8010_ & new_n8017_;
  assign new_n8020_ = ~new_n8018_ & ~new_n8019_;
  assign new_n8021_ = ~new_n4466_ & ~new_n4476_;
  assign new_n8022_ = ~new_n4469_ & ~new_n8021_;
  assign new_n8023_ = new_n4469_ & ~new_n8022_;
  assign new_n8024_ = new_n4469_ & new_n8021_;
  assign new_n8025_ = new_n8023_ & ~new_n8024_;
  assign new_n8026_ = ~new_n4476_ & ~new_n8025_;
  assign new_n8027_ = ~new_n4493_ & ~new_n8026_;
  assign new_n8028_ = ~new_n4511_ & ~new_n4521_;
  assign new_n8029_ = ~new_n4514_ & ~new_n8028_;
  assign new_n8030_ = new_n4514_ & ~new_n8029_;
  assign new_n8031_ = new_n4514_ & new_n8028_;
  assign new_n8032_ = new_n8030_ & ~new_n8031_;
  assign new_n8033_ = ~new_n4521_ & ~new_n8032_;
  assign new_n8034_ = ~new_n4538_ & ~new_n8033_;
  assign new_n8035_ = new_n8020_ & new_n8034_;
  assign new_n8036_ = ~new_n4557_ & ~new_n4567_;
  assign new_n8037_ = ~new_n4560_ & ~new_n8036_;
  assign new_n8038_ = new_n4560_ & ~new_n8037_;
  assign new_n8039_ = new_n4560_ & new_n8036_;
  assign new_n8040_ = new_n8038_ & ~new_n8039_;
  assign new_n8041_ = ~new_n4567_ & ~new_n8040_;
  assign new_n8042_ = ~new_n4584_ & ~new_n8041_;
  assign new_n8043_ = new_n8034_ & new_n8042_;
  assign new_n8044_ = ~new_n8035_ & ~new_n8043_;
  assign new_n8045_ = ~new_n8027_ & new_n8044_;
  assign new_n8046_ = new_n8027_ & ~new_n8044_;
  assign new_n8047_ = ~new_n8045_ & ~new_n8046_;
  assign new_n8048_ = ~new_n8020_ & ~new_n8047_;
  assign new_n8049_ = ~new_n8002_ & ~new_n8048_;
  assign new_n8050_ = ~new_n8003_ & ~new_n8049_;
  assign new_n8051_ = new_n7957_ & new_n8050_;
  assign new_n8052_ = ~new_n7957_ & ~new_n8050_;
  assign new_n8053_ = ~new_n8051_ & ~new_n8052_;
  assign A6511 = ~new_n7912_ & ~new_n8053_;
  assign new_n8055_ = ~new_n7909_ & ~new_n8051_;
  assign A6510 = ~new_n7912_ & ~new_n8055_;
  assign new_n8057_ = new_n7909_ & new_n7957_;
  assign new_n8058_ = ~new_n7912_ & ~new_n8057_;
  assign new_n8059_ = new_n7912_ & ~new_n8058_;
  assign new_n8060_ = new_n7912_ & new_n8057_;
  assign new_n8061_ = new_n8059_ & ~new_n8060_;
  assign new_n8062_ = new_n7957_ & ~new_n8061_;
  assign A6509 = new_n8050_ | new_n8062_;
  assign new_n8064_ = new_n8002_ & new_n8048_;
  assign new_n8065_ = ~new_n8049_ & ~new_n8064_;
  assign new_n8066_ = ~new_n7912_ & ~new_n8002_;
  assign new_n8067_ = new_n7912_ & new_n8002_;
  assign new_n8068_ = ~new_n8066_ & ~new_n8067_;
  assign new_n8069_ = new_n8065_ & ~new_n8068_;
  assign A6508 = new_n8062_ | new_n8069_;
  assign new_n8071_ = new_n7957_ & ~new_n8069_;
  assign new_n8072_ = ~new_n7957_ & new_n8069_;
  assign new_n8073_ = ~new_n8071_ & ~new_n8072_;
  assign A6507 = ~new_n7912_ & ~new_n8073_;
  assign new_n8075_ = ~new_n4630_ & ~new_n4640_;
  assign new_n8076_ = ~new_n4633_ & ~new_n8075_;
  assign new_n8077_ = new_n4633_ & ~new_n8076_;
  assign new_n8078_ = new_n4633_ & new_n8075_;
  assign new_n8079_ = new_n8077_ & ~new_n8078_;
  assign new_n8080_ = ~new_n4640_ & ~new_n8079_;
  assign new_n8081_ = ~new_n4657_ & ~new_n8080_;
  assign new_n8082_ = ~new_n4675_ & ~new_n4685_;
  assign new_n8083_ = ~new_n4678_ & ~new_n8082_;
  assign new_n8084_ = new_n4678_ & ~new_n8083_;
  assign new_n8085_ = new_n4678_ & new_n8082_;
  assign new_n8086_ = new_n8084_ & ~new_n8085_;
  assign new_n8087_ = ~new_n4685_ & ~new_n8086_;
  assign new_n8088_ = ~new_n4702_ & ~new_n8087_;
  assign new_n8089_ = new_n8081_ & ~new_n8088_;
  assign new_n8090_ = ~new_n8081_ & new_n8088_;
  assign new_n8091_ = ~new_n8089_ & ~new_n8090_;
  assign new_n8092_ = ~new_n4723_ & ~new_n4733_;
  assign new_n8093_ = ~new_n4726_ & ~new_n8092_;
  assign new_n8094_ = new_n4726_ & ~new_n8093_;
  assign new_n8095_ = new_n4726_ & new_n8092_;
  assign new_n8096_ = new_n8094_ & ~new_n8095_;
  assign new_n8097_ = ~new_n4733_ & ~new_n8096_;
  assign new_n8098_ = ~new_n4750_ & ~new_n8097_;
  assign new_n8099_ = ~new_n4768_ & ~new_n4778_;
  assign new_n8100_ = ~new_n4771_ & ~new_n8099_;
  assign new_n8101_ = new_n4771_ & ~new_n8100_;
  assign new_n8102_ = new_n4771_ & new_n8099_;
  assign new_n8103_ = new_n8101_ & ~new_n8102_;
  assign new_n8104_ = ~new_n4778_ & ~new_n8103_;
  assign new_n8105_ = ~new_n4795_ & ~new_n8104_;
  assign new_n8106_ = new_n8091_ & new_n8105_;
  assign new_n8107_ = ~new_n4814_ & ~new_n4824_;
  assign new_n8108_ = ~new_n4817_ & ~new_n8107_;
  assign new_n8109_ = new_n4817_ & ~new_n8108_;
  assign new_n8110_ = new_n4817_ & new_n8107_;
  assign new_n8111_ = new_n8109_ & ~new_n8110_;
  assign new_n8112_ = ~new_n4824_ & ~new_n8111_;
  assign new_n8113_ = ~new_n4841_ & ~new_n8112_;
  assign new_n8114_ = new_n8105_ & new_n8113_;
  assign new_n8115_ = ~new_n8106_ & ~new_n8114_;
  assign new_n8116_ = ~new_n8098_ & new_n8115_;
  assign new_n8117_ = new_n8098_ & ~new_n8115_;
  assign new_n8118_ = ~new_n8116_ & ~new_n8117_;
  assign new_n8119_ = ~new_n8091_ & ~new_n8118_;
  assign new_n8120_ = ~new_n4865_ & ~new_n4875_;
  assign new_n8121_ = ~new_n4868_ & ~new_n8120_;
  assign new_n8122_ = new_n4868_ & ~new_n8121_;
  assign new_n8123_ = new_n4868_ & new_n8120_;
  assign new_n8124_ = new_n8122_ & ~new_n8123_;
  assign new_n8125_ = ~new_n4875_ & ~new_n8124_;
  assign new_n8126_ = ~new_n4892_ & ~new_n8125_;
  assign new_n8127_ = ~new_n4910_ & ~new_n4920_;
  assign new_n8128_ = ~new_n4913_ & ~new_n8127_;
  assign new_n8129_ = new_n4913_ & ~new_n8128_;
  assign new_n8130_ = new_n4913_ & new_n8127_;
  assign new_n8131_ = new_n8129_ & ~new_n8130_;
  assign new_n8132_ = ~new_n4920_ & ~new_n8131_;
  assign new_n8133_ = ~new_n4937_ & ~new_n8132_;
  assign new_n8134_ = new_n8126_ & ~new_n8133_;
  assign new_n8135_ = ~new_n8126_ & new_n8133_;
  assign new_n8136_ = ~new_n8134_ & ~new_n8135_;
  assign new_n8137_ = ~new_n4958_ & ~new_n4968_;
  assign new_n8138_ = ~new_n4961_ & ~new_n8137_;
  assign new_n8139_ = new_n4961_ & ~new_n8138_;
  assign new_n8140_ = new_n4961_ & new_n8137_;
  assign new_n8141_ = new_n8139_ & ~new_n8140_;
  assign new_n8142_ = ~new_n4968_ & ~new_n8141_;
  assign new_n8143_ = ~new_n4985_ & ~new_n8142_;
  assign new_n8144_ = ~new_n5003_ & ~new_n5013_;
  assign new_n8145_ = ~new_n5006_ & ~new_n8144_;
  assign new_n8146_ = new_n5006_ & ~new_n8145_;
  assign new_n8147_ = new_n5006_ & new_n8144_;
  assign new_n8148_ = new_n8146_ & ~new_n8147_;
  assign new_n8149_ = ~new_n5013_ & ~new_n8148_;
  assign new_n8150_ = ~new_n5030_ & ~new_n8149_;
  assign new_n8151_ = new_n8136_ & new_n8150_;
  assign new_n8152_ = ~new_n5049_ & ~new_n5059_;
  assign new_n8153_ = ~new_n5052_ & ~new_n8152_;
  assign new_n8154_ = new_n5052_ & ~new_n8153_;
  assign new_n8155_ = new_n5052_ & new_n8152_;
  assign new_n8156_ = new_n8154_ & ~new_n8155_;
  assign new_n8157_ = ~new_n5059_ & ~new_n8156_;
  assign new_n8158_ = ~new_n5076_ & ~new_n8157_;
  assign new_n8159_ = new_n8150_ & new_n8158_;
  assign new_n8160_ = ~new_n8151_ & ~new_n8159_;
  assign new_n8161_ = ~new_n8143_ & new_n8160_;
  assign new_n8162_ = new_n8143_ & ~new_n8160_;
  assign new_n8163_ = ~new_n8161_ & ~new_n8162_;
  assign new_n8164_ = ~new_n8136_ & ~new_n8163_;
  assign new_n8165_ = ~new_n8119_ & new_n8164_;
  assign new_n8166_ = new_n8119_ & ~new_n8164_;
  assign new_n8167_ = ~new_n8165_ & ~new_n8166_;
  assign new_n8168_ = ~new_n5103_ & ~new_n5113_;
  assign new_n8169_ = ~new_n5106_ & ~new_n8168_;
  assign new_n8170_ = new_n5106_ & ~new_n8169_;
  assign new_n8171_ = new_n5106_ & new_n8168_;
  assign new_n8172_ = new_n8170_ & ~new_n8171_;
  assign new_n8173_ = ~new_n5113_ & ~new_n8172_;
  assign new_n8174_ = ~new_n5130_ & ~new_n8173_;
  assign new_n8175_ = ~new_n5148_ & ~new_n5158_;
  assign new_n8176_ = ~new_n5151_ & ~new_n8175_;
  assign new_n8177_ = new_n5151_ & ~new_n8176_;
  assign new_n8178_ = new_n5151_ & new_n8175_;
  assign new_n8179_ = new_n8177_ & ~new_n8178_;
  assign new_n8180_ = ~new_n5158_ & ~new_n8179_;
  assign new_n8181_ = ~new_n5175_ & ~new_n8180_;
  assign new_n8182_ = new_n8174_ & ~new_n8181_;
  assign new_n8183_ = ~new_n8174_ & new_n8181_;
  assign new_n8184_ = ~new_n8182_ & ~new_n8183_;
  assign new_n8185_ = ~new_n5196_ & ~new_n5206_;
  assign new_n8186_ = ~new_n5199_ & ~new_n8185_;
  assign new_n8187_ = new_n5199_ & ~new_n8186_;
  assign new_n8188_ = new_n5199_ & new_n8185_;
  assign new_n8189_ = new_n8187_ & ~new_n8188_;
  assign new_n8190_ = ~new_n5206_ & ~new_n8189_;
  assign new_n8191_ = ~new_n5223_ & ~new_n8190_;
  assign new_n8192_ = ~new_n5241_ & ~new_n5251_;
  assign new_n8193_ = ~new_n5244_ & ~new_n8192_;
  assign new_n8194_ = new_n5244_ & ~new_n8193_;
  assign new_n8195_ = new_n5244_ & new_n8192_;
  assign new_n8196_ = new_n8194_ & ~new_n8195_;
  assign new_n8197_ = ~new_n5251_ & ~new_n8196_;
  assign new_n8198_ = ~new_n5268_ & ~new_n8197_;
  assign new_n8199_ = new_n8184_ & new_n8198_;
  assign new_n8200_ = ~new_n5287_ & ~new_n5297_;
  assign new_n8201_ = ~new_n5290_ & ~new_n8200_;
  assign new_n8202_ = new_n5290_ & ~new_n8201_;
  assign new_n8203_ = new_n5290_ & new_n8200_;
  assign new_n8204_ = new_n8202_ & ~new_n8203_;
  assign new_n8205_ = ~new_n5297_ & ~new_n8204_;
  assign new_n8206_ = ~new_n5314_ & ~new_n8205_;
  assign new_n8207_ = new_n8198_ & new_n8206_;
  assign new_n8208_ = ~new_n8199_ & ~new_n8207_;
  assign new_n8209_ = ~new_n8191_ & new_n8208_;
  assign new_n8210_ = new_n8191_ & ~new_n8208_;
  assign new_n8211_ = ~new_n8209_ & ~new_n8210_;
  assign new_n8212_ = ~new_n8184_ & ~new_n8211_;
  assign new_n8213_ = ~new_n5338_ & ~new_n5348_;
  assign new_n8214_ = ~new_n5341_ & ~new_n8213_;
  assign new_n8215_ = new_n5341_ & ~new_n8214_;
  assign new_n8216_ = new_n5341_ & new_n8213_;
  assign new_n8217_ = new_n8215_ & ~new_n8216_;
  assign new_n8218_ = ~new_n5348_ & ~new_n8217_;
  assign new_n8219_ = ~new_n5365_ & ~new_n8218_;
  assign new_n8220_ = ~new_n5383_ & ~new_n5393_;
  assign new_n8221_ = ~new_n5386_ & ~new_n8220_;
  assign new_n8222_ = new_n5386_ & ~new_n8221_;
  assign new_n8223_ = new_n5386_ & new_n8220_;
  assign new_n8224_ = new_n8222_ & ~new_n8223_;
  assign new_n8225_ = ~new_n5393_ & ~new_n8224_;
  assign new_n8226_ = ~new_n5410_ & ~new_n8225_;
  assign new_n8227_ = new_n8219_ & ~new_n8226_;
  assign new_n8228_ = ~new_n8219_ & new_n8226_;
  assign new_n8229_ = ~new_n8227_ & ~new_n8228_;
  assign new_n8230_ = ~new_n5431_ & ~new_n5441_;
  assign new_n8231_ = ~new_n5434_ & ~new_n8230_;
  assign new_n8232_ = new_n5434_ & ~new_n8231_;
  assign new_n8233_ = new_n5434_ & new_n8230_;
  assign new_n8234_ = new_n8232_ & ~new_n8233_;
  assign new_n8235_ = ~new_n5441_ & ~new_n8234_;
  assign new_n8236_ = ~new_n5458_ & ~new_n8235_;
  assign new_n8237_ = ~new_n5476_ & ~new_n5486_;
  assign new_n8238_ = ~new_n5479_ & ~new_n8237_;
  assign new_n8239_ = new_n5479_ & ~new_n8238_;
  assign new_n8240_ = new_n5479_ & new_n8237_;
  assign new_n8241_ = new_n8239_ & ~new_n8240_;
  assign new_n8242_ = ~new_n5486_ & ~new_n8241_;
  assign new_n8243_ = ~new_n5503_ & ~new_n8242_;
  assign new_n8244_ = new_n8229_ & new_n8243_;
  assign new_n8245_ = ~new_n5522_ & ~new_n5532_;
  assign new_n8246_ = ~new_n5525_ & ~new_n8245_;
  assign new_n8247_ = new_n5525_ & ~new_n8246_;
  assign new_n8248_ = new_n5525_ & new_n8245_;
  assign new_n8249_ = new_n8247_ & ~new_n8248_;
  assign new_n8250_ = ~new_n5532_ & ~new_n8249_;
  assign new_n8251_ = ~new_n5549_ & ~new_n8250_;
  assign new_n8252_ = new_n8243_ & new_n8251_;
  assign new_n8253_ = ~new_n8244_ & ~new_n8252_;
  assign new_n8254_ = ~new_n8236_ & new_n8253_;
  assign new_n8255_ = new_n8236_ & ~new_n8253_;
  assign new_n8256_ = ~new_n8254_ & ~new_n8255_;
  assign new_n8257_ = ~new_n8229_ & ~new_n8256_;
  assign new_n8258_ = new_n8167_ & ~new_n8257_;
  assign new_n8259_ = ~new_n5574_ & ~new_n5584_;
  assign new_n8260_ = ~new_n5577_ & ~new_n8259_;
  assign new_n8261_ = new_n5577_ & ~new_n8260_;
  assign new_n8262_ = new_n5577_ & new_n8259_;
  assign new_n8263_ = new_n8261_ & ~new_n8262_;
  assign new_n8264_ = ~new_n5584_ & ~new_n8263_;
  assign new_n8265_ = ~new_n5601_ & ~new_n8264_;
  assign new_n8266_ = ~new_n5619_ & ~new_n5629_;
  assign new_n8267_ = ~new_n5622_ & ~new_n8266_;
  assign new_n8268_ = new_n5622_ & ~new_n8267_;
  assign new_n8269_ = new_n5622_ & new_n8266_;
  assign new_n8270_ = new_n8268_ & ~new_n8269_;
  assign new_n8271_ = ~new_n5629_ & ~new_n8270_;
  assign new_n8272_ = ~new_n5646_ & ~new_n8271_;
  assign new_n8273_ = new_n8265_ & ~new_n8272_;
  assign new_n8274_ = ~new_n8265_ & new_n8272_;
  assign new_n8275_ = ~new_n8273_ & ~new_n8274_;
  assign new_n8276_ = ~new_n5667_ & ~new_n5677_;
  assign new_n8277_ = ~new_n5670_ & ~new_n8276_;
  assign new_n8278_ = new_n5670_ & ~new_n8277_;
  assign new_n8279_ = new_n5670_ & new_n8276_;
  assign new_n8280_ = new_n8278_ & ~new_n8279_;
  assign new_n8281_ = ~new_n5677_ & ~new_n8280_;
  assign new_n8282_ = ~new_n5694_ & ~new_n8281_;
  assign new_n8283_ = ~new_n5712_ & ~new_n5722_;
  assign new_n8284_ = ~new_n5715_ & ~new_n8283_;
  assign new_n8285_ = new_n5715_ & ~new_n8284_;
  assign new_n8286_ = new_n5715_ & new_n8283_;
  assign new_n8287_ = new_n8285_ & ~new_n8286_;
  assign new_n8288_ = ~new_n5722_ & ~new_n8287_;
  assign new_n8289_ = ~new_n5739_ & ~new_n8288_;
  assign new_n8290_ = new_n8275_ & new_n8289_;
  assign new_n8291_ = ~new_n5758_ & ~new_n5768_;
  assign new_n8292_ = ~new_n5761_ & ~new_n8291_;
  assign new_n8293_ = new_n5761_ & ~new_n8292_;
  assign new_n8294_ = new_n5761_ & new_n8291_;
  assign new_n8295_ = new_n8293_ & ~new_n8294_;
  assign new_n8296_ = ~new_n5768_ & ~new_n8295_;
  assign new_n8297_ = ~new_n5785_ & ~new_n8296_;
  assign new_n8298_ = new_n8289_ & new_n8297_;
  assign new_n8299_ = ~new_n8290_ & ~new_n8298_;
  assign new_n8300_ = ~new_n8282_ & new_n8299_;
  assign new_n8301_ = new_n8282_ & ~new_n8299_;
  assign new_n8302_ = ~new_n8300_ & ~new_n8301_;
  assign new_n8303_ = ~new_n8275_ & ~new_n8302_;
  assign new_n8304_ = ~new_n8257_ & ~new_n8303_;
  assign new_n8305_ = ~new_n8258_ & ~new_n8304_;
  assign new_n8306_ = new_n8212_ & new_n8305_;
  assign new_n8307_ = ~new_n8212_ & ~new_n8305_;
  assign new_n8308_ = ~new_n8306_ & ~new_n8307_;
  assign A6478 = ~new_n8167_ & ~new_n8308_;
  assign new_n8310_ = ~new_n8164_ & ~new_n8306_;
  assign A6477 = ~new_n8167_ & ~new_n8310_;
  assign new_n8312_ = new_n8164_ & new_n8212_;
  assign new_n8313_ = ~new_n8167_ & ~new_n8312_;
  assign new_n8314_ = new_n8167_ & ~new_n8313_;
  assign new_n8315_ = new_n8167_ & new_n8312_;
  assign new_n8316_ = new_n8314_ & ~new_n8315_;
  assign new_n8317_ = new_n8212_ & ~new_n8316_;
  assign A6476 = new_n8305_ | new_n8317_;
  assign new_n8319_ = new_n8257_ & new_n8303_;
  assign new_n8320_ = ~new_n8304_ & ~new_n8319_;
  assign new_n8321_ = ~new_n8167_ & ~new_n8257_;
  assign new_n8322_ = new_n8167_ & new_n8257_;
  assign new_n8323_ = ~new_n8321_ & ~new_n8322_;
  assign new_n8324_ = new_n8320_ & ~new_n8323_;
  assign A6475 = new_n8317_ | new_n8324_;
  assign new_n8326_ = new_n8212_ & ~new_n8324_;
  assign new_n8327_ = ~new_n8212_ & new_n8324_;
  assign new_n8328_ = ~new_n8326_ & ~new_n8327_;
  assign A6474 = ~new_n8167_ & ~new_n8328_;
  assign new_n8330_ = ~new_n5825_ & new_n5842_;
  assign new_n8331_ = ~new_n5830_ & ~new_n8330_;
  assign new_n8332_ = ~new_n7180_ & ~new_n8331_;
  assign new_n8333_ = new_n5862_ & new_n5869_;
  assign new_n8334_ = ~new_n5865_ & ~new_n8333_;
  assign new_n8335_ = new_n5865_ & ~new_n8334_;
  assign new_n8336_ = new_n5865_ & new_n8333_;
  assign new_n8337_ = new_n8335_ & ~new_n8336_;
  assign new_n8338_ = new_n5869_ & ~new_n8337_;
  assign new_n8339_ = ~new_n5880_ & ~new_n8338_;
  assign new_n8340_ = new_n8332_ & ~new_n8339_;
  assign new_n8341_ = ~new_n8332_ & new_n8339_;
  assign new_n8342_ = ~new_n8340_ & ~new_n8341_;
  assign new_n8343_ = new_n5895_ & new_n5902_;
  assign new_n8344_ = ~new_n5898_ & ~new_n8343_;
  assign new_n8345_ = new_n5898_ & ~new_n8344_;
  assign new_n8346_ = new_n5898_ & new_n8343_;
  assign new_n8347_ = new_n8345_ & ~new_n8346_;
  assign new_n8348_ = new_n5902_ & ~new_n8347_;
  assign new_n8349_ = ~new_n5913_ & ~new_n8348_;
  assign new_n8350_ = new_n5925_ & new_n5932_;
  assign new_n8351_ = ~new_n5928_ & ~new_n8350_;
  assign new_n8352_ = new_n5928_ & ~new_n8351_;
  assign new_n8353_ = new_n5928_ & new_n8350_;
  assign new_n8354_ = new_n8352_ & ~new_n8353_;
  assign new_n8355_ = new_n5932_ & ~new_n8354_;
  assign new_n8356_ = ~new_n5943_ & ~new_n8355_;
  assign new_n8357_ = new_n8342_ & new_n8356_;
  assign new_n8358_ = new_n5956_ & new_n5963_;
  assign new_n8359_ = ~new_n5959_ & ~new_n8358_;
  assign new_n8360_ = new_n5959_ & ~new_n8359_;
  assign new_n8361_ = new_n5959_ & new_n8358_;
  assign new_n8362_ = new_n8360_ & ~new_n8361_;
  assign new_n8363_ = new_n5963_ & ~new_n8362_;
  assign new_n8364_ = ~new_n5974_ & ~new_n8363_;
  assign new_n8365_ = new_n8356_ & new_n8364_;
  assign new_n8366_ = ~new_n8357_ & ~new_n8365_;
  assign new_n8367_ = ~new_n8349_ & new_n8366_;
  assign new_n8368_ = new_n8349_ & ~new_n8366_;
  assign new_n8369_ = ~new_n8367_ & ~new_n8368_;
  assign new_n8370_ = ~new_n8342_ & ~new_n8369_;
  assign new_n8371_ = new_n5992_ & new_n5999_;
  assign new_n8372_ = ~new_n5995_ & ~new_n8371_;
  assign new_n8373_ = new_n5995_ & ~new_n8372_;
  assign new_n8374_ = new_n5995_ & new_n8371_;
  assign new_n8375_ = new_n8373_ & ~new_n8374_;
  assign new_n8376_ = new_n5999_ & ~new_n8375_;
  assign new_n8377_ = ~new_n6010_ & ~new_n8376_;
  assign new_n8378_ = new_n6022_ & new_n6029_;
  assign new_n8379_ = ~new_n6025_ & ~new_n8378_;
  assign new_n8380_ = new_n6025_ & ~new_n8379_;
  assign new_n8381_ = new_n6025_ & new_n8378_;
  assign new_n8382_ = new_n8380_ & ~new_n8381_;
  assign new_n8383_ = new_n6029_ & ~new_n8382_;
  assign new_n8384_ = ~new_n6040_ & ~new_n8383_;
  assign new_n8385_ = new_n8377_ & ~new_n8384_;
  assign new_n8386_ = ~new_n8377_ & new_n8384_;
  assign new_n8387_ = ~new_n8385_ & ~new_n8386_;
  assign new_n8388_ = new_n6055_ & new_n6062_;
  assign new_n8389_ = ~new_n6058_ & ~new_n8388_;
  assign new_n8390_ = new_n6058_ & ~new_n8389_;
  assign new_n8391_ = new_n6058_ & new_n8388_;
  assign new_n8392_ = new_n8390_ & ~new_n8391_;
  assign new_n8393_ = new_n6062_ & ~new_n8392_;
  assign new_n8394_ = ~new_n6073_ & ~new_n8393_;
  assign new_n8395_ = new_n6085_ & new_n6092_;
  assign new_n8396_ = ~new_n6088_ & ~new_n8395_;
  assign new_n8397_ = new_n6088_ & ~new_n8396_;
  assign new_n8398_ = new_n6088_ & new_n8395_;
  assign new_n8399_ = new_n8397_ & ~new_n8398_;
  assign new_n8400_ = new_n6092_ & ~new_n8399_;
  assign new_n8401_ = ~new_n6103_ & ~new_n8400_;
  assign new_n8402_ = new_n8387_ & new_n8401_;
  assign new_n8403_ = new_n6116_ & new_n6123_;
  assign new_n8404_ = ~new_n6119_ & ~new_n8403_;
  assign new_n8405_ = new_n6119_ & ~new_n8404_;
  assign new_n8406_ = new_n6119_ & new_n8403_;
  assign new_n8407_ = new_n8405_ & ~new_n8406_;
  assign new_n8408_ = new_n6123_ & ~new_n8407_;
  assign new_n8409_ = ~new_n6134_ & ~new_n8408_;
  assign new_n8410_ = new_n8401_ & new_n8409_;
  assign new_n8411_ = ~new_n8402_ & ~new_n8410_;
  assign new_n8412_ = ~new_n8394_ & new_n8411_;
  assign new_n8413_ = new_n8394_ & ~new_n8411_;
  assign new_n8414_ = ~new_n8412_ & ~new_n8413_;
  assign new_n8415_ = ~new_n8387_ & ~new_n8414_;
  assign new_n8416_ = ~new_n8370_ & new_n8415_;
  assign new_n8417_ = new_n8370_ & ~new_n8415_;
  assign new_n8418_ = ~new_n8416_ & ~new_n8417_;
  assign new_n8419_ = new_n6155_ & new_n6162_;
  assign new_n8420_ = ~new_n6158_ & ~new_n8419_;
  assign new_n8421_ = new_n6158_ & ~new_n8420_;
  assign new_n8422_ = new_n6158_ & new_n8419_;
  assign new_n8423_ = new_n8421_ & ~new_n8422_;
  assign new_n8424_ = new_n6162_ & ~new_n8423_;
  assign new_n8425_ = ~new_n6173_ & ~new_n8424_;
  assign new_n8426_ = new_n6185_ & new_n6192_;
  assign new_n8427_ = ~new_n6188_ & ~new_n8426_;
  assign new_n8428_ = new_n6188_ & ~new_n8427_;
  assign new_n8429_ = new_n6188_ & new_n8426_;
  assign new_n8430_ = new_n8428_ & ~new_n8429_;
  assign new_n8431_ = new_n6192_ & ~new_n8430_;
  assign new_n8432_ = ~new_n6203_ & ~new_n8431_;
  assign new_n8433_ = new_n8425_ & ~new_n8432_;
  assign new_n8434_ = ~new_n8425_ & new_n8432_;
  assign new_n8435_ = ~new_n8433_ & ~new_n8434_;
  assign new_n8436_ = new_n6218_ & new_n6225_;
  assign new_n8437_ = ~new_n6221_ & ~new_n8436_;
  assign new_n8438_ = new_n6221_ & ~new_n8437_;
  assign new_n8439_ = new_n6221_ & new_n8436_;
  assign new_n8440_ = new_n8438_ & ~new_n8439_;
  assign new_n8441_ = new_n6225_ & ~new_n8440_;
  assign new_n8442_ = ~new_n6236_ & ~new_n8441_;
  assign new_n8443_ = new_n6248_ & new_n6255_;
  assign new_n8444_ = ~new_n6251_ & ~new_n8443_;
  assign new_n8445_ = new_n6251_ & ~new_n8444_;
  assign new_n8446_ = new_n6251_ & new_n8443_;
  assign new_n8447_ = new_n8445_ & ~new_n8446_;
  assign new_n8448_ = new_n6255_ & ~new_n8447_;
  assign new_n8449_ = ~new_n6266_ & ~new_n8448_;
  assign new_n8450_ = new_n8435_ & new_n8449_;
  assign new_n8451_ = new_n6279_ & new_n6286_;
  assign new_n8452_ = ~new_n6282_ & ~new_n8451_;
  assign new_n8453_ = new_n6282_ & ~new_n8452_;
  assign new_n8454_ = new_n6282_ & new_n8451_;
  assign new_n8455_ = new_n8453_ & ~new_n8454_;
  assign new_n8456_ = new_n6286_ & ~new_n8455_;
  assign new_n8457_ = ~new_n6297_ & ~new_n8456_;
  assign new_n8458_ = new_n8449_ & new_n8457_;
  assign new_n8459_ = ~new_n8450_ & ~new_n8458_;
  assign new_n8460_ = ~new_n8442_ & new_n8459_;
  assign new_n8461_ = new_n8442_ & ~new_n8459_;
  assign new_n8462_ = ~new_n8460_ & ~new_n8461_;
  assign new_n8463_ = ~new_n8435_ & ~new_n8462_;
  assign new_n8464_ = new_n6315_ & new_n6322_;
  assign new_n8465_ = ~new_n6318_ & ~new_n8464_;
  assign new_n8466_ = new_n6318_ & ~new_n8465_;
  assign new_n8467_ = new_n6318_ & new_n8464_;
  assign new_n8468_ = new_n8466_ & ~new_n8467_;
  assign new_n8469_ = new_n6322_ & ~new_n8468_;
  assign new_n8470_ = ~new_n6333_ & ~new_n8469_;
  assign new_n8471_ = new_n6345_ & new_n6352_;
  assign new_n8472_ = ~new_n6348_ & ~new_n8471_;
  assign new_n8473_ = new_n6348_ & ~new_n8472_;
  assign new_n8474_ = new_n6348_ & new_n8471_;
  assign new_n8475_ = new_n8473_ & ~new_n8474_;
  assign new_n8476_ = new_n6352_ & ~new_n8475_;
  assign new_n8477_ = ~new_n6363_ & ~new_n8476_;
  assign new_n8478_ = new_n8470_ & ~new_n8477_;
  assign new_n8479_ = ~new_n8470_ & new_n8477_;
  assign new_n8480_ = ~new_n8478_ & ~new_n8479_;
  assign new_n8481_ = new_n6378_ & new_n6385_;
  assign new_n8482_ = ~new_n6381_ & ~new_n8481_;
  assign new_n8483_ = new_n6381_ & ~new_n8482_;
  assign new_n8484_ = new_n6381_ & new_n8481_;
  assign new_n8485_ = new_n8483_ & ~new_n8484_;
  assign new_n8486_ = new_n6385_ & ~new_n8485_;
  assign new_n8487_ = ~new_n6396_ & ~new_n8486_;
  assign new_n8488_ = new_n6408_ & new_n6415_;
  assign new_n8489_ = ~new_n6411_ & ~new_n8488_;
  assign new_n8490_ = new_n6411_ & ~new_n8489_;
  assign new_n8491_ = new_n6411_ & new_n8488_;
  assign new_n8492_ = new_n8490_ & ~new_n8491_;
  assign new_n8493_ = new_n6415_ & ~new_n8492_;
  assign new_n8494_ = ~new_n6426_ & ~new_n8493_;
  assign new_n8495_ = new_n8480_ & new_n8494_;
  assign new_n8496_ = new_n6439_ & new_n6446_;
  assign new_n8497_ = ~new_n6442_ & ~new_n8496_;
  assign new_n8498_ = new_n6442_ & ~new_n8497_;
  assign new_n8499_ = new_n6442_ & new_n8496_;
  assign new_n8500_ = new_n8498_ & ~new_n8499_;
  assign new_n8501_ = new_n6446_ & ~new_n8500_;
  assign new_n8502_ = ~new_n6457_ & ~new_n8501_;
  assign new_n8503_ = new_n8494_ & new_n8502_;
  assign new_n8504_ = ~new_n8495_ & ~new_n8503_;
  assign new_n8505_ = ~new_n8487_ & new_n8504_;
  assign new_n8506_ = new_n8487_ & ~new_n8504_;
  assign new_n8507_ = ~new_n8505_ & ~new_n8506_;
  assign new_n8508_ = ~new_n8480_ & ~new_n8507_;
  assign new_n8509_ = new_n8418_ & ~new_n8508_;
  assign new_n8510_ = new_n6476_ & new_n6483_;
  assign new_n8511_ = ~new_n6479_ & ~new_n8510_;
  assign new_n8512_ = new_n6479_ & ~new_n8511_;
  assign new_n8513_ = new_n6479_ & new_n8510_;
  assign new_n8514_ = new_n8512_ & ~new_n8513_;
  assign new_n8515_ = new_n6483_ & ~new_n8514_;
  assign new_n8516_ = ~new_n6494_ & ~new_n8515_;
  assign new_n8517_ = new_n6506_ & new_n6513_;
  assign new_n8518_ = ~new_n6509_ & ~new_n8517_;
  assign new_n8519_ = new_n6509_ & ~new_n8518_;
  assign new_n8520_ = new_n6509_ & new_n8517_;
  assign new_n8521_ = new_n8519_ & ~new_n8520_;
  assign new_n8522_ = new_n6513_ & ~new_n8521_;
  assign new_n8523_ = ~new_n6524_ & ~new_n8522_;
  assign new_n8524_ = new_n8516_ & ~new_n8523_;
  assign new_n8525_ = ~new_n8516_ & new_n8523_;
  assign new_n8526_ = ~new_n8524_ & ~new_n8525_;
  assign new_n8527_ = new_n6539_ & new_n6546_;
  assign new_n8528_ = ~new_n6542_ & ~new_n8527_;
  assign new_n8529_ = new_n6542_ & ~new_n8528_;
  assign new_n8530_ = new_n6542_ & new_n8527_;
  assign new_n8531_ = new_n8529_ & ~new_n8530_;
  assign new_n8532_ = new_n6546_ & ~new_n8531_;
  assign new_n8533_ = ~new_n6557_ & ~new_n8532_;
  assign new_n8534_ = new_n6569_ & new_n6576_;
  assign new_n8535_ = ~new_n6572_ & ~new_n8534_;
  assign new_n8536_ = new_n6572_ & ~new_n8535_;
  assign new_n8537_ = new_n6572_ & new_n8534_;
  assign new_n8538_ = new_n8536_ & ~new_n8537_;
  assign new_n8539_ = new_n6576_ & ~new_n8538_;
  assign new_n8540_ = ~new_n6587_ & ~new_n8539_;
  assign new_n8541_ = new_n8526_ & new_n8540_;
  assign new_n8542_ = new_n6600_ & new_n6607_;
  assign new_n8543_ = ~new_n6603_ & ~new_n8542_;
  assign new_n8544_ = new_n6603_ & ~new_n8543_;
  assign new_n8545_ = new_n6603_ & new_n8542_;
  assign new_n8546_ = new_n8544_ & ~new_n8545_;
  assign new_n8547_ = new_n6607_ & ~new_n8546_;
  assign new_n8548_ = ~new_n6618_ & ~new_n8547_;
  assign new_n8549_ = new_n8540_ & new_n8548_;
  assign new_n8550_ = ~new_n8541_ & ~new_n8549_;
  assign new_n8551_ = ~new_n8533_ & new_n8550_;
  assign new_n8552_ = new_n8533_ & ~new_n8550_;
  assign new_n8553_ = ~new_n8551_ & ~new_n8552_;
  assign new_n8554_ = ~new_n8526_ & ~new_n8553_;
  assign new_n8555_ = ~new_n8508_ & ~new_n8554_;
  assign new_n8556_ = ~new_n8509_ & ~new_n8555_;
  assign new_n8557_ = new_n8463_ & new_n8556_;
  assign new_n8558_ = ~new_n8463_ & ~new_n8556_;
  assign new_n8559_ = ~new_n8557_ & ~new_n8558_;
  assign A6445 = ~new_n8418_ & ~new_n8559_;
  assign new_n8561_ = ~new_n8415_ & ~new_n8557_;
  assign A6444 = ~new_n8418_ & ~new_n8561_;
  assign new_n8563_ = new_n8415_ & new_n8463_;
  assign new_n8564_ = ~new_n8418_ & ~new_n8563_;
  assign new_n8565_ = new_n8418_ & ~new_n8564_;
  assign new_n8566_ = new_n8418_ & new_n8563_;
  assign new_n8567_ = new_n8565_ & ~new_n8566_;
  assign new_n8568_ = new_n8463_ & ~new_n8567_;
  assign A6443 = new_n8556_ | new_n8568_;
  assign new_n8570_ = new_n8508_ & new_n8554_;
  assign new_n8571_ = ~new_n8555_ & ~new_n8570_;
  assign new_n8572_ = ~new_n8418_ & ~new_n8508_;
  assign new_n8573_ = new_n8418_ & new_n8508_;
  assign new_n8574_ = ~new_n8572_ & ~new_n8573_;
  assign new_n8575_ = new_n8571_ & ~new_n8574_;
  assign A6442 = new_n8568_ | new_n8575_;
  assign new_n8577_ = new_n8463_ & ~new_n8575_;
  assign new_n8578_ = ~new_n8463_ & new_n8575_;
  assign new_n8579_ = ~new_n8577_ & ~new_n8578_;
  assign A6441 = ~new_n8418_ & ~new_n8579_;
  assign new_n8581_ = new_n1297_ & new_n1308_;
  assign new_n8582_ = ~new_n1309_ & ~new_n8581_;
  assign new_n8583_ = ~new_n1277_ & ~new_n1297_;
  assign new_n8584_ = new_n1277_ & new_n1297_;
  assign new_n8585_ = ~new_n8583_ & ~new_n8584_;
  assign new_n8586_ = new_n8582_ & ~new_n8585_;
  assign new_n8587_ = ~new_n7315_ & ~new_n8586_;
  assign new_n8588_ = new_n1357_ & new_n1368_;
  assign new_n8589_ = ~new_n1369_ & ~new_n8588_;
  assign new_n8590_ = ~new_n1337_ & ~new_n1357_;
  assign new_n8591_ = new_n1337_ & new_n1357_;
  assign new_n8592_ = ~new_n8590_ & ~new_n8591_;
  assign new_n8593_ = new_n8589_ & ~new_n8592_;
  assign new_n8594_ = ~new_n7322_ & ~new_n8593_;
  assign new_n8595_ = new_n8587_ & ~new_n8594_;
  assign new_n8596_ = ~new_n8587_ & new_n8594_;
  assign new_n8597_ = ~new_n8595_ & ~new_n8596_;
  assign new_n8598_ = new_n1420_ & new_n1431_;
  assign new_n8599_ = ~new_n1432_ & ~new_n8598_;
  assign new_n8600_ = ~new_n1400_ & ~new_n1420_;
  assign new_n8601_ = new_n1400_ & new_n1420_;
  assign new_n8602_ = ~new_n8600_ & ~new_n8601_;
  assign new_n8603_ = new_n8599_ & ~new_n8602_;
  assign new_n8604_ = ~new_n7332_ & ~new_n8603_;
  assign new_n8605_ = new_n1480_ & new_n1491_;
  assign new_n8606_ = ~new_n1492_ & ~new_n8605_;
  assign new_n8607_ = ~new_n1460_ & ~new_n1480_;
  assign new_n8608_ = new_n1460_ & new_n1480_;
  assign new_n8609_ = ~new_n8607_ & ~new_n8608_;
  assign new_n8610_ = new_n8606_ & ~new_n8609_;
  assign new_n8611_ = ~new_n7339_ & ~new_n8610_;
  assign new_n8612_ = new_n8597_ & new_n8611_;
  assign new_n8613_ = new_n1541_ & new_n1552_;
  assign new_n8614_ = ~new_n1553_ & ~new_n8613_;
  assign new_n8615_ = ~new_n1521_ & ~new_n1541_;
  assign new_n8616_ = new_n1521_ & new_n1541_;
  assign new_n8617_ = ~new_n8615_ & ~new_n8616_;
  assign new_n8618_ = new_n8614_ & ~new_n8617_;
  assign new_n8619_ = ~new_n7347_ & ~new_n8618_;
  assign new_n8620_ = new_n8611_ & new_n8619_;
  assign new_n8621_ = ~new_n8612_ & ~new_n8620_;
  assign new_n8622_ = ~new_n8604_ & new_n8621_;
  assign new_n8623_ = new_n8604_ & ~new_n8621_;
  assign new_n8624_ = ~new_n8622_ & ~new_n8623_;
  assign new_n8625_ = ~new_n8597_ & ~new_n8624_;
  assign new_n8626_ = new_n1607_ & new_n1618_;
  assign new_n8627_ = ~new_n1619_ & ~new_n8626_;
  assign new_n8628_ = ~new_n1587_ & ~new_n1607_;
  assign new_n8629_ = new_n1587_ & new_n1607_;
  assign new_n8630_ = ~new_n8628_ & ~new_n8629_;
  assign new_n8631_ = new_n8627_ & ~new_n8630_;
  assign new_n8632_ = ~new_n7360_ & ~new_n8631_;
  assign new_n8633_ = new_n1667_ & new_n1678_;
  assign new_n8634_ = ~new_n1679_ & ~new_n8633_;
  assign new_n8635_ = ~new_n1647_ & ~new_n1667_;
  assign new_n8636_ = new_n1647_ & new_n1667_;
  assign new_n8637_ = ~new_n8635_ & ~new_n8636_;
  assign new_n8638_ = new_n8634_ & ~new_n8637_;
  assign new_n8639_ = ~new_n7367_ & ~new_n8638_;
  assign new_n8640_ = new_n8632_ & ~new_n8639_;
  assign new_n8641_ = ~new_n8632_ & new_n8639_;
  assign new_n8642_ = ~new_n8640_ & ~new_n8641_;
  assign new_n8643_ = new_n1730_ & new_n1741_;
  assign new_n8644_ = ~new_n1742_ & ~new_n8643_;
  assign new_n8645_ = ~new_n1710_ & ~new_n1730_;
  assign new_n8646_ = new_n1710_ & new_n1730_;
  assign new_n8647_ = ~new_n8645_ & ~new_n8646_;
  assign new_n8648_ = new_n8644_ & ~new_n8647_;
  assign new_n8649_ = ~new_n7377_ & ~new_n8648_;
  assign new_n8650_ = new_n1790_ & new_n1801_;
  assign new_n8651_ = ~new_n1802_ & ~new_n8650_;
  assign new_n8652_ = ~new_n1770_ & ~new_n1790_;
  assign new_n8653_ = new_n1770_ & new_n1790_;
  assign new_n8654_ = ~new_n8652_ & ~new_n8653_;
  assign new_n8655_ = new_n8651_ & ~new_n8654_;
  assign new_n8656_ = ~new_n7384_ & ~new_n8655_;
  assign new_n8657_ = new_n8642_ & new_n8656_;
  assign new_n8658_ = new_n1851_ & new_n1862_;
  assign new_n8659_ = ~new_n1863_ & ~new_n8658_;
  assign new_n8660_ = ~new_n1831_ & ~new_n1851_;
  assign new_n8661_ = new_n1831_ & new_n1851_;
  assign new_n8662_ = ~new_n8660_ & ~new_n8661_;
  assign new_n8663_ = new_n8659_ & ~new_n8662_;
  assign new_n8664_ = ~new_n7392_ & ~new_n8663_;
  assign new_n8665_ = new_n8656_ & new_n8664_;
  assign new_n8666_ = ~new_n8657_ & ~new_n8665_;
  assign new_n8667_ = ~new_n8649_ & new_n8666_;
  assign new_n8668_ = new_n8649_ & ~new_n8666_;
  assign new_n8669_ = ~new_n8667_ & ~new_n8668_;
  assign new_n8670_ = ~new_n8642_ & ~new_n8669_;
  assign new_n8671_ = ~new_n8625_ & new_n8670_;
  assign new_n8672_ = new_n8625_ & ~new_n8670_;
  assign new_n8673_ = ~new_n8671_ & ~new_n8672_;
  assign new_n8674_ = new_n1920_ & new_n1931_;
  assign new_n8675_ = ~new_n1932_ & ~new_n8674_;
  assign new_n8676_ = ~new_n1900_ & ~new_n1920_;
  assign new_n8677_ = new_n1900_ & new_n1920_;
  assign new_n8678_ = ~new_n8676_ & ~new_n8677_;
  assign new_n8679_ = new_n8675_ & ~new_n8678_;
  assign new_n8680_ = ~new_n7408_ & ~new_n8679_;
  assign new_n8681_ = new_n1980_ & new_n1991_;
  assign new_n8682_ = ~new_n1992_ & ~new_n8681_;
  assign new_n8683_ = ~new_n1960_ & ~new_n1980_;
  assign new_n8684_ = new_n1960_ & new_n1980_;
  assign new_n8685_ = ~new_n8683_ & ~new_n8684_;
  assign new_n8686_ = new_n8682_ & ~new_n8685_;
  assign new_n8687_ = ~new_n7415_ & ~new_n8686_;
  assign new_n8688_ = new_n8680_ & ~new_n8687_;
  assign new_n8689_ = ~new_n8680_ & new_n8687_;
  assign new_n8690_ = ~new_n8688_ & ~new_n8689_;
  assign new_n8691_ = new_n2043_ & new_n2054_;
  assign new_n8692_ = ~new_n2055_ & ~new_n8691_;
  assign new_n8693_ = ~new_n2023_ & ~new_n2043_;
  assign new_n8694_ = new_n2023_ & new_n2043_;
  assign new_n8695_ = ~new_n8693_ & ~new_n8694_;
  assign new_n8696_ = new_n8692_ & ~new_n8695_;
  assign new_n8697_ = ~new_n7425_ & ~new_n8696_;
  assign new_n8698_ = new_n2103_ & new_n2114_;
  assign new_n8699_ = ~new_n2115_ & ~new_n8698_;
  assign new_n8700_ = ~new_n2083_ & ~new_n2103_;
  assign new_n8701_ = new_n2083_ & new_n2103_;
  assign new_n8702_ = ~new_n8700_ & ~new_n8701_;
  assign new_n8703_ = new_n8699_ & ~new_n8702_;
  assign new_n8704_ = ~new_n7432_ & ~new_n8703_;
  assign new_n8705_ = new_n8690_ & new_n8704_;
  assign new_n8706_ = new_n2164_ & new_n2175_;
  assign new_n8707_ = ~new_n2176_ & ~new_n8706_;
  assign new_n8708_ = ~new_n2144_ & ~new_n2164_;
  assign new_n8709_ = new_n2144_ & new_n2164_;
  assign new_n8710_ = ~new_n8708_ & ~new_n8709_;
  assign new_n8711_ = new_n8707_ & ~new_n8710_;
  assign new_n8712_ = ~new_n7440_ & ~new_n8711_;
  assign new_n8713_ = new_n8704_ & new_n8712_;
  assign new_n8714_ = ~new_n8705_ & ~new_n8713_;
  assign new_n8715_ = ~new_n8697_ & new_n8714_;
  assign new_n8716_ = new_n8697_ & ~new_n8714_;
  assign new_n8717_ = ~new_n8715_ & ~new_n8716_;
  assign new_n8718_ = ~new_n8690_ & ~new_n8717_;
  assign new_n8719_ = new_n2230_ & new_n2241_;
  assign new_n8720_ = ~new_n2242_ & ~new_n8719_;
  assign new_n8721_ = ~new_n2210_ & ~new_n2230_;
  assign new_n8722_ = new_n2210_ & new_n2230_;
  assign new_n8723_ = ~new_n8721_ & ~new_n8722_;
  assign new_n8724_ = new_n8720_ & ~new_n8723_;
  assign new_n8725_ = ~new_n7453_ & ~new_n8724_;
  assign new_n8726_ = new_n2290_ & new_n2301_;
  assign new_n8727_ = ~new_n2302_ & ~new_n8726_;
  assign new_n8728_ = ~new_n2270_ & ~new_n2290_;
  assign new_n8729_ = new_n2270_ & new_n2290_;
  assign new_n8730_ = ~new_n8728_ & ~new_n8729_;
  assign new_n8731_ = new_n8727_ & ~new_n8730_;
  assign new_n8732_ = ~new_n7460_ & ~new_n8731_;
  assign new_n8733_ = new_n8725_ & ~new_n8732_;
  assign new_n8734_ = ~new_n8725_ & new_n8732_;
  assign new_n8735_ = ~new_n8733_ & ~new_n8734_;
  assign new_n8736_ = new_n2353_ & new_n2364_;
  assign new_n8737_ = ~new_n2365_ & ~new_n8736_;
  assign new_n8738_ = ~new_n2333_ & ~new_n2353_;
  assign new_n8739_ = new_n2333_ & new_n2353_;
  assign new_n8740_ = ~new_n8738_ & ~new_n8739_;
  assign new_n8741_ = new_n8737_ & ~new_n8740_;
  assign new_n8742_ = ~new_n7470_ & ~new_n8741_;
  assign new_n8743_ = new_n2413_ & new_n2424_;
  assign new_n8744_ = ~new_n2425_ & ~new_n8743_;
  assign new_n8745_ = ~new_n2393_ & ~new_n2413_;
  assign new_n8746_ = new_n2393_ & new_n2413_;
  assign new_n8747_ = ~new_n8745_ & ~new_n8746_;
  assign new_n8748_ = new_n8744_ & ~new_n8747_;
  assign new_n8749_ = ~new_n7477_ & ~new_n8748_;
  assign new_n8750_ = new_n8735_ & new_n8749_;
  assign new_n8751_ = new_n2474_ & new_n2485_;
  assign new_n8752_ = ~new_n2486_ & ~new_n8751_;
  assign new_n8753_ = ~new_n2454_ & ~new_n2474_;
  assign new_n8754_ = new_n2454_ & new_n2474_;
  assign new_n8755_ = ~new_n8753_ & ~new_n8754_;
  assign new_n8756_ = new_n8752_ & ~new_n8755_;
  assign new_n8757_ = ~new_n7485_ & ~new_n8756_;
  assign new_n8758_ = new_n8749_ & new_n8757_;
  assign new_n8759_ = ~new_n8750_ & ~new_n8758_;
  assign new_n8760_ = ~new_n8742_ & new_n8759_;
  assign new_n8761_ = new_n8742_ & ~new_n8759_;
  assign new_n8762_ = ~new_n8760_ & ~new_n8761_;
  assign new_n8763_ = ~new_n8735_ & ~new_n8762_;
  assign new_n8764_ = new_n8673_ & ~new_n8763_;
  assign new_n8765_ = new_n2541_ & new_n2552_;
  assign new_n8766_ = ~new_n2553_ & ~new_n8765_;
  assign new_n8767_ = ~new_n2521_ & ~new_n2541_;
  assign new_n8768_ = new_n2521_ & new_n2541_;
  assign new_n8769_ = ~new_n8767_ & ~new_n8768_;
  assign new_n8770_ = new_n8766_ & ~new_n8769_;
  assign new_n8771_ = ~new_n7499_ & ~new_n8770_;
  assign new_n8772_ = new_n2601_ & new_n2612_;
  assign new_n8773_ = ~new_n2613_ & ~new_n8772_;
  assign new_n8774_ = ~new_n2581_ & ~new_n2601_;
  assign new_n8775_ = new_n2581_ & new_n2601_;
  assign new_n8776_ = ~new_n8774_ & ~new_n8775_;
  assign new_n8777_ = new_n8773_ & ~new_n8776_;
  assign new_n8778_ = ~new_n7506_ & ~new_n8777_;
  assign new_n8779_ = new_n8771_ & ~new_n8778_;
  assign new_n8780_ = ~new_n8771_ & new_n8778_;
  assign new_n8781_ = ~new_n8779_ & ~new_n8780_;
  assign new_n8782_ = new_n2664_ & new_n2675_;
  assign new_n8783_ = ~new_n2676_ & ~new_n8782_;
  assign new_n8784_ = ~new_n2644_ & ~new_n2664_;
  assign new_n8785_ = new_n2644_ & new_n2664_;
  assign new_n8786_ = ~new_n8784_ & ~new_n8785_;
  assign new_n8787_ = new_n8783_ & ~new_n8786_;
  assign new_n8788_ = ~new_n7516_ & ~new_n8787_;
  assign new_n8789_ = new_n2724_ & new_n2735_;
  assign new_n8790_ = ~new_n2736_ & ~new_n8789_;
  assign new_n8791_ = ~new_n2704_ & ~new_n2724_;
  assign new_n8792_ = new_n2704_ & new_n2724_;
  assign new_n8793_ = ~new_n8791_ & ~new_n8792_;
  assign new_n8794_ = new_n8790_ & ~new_n8793_;
  assign new_n8795_ = ~new_n7523_ & ~new_n8794_;
  assign new_n8796_ = new_n8781_ & new_n8795_;
  assign new_n8797_ = new_n2785_ & new_n2796_;
  assign new_n8798_ = ~new_n2797_ & ~new_n8797_;
  assign new_n8799_ = ~new_n2765_ & ~new_n2785_;
  assign new_n8800_ = new_n2765_ & new_n2785_;
  assign new_n8801_ = ~new_n8799_ & ~new_n8800_;
  assign new_n8802_ = new_n8798_ & ~new_n8801_;
  assign new_n8803_ = ~new_n7531_ & ~new_n8802_;
  assign new_n8804_ = new_n8795_ & new_n8803_;
  assign new_n8805_ = ~new_n8796_ & ~new_n8804_;
  assign new_n8806_ = ~new_n8788_ & new_n8805_;
  assign new_n8807_ = new_n8788_ & ~new_n8805_;
  assign new_n8808_ = ~new_n8806_ & ~new_n8807_;
  assign new_n8809_ = ~new_n8781_ & ~new_n8808_;
  assign new_n8810_ = ~new_n8763_ & ~new_n8809_;
  assign new_n8811_ = ~new_n8764_ & ~new_n8810_;
  assign new_n8812_ = new_n8718_ & new_n8811_;
  assign new_n8813_ = ~new_n8718_ & ~new_n8811_;
  assign new_n8814_ = ~new_n8812_ & ~new_n8813_;
  assign A6412 = ~new_n8673_ & ~new_n8814_;
  assign new_n8816_ = ~new_n8670_ & ~new_n8812_;
  assign A6411 = ~new_n8673_ & ~new_n8816_;
  assign new_n8818_ = new_n8670_ & new_n8718_;
  assign new_n8819_ = ~new_n8673_ & ~new_n8818_;
  assign new_n8820_ = new_n8673_ & ~new_n8819_;
  assign new_n8821_ = new_n8673_ & new_n8818_;
  assign new_n8822_ = new_n8820_ & ~new_n8821_;
  assign new_n8823_ = new_n8718_ & ~new_n8822_;
  assign A6410 = new_n8811_ | new_n8823_;
  assign new_n8825_ = new_n8763_ & new_n8809_;
  assign new_n8826_ = ~new_n8810_ & ~new_n8825_;
  assign new_n8827_ = ~new_n8673_ & ~new_n8763_;
  assign new_n8828_ = new_n8673_ & new_n8763_;
  assign new_n8829_ = ~new_n8827_ & ~new_n8828_;
  assign new_n8830_ = new_n8826_ & ~new_n8829_;
  assign A6409 = new_n8823_ | new_n8830_;
  assign new_n8832_ = new_n8718_ & ~new_n8830_;
  assign new_n8833_ = ~new_n8718_ & new_n8830_;
  assign new_n8834_ = ~new_n8832_ & ~new_n8833_;
  assign A6408 = ~new_n8673_ & ~new_n8834_;
  assign new_n8836_ = new_n2850_ & new_n2853_;
  assign new_n8837_ = ~new_n2854_ & ~new_n8836_;
  assign new_n8838_ = ~new_n2846_ & ~new_n2850_;
  assign new_n8839_ = new_n2846_ & new_n2850_;
  assign new_n8840_ = ~new_n8838_ & ~new_n8839_;
  assign new_n8841_ = new_n8837_ & ~new_n8840_;
  assign new_n8842_ = ~new_n7570_ & ~new_n8841_;
  assign new_n8843_ = new_n2870_ & new_n2873_;
  assign new_n8844_ = ~new_n2874_ & ~new_n8843_;
  assign new_n8845_ = ~new_n2866_ & ~new_n2870_;
  assign new_n8846_ = new_n2866_ & new_n2870_;
  assign new_n8847_ = ~new_n8845_ & ~new_n8846_;
  assign new_n8848_ = new_n8844_ & ~new_n8847_;
  assign new_n8849_ = ~new_n7577_ & ~new_n8848_;
  assign new_n8850_ = new_n8842_ & ~new_n8849_;
  assign new_n8851_ = ~new_n8842_ & new_n8849_;
  assign new_n8852_ = ~new_n8850_ & ~new_n8851_;
  assign new_n8853_ = new_n2893_ & new_n2896_;
  assign new_n8854_ = ~new_n2897_ & ~new_n8853_;
  assign new_n8855_ = ~new_n2889_ & ~new_n2893_;
  assign new_n8856_ = new_n2889_ & new_n2893_;
  assign new_n8857_ = ~new_n8855_ & ~new_n8856_;
  assign new_n8858_ = new_n8854_ & ~new_n8857_;
  assign new_n8859_ = ~new_n7587_ & ~new_n8858_;
  assign new_n8860_ = new_n2913_ & new_n2916_;
  assign new_n8861_ = ~new_n2917_ & ~new_n8860_;
  assign new_n8862_ = ~new_n2909_ & ~new_n2913_;
  assign new_n8863_ = new_n2909_ & new_n2913_;
  assign new_n8864_ = ~new_n8862_ & ~new_n8863_;
  assign new_n8865_ = new_n8861_ & ~new_n8864_;
  assign new_n8866_ = ~new_n7594_ & ~new_n8865_;
  assign new_n8867_ = new_n8852_ & new_n8866_;
  assign new_n8868_ = new_n2934_ & new_n2937_;
  assign new_n8869_ = ~new_n2938_ & ~new_n8868_;
  assign new_n8870_ = ~new_n2930_ & ~new_n2934_;
  assign new_n8871_ = new_n2930_ & new_n2934_;
  assign new_n8872_ = ~new_n8870_ & ~new_n8871_;
  assign new_n8873_ = new_n8869_ & ~new_n8872_;
  assign new_n8874_ = ~new_n7602_ & ~new_n8873_;
  assign new_n8875_ = new_n8866_ & new_n8874_;
  assign new_n8876_ = ~new_n8867_ & ~new_n8875_;
  assign new_n8877_ = ~new_n8859_ & new_n8876_;
  assign new_n8878_ = new_n8859_ & ~new_n8876_;
  assign new_n8879_ = ~new_n8877_ & ~new_n8878_;
  assign new_n8880_ = ~new_n8852_ & ~new_n8879_;
  assign new_n8881_ = new_n2960_ & new_n2963_;
  assign new_n8882_ = ~new_n2964_ & ~new_n8881_;
  assign new_n8883_ = ~new_n2956_ & ~new_n2960_;
  assign new_n8884_ = new_n2956_ & new_n2960_;
  assign new_n8885_ = ~new_n8883_ & ~new_n8884_;
  assign new_n8886_ = new_n8882_ & ~new_n8885_;
  assign new_n8887_ = ~new_n7615_ & ~new_n8886_;
  assign new_n8888_ = new_n2980_ & new_n2983_;
  assign new_n8889_ = ~new_n2984_ & ~new_n8888_;
  assign new_n8890_ = ~new_n2976_ & ~new_n2980_;
  assign new_n8891_ = new_n2976_ & new_n2980_;
  assign new_n8892_ = ~new_n8890_ & ~new_n8891_;
  assign new_n8893_ = new_n8889_ & ~new_n8892_;
  assign new_n8894_ = ~new_n7622_ & ~new_n8893_;
  assign new_n8895_ = new_n8887_ & ~new_n8894_;
  assign new_n8896_ = ~new_n8887_ & new_n8894_;
  assign new_n8897_ = ~new_n8895_ & ~new_n8896_;
  assign new_n8898_ = new_n3003_ & new_n3006_;
  assign new_n8899_ = ~new_n3007_ & ~new_n8898_;
  assign new_n8900_ = ~new_n2999_ & ~new_n3003_;
  assign new_n8901_ = new_n2999_ & new_n3003_;
  assign new_n8902_ = ~new_n8900_ & ~new_n8901_;
  assign new_n8903_ = new_n8899_ & ~new_n8902_;
  assign new_n8904_ = ~new_n7632_ & ~new_n8903_;
  assign new_n8905_ = new_n3023_ & new_n3026_;
  assign new_n8906_ = ~new_n3027_ & ~new_n8905_;
  assign new_n8907_ = ~new_n3019_ & ~new_n3023_;
  assign new_n8908_ = new_n3019_ & new_n3023_;
  assign new_n8909_ = ~new_n8907_ & ~new_n8908_;
  assign new_n8910_ = new_n8906_ & ~new_n8909_;
  assign new_n8911_ = ~new_n7639_ & ~new_n8910_;
  assign new_n8912_ = new_n8897_ & new_n8911_;
  assign new_n8913_ = new_n3044_ & new_n3047_;
  assign new_n8914_ = ~new_n3048_ & ~new_n8913_;
  assign new_n8915_ = ~new_n3040_ & ~new_n3044_;
  assign new_n8916_ = new_n3040_ & new_n3044_;
  assign new_n8917_ = ~new_n8915_ & ~new_n8916_;
  assign new_n8918_ = new_n8914_ & ~new_n8917_;
  assign new_n8919_ = ~new_n7647_ & ~new_n8918_;
  assign new_n8920_ = new_n8911_ & new_n8919_;
  assign new_n8921_ = ~new_n8912_ & ~new_n8920_;
  assign new_n8922_ = ~new_n8904_ & new_n8921_;
  assign new_n8923_ = new_n8904_ & ~new_n8921_;
  assign new_n8924_ = ~new_n8922_ & ~new_n8923_;
  assign new_n8925_ = ~new_n8897_ & ~new_n8924_;
  assign new_n8926_ = ~new_n8880_ & new_n8925_;
  assign new_n8927_ = new_n8880_ & ~new_n8925_;
  assign new_n8928_ = ~new_n8926_ & ~new_n8927_;
  assign new_n8929_ = new_n3073_ & new_n3076_;
  assign new_n8930_ = ~new_n3077_ & ~new_n8929_;
  assign new_n8931_ = ~new_n3069_ & ~new_n3073_;
  assign new_n8932_ = new_n3069_ & new_n3073_;
  assign new_n8933_ = ~new_n8931_ & ~new_n8932_;
  assign new_n8934_ = new_n8930_ & ~new_n8933_;
  assign new_n8935_ = ~new_n7663_ & ~new_n8934_;
  assign new_n8936_ = new_n3093_ & new_n3096_;
  assign new_n8937_ = ~new_n3097_ & ~new_n8936_;
  assign new_n8938_ = ~new_n3089_ & ~new_n3093_;
  assign new_n8939_ = new_n3089_ & new_n3093_;
  assign new_n8940_ = ~new_n8938_ & ~new_n8939_;
  assign new_n8941_ = new_n8937_ & ~new_n8940_;
  assign new_n8942_ = ~new_n7670_ & ~new_n8941_;
  assign new_n8943_ = new_n8935_ & ~new_n8942_;
  assign new_n8944_ = ~new_n8935_ & new_n8942_;
  assign new_n8945_ = ~new_n8943_ & ~new_n8944_;
  assign new_n8946_ = new_n3116_ & new_n3119_;
  assign new_n8947_ = ~new_n3120_ & ~new_n8946_;
  assign new_n8948_ = ~new_n3112_ & ~new_n3116_;
  assign new_n8949_ = new_n3112_ & new_n3116_;
  assign new_n8950_ = ~new_n8948_ & ~new_n8949_;
  assign new_n8951_ = new_n8947_ & ~new_n8950_;
  assign new_n8952_ = ~new_n7680_ & ~new_n8951_;
  assign new_n8953_ = new_n3136_ & new_n3139_;
  assign new_n8954_ = ~new_n3140_ & ~new_n8953_;
  assign new_n8955_ = ~new_n3132_ & ~new_n3136_;
  assign new_n8956_ = new_n3132_ & new_n3136_;
  assign new_n8957_ = ~new_n8955_ & ~new_n8956_;
  assign new_n8958_ = new_n8954_ & ~new_n8957_;
  assign new_n8959_ = ~new_n7687_ & ~new_n8958_;
  assign new_n8960_ = new_n8945_ & new_n8959_;
  assign new_n8961_ = new_n3157_ & new_n3160_;
  assign new_n8962_ = ~new_n3161_ & ~new_n8961_;
  assign new_n8963_ = ~new_n3153_ & ~new_n3157_;
  assign new_n8964_ = new_n3153_ & new_n3157_;
  assign new_n8965_ = ~new_n8963_ & ~new_n8964_;
  assign new_n8966_ = new_n8962_ & ~new_n8965_;
  assign new_n8967_ = ~new_n7695_ & ~new_n8966_;
  assign new_n8968_ = new_n8959_ & new_n8967_;
  assign new_n8969_ = ~new_n8960_ & ~new_n8968_;
  assign new_n8970_ = ~new_n8952_ & new_n8969_;
  assign new_n8971_ = new_n8952_ & ~new_n8969_;
  assign new_n8972_ = ~new_n8970_ & ~new_n8971_;
  assign new_n8973_ = ~new_n8945_ & ~new_n8972_;
  assign new_n8974_ = new_n3183_ & new_n3186_;
  assign new_n8975_ = ~new_n3187_ & ~new_n8974_;
  assign new_n8976_ = ~new_n3179_ & ~new_n3183_;
  assign new_n8977_ = new_n3179_ & new_n3183_;
  assign new_n8978_ = ~new_n8976_ & ~new_n8977_;
  assign new_n8979_ = new_n8975_ & ~new_n8978_;
  assign new_n8980_ = ~new_n7708_ & ~new_n8979_;
  assign new_n8981_ = new_n3203_ & new_n3206_;
  assign new_n8982_ = ~new_n3207_ & ~new_n8981_;
  assign new_n8983_ = ~new_n3199_ & ~new_n3203_;
  assign new_n8984_ = new_n3199_ & new_n3203_;
  assign new_n8985_ = ~new_n8983_ & ~new_n8984_;
  assign new_n8986_ = new_n8982_ & ~new_n8985_;
  assign new_n8987_ = ~new_n7715_ & ~new_n8986_;
  assign new_n8988_ = new_n8980_ & ~new_n8987_;
  assign new_n8989_ = ~new_n8980_ & new_n8987_;
  assign new_n8990_ = ~new_n8988_ & ~new_n8989_;
  assign new_n8991_ = new_n3226_ & new_n3229_;
  assign new_n8992_ = ~new_n3230_ & ~new_n8991_;
  assign new_n8993_ = ~new_n3222_ & ~new_n3226_;
  assign new_n8994_ = new_n3222_ & new_n3226_;
  assign new_n8995_ = ~new_n8993_ & ~new_n8994_;
  assign new_n8996_ = new_n8992_ & ~new_n8995_;
  assign new_n8997_ = ~new_n7725_ & ~new_n8996_;
  assign new_n8998_ = new_n3246_ & new_n3249_;
  assign new_n8999_ = ~new_n3250_ & ~new_n8998_;
  assign new_n9000_ = ~new_n3242_ & ~new_n3246_;
  assign new_n9001_ = new_n3242_ & new_n3246_;
  assign new_n9002_ = ~new_n9000_ & ~new_n9001_;
  assign new_n9003_ = new_n8999_ & ~new_n9002_;
  assign new_n9004_ = ~new_n7732_ & ~new_n9003_;
  assign new_n9005_ = new_n8990_ & new_n9004_;
  assign new_n9006_ = new_n3267_ & new_n3270_;
  assign new_n9007_ = ~new_n3271_ & ~new_n9006_;
  assign new_n9008_ = ~new_n3263_ & ~new_n3267_;
  assign new_n9009_ = new_n3263_ & new_n3267_;
  assign new_n9010_ = ~new_n9008_ & ~new_n9009_;
  assign new_n9011_ = new_n9007_ & ~new_n9010_;
  assign new_n9012_ = ~new_n7740_ & ~new_n9011_;
  assign new_n9013_ = new_n9004_ & new_n9012_;
  assign new_n9014_ = ~new_n9005_ & ~new_n9013_;
  assign new_n9015_ = ~new_n8997_ & new_n9014_;
  assign new_n9016_ = new_n8997_ & ~new_n9014_;
  assign new_n9017_ = ~new_n9015_ & ~new_n9016_;
  assign new_n9018_ = ~new_n8990_ & ~new_n9017_;
  assign new_n9019_ = new_n8928_ & ~new_n9018_;
  assign new_n9020_ = new_n3294_ & new_n3297_;
  assign new_n9021_ = ~new_n3298_ & ~new_n9020_;
  assign new_n9022_ = ~new_n3290_ & ~new_n3294_;
  assign new_n9023_ = new_n3290_ & new_n3294_;
  assign new_n9024_ = ~new_n9022_ & ~new_n9023_;
  assign new_n9025_ = new_n9021_ & ~new_n9024_;
  assign new_n9026_ = ~new_n7754_ & ~new_n9025_;
  assign new_n9027_ = new_n3314_ & new_n3317_;
  assign new_n9028_ = ~new_n3318_ & ~new_n9027_;
  assign new_n9029_ = ~new_n3310_ & ~new_n3314_;
  assign new_n9030_ = new_n3310_ & new_n3314_;
  assign new_n9031_ = ~new_n9029_ & ~new_n9030_;
  assign new_n9032_ = new_n9028_ & ~new_n9031_;
  assign new_n9033_ = ~new_n7761_ & ~new_n9032_;
  assign new_n9034_ = new_n9026_ & ~new_n9033_;
  assign new_n9035_ = ~new_n9026_ & new_n9033_;
  assign new_n9036_ = ~new_n9034_ & ~new_n9035_;
  assign new_n9037_ = new_n3337_ & new_n3340_;
  assign new_n9038_ = ~new_n3341_ & ~new_n9037_;
  assign new_n9039_ = ~new_n3333_ & ~new_n3337_;
  assign new_n9040_ = new_n3333_ & new_n3337_;
  assign new_n9041_ = ~new_n9039_ & ~new_n9040_;
  assign new_n9042_ = new_n9038_ & ~new_n9041_;
  assign new_n9043_ = ~new_n7771_ & ~new_n9042_;
  assign new_n9044_ = new_n3357_ & new_n3360_;
  assign new_n9045_ = ~new_n3361_ & ~new_n9044_;
  assign new_n9046_ = ~new_n3353_ & ~new_n3357_;
  assign new_n9047_ = new_n3353_ & new_n3357_;
  assign new_n9048_ = ~new_n9046_ & ~new_n9047_;
  assign new_n9049_ = new_n9045_ & ~new_n9048_;
  assign new_n9050_ = ~new_n7778_ & ~new_n9049_;
  assign new_n9051_ = new_n9036_ & new_n9050_;
  assign new_n9052_ = new_n3378_ & new_n3381_;
  assign new_n9053_ = ~new_n3382_ & ~new_n9052_;
  assign new_n9054_ = ~new_n3374_ & ~new_n3378_;
  assign new_n9055_ = new_n3374_ & new_n3378_;
  assign new_n9056_ = ~new_n9054_ & ~new_n9055_;
  assign new_n9057_ = new_n9053_ & ~new_n9056_;
  assign new_n9058_ = ~new_n7786_ & ~new_n9057_;
  assign new_n9059_ = new_n9050_ & new_n9058_;
  assign new_n9060_ = ~new_n9051_ & ~new_n9059_;
  assign new_n9061_ = ~new_n9043_ & new_n9060_;
  assign new_n9062_ = new_n9043_ & ~new_n9060_;
  assign new_n9063_ = ~new_n9061_ & ~new_n9062_;
  assign new_n9064_ = ~new_n9036_ & ~new_n9063_;
  assign new_n9065_ = ~new_n9018_ & ~new_n9064_;
  assign new_n9066_ = ~new_n9019_ & ~new_n9065_;
  assign new_n9067_ = new_n8973_ & new_n9066_;
  assign new_n9068_ = ~new_n8973_ & ~new_n9066_;
  assign new_n9069_ = ~new_n9067_ & ~new_n9068_;
  assign A6379 = ~new_n8928_ & ~new_n9069_;
  assign new_n9071_ = ~new_n8925_ & ~new_n9067_;
  assign A6378 = ~new_n8928_ & ~new_n9071_;
  assign new_n9073_ = new_n8925_ & new_n8973_;
  assign new_n9074_ = ~new_n8928_ & ~new_n9073_;
  assign new_n9075_ = new_n8928_ & ~new_n9074_;
  assign new_n9076_ = new_n8928_ & new_n9073_;
  assign new_n9077_ = new_n9075_ & ~new_n9076_;
  assign new_n9078_ = new_n8973_ & ~new_n9077_;
  assign A6377 = new_n9066_ | new_n9078_;
  assign new_n9080_ = new_n9018_ & new_n9064_;
  assign new_n9081_ = ~new_n9065_ & ~new_n9080_;
  assign new_n9082_ = ~new_n8928_ & ~new_n9018_;
  assign new_n9083_ = new_n8928_ & new_n9018_;
  assign new_n9084_ = ~new_n9082_ & ~new_n9083_;
  assign new_n9085_ = new_n9081_ & ~new_n9084_;
  assign A6376 = new_n9078_ | new_n9085_;
  assign new_n9087_ = new_n8973_ & ~new_n9085_;
  assign new_n9088_ = ~new_n8973_ & new_n9085_;
  assign new_n9089_ = ~new_n9087_ & ~new_n9088_;
  assign A6375 = ~new_n8928_ & ~new_n9089_;
  assign new_n9091_ = ~new_n3446_ & ~new_n3454_;
  assign new_n9092_ = ~new_n3455_ & ~new_n9091_;
  assign new_n9093_ = ~new_n3432_ & new_n3446_;
  assign new_n9094_ = new_n3432_ & ~new_n3446_;
  assign new_n9095_ = ~new_n9093_ & ~new_n9094_;
  assign new_n9096_ = new_n9092_ & ~new_n9095_;
  assign new_n9097_ = ~new_n7825_ & ~new_n9096_;
  assign new_n9098_ = ~new_n3491_ & ~new_n3499_;
  assign new_n9099_ = ~new_n3500_ & ~new_n9098_;
  assign new_n9100_ = ~new_n3477_ & new_n3491_;
  assign new_n9101_ = new_n3477_ & ~new_n3491_;
  assign new_n9102_ = ~new_n9100_ & ~new_n9101_;
  assign new_n9103_ = new_n9099_ & ~new_n9102_;
  assign new_n9104_ = ~new_n7832_ & ~new_n9103_;
  assign new_n9105_ = new_n9097_ & ~new_n9104_;
  assign new_n9106_ = ~new_n9097_ & new_n9104_;
  assign new_n9107_ = ~new_n9105_ & ~new_n9106_;
  assign new_n9108_ = ~new_n3539_ & ~new_n3547_;
  assign new_n9109_ = ~new_n3548_ & ~new_n9108_;
  assign new_n9110_ = ~new_n3525_ & new_n3539_;
  assign new_n9111_ = new_n3525_ & ~new_n3539_;
  assign new_n9112_ = ~new_n9110_ & ~new_n9111_;
  assign new_n9113_ = new_n9109_ & ~new_n9112_;
  assign new_n9114_ = ~new_n7842_ & ~new_n9113_;
  assign new_n9115_ = ~new_n3584_ & ~new_n3592_;
  assign new_n9116_ = ~new_n3593_ & ~new_n9115_;
  assign new_n9117_ = ~new_n3570_ & new_n3584_;
  assign new_n9118_ = new_n3570_ & ~new_n3584_;
  assign new_n9119_ = ~new_n9117_ & ~new_n9118_;
  assign new_n9120_ = new_n9116_ & ~new_n9119_;
  assign new_n9121_ = ~new_n7849_ & ~new_n9120_;
  assign new_n9122_ = new_n9107_ & new_n9121_;
  assign new_n9123_ = ~new_n3630_ & ~new_n3638_;
  assign new_n9124_ = ~new_n3639_ & ~new_n9123_;
  assign new_n9125_ = ~new_n3616_ & new_n3630_;
  assign new_n9126_ = new_n3616_ & ~new_n3630_;
  assign new_n9127_ = ~new_n9125_ & ~new_n9126_;
  assign new_n9128_ = new_n9124_ & ~new_n9127_;
  assign new_n9129_ = ~new_n7857_ & ~new_n9128_;
  assign new_n9130_ = new_n9121_ & new_n9129_;
  assign new_n9131_ = ~new_n9122_ & ~new_n9130_;
  assign new_n9132_ = ~new_n9114_ & new_n9131_;
  assign new_n9133_ = new_n9114_ & ~new_n9131_;
  assign new_n9134_ = ~new_n9132_ & ~new_n9133_;
  assign new_n9135_ = ~new_n9107_ & ~new_n9134_;
  assign new_n9136_ = ~new_n3681_ & ~new_n3689_;
  assign new_n9137_ = ~new_n3690_ & ~new_n9136_;
  assign new_n9138_ = ~new_n3667_ & new_n3681_;
  assign new_n9139_ = new_n3667_ & ~new_n3681_;
  assign new_n9140_ = ~new_n9138_ & ~new_n9139_;
  assign new_n9141_ = new_n9137_ & ~new_n9140_;
  assign new_n9142_ = ~new_n7870_ & ~new_n9141_;
  assign new_n9143_ = ~new_n3726_ & ~new_n3734_;
  assign new_n9144_ = ~new_n3735_ & ~new_n9143_;
  assign new_n9145_ = ~new_n3712_ & new_n3726_;
  assign new_n9146_ = new_n3712_ & ~new_n3726_;
  assign new_n9147_ = ~new_n9145_ & ~new_n9146_;
  assign new_n9148_ = new_n9144_ & ~new_n9147_;
  assign new_n9149_ = ~new_n7877_ & ~new_n9148_;
  assign new_n9150_ = new_n9142_ & ~new_n9149_;
  assign new_n9151_ = ~new_n9142_ & new_n9149_;
  assign new_n9152_ = ~new_n9150_ & ~new_n9151_;
  assign new_n9153_ = ~new_n3774_ & ~new_n3782_;
  assign new_n9154_ = ~new_n3783_ & ~new_n9153_;
  assign new_n9155_ = ~new_n3760_ & new_n3774_;
  assign new_n9156_ = new_n3760_ & ~new_n3774_;
  assign new_n9157_ = ~new_n9155_ & ~new_n9156_;
  assign new_n9158_ = new_n9154_ & ~new_n9157_;
  assign new_n9159_ = ~new_n7887_ & ~new_n9158_;
  assign new_n9160_ = ~new_n3819_ & ~new_n3827_;
  assign new_n9161_ = ~new_n3828_ & ~new_n9160_;
  assign new_n9162_ = ~new_n3805_ & new_n3819_;
  assign new_n9163_ = new_n3805_ & ~new_n3819_;
  assign new_n9164_ = ~new_n9162_ & ~new_n9163_;
  assign new_n9165_ = new_n9161_ & ~new_n9164_;
  assign new_n9166_ = ~new_n7894_ & ~new_n9165_;
  assign new_n9167_ = new_n9152_ & new_n9166_;
  assign new_n9168_ = ~new_n3865_ & ~new_n3873_;
  assign new_n9169_ = ~new_n3874_ & ~new_n9168_;
  assign new_n9170_ = ~new_n3851_ & new_n3865_;
  assign new_n9171_ = new_n3851_ & ~new_n3865_;
  assign new_n9172_ = ~new_n9170_ & ~new_n9171_;
  assign new_n9173_ = new_n9169_ & ~new_n9172_;
  assign new_n9174_ = ~new_n7902_ & ~new_n9173_;
  assign new_n9175_ = new_n9166_ & new_n9174_;
  assign new_n9176_ = ~new_n9167_ & ~new_n9175_;
  assign new_n9177_ = ~new_n9159_ & new_n9176_;
  assign new_n9178_ = new_n9159_ & ~new_n9176_;
  assign new_n9179_ = ~new_n9177_ & ~new_n9178_;
  assign new_n9180_ = ~new_n9152_ & ~new_n9179_;
  assign new_n9181_ = ~new_n9135_ & new_n9180_;
  assign new_n9182_ = new_n9135_ & ~new_n9180_;
  assign new_n9183_ = ~new_n9181_ & ~new_n9182_;
  assign new_n9184_ = ~new_n3919_ & ~new_n3927_;
  assign new_n9185_ = ~new_n3928_ & ~new_n9184_;
  assign new_n9186_ = ~new_n3905_ & new_n3919_;
  assign new_n9187_ = new_n3905_ & ~new_n3919_;
  assign new_n9188_ = ~new_n9186_ & ~new_n9187_;
  assign new_n9189_ = new_n9185_ & ~new_n9188_;
  assign new_n9190_ = ~new_n7918_ & ~new_n9189_;
  assign new_n9191_ = ~new_n3964_ & ~new_n3972_;
  assign new_n9192_ = ~new_n3973_ & ~new_n9191_;
  assign new_n9193_ = ~new_n3950_ & new_n3964_;
  assign new_n9194_ = new_n3950_ & ~new_n3964_;
  assign new_n9195_ = ~new_n9193_ & ~new_n9194_;
  assign new_n9196_ = new_n9192_ & ~new_n9195_;
  assign new_n9197_ = ~new_n7925_ & ~new_n9196_;
  assign new_n9198_ = new_n9190_ & ~new_n9197_;
  assign new_n9199_ = ~new_n9190_ & new_n9197_;
  assign new_n9200_ = ~new_n9198_ & ~new_n9199_;
  assign new_n9201_ = ~new_n4012_ & ~new_n4020_;
  assign new_n9202_ = ~new_n4021_ & ~new_n9201_;
  assign new_n9203_ = ~new_n3998_ & new_n4012_;
  assign new_n9204_ = new_n3998_ & ~new_n4012_;
  assign new_n9205_ = ~new_n9203_ & ~new_n9204_;
  assign new_n9206_ = new_n9202_ & ~new_n9205_;
  assign new_n9207_ = ~new_n7935_ & ~new_n9206_;
  assign new_n9208_ = ~new_n4057_ & ~new_n4065_;
  assign new_n9209_ = ~new_n4066_ & ~new_n9208_;
  assign new_n9210_ = ~new_n4043_ & new_n4057_;
  assign new_n9211_ = new_n4043_ & ~new_n4057_;
  assign new_n9212_ = ~new_n9210_ & ~new_n9211_;
  assign new_n9213_ = new_n9209_ & ~new_n9212_;
  assign new_n9214_ = ~new_n7942_ & ~new_n9213_;
  assign new_n9215_ = new_n9200_ & new_n9214_;
  assign new_n9216_ = ~new_n4103_ & ~new_n4111_;
  assign new_n9217_ = ~new_n4112_ & ~new_n9216_;
  assign new_n9218_ = ~new_n4089_ & new_n4103_;
  assign new_n9219_ = new_n4089_ & ~new_n4103_;
  assign new_n9220_ = ~new_n9218_ & ~new_n9219_;
  assign new_n9221_ = new_n9217_ & ~new_n9220_;
  assign new_n9222_ = ~new_n7950_ & ~new_n9221_;
  assign new_n9223_ = new_n9214_ & new_n9222_;
  assign new_n9224_ = ~new_n9215_ & ~new_n9223_;
  assign new_n9225_ = ~new_n9207_ & new_n9224_;
  assign new_n9226_ = new_n9207_ & ~new_n9224_;
  assign new_n9227_ = ~new_n9225_ & ~new_n9226_;
  assign new_n9228_ = ~new_n9200_ & ~new_n9227_;
  assign new_n9229_ = ~new_n4154_ & ~new_n4162_;
  assign new_n9230_ = ~new_n4163_ & ~new_n9229_;
  assign new_n9231_ = ~new_n4140_ & new_n4154_;
  assign new_n9232_ = new_n4140_ & ~new_n4154_;
  assign new_n9233_ = ~new_n9231_ & ~new_n9232_;
  assign new_n9234_ = new_n9230_ & ~new_n9233_;
  assign new_n9235_ = ~new_n7963_ & ~new_n9234_;
  assign new_n9236_ = ~new_n4199_ & ~new_n4207_;
  assign new_n9237_ = ~new_n4208_ & ~new_n9236_;
  assign new_n9238_ = ~new_n4185_ & new_n4199_;
  assign new_n9239_ = new_n4185_ & ~new_n4199_;
  assign new_n9240_ = ~new_n9238_ & ~new_n9239_;
  assign new_n9241_ = new_n9237_ & ~new_n9240_;
  assign new_n9242_ = ~new_n7970_ & ~new_n9241_;
  assign new_n9243_ = new_n9235_ & ~new_n9242_;
  assign new_n9244_ = ~new_n9235_ & new_n9242_;
  assign new_n9245_ = ~new_n9243_ & ~new_n9244_;
  assign new_n9246_ = ~new_n4247_ & ~new_n4255_;
  assign new_n9247_ = ~new_n4256_ & ~new_n9246_;
  assign new_n9248_ = ~new_n4233_ & new_n4247_;
  assign new_n9249_ = new_n4233_ & ~new_n4247_;
  assign new_n9250_ = ~new_n9248_ & ~new_n9249_;
  assign new_n9251_ = new_n9247_ & ~new_n9250_;
  assign new_n9252_ = ~new_n7980_ & ~new_n9251_;
  assign new_n9253_ = ~new_n4292_ & ~new_n4300_;
  assign new_n9254_ = ~new_n4301_ & ~new_n9253_;
  assign new_n9255_ = ~new_n4278_ & new_n4292_;
  assign new_n9256_ = new_n4278_ & ~new_n4292_;
  assign new_n9257_ = ~new_n9255_ & ~new_n9256_;
  assign new_n9258_ = new_n9254_ & ~new_n9257_;
  assign new_n9259_ = ~new_n7987_ & ~new_n9258_;
  assign new_n9260_ = new_n9245_ & new_n9259_;
  assign new_n9261_ = ~new_n4338_ & ~new_n4346_;
  assign new_n9262_ = ~new_n4347_ & ~new_n9261_;
  assign new_n9263_ = ~new_n4324_ & new_n4338_;
  assign new_n9264_ = new_n4324_ & ~new_n4338_;
  assign new_n9265_ = ~new_n9263_ & ~new_n9264_;
  assign new_n9266_ = new_n9262_ & ~new_n9265_;
  assign new_n9267_ = ~new_n7995_ & ~new_n9266_;
  assign new_n9268_ = new_n9259_ & new_n9267_;
  assign new_n9269_ = ~new_n9260_ & ~new_n9268_;
  assign new_n9270_ = ~new_n9252_ & new_n9269_;
  assign new_n9271_ = new_n9252_ & ~new_n9269_;
  assign new_n9272_ = ~new_n9270_ & ~new_n9271_;
  assign new_n9273_ = ~new_n9245_ & ~new_n9272_;
  assign new_n9274_ = new_n9183_ & ~new_n9273_;
  assign new_n9275_ = ~new_n4390_ & ~new_n4398_;
  assign new_n9276_ = ~new_n4399_ & ~new_n9275_;
  assign new_n9277_ = ~new_n4376_ & new_n4390_;
  assign new_n9278_ = new_n4376_ & ~new_n4390_;
  assign new_n9279_ = ~new_n9277_ & ~new_n9278_;
  assign new_n9280_ = new_n9276_ & ~new_n9279_;
  assign new_n9281_ = ~new_n8009_ & ~new_n9280_;
  assign new_n9282_ = ~new_n4435_ & ~new_n4443_;
  assign new_n9283_ = ~new_n4444_ & ~new_n9282_;
  assign new_n9284_ = ~new_n4421_ & new_n4435_;
  assign new_n9285_ = new_n4421_ & ~new_n4435_;
  assign new_n9286_ = ~new_n9284_ & ~new_n9285_;
  assign new_n9287_ = new_n9283_ & ~new_n9286_;
  assign new_n9288_ = ~new_n8016_ & ~new_n9287_;
  assign new_n9289_ = new_n9281_ & ~new_n9288_;
  assign new_n9290_ = ~new_n9281_ & new_n9288_;
  assign new_n9291_ = ~new_n9289_ & ~new_n9290_;
  assign new_n9292_ = ~new_n4483_ & ~new_n4491_;
  assign new_n9293_ = ~new_n4492_ & ~new_n9292_;
  assign new_n9294_ = ~new_n4469_ & new_n4483_;
  assign new_n9295_ = new_n4469_ & ~new_n4483_;
  assign new_n9296_ = ~new_n9294_ & ~new_n9295_;
  assign new_n9297_ = new_n9293_ & ~new_n9296_;
  assign new_n9298_ = ~new_n8026_ & ~new_n9297_;
  assign new_n9299_ = ~new_n4528_ & ~new_n4536_;
  assign new_n9300_ = ~new_n4537_ & ~new_n9299_;
  assign new_n9301_ = ~new_n4514_ & new_n4528_;
  assign new_n9302_ = new_n4514_ & ~new_n4528_;
  assign new_n9303_ = ~new_n9301_ & ~new_n9302_;
  assign new_n9304_ = new_n9300_ & ~new_n9303_;
  assign new_n9305_ = ~new_n8033_ & ~new_n9304_;
  assign new_n9306_ = new_n9291_ & new_n9305_;
  assign new_n9307_ = ~new_n4574_ & ~new_n4582_;
  assign new_n9308_ = ~new_n4583_ & ~new_n9307_;
  assign new_n9309_ = ~new_n4560_ & new_n4574_;
  assign new_n9310_ = new_n4560_ & ~new_n4574_;
  assign new_n9311_ = ~new_n9309_ & ~new_n9310_;
  assign new_n9312_ = new_n9308_ & ~new_n9311_;
  assign new_n9313_ = ~new_n8041_ & ~new_n9312_;
  assign new_n9314_ = new_n9305_ & new_n9313_;
  assign new_n9315_ = ~new_n9306_ & ~new_n9314_;
  assign new_n9316_ = ~new_n9298_ & new_n9315_;
  assign new_n9317_ = new_n9298_ & ~new_n9315_;
  assign new_n9318_ = ~new_n9316_ & ~new_n9317_;
  assign new_n9319_ = ~new_n9291_ & ~new_n9318_;
  assign new_n9320_ = ~new_n9273_ & ~new_n9319_;
  assign new_n9321_ = ~new_n9274_ & ~new_n9320_;
  assign new_n9322_ = new_n9228_ & new_n9321_;
  assign new_n9323_ = ~new_n9228_ & ~new_n9321_;
  assign new_n9324_ = ~new_n9322_ & ~new_n9323_;
  assign A6346 = ~new_n9183_ & ~new_n9324_;
  assign new_n9326_ = ~new_n9180_ & ~new_n9322_;
  assign A6345 = ~new_n9183_ & ~new_n9326_;
  assign new_n9328_ = new_n9180_ & new_n9228_;
  assign new_n9329_ = ~new_n9183_ & ~new_n9328_;
  assign new_n9330_ = new_n9183_ & ~new_n9329_;
  assign new_n9331_ = new_n9183_ & new_n9328_;
  assign new_n9332_ = new_n9330_ & ~new_n9331_;
  assign new_n9333_ = new_n9228_ & ~new_n9332_;
  assign A6344 = new_n9321_ | new_n9333_;
  assign new_n9335_ = new_n9273_ & new_n9319_;
  assign new_n9336_ = ~new_n9320_ & ~new_n9335_;
  assign new_n9337_ = ~new_n9183_ & ~new_n9273_;
  assign new_n9338_ = new_n9183_ & new_n9273_;
  assign new_n9339_ = ~new_n9337_ & ~new_n9338_;
  assign new_n9340_ = new_n9336_ & ~new_n9339_;
  assign A6343 = new_n9333_ | new_n9340_;
  assign new_n9342_ = new_n9228_ & ~new_n9340_;
  assign new_n9343_ = ~new_n9228_ & new_n9340_;
  assign new_n9344_ = ~new_n9342_ & ~new_n9343_;
  assign A6342 = ~new_n9183_ & ~new_n9344_;
  assign new_n9346_ = ~new_n4647_ & ~new_n4655_;
  assign new_n9347_ = ~new_n4656_ & ~new_n9346_;
  assign new_n9348_ = ~new_n4633_ & new_n4647_;
  assign new_n9349_ = new_n4633_ & ~new_n4647_;
  assign new_n9350_ = ~new_n9348_ & ~new_n9349_;
  assign new_n9351_ = new_n9347_ & ~new_n9350_;
  assign new_n9352_ = ~new_n8080_ & ~new_n9351_;
  assign new_n9353_ = ~new_n4692_ & ~new_n4700_;
  assign new_n9354_ = ~new_n4701_ & ~new_n9353_;
  assign new_n9355_ = ~new_n4678_ & new_n4692_;
  assign new_n9356_ = new_n4678_ & ~new_n4692_;
  assign new_n9357_ = ~new_n9355_ & ~new_n9356_;
  assign new_n9358_ = new_n9354_ & ~new_n9357_;
  assign new_n9359_ = ~new_n8087_ & ~new_n9358_;
  assign new_n9360_ = new_n9352_ & ~new_n9359_;
  assign new_n9361_ = ~new_n9352_ & new_n9359_;
  assign new_n9362_ = ~new_n9360_ & ~new_n9361_;
  assign new_n9363_ = ~new_n4740_ & ~new_n4748_;
  assign new_n9364_ = ~new_n4749_ & ~new_n9363_;
  assign new_n9365_ = ~new_n4726_ & new_n4740_;
  assign new_n9366_ = new_n4726_ & ~new_n4740_;
  assign new_n9367_ = ~new_n9365_ & ~new_n9366_;
  assign new_n9368_ = new_n9364_ & ~new_n9367_;
  assign new_n9369_ = ~new_n8097_ & ~new_n9368_;
  assign new_n9370_ = ~new_n4785_ & ~new_n4793_;
  assign new_n9371_ = ~new_n4794_ & ~new_n9370_;
  assign new_n9372_ = ~new_n4771_ & new_n4785_;
  assign new_n9373_ = new_n4771_ & ~new_n4785_;
  assign new_n9374_ = ~new_n9372_ & ~new_n9373_;
  assign new_n9375_ = new_n9371_ & ~new_n9374_;
  assign new_n9376_ = ~new_n8104_ & ~new_n9375_;
  assign new_n9377_ = new_n9362_ & new_n9376_;
  assign new_n9378_ = ~new_n4831_ & ~new_n4839_;
  assign new_n9379_ = ~new_n4840_ & ~new_n9378_;
  assign new_n9380_ = ~new_n4817_ & new_n4831_;
  assign new_n9381_ = new_n4817_ & ~new_n4831_;
  assign new_n9382_ = ~new_n9380_ & ~new_n9381_;
  assign new_n9383_ = new_n9379_ & ~new_n9382_;
  assign new_n9384_ = ~new_n8112_ & ~new_n9383_;
  assign new_n9385_ = new_n9376_ & new_n9384_;
  assign new_n9386_ = ~new_n9377_ & ~new_n9385_;
  assign new_n9387_ = ~new_n9369_ & new_n9386_;
  assign new_n9388_ = new_n9369_ & ~new_n9386_;
  assign new_n9389_ = ~new_n9387_ & ~new_n9388_;
  assign new_n9390_ = ~new_n9362_ & ~new_n9389_;
  assign new_n9391_ = ~new_n4882_ & ~new_n4890_;
  assign new_n9392_ = ~new_n4891_ & ~new_n9391_;
  assign new_n9393_ = ~new_n4868_ & new_n4882_;
  assign new_n9394_ = new_n4868_ & ~new_n4882_;
  assign new_n9395_ = ~new_n9393_ & ~new_n9394_;
  assign new_n9396_ = new_n9392_ & ~new_n9395_;
  assign new_n9397_ = ~new_n8125_ & ~new_n9396_;
  assign new_n9398_ = ~new_n4927_ & ~new_n4935_;
  assign new_n9399_ = ~new_n4936_ & ~new_n9398_;
  assign new_n9400_ = ~new_n4913_ & new_n4927_;
  assign new_n9401_ = new_n4913_ & ~new_n4927_;
  assign new_n9402_ = ~new_n9400_ & ~new_n9401_;
  assign new_n9403_ = new_n9399_ & ~new_n9402_;
  assign new_n9404_ = ~new_n8132_ & ~new_n9403_;
  assign new_n9405_ = new_n9397_ & ~new_n9404_;
  assign new_n9406_ = ~new_n9397_ & new_n9404_;
  assign new_n9407_ = ~new_n9405_ & ~new_n9406_;
  assign new_n9408_ = ~new_n4975_ & ~new_n4983_;
  assign new_n9409_ = ~new_n4984_ & ~new_n9408_;
  assign new_n9410_ = ~new_n4961_ & new_n4975_;
  assign new_n9411_ = new_n4961_ & ~new_n4975_;
  assign new_n9412_ = ~new_n9410_ & ~new_n9411_;
  assign new_n9413_ = new_n9409_ & ~new_n9412_;
  assign new_n9414_ = ~new_n8142_ & ~new_n9413_;
  assign new_n9415_ = ~new_n5020_ & ~new_n5028_;
  assign new_n9416_ = ~new_n5029_ & ~new_n9415_;
  assign new_n9417_ = ~new_n5006_ & new_n5020_;
  assign new_n9418_ = new_n5006_ & ~new_n5020_;
  assign new_n9419_ = ~new_n9417_ & ~new_n9418_;
  assign new_n9420_ = new_n9416_ & ~new_n9419_;
  assign new_n9421_ = ~new_n8149_ & ~new_n9420_;
  assign new_n9422_ = new_n9407_ & new_n9421_;
  assign new_n9423_ = ~new_n5066_ & ~new_n5074_;
  assign new_n9424_ = ~new_n5075_ & ~new_n9423_;
  assign new_n9425_ = ~new_n5052_ & new_n5066_;
  assign new_n9426_ = new_n5052_ & ~new_n5066_;
  assign new_n9427_ = ~new_n9425_ & ~new_n9426_;
  assign new_n9428_ = new_n9424_ & ~new_n9427_;
  assign new_n9429_ = ~new_n8157_ & ~new_n9428_;
  assign new_n9430_ = new_n9421_ & new_n9429_;
  assign new_n9431_ = ~new_n9422_ & ~new_n9430_;
  assign new_n9432_ = ~new_n9414_ & new_n9431_;
  assign new_n9433_ = new_n9414_ & ~new_n9431_;
  assign new_n9434_ = ~new_n9432_ & ~new_n9433_;
  assign new_n9435_ = ~new_n9407_ & ~new_n9434_;
  assign new_n9436_ = ~new_n9390_ & new_n9435_;
  assign new_n9437_ = new_n9390_ & ~new_n9435_;
  assign new_n9438_ = ~new_n9436_ & ~new_n9437_;
  assign new_n9439_ = ~new_n5120_ & ~new_n5128_;
  assign new_n9440_ = ~new_n5129_ & ~new_n9439_;
  assign new_n9441_ = ~new_n5106_ & new_n5120_;
  assign new_n9442_ = new_n5106_ & ~new_n5120_;
  assign new_n9443_ = ~new_n9441_ & ~new_n9442_;
  assign new_n9444_ = new_n9440_ & ~new_n9443_;
  assign new_n9445_ = ~new_n8173_ & ~new_n9444_;
  assign new_n9446_ = ~new_n5165_ & ~new_n5173_;
  assign new_n9447_ = ~new_n5174_ & ~new_n9446_;
  assign new_n9448_ = ~new_n5151_ & new_n5165_;
  assign new_n9449_ = new_n5151_ & ~new_n5165_;
  assign new_n9450_ = ~new_n9448_ & ~new_n9449_;
  assign new_n9451_ = new_n9447_ & ~new_n9450_;
  assign new_n9452_ = ~new_n8180_ & ~new_n9451_;
  assign new_n9453_ = new_n9445_ & ~new_n9452_;
  assign new_n9454_ = ~new_n9445_ & new_n9452_;
  assign new_n9455_ = ~new_n9453_ & ~new_n9454_;
  assign new_n9456_ = ~new_n5213_ & ~new_n5221_;
  assign new_n9457_ = ~new_n5222_ & ~new_n9456_;
  assign new_n9458_ = ~new_n5199_ & new_n5213_;
  assign new_n9459_ = new_n5199_ & ~new_n5213_;
  assign new_n9460_ = ~new_n9458_ & ~new_n9459_;
  assign new_n9461_ = new_n9457_ & ~new_n9460_;
  assign new_n9462_ = ~new_n8190_ & ~new_n9461_;
  assign new_n9463_ = ~new_n5258_ & ~new_n5266_;
  assign new_n9464_ = ~new_n5267_ & ~new_n9463_;
  assign new_n9465_ = ~new_n5244_ & new_n5258_;
  assign new_n9466_ = new_n5244_ & ~new_n5258_;
  assign new_n9467_ = ~new_n9465_ & ~new_n9466_;
  assign new_n9468_ = new_n9464_ & ~new_n9467_;
  assign new_n9469_ = ~new_n8197_ & ~new_n9468_;
  assign new_n9470_ = new_n9455_ & new_n9469_;
  assign new_n9471_ = ~new_n5304_ & ~new_n5312_;
  assign new_n9472_ = ~new_n5313_ & ~new_n9471_;
  assign new_n9473_ = ~new_n5290_ & new_n5304_;
  assign new_n9474_ = new_n5290_ & ~new_n5304_;
  assign new_n9475_ = ~new_n9473_ & ~new_n9474_;
  assign new_n9476_ = new_n9472_ & ~new_n9475_;
  assign new_n9477_ = ~new_n8205_ & ~new_n9476_;
  assign new_n9478_ = new_n9469_ & new_n9477_;
  assign new_n9479_ = ~new_n9470_ & ~new_n9478_;
  assign new_n9480_ = ~new_n9462_ & new_n9479_;
  assign new_n9481_ = new_n9462_ & ~new_n9479_;
  assign new_n9482_ = ~new_n9480_ & ~new_n9481_;
  assign new_n9483_ = ~new_n9455_ & ~new_n9482_;
  assign new_n9484_ = ~new_n5355_ & ~new_n5363_;
  assign new_n9485_ = ~new_n5364_ & ~new_n9484_;
  assign new_n9486_ = ~new_n5341_ & new_n5355_;
  assign new_n9487_ = new_n5341_ & ~new_n5355_;
  assign new_n9488_ = ~new_n9486_ & ~new_n9487_;
  assign new_n9489_ = new_n9485_ & ~new_n9488_;
  assign new_n9490_ = ~new_n8218_ & ~new_n9489_;
  assign new_n9491_ = ~new_n5400_ & ~new_n5408_;
  assign new_n9492_ = ~new_n5409_ & ~new_n9491_;
  assign new_n9493_ = ~new_n5386_ & new_n5400_;
  assign new_n9494_ = new_n5386_ & ~new_n5400_;
  assign new_n9495_ = ~new_n9493_ & ~new_n9494_;
  assign new_n9496_ = new_n9492_ & ~new_n9495_;
  assign new_n9497_ = ~new_n8225_ & ~new_n9496_;
  assign new_n9498_ = new_n9490_ & ~new_n9497_;
  assign new_n9499_ = ~new_n9490_ & new_n9497_;
  assign new_n9500_ = ~new_n9498_ & ~new_n9499_;
  assign new_n9501_ = ~new_n5448_ & ~new_n5456_;
  assign new_n9502_ = ~new_n5457_ & ~new_n9501_;
  assign new_n9503_ = ~new_n5434_ & new_n5448_;
  assign new_n9504_ = new_n5434_ & ~new_n5448_;
  assign new_n9505_ = ~new_n9503_ & ~new_n9504_;
  assign new_n9506_ = new_n9502_ & ~new_n9505_;
  assign new_n9507_ = ~new_n8235_ & ~new_n9506_;
  assign new_n9508_ = ~new_n5493_ & ~new_n5501_;
  assign new_n9509_ = ~new_n5502_ & ~new_n9508_;
  assign new_n9510_ = ~new_n5479_ & new_n5493_;
  assign new_n9511_ = new_n5479_ & ~new_n5493_;
  assign new_n9512_ = ~new_n9510_ & ~new_n9511_;
  assign new_n9513_ = new_n9509_ & ~new_n9512_;
  assign new_n9514_ = ~new_n8242_ & ~new_n9513_;
  assign new_n9515_ = new_n9500_ & new_n9514_;
  assign new_n9516_ = ~new_n5539_ & ~new_n5547_;
  assign new_n9517_ = ~new_n5548_ & ~new_n9516_;
  assign new_n9518_ = ~new_n5525_ & new_n5539_;
  assign new_n9519_ = new_n5525_ & ~new_n5539_;
  assign new_n9520_ = ~new_n9518_ & ~new_n9519_;
  assign new_n9521_ = new_n9517_ & ~new_n9520_;
  assign new_n9522_ = ~new_n8250_ & ~new_n9521_;
  assign new_n9523_ = new_n9514_ & new_n9522_;
  assign new_n9524_ = ~new_n9515_ & ~new_n9523_;
  assign new_n9525_ = ~new_n9507_ & new_n9524_;
  assign new_n9526_ = new_n9507_ & ~new_n9524_;
  assign new_n9527_ = ~new_n9525_ & ~new_n9526_;
  assign new_n9528_ = ~new_n9500_ & ~new_n9527_;
  assign new_n9529_ = new_n9438_ & ~new_n9528_;
  assign new_n9530_ = ~new_n5591_ & ~new_n5599_;
  assign new_n9531_ = ~new_n5600_ & ~new_n9530_;
  assign new_n9532_ = ~new_n5577_ & new_n5591_;
  assign new_n9533_ = new_n5577_ & ~new_n5591_;
  assign new_n9534_ = ~new_n9532_ & ~new_n9533_;
  assign new_n9535_ = new_n9531_ & ~new_n9534_;
  assign new_n9536_ = ~new_n8264_ & ~new_n9535_;
  assign new_n9537_ = ~new_n5636_ & ~new_n5644_;
  assign new_n9538_ = ~new_n5645_ & ~new_n9537_;
  assign new_n9539_ = ~new_n5622_ & new_n5636_;
  assign new_n9540_ = new_n5622_ & ~new_n5636_;
  assign new_n9541_ = ~new_n9539_ & ~new_n9540_;
  assign new_n9542_ = new_n9538_ & ~new_n9541_;
  assign new_n9543_ = ~new_n8271_ & ~new_n9542_;
  assign new_n9544_ = new_n9536_ & ~new_n9543_;
  assign new_n9545_ = ~new_n9536_ & new_n9543_;
  assign new_n9546_ = ~new_n9544_ & ~new_n9545_;
  assign new_n9547_ = ~new_n5684_ & ~new_n5692_;
  assign new_n9548_ = ~new_n5693_ & ~new_n9547_;
  assign new_n9549_ = ~new_n5670_ & new_n5684_;
  assign new_n9550_ = new_n5670_ & ~new_n5684_;
  assign new_n9551_ = ~new_n9549_ & ~new_n9550_;
  assign new_n9552_ = new_n9548_ & ~new_n9551_;
  assign new_n9553_ = ~new_n8281_ & ~new_n9552_;
  assign new_n9554_ = ~new_n5729_ & ~new_n5737_;
  assign new_n9555_ = ~new_n5738_ & ~new_n9554_;
  assign new_n9556_ = ~new_n5715_ & new_n5729_;
  assign new_n9557_ = new_n5715_ & ~new_n5729_;
  assign new_n9558_ = ~new_n9556_ & ~new_n9557_;
  assign new_n9559_ = new_n9555_ & ~new_n9558_;
  assign new_n9560_ = ~new_n8288_ & ~new_n9559_;
  assign new_n9561_ = new_n9546_ & new_n9560_;
  assign new_n9562_ = ~new_n5775_ & ~new_n5783_;
  assign new_n9563_ = ~new_n5784_ & ~new_n9562_;
  assign new_n9564_ = ~new_n5761_ & new_n5775_;
  assign new_n9565_ = new_n5761_ & ~new_n5775_;
  assign new_n9566_ = ~new_n9564_ & ~new_n9565_;
  assign new_n9567_ = new_n9563_ & ~new_n9566_;
  assign new_n9568_ = ~new_n8296_ & ~new_n9567_;
  assign new_n9569_ = new_n9560_ & new_n9568_;
  assign new_n9570_ = ~new_n9561_ & ~new_n9569_;
  assign new_n9571_ = ~new_n9553_ & new_n9570_;
  assign new_n9572_ = new_n9553_ & ~new_n9570_;
  assign new_n9573_ = ~new_n9571_ & ~new_n9572_;
  assign new_n9574_ = ~new_n9546_ & ~new_n9573_;
  assign new_n9575_ = ~new_n9528_ & ~new_n9574_;
  assign new_n9576_ = ~new_n9529_ & ~new_n9575_;
  assign new_n9577_ = new_n9483_ & new_n9576_;
  assign new_n9578_ = ~new_n9483_ & ~new_n9576_;
  assign new_n9579_ = ~new_n9577_ & ~new_n9578_;
  assign A6313 = ~new_n9438_ & ~new_n9579_;
  assign new_n9581_ = ~new_n9435_ & ~new_n9577_;
  assign A6312 = ~new_n9438_ & ~new_n9581_;
  assign new_n9583_ = new_n9435_ & new_n9483_;
  assign new_n9584_ = ~new_n9438_ & ~new_n9583_;
  assign new_n9585_ = new_n9438_ & ~new_n9584_;
  assign new_n9586_ = new_n9438_ & new_n9583_;
  assign new_n9587_ = new_n9585_ & ~new_n9586_;
  assign new_n9588_ = new_n9483_ & ~new_n9587_;
  assign A6311 = new_n9576_ | new_n9588_;
  assign new_n9590_ = new_n9528_ & new_n9574_;
  assign new_n9591_ = ~new_n9575_ & ~new_n9590_;
  assign new_n9592_ = ~new_n9438_ & ~new_n9528_;
  assign new_n9593_ = new_n9438_ & new_n9528_;
  assign new_n9594_ = ~new_n9592_ & ~new_n9593_;
  assign new_n9595_ = new_n9591_ & ~new_n9594_;
  assign A6310 = new_n9588_ | new_n9595_;
  assign new_n9597_ = new_n9483_ & ~new_n9595_;
  assign new_n9598_ = ~new_n9483_ & new_n9595_;
  assign new_n9599_ = ~new_n9597_ & ~new_n9598_;
  assign A6309 = ~new_n9438_ & ~new_n9599_;
  assign new_n9601_ = new_n5850_ & new_n8331_;
  assign new_n9602_ = ~new_n5839_ & ~new_n9601_;
  assign new_n9603_ = ~new_n5842_ & ~new_n9602_;
  assign new_n9604_ = new_n5873_ & new_n5878_;
  assign new_n9605_ = ~new_n5879_ & ~new_n9604_;
  assign new_n9606_ = ~new_n5865_ & ~new_n5873_;
  assign new_n9607_ = new_n5865_ & new_n5873_;
  assign new_n9608_ = ~new_n9606_ & ~new_n9607_;
  assign new_n9609_ = new_n9605_ & ~new_n9608_;
  assign new_n9610_ = ~new_n8338_ & ~new_n9609_;
  assign new_n9611_ = ~new_n9603_ & ~new_n9610_;
  assign new_n9612_ = new_n9603_ & new_n9610_;
  assign new_n9613_ = ~new_n9611_ & ~new_n9612_;
  assign new_n9614_ = new_n5906_ & new_n5911_;
  assign new_n9615_ = ~new_n5912_ & ~new_n9614_;
  assign new_n9616_ = ~new_n5898_ & ~new_n5906_;
  assign new_n9617_ = new_n5898_ & new_n5906_;
  assign new_n9618_ = ~new_n9616_ & ~new_n9617_;
  assign new_n9619_ = new_n9615_ & ~new_n9618_;
  assign new_n9620_ = ~new_n8348_ & ~new_n9619_;
  assign new_n9621_ = new_n5936_ & new_n5941_;
  assign new_n9622_ = ~new_n5942_ & ~new_n9621_;
  assign new_n9623_ = ~new_n5928_ & ~new_n5936_;
  assign new_n9624_ = new_n5928_ & new_n5936_;
  assign new_n9625_ = ~new_n9623_ & ~new_n9624_;
  assign new_n9626_ = new_n9622_ & ~new_n9625_;
  assign new_n9627_ = ~new_n8355_ & ~new_n9626_;
  assign new_n9628_ = new_n9613_ & new_n9627_;
  assign new_n9629_ = new_n5967_ & new_n5972_;
  assign new_n9630_ = ~new_n5973_ & ~new_n9629_;
  assign new_n9631_ = ~new_n5959_ & ~new_n5967_;
  assign new_n9632_ = new_n5959_ & new_n5967_;
  assign new_n9633_ = ~new_n9631_ & ~new_n9632_;
  assign new_n9634_ = new_n9630_ & ~new_n9633_;
  assign new_n9635_ = ~new_n8363_ & ~new_n9634_;
  assign new_n9636_ = new_n9627_ & new_n9635_;
  assign new_n9637_ = ~new_n9628_ & ~new_n9636_;
  assign new_n9638_ = ~new_n9620_ & new_n9637_;
  assign new_n9639_ = new_n9620_ & ~new_n9637_;
  assign new_n9640_ = ~new_n9638_ & ~new_n9639_;
  assign new_n9641_ = ~new_n9613_ & ~new_n9640_;
  assign new_n9642_ = new_n6003_ & new_n6008_;
  assign new_n9643_ = ~new_n6009_ & ~new_n9642_;
  assign new_n9644_ = ~new_n5995_ & ~new_n6003_;
  assign new_n9645_ = new_n5995_ & new_n6003_;
  assign new_n9646_ = ~new_n9644_ & ~new_n9645_;
  assign new_n9647_ = new_n9643_ & ~new_n9646_;
  assign new_n9648_ = ~new_n8376_ & ~new_n9647_;
  assign new_n9649_ = new_n6033_ & new_n6038_;
  assign new_n9650_ = ~new_n6039_ & ~new_n9649_;
  assign new_n9651_ = ~new_n6025_ & ~new_n6033_;
  assign new_n9652_ = new_n6025_ & new_n6033_;
  assign new_n9653_ = ~new_n9651_ & ~new_n9652_;
  assign new_n9654_ = new_n9650_ & ~new_n9653_;
  assign new_n9655_ = ~new_n8383_ & ~new_n9654_;
  assign new_n9656_ = new_n9648_ & ~new_n9655_;
  assign new_n9657_ = ~new_n9648_ & new_n9655_;
  assign new_n9658_ = ~new_n9656_ & ~new_n9657_;
  assign new_n9659_ = new_n6066_ & new_n6071_;
  assign new_n9660_ = ~new_n6072_ & ~new_n9659_;
  assign new_n9661_ = ~new_n6058_ & ~new_n6066_;
  assign new_n9662_ = new_n6058_ & new_n6066_;
  assign new_n9663_ = ~new_n9661_ & ~new_n9662_;
  assign new_n9664_ = new_n9660_ & ~new_n9663_;
  assign new_n9665_ = ~new_n8393_ & ~new_n9664_;
  assign new_n9666_ = new_n6096_ & new_n6101_;
  assign new_n9667_ = ~new_n6102_ & ~new_n9666_;
  assign new_n9668_ = ~new_n6088_ & ~new_n6096_;
  assign new_n9669_ = new_n6088_ & new_n6096_;
  assign new_n9670_ = ~new_n9668_ & ~new_n9669_;
  assign new_n9671_ = new_n9667_ & ~new_n9670_;
  assign new_n9672_ = ~new_n8400_ & ~new_n9671_;
  assign new_n9673_ = new_n9658_ & new_n9672_;
  assign new_n9674_ = new_n6127_ & new_n6132_;
  assign new_n9675_ = ~new_n6133_ & ~new_n9674_;
  assign new_n9676_ = ~new_n6119_ & ~new_n6127_;
  assign new_n9677_ = new_n6119_ & new_n6127_;
  assign new_n9678_ = ~new_n9676_ & ~new_n9677_;
  assign new_n9679_ = new_n9675_ & ~new_n9678_;
  assign new_n9680_ = ~new_n8408_ & ~new_n9679_;
  assign new_n9681_ = new_n9672_ & new_n9680_;
  assign new_n9682_ = ~new_n9673_ & ~new_n9681_;
  assign new_n9683_ = ~new_n9665_ & new_n9682_;
  assign new_n9684_ = new_n9665_ & ~new_n9682_;
  assign new_n9685_ = ~new_n9683_ & ~new_n9684_;
  assign new_n9686_ = ~new_n9658_ & ~new_n9685_;
  assign new_n9687_ = ~new_n9641_ & new_n9686_;
  assign new_n9688_ = new_n9641_ & ~new_n9686_;
  assign new_n9689_ = ~new_n9687_ & ~new_n9688_;
  assign new_n9690_ = new_n6166_ & new_n6171_;
  assign new_n9691_ = ~new_n6172_ & ~new_n9690_;
  assign new_n9692_ = ~new_n6158_ & ~new_n6166_;
  assign new_n9693_ = new_n6158_ & new_n6166_;
  assign new_n9694_ = ~new_n9692_ & ~new_n9693_;
  assign new_n9695_ = new_n9691_ & ~new_n9694_;
  assign new_n9696_ = ~new_n8424_ & ~new_n9695_;
  assign new_n9697_ = new_n6196_ & new_n6201_;
  assign new_n9698_ = ~new_n6202_ & ~new_n9697_;
  assign new_n9699_ = ~new_n6188_ & ~new_n6196_;
  assign new_n9700_ = new_n6188_ & new_n6196_;
  assign new_n9701_ = ~new_n9699_ & ~new_n9700_;
  assign new_n9702_ = new_n9698_ & ~new_n9701_;
  assign new_n9703_ = ~new_n8431_ & ~new_n9702_;
  assign new_n9704_ = new_n9696_ & ~new_n9703_;
  assign new_n9705_ = ~new_n9696_ & new_n9703_;
  assign new_n9706_ = ~new_n9704_ & ~new_n9705_;
  assign new_n9707_ = new_n6229_ & new_n6234_;
  assign new_n9708_ = ~new_n6235_ & ~new_n9707_;
  assign new_n9709_ = ~new_n6221_ & ~new_n6229_;
  assign new_n9710_ = new_n6221_ & new_n6229_;
  assign new_n9711_ = ~new_n9709_ & ~new_n9710_;
  assign new_n9712_ = new_n9708_ & ~new_n9711_;
  assign new_n9713_ = ~new_n8441_ & ~new_n9712_;
  assign new_n9714_ = new_n6259_ & new_n6264_;
  assign new_n9715_ = ~new_n6265_ & ~new_n9714_;
  assign new_n9716_ = ~new_n6251_ & ~new_n6259_;
  assign new_n9717_ = new_n6251_ & new_n6259_;
  assign new_n9718_ = ~new_n9716_ & ~new_n9717_;
  assign new_n9719_ = new_n9715_ & ~new_n9718_;
  assign new_n9720_ = ~new_n8448_ & ~new_n9719_;
  assign new_n9721_ = new_n9706_ & new_n9720_;
  assign new_n9722_ = new_n6290_ & new_n6295_;
  assign new_n9723_ = ~new_n6296_ & ~new_n9722_;
  assign new_n9724_ = ~new_n6282_ & ~new_n6290_;
  assign new_n9725_ = new_n6282_ & new_n6290_;
  assign new_n9726_ = ~new_n9724_ & ~new_n9725_;
  assign new_n9727_ = new_n9723_ & ~new_n9726_;
  assign new_n9728_ = ~new_n8456_ & ~new_n9727_;
  assign new_n9729_ = new_n9720_ & new_n9728_;
  assign new_n9730_ = ~new_n9721_ & ~new_n9729_;
  assign new_n9731_ = ~new_n9713_ & new_n9730_;
  assign new_n9732_ = new_n9713_ & ~new_n9730_;
  assign new_n9733_ = ~new_n9731_ & ~new_n9732_;
  assign new_n9734_ = ~new_n9706_ & ~new_n9733_;
  assign new_n9735_ = new_n6326_ & new_n6331_;
  assign new_n9736_ = ~new_n6332_ & ~new_n9735_;
  assign new_n9737_ = ~new_n6318_ & ~new_n6326_;
  assign new_n9738_ = new_n6318_ & new_n6326_;
  assign new_n9739_ = ~new_n9737_ & ~new_n9738_;
  assign new_n9740_ = new_n9736_ & ~new_n9739_;
  assign new_n9741_ = ~new_n8469_ & ~new_n9740_;
  assign new_n9742_ = new_n6356_ & new_n6361_;
  assign new_n9743_ = ~new_n6362_ & ~new_n9742_;
  assign new_n9744_ = ~new_n6348_ & ~new_n6356_;
  assign new_n9745_ = new_n6348_ & new_n6356_;
  assign new_n9746_ = ~new_n9744_ & ~new_n9745_;
  assign new_n9747_ = new_n9743_ & ~new_n9746_;
  assign new_n9748_ = ~new_n8476_ & ~new_n9747_;
  assign new_n9749_ = new_n9741_ & ~new_n9748_;
  assign new_n9750_ = ~new_n9741_ & new_n9748_;
  assign new_n9751_ = ~new_n9749_ & ~new_n9750_;
  assign new_n9752_ = new_n6389_ & new_n6394_;
  assign new_n9753_ = ~new_n6395_ & ~new_n9752_;
  assign new_n9754_ = ~new_n6381_ & ~new_n6389_;
  assign new_n9755_ = new_n6381_ & new_n6389_;
  assign new_n9756_ = ~new_n9754_ & ~new_n9755_;
  assign new_n9757_ = new_n9753_ & ~new_n9756_;
  assign new_n9758_ = ~new_n8486_ & ~new_n9757_;
  assign new_n9759_ = new_n6419_ & new_n6424_;
  assign new_n9760_ = ~new_n6425_ & ~new_n9759_;
  assign new_n9761_ = ~new_n6411_ & ~new_n6419_;
  assign new_n9762_ = new_n6411_ & new_n6419_;
  assign new_n9763_ = ~new_n9761_ & ~new_n9762_;
  assign new_n9764_ = new_n9760_ & ~new_n9763_;
  assign new_n9765_ = ~new_n8493_ & ~new_n9764_;
  assign new_n9766_ = new_n9751_ & new_n9765_;
  assign new_n9767_ = new_n6450_ & new_n6455_;
  assign new_n9768_ = ~new_n6456_ & ~new_n9767_;
  assign new_n9769_ = ~new_n6442_ & ~new_n6450_;
  assign new_n9770_ = new_n6442_ & new_n6450_;
  assign new_n9771_ = ~new_n9769_ & ~new_n9770_;
  assign new_n9772_ = new_n9768_ & ~new_n9771_;
  assign new_n9773_ = ~new_n8501_ & ~new_n9772_;
  assign new_n9774_ = new_n9765_ & new_n9773_;
  assign new_n9775_ = ~new_n9766_ & ~new_n9774_;
  assign new_n9776_ = ~new_n9758_ & new_n9775_;
  assign new_n9777_ = new_n9758_ & ~new_n9775_;
  assign new_n9778_ = ~new_n9776_ & ~new_n9777_;
  assign new_n9779_ = ~new_n9751_ & ~new_n9778_;
  assign new_n9780_ = new_n9689_ & ~new_n9779_;
  assign new_n9781_ = new_n6487_ & new_n6492_;
  assign new_n9782_ = ~new_n6493_ & ~new_n9781_;
  assign new_n9783_ = ~new_n6479_ & ~new_n6487_;
  assign new_n9784_ = new_n6479_ & new_n6487_;
  assign new_n9785_ = ~new_n9783_ & ~new_n9784_;
  assign new_n9786_ = new_n9782_ & ~new_n9785_;
  assign new_n9787_ = ~new_n8515_ & ~new_n9786_;
  assign new_n9788_ = new_n6517_ & new_n6522_;
  assign new_n9789_ = ~new_n6523_ & ~new_n9788_;
  assign new_n9790_ = ~new_n6509_ & ~new_n6517_;
  assign new_n9791_ = new_n6509_ & new_n6517_;
  assign new_n9792_ = ~new_n9790_ & ~new_n9791_;
  assign new_n9793_ = new_n9789_ & ~new_n9792_;
  assign new_n9794_ = ~new_n8522_ & ~new_n9793_;
  assign new_n9795_ = new_n9787_ & ~new_n9794_;
  assign new_n9796_ = ~new_n9787_ & new_n9794_;
  assign new_n9797_ = ~new_n9795_ & ~new_n9796_;
  assign new_n9798_ = new_n6550_ & new_n6555_;
  assign new_n9799_ = ~new_n6556_ & ~new_n9798_;
  assign new_n9800_ = ~new_n6542_ & ~new_n6550_;
  assign new_n9801_ = new_n6542_ & new_n6550_;
  assign new_n9802_ = ~new_n9800_ & ~new_n9801_;
  assign new_n9803_ = new_n9799_ & ~new_n9802_;
  assign new_n9804_ = ~new_n8532_ & ~new_n9803_;
  assign new_n9805_ = new_n6580_ & new_n6585_;
  assign new_n9806_ = ~new_n6586_ & ~new_n9805_;
  assign new_n9807_ = ~new_n6572_ & ~new_n6580_;
  assign new_n9808_ = new_n6572_ & new_n6580_;
  assign new_n9809_ = ~new_n9807_ & ~new_n9808_;
  assign new_n9810_ = new_n9806_ & ~new_n9809_;
  assign new_n9811_ = ~new_n8539_ & ~new_n9810_;
  assign new_n9812_ = new_n9797_ & new_n9811_;
  assign new_n9813_ = new_n6611_ & new_n6616_;
  assign new_n9814_ = ~new_n6617_ & ~new_n9813_;
  assign new_n9815_ = ~new_n6603_ & ~new_n6611_;
  assign new_n9816_ = new_n6603_ & new_n6611_;
  assign new_n9817_ = ~new_n9815_ & ~new_n9816_;
  assign new_n9818_ = new_n9814_ & ~new_n9817_;
  assign new_n9819_ = ~new_n8547_ & ~new_n9818_;
  assign new_n9820_ = new_n9811_ & new_n9819_;
  assign new_n9821_ = ~new_n9812_ & ~new_n9820_;
  assign new_n9822_ = ~new_n9804_ & new_n9821_;
  assign new_n9823_ = new_n9804_ & ~new_n9821_;
  assign new_n9824_ = ~new_n9822_ & ~new_n9823_;
  assign new_n9825_ = ~new_n9797_ & ~new_n9824_;
  assign new_n9826_ = ~new_n9779_ & ~new_n9825_;
  assign new_n9827_ = ~new_n9780_ & ~new_n9826_;
  assign new_n9828_ = new_n9734_ & new_n9827_;
  assign new_n9829_ = ~new_n9734_ & ~new_n9827_;
  assign new_n9830_ = ~new_n9828_ & ~new_n9829_;
  assign A6280 = ~new_n9689_ & ~new_n9830_;
  assign new_n9832_ = ~new_n9686_ & ~new_n9828_;
  assign A6279 = ~new_n9689_ & ~new_n9832_;
  assign new_n9834_ = new_n9686_ & new_n9734_;
  assign new_n9835_ = ~new_n9689_ & ~new_n9834_;
  assign new_n9836_ = new_n9689_ & ~new_n9835_;
  assign new_n9837_ = new_n9689_ & new_n9834_;
  assign new_n9838_ = new_n9836_ & ~new_n9837_;
  assign new_n9839_ = new_n9734_ & ~new_n9838_;
  assign A6278 = new_n9827_ | new_n9839_;
  assign new_n9841_ = new_n9779_ & new_n9825_;
  assign new_n9842_ = ~new_n9826_ & ~new_n9841_;
  assign new_n9843_ = ~new_n9689_ & ~new_n9779_;
  assign new_n9844_ = new_n9689_ & new_n9779_;
  assign new_n9845_ = ~new_n9843_ & ~new_n9844_;
  assign new_n9846_ = new_n9842_ & ~new_n9845_;
  assign A6277 = new_n9839_ | new_n9846_;
  assign new_n9848_ = new_n9734_ & ~new_n9846_;
  assign new_n9849_ = ~new_n9734_ & new_n9846_;
  assign new_n9850_ = ~new_n9848_ & ~new_n9849_;
  assign A6276 = ~new_n9689_ & ~new_n9850_;
  assign new_n9852_ = new_n1287_ & ~new_n8586_;
  assign new_n9853_ = ~new_n1287_ & new_n8586_;
  assign new_n9854_ = ~new_n9852_ & ~new_n9853_;
  assign new_n9855_ = ~new_n1277_ & ~new_n9854_;
  assign new_n9856_ = new_n1347_ & ~new_n8593_;
  assign new_n9857_ = ~new_n1347_ & new_n8593_;
  assign new_n9858_ = ~new_n9856_ & ~new_n9857_;
  assign new_n9859_ = ~new_n1337_ & ~new_n9858_;
  assign new_n9860_ = ~new_n9855_ & new_n9859_;
  assign new_n9861_ = new_n9855_ & ~new_n9859_;
  assign new_n9862_ = ~new_n9860_ & ~new_n9861_;
  assign new_n9863_ = new_n1410_ & ~new_n8603_;
  assign new_n9864_ = ~new_n1410_ & new_n8603_;
  assign new_n9865_ = ~new_n9863_ & ~new_n9864_;
  assign new_n9866_ = ~new_n1400_ & ~new_n9865_;
  assign new_n9867_ = new_n1470_ & ~new_n8610_;
  assign new_n9868_ = ~new_n1470_ & new_n8610_;
  assign new_n9869_ = ~new_n9867_ & ~new_n9868_;
  assign new_n9870_ = ~new_n1460_ & ~new_n9869_;
  assign new_n9871_ = new_n9862_ & ~new_n9870_;
  assign new_n9872_ = new_n1531_ & ~new_n8618_;
  assign new_n9873_ = ~new_n1531_ & new_n8618_;
  assign new_n9874_ = ~new_n9872_ & ~new_n9873_;
  assign new_n9875_ = ~new_n1521_ & ~new_n9874_;
  assign new_n9876_ = ~new_n9870_ & ~new_n9875_;
  assign new_n9877_ = ~new_n9871_ & ~new_n9876_;
  assign new_n9878_ = new_n9866_ & new_n9877_;
  assign new_n9879_ = ~new_n9866_ & ~new_n9877_;
  assign new_n9880_ = ~new_n9878_ & ~new_n9879_;
  assign new_n9881_ = ~new_n9862_ & ~new_n9880_;
  assign new_n9882_ = new_n1597_ & ~new_n8631_;
  assign new_n9883_ = ~new_n1597_ & new_n8631_;
  assign new_n9884_ = ~new_n9882_ & ~new_n9883_;
  assign new_n9885_ = ~new_n1587_ & ~new_n9884_;
  assign new_n9886_ = new_n1657_ & ~new_n8638_;
  assign new_n9887_ = ~new_n1657_ & new_n8638_;
  assign new_n9888_ = ~new_n9886_ & ~new_n9887_;
  assign new_n9889_ = ~new_n1647_ & ~new_n9888_;
  assign new_n9890_ = ~new_n9885_ & new_n9889_;
  assign new_n9891_ = new_n9885_ & ~new_n9889_;
  assign new_n9892_ = ~new_n9890_ & ~new_n9891_;
  assign new_n9893_ = new_n1720_ & ~new_n8648_;
  assign new_n9894_ = ~new_n1720_ & new_n8648_;
  assign new_n9895_ = ~new_n9893_ & ~new_n9894_;
  assign new_n9896_ = ~new_n1710_ & ~new_n9895_;
  assign new_n9897_ = new_n1780_ & ~new_n8655_;
  assign new_n9898_ = ~new_n1780_ & new_n8655_;
  assign new_n9899_ = ~new_n9897_ & ~new_n9898_;
  assign new_n9900_ = ~new_n1770_ & ~new_n9899_;
  assign new_n9901_ = new_n9892_ & ~new_n9900_;
  assign new_n9902_ = new_n1841_ & ~new_n8663_;
  assign new_n9903_ = ~new_n1841_ & new_n8663_;
  assign new_n9904_ = ~new_n9902_ & ~new_n9903_;
  assign new_n9905_ = ~new_n1831_ & ~new_n9904_;
  assign new_n9906_ = ~new_n9900_ & ~new_n9905_;
  assign new_n9907_ = ~new_n9901_ & ~new_n9906_;
  assign new_n9908_ = new_n9896_ & new_n9907_;
  assign new_n9909_ = ~new_n9896_ & ~new_n9907_;
  assign new_n9910_ = ~new_n9908_ & ~new_n9909_;
  assign new_n9911_ = ~new_n9892_ & ~new_n9910_;
  assign new_n9912_ = ~new_n9881_ & new_n9911_;
  assign new_n9913_ = new_n9881_ & ~new_n9911_;
  assign new_n9914_ = ~new_n9912_ & ~new_n9913_;
  assign new_n9915_ = new_n1910_ & ~new_n8679_;
  assign new_n9916_ = ~new_n1910_ & new_n8679_;
  assign new_n9917_ = ~new_n9915_ & ~new_n9916_;
  assign new_n9918_ = ~new_n1900_ & ~new_n9917_;
  assign new_n9919_ = new_n1970_ & ~new_n8686_;
  assign new_n9920_ = ~new_n1970_ & new_n8686_;
  assign new_n9921_ = ~new_n9919_ & ~new_n9920_;
  assign new_n9922_ = ~new_n1960_ & ~new_n9921_;
  assign new_n9923_ = ~new_n9918_ & new_n9922_;
  assign new_n9924_ = new_n9918_ & ~new_n9922_;
  assign new_n9925_ = ~new_n9923_ & ~new_n9924_;
  assign new_n9926_ = new_n2033_ & ~new_n8696_;
  assign new_n9927_ = ~new_n2033_ & new_n8696_;
  assign new_n9928_ = ~new_n9926_ & ~new_n9927_;
  assign new_n9929_ = ~new_n2023_ & ~new_n9928_;
  assign new_n9930_ = new_n2093_ & ~new_n8703_;
  assign new_n9931_ = ~new_n2093_ & new_n8703_;
  assign new_n9932_ = ~new_n9930_ & ~new_n9931_;
  assign new_n9933_ = ~new_n2083_ & ~new_n9932_;
  assign new_n9934_ = new_n9925_ & ~new_n9933_;
  assign new_n9935_ = new_n2154_ & ~new_n8711_;
  assign new_n9936_ = ~new_n2154_ & new_n8711_;
  assign new_n9937_ = ~new_n9935_ & ~new_n9936_;
  assign new_n9938_ = ~new_n2144_ & ~new_n9937_;
  assign new_n9939_ = ~new_n9933_ & ~new_n9938_;
  assign new_n9940_ = ~new_n9934_ & ~new_n9939_;
  assign new_n9941_ = new_n9929_ & new_n9940_;
  assign new_n9942_ = ~new_n9929_ & ~new_n9940_;
  assign new_n9943_ = ~new_n9941_ & ~new_n9942_;
  assign new_n9944_ = ~new_n9925_ & ~new_n9943_;
  assign new_n9945_ = new_n2220_ & ~new_n8724_;
  assign new_n9946_ = ~new_n2220_ & new_n8724_;
  assign new_n9947_ = ~new_n9945_ & ~new_n9946_;
  assign new_n9948_ = ~new_n2210_ & ~new_n9947_;
  assign new_n9949_ = new_n2280_ & ~new_n8731_;
  assign new_n9950_ = ~new_n2280_ & new_n8731_;
  assign new_n9951_ = ~new_n9949_ & ~new_n9950_;
  assign new_n9952_ = ~new_n2270_ & ~new_n9951_;
  assign new_n9953_ = ~new_n9948_ & new_n9952_;
  assign new_n9954_ = new_n9948_ & ~new_n9952_;
  assign new_n9955_ = ~new_n9953_ & ~new_n9954_;
  assign new_n9956_ = new_n2343_ & ~new_n8741_;
  assign new_n9957_ = ~new_n2343_ & new_n8741_;
  assign new_n9958_ = ~new_n9956_ & ~new_n9957_;
  assign new_n9959_ = ~new_n2333_ & ~new_n9958_;
  assign new_n9960_ = new_n2403_ & ~new_n8748_;
  assign new_n9961_ = ~new_n2403_ & new_n8748_;
  assign new_n9962_ = ~new_n9960_ & ~new_n9961_;
  assign new_n9963_ = ~new_n2393_ & ~new_n9962_;
  assign new_n9964_ = new_n9955_ & ~new_n9963_;
  assign new_n9965_ = new_n2464_ & ~new_n8756_;
  assign new_n9966_ = ~new_n2464_ & new_n8756_;
  assign new_n9967_ = ~new_n9965_ & ~new_n9966_;
  assign new_n9968_ = ~new_n2454_ & ~new_n9967_;
  assign new_n9969_ = ~new_n9963_ & ~new_n9968_;
  assign new_n9970_ = ~new_n9964_ & ~new_n9969_;
  assign new_n9971_ = new_n9959_ & new_n9970_;
  assign new_n9972_ = ~new_n9959_ & ~new_n9970_;
  assign new_n9973_ = ~new_n9971_ & ~new_n9972_;
  assign new_n9974_ = ~new_n9955_ & ~new_n9973_;
  assign new_n9975_ = new_n9914_ & ~new_n9974_;
  assign new_n9976_ = new_n2531_ & ~new_n8770_;
  assign new_n9977_ = ~new_n2531_ & new_n8770_;
  assign new_n9978_ = ~new_n9976_ & ~new_n9977_;
  assign new_n9979_ = ~new_n2521_ & ~new_n9978_;
  assign new_n9980_ = new_n2591_ & ~new_n8777_;
  assign new_n9981_ = ~new_n2591_ & new_n8777_;
  assign new_n9982_ = ~new_n9980_ & ~new_n9981_;
  assign new_n9983_ = ~new_n2581_ & ~new_n9982_;
  assign new_n9984_ = ~new_n9979_ & new_n9983_;
  assign new_n9985_ = new_n9979_ & ~new_n9983_;
  assign new_n9986_ = ~new_n9984_ & ~new_n9985_;
  assign new_n9987_ = new_n2654_ & ~new_n8787_;
  assign new_n9988_ = ~new_n2654_ & new_n8787_;
  assign new_n9989_ = ~new_n9987_ & ~new_n9988_;
  assign new_n9990_ = ~new_n2644_ & ~new_n9989_;
  assign new_n9991_ = new_n2714_ & ~new_n8794_;
  assign new_n9992_ = ~new_n2714_ & new_n8794_;
  assign new_n9993_ = ~new_n9991_ & ~new_n9992_;
  assign new_n9994_ = ~new_n2704_ & ~new_n9993_;
  assign new_n9995_ = new_n9986_ & ~new_n9994_;
  assign new_n9996_ = new_n2775_ & ~new_n8802_;
  assign new_n9997_ = ~new_n2775_ & new_n8802_;
  assign new_n9998_ = ~new_n9996_ & ~new_n9997_;
  assign new_n9999_ = ~new_n2765_ & ~new_n9998_;
  assign new_n10000_ = ~new_n9994_ & ~new_n9999_;
  assign new_n10001_ = ~new_n9995_ & ~new_n10000_;
  assign new_n10002_ = new_n9990_ & new_n10001_;
  assign new_n10003_ = ~new_n9990_ & ~new_n10001_;
  assign new_n10004_ = ~new_n10002_ & ~new_n10003_;
  assign new_n10005_ = ~new_n9986_ & ~new_n10004_;
  assign new_n10006_ = ~new_n9974_ & ~new_n10005_;
  assign new_n10007_ = ~new_n9975_ & ~new_n10006_;
  assign new_n10008_ = new_n9944_ & new_n10007_;
  assign new_n10009_ = ~new_n9944_ & ~new_n10007_;
  assign new_n10010_ = ~new_n10008_ & ~new_n10009_;
  assign A6247 = ~new_n9914_ & ~new_n10010_;
  assign new_n10012_ = ~new_n9911_ & ~new_n10008_;
  assign A6246 = ~new_n9914_ & ~new_n10012_;
  assign new_n10014_ = new_n9911_ & new_n9944_;
  assign new_n10015_ = ~new_n9914_ & ~new_n10014_;
  assign new_n10016_ = new_n9914_ & ~new_n10015_;
  assign new_n10017_ = new_n9914_ & new_n10014_;
  assign new_n10018_ = new_n10016_ & ~new_n10017_;
  assign new_n10019_ = new_n9944_ & ~new_n10018_;
  assign A6245 = new_n10007_ | new_n10019_;
  assign new_n10021_ = new_n9974_ & new_n10005_;
  assign new_n10022_ = ~new_n10006_ & ~new_n10021_;
  assign new_n10023_ = ~new_n9914_ & ~new_n9974_;
  assign new_n10024_ = new_n9914_ & new_n9974_;
  assign new_n10025_ = ~new_n10023_ & ~new_n10024_;
  assign new_n10026_ = new_n10022_ & ~new_n10025_;
  assign A6244 = new_n10019_ | new_n10026_;
  assign new_n10028_ = new_n9944_ & ~new_n10026_;
  assign new_n10029_ = ~new_n9944_ & new_n10026_;
  assign new_n10030_ = ~new_n10028_ & ~new_n10029_;
  assign A6243 = ~new_n9914_ & ~new_n10030_;
  assign new_n10032_ = new_n2848_ & ~new_n8841_;
  assign new_n10033_ = ~new_n2848_ & new_n8841_;
  assign new_n10034_ = ~new_n10032_ & ~new_n10033_;
  assign new_n10035_ = ~new_n2846_ & ~new_n10034_;
  assign new_n10036_ = new_n2868_ & ~new_n8848_;
  assign new_n10037_ = ~new_n2868_ & new_n8848_;
  assign new_n10038_ = ~new_n10036_ & ~new_n10037_;
  assign new_n10039_ = ~new_n2866_ & ~new_n10038_;
  assign new_n10040_ = ~new_n10035_ & new_n10039_;
  assign new_n10041_ = new_n10035_ & ~new_n10039_;
  assign new_n10042_ = ~new_n10040_ & ~new_n10041_;
  assign new_n10043_ = new_n2891_ & ~new_n8858_;
  assign new_n10044_ = ~new_n2891_ & new_n8858_;
  assign new_n10045_ = ~new_n10043_ & ~new_n10044_;
  assign new_n10046_ = ~new_n2889_ & ~new_n10045_;
  assign new_n10047_ = new_n2911_ & ~new_n8865_;
  assign new_n10048_ = ~new_n2911_ & new_n8865_;
  assign new_n10049_ = ~new_n10047_ & ~new_n10048_;
  assign new_n10050_ = ~new_n2909_ & ~new_n10049_;
  assign new_n10051_ = new_n10042_ & ~new_n10050_;
  assign new_n10052_ = new_n2932_ & ~new_n8873_;
  assign new_n10053_ = ~new_n2932_ & new_n8873_;
  assign new_n10054_ = ~new_n10052_ & ~new_n10053_;
  assign new_n10055_ = ~new_n2930_ & ~new_n10054_;
  assign new_n10056_ = ~new_n10050_ & ~new_n10055_;
  assign new_n10057_ = ~new_n10051_ & ~new_n10056_;
  assign new_n10058_ = new_n10046_ & new_n10057_;
  assign new_n10059_ = ~new_n10046_ & ~new_n10057_;
  assign new_n10060_ = ~new_n10058_ & ~new_n10059_;
  assign new_n10061_ = ~new_n10042_ & ~new_n10060_;
  assign new_n10062_ = new_n2958_ & ~new_n8886_;
  assign new_n10063_ = ~new_n2958_ & new_n8886_;
  assign new_n10064_ = ~new_n10062_ & ~new_n10063_;
  assign new_n10065_ = ~new_n2956_ & ~new_n10064_;
  assign new_n10066_ = new_n2978_ & ~new_n8893_;
  assign new_n10067_ = ~new_n2978_ & new_n8893_;
  assign new_n10068_ = ~new_n10066_ & ~new_n10067_;
  assign new_n10069_ = ~new_n2976_ & ~new_n10068_;
  assign new_n10070_ = ~new_n10065_ & new_n10069_;
  assign new_n10071_ = new_n10065_ & ~new_n10069_;
  assign new_n10072_ = ~new_n10070_ & ~new_n10071_;
  assign new_n10073_ = new_n3001_ & ~new_n8903_;
  assign new_n10074_ = ~new_n3001_ & new_n8903_;
  assign new_n10075_ = ~new_n10073_ & ~new_n10074_;
  assign new_n10076_ = ~new_n2999_ & ~new_n10075_;
  assign new_n10077_ = new_n3021_ & ~new_n8910_;
  assign new_n10078_ = ~new_n3021_ & new_n8910_;
  assign new_n10079_ = ~new_n10077_ & ~new_n10078_;
  assign new_n10080_ = ~new_n3019_ & ~new_n10079_;
  assign new_n10081_ = new_n10072_ & ~new_n10080_;
  assign new_n10082_ = new_n3042_ & ~new_n8918_;
  assign new_n10083_ = ~new_n3042_ & new_n8918_;
  assign new_n10084_ = ~new_n10082_ & ~new_n10083_;
  assign new_n10085_ = ~new_n3040_ & ~new_n10084_;
  assign new_n10086_ = ~new_n10080_ & ~new_n10085_;
  assign new_n10087_ = ~new_n10081_ & ~new_n10086_;
  assign new_n10088_ = new_n10076_ & new_n10087_;
  assign new_n10089_ = ~new_n10076_ & ~new_n10087_;
  assign new_n10090_ = ~new_n10088_ & ~new_n10089_;
  assign new_n10091_ = ~new_n10072_ & ~new_n10090_;
  assign new_n10092_ = ~new_n10061_ & new_n10091_;
  assign new_n10093_ = new_n10061_ & ~new_n10091_;
  assign new_n10094_ = ~new_n10092_ & ~new_n10093_;
  assign new_n10095_ = new_n3071_ & ~new_n8934_;
  assign new_n10096_ = ~new_n3071_ & new_n8934_;
  assign new_n10097_ = ~new_n10095_ & ~new_n10096_;
  assign new_n10098_ = ~new_n3069_ & ~new_n10097_;
  assign new_n10099_ = new_n3091_ & ~new_n8941_;
  assign new_n10100_ = ~new_n3091_ & new_n8941_;
  assign new_n10101_ = ~new_n10099_ & ~new_n10100_;
  assign new_n10102_ = ~new_n3089_ & ~new_n10101_;
  assign new_n10103_ = ~new_n10098_ & new_n10102_;
  assign new_n10104_ = new_n10098_ & ~new_n10102_;
  assign new_n10105_ = ~new_n10103_ & ~new_n10104_;
  assign new_n10106_ = new_n3114_ & ~new_n8951_;
  assign new_n10107_ = ~new_n3114_ & new_n8951_;
  assign new_n10108_ = ~new_n10106_ & ~new_n10107_;
  assign new_n10109_ = ~new_n3112_ & ~new_n10108_;
  assign new_n10110_ = new_n3134_ & ~new_n8958_;
  assign new_n10111_ = ~new_n3134_ & new_n8958_;
  assign new_n10112_ = ~new_n10110_ & ~new_n10111_;
  assign new_n10113_ = ~new_n3132_ & ~new_n10112_;
  assign new_n10114_ = new_n10105_ & ~new_n10113_;
  assign new_n10115_ = new_n3155_ & ~new_n8966_;
  assign new_n10116_ = ~new_n3155_ & new_n8966_;
  assign new_n10117_ = ~new_n10115_ & ~new_n10116_;
  assign new_n10118_ = ~new_n3153_ & ~new_n10117_;
  assign new_n10119_ = ~new_n10113_ & ~new_n10118_;
  assign new_n10120_ = ~new_n10114_ & ~new_n10119_;
  assign new_n10121_ = new_n10109_ & new_n10120_;
  assign new_n10122_ = ~new_n10109_ & ~new_n10120_;
  assign new_n10123_ = ~new_n10121_ & ~new_n10122_;
  assign new_n10124_ = ~new_n10105_ & ~new_n10123_;
  assign new_n10125_ = new_n3181_ & ~new_n8979_;
  assign new_n10126_ = ~new_n3181_ & new_n8979_;
  assign new_n10127_ = ~new_n10125_ & ~new_n10126_;
  assign new_n10128_ = ~new_n3179_ & ~new_n10127_;
  assign new_n10129_ = new_n3201_ & ~new_n8986_;
  assign new_n10130_ = ~new_n3201_ & new_n8986_;
  assign new_n10131_ = ~new_n10129_ & ~new_n10130_;
  assign new_n10132_ = ~new_n3199_ & ~new_n10131_;
  assign new_n10133_ = ~new_n10128_ & new_n10132_;
  assign new_n10134_ = new_n10128_ & ~new_n10132_;
  assign new_n10135_ = ~new_n10133_ & ~new_n10134_;
  assign new_n10136_ = new_n3224_ & ~new_n8996_;
  assign new_n10137_ = ~new_n3224_ & new_n8996_;
  assign new_n10138_ = ~new_n10136_ & ~new_n10137_;
  assign new_n10139_ = ~new_n3222_ & ~new_n10138_;
  assign new_n10140_ = new_n3244_ & ~new_n9003_;
  assign new_n10141_ = ~new_n3244_ & new_n9003_;
  assign new_n10142_ = ~new_n10140_ & ~new_n10141_;
  assign new_n10143_ = ~new_n3242_ & ~new_n10142_;
  assign new_n10144_ = new_n10135_ & ~new_n10143_;
  assign new_n10145_ = new_n3265_ & ~new_n9011_;
  assign new_n10146_ = ~new_n3265_ & new_n9011_;
  assign new_n10147_ = ~new_n10145_ & ~new_n10146_;
  assign new_n10148_ = ~new_n3263_ & ~new_n10147_;
  assign new_n10149_ = ~new_n10143_ & ~new_n10148_;
  assign new_n10150_ = ~new_n10144_ & ~new_n10149_;
  assign new_n10151_ = new_n10139_ & new_n10150_;
  assign new_n10152_ = ~new_n10139_ & ~new_n10150_;
  assign new_n10153_ = ~new_n10151_ & ~new_n10152_;
  assign new_n10154_ = ~new_n10135_ & ~new_n10153_;
  assign new_n10155_ = new_n10094_ & ~new_n10154_;
  assign new_n10156_ = new_n3292_ & ~new_n9025_;
  assign new_n10157_ = ~new_n3292_ & new_n9025_;
  assign new_n10158_ = ~new_n10156_ & ~new_n10157_;
  assign new_n10159_ = ~new_n3290_ & ~new_n10158_;
  assign new_n10160_ = new_n3312_ & ~new_n9032_;
  assign new_n10161_ = ~new_n3312_ & new_n9032_;
  assign new_n10162_ = ~new_n10160_ & ~new_n10161_;
  assign new_n10163_ = ~new_n3310_ & ~new_n10162_;
  assign new_n10164_ = ~new_n10159_ & new_n10163_;
  assign new_n10165_ = new_n10159_ & ~new_n10163_;
  assign new_n10166_ = ~new_n10164_ & ~new_n10165_;
  assign new_n10167_ = new_n3335_ & ~new_n9042_;
  assign new_n10168_ = ~new_n3335_ & new_n9042_;
  assign new_n10169_ = ~new_n10167_ & ~new_n10168_;
  assign new_n10170_ = ~new_n3333_ & ~new_n10169_;
  assign new_n10171_ = new_n3355_ & ~new_n9049_;
  assign new_n10172_ = ~new_n3355_ & new_n9049_;
  assign new_n10173_ = ~new_n10171_ & ~new_n10172_;
  assign new_n10174_ = ~new_n3353_ & ~new_n10173_;
  assign new_n10175_ = new_n10166_ & ~new_n10174_;
  assign new_n10176_ = new_n3376_ & ~new_n9057_;
  assign new_n10177_ = ~new_n3376_ & new_n9057_;
  assign new_n10178_ = ~new_n10176_ & ~new_n10177_;
  assign new_n10179_ = ~new_n3374_ & ~new_n10178_;
  assign new_n10180_ = ~new_n10174_ & ~new_n10179_;
  assign new_n10181_ = ~new_n10175_ & ~new_n10180_;
  assign new_n10182_ = new_n10170_ & new_n10181_;
  assign new_n10183_ = ~new_n10170_ & ~new_n10181_;
  assign new_n10184_ = ~new_n10182_ & ~new_n10183_;
  assign new_n10185_ = ~new_n10166_ & ~new_n10184_;
  assign new_n10186_ = ~new_n10154_ & ~new_n10185_;
  assign new_n10187_ = ~new_n10155_ & ~new_n10186_;
  assign new_n10188_ = new_n10124_ & new_n10187_;
  assign new_n10189_ = ~new_n10124_ & ~new_n10187_;
  assign new_n10190_ = ~new_n10188_ & ~new_n10189_;
  assign A6214 = ~new_n10094_ & ~new_n10190_;
  assign new_n10192_ = ~new_n10091_ & ~new_n10188_;
  assign A6213 = ~new_n10094_ & ~new_n10192_;
  assign new_n10194_ = new_n10091_ & new_n10124_;
  assign new_n10195_ = ~new_n10094_ & ~new_n10194_;
  assign new_n10196_ = new_n10094_ & ~new_n10195_;
  assign new_n10197_ = new_n10094_ & new_n10194_;
  assign new_n10198_ = new_n10196_ & ~new_n10197_;
  assign new_n10199_ = new_n10124_ & ~new_n10198_;
  assign A6212 = new_n10187_ | new_n10199_;
  assign new_n10201_ = new_n10154_ & new_n10185_;
  assign new_n10202_ = ~new_n10186_ & ~new_n10201_;
  assign new_n10203_ = ~new_n10094_ & ~new_n10154_;
  assign new_n10204_ = new_n10094_ & new_n10154_;
  assign new_n10205_ = ~new_n10203_ & ~new_n10204_;
  assign new_n10206_ = new_n10202_ & ~new_n10205_;
  assign A6211 = new_n10199_ | new_n10206_;
  assign new_n10208_ = new_n10124_ & ~new_n10206_;
  assign new_n10209_ = ~new_n10124_ & new_n10206_;
  assign new_n10210_ = ~new_n10208_ & ~new_n10209_;
  assign A6210 = ~new_n10094_ & ~new_n10210_;
  assign new_n10212_ = ~new_n3439_ & ~new_n9096_;
  assign new_n10213_ = new_n3439_ & new_n9096_;
  assign new_n10214_ = ~new_n10212_ & ~new_n10213_;
  assign new_n10215_ = ~new_n3432_ & ~new_n10214_;
  assign new_n10216_ = ~new_n3484_ & ~new_n9103_;
  assign new_n10217_ = new_n3484_ & new_n9103_;
  assign new_n10218_ = ~new_n10216_ & ~new_n10217_;
  assign new_n10219_ = ~new_n3477_ & ~new_n10218_;
  assign new_n10220_ = ~new_n10215_ & new_n10219_;
  assign new_n10221_ = new_n10215_ & ~new_n10219_;
  assign new_n10222_ = ~new_n10220_ & ~new_n10221_;
  assign new_n10223_ = ~new_n3532_ & ~new_n9113_;
  assign new_n10224_ = new_n3532_ & new_n9113_;
  assign new_n10225_ = ~new_n10223_ & ~new_n10224_;
  assign new_n10226_ = ~new_n3525_ & ~new_n10225_;
  assign new_n10227_ = ~new_n3577_ & ~new_n9120_;
  assign new_n10228_ = new_n3577_ & new_n9120_;
  assign new_n10229_ = ~new_n10227_ & ~new_n10228_;
  assign new_n10230_ = ~new_n3570_ & ~new_n10229_;
  assign new_n10231_ = new_n10222_ & ~new_n10230_;
  assign new_n10232_ = ~new_n3623_ & ~new_n9128_;
  assign new_n10233_ = new_n3623_ & new_n9128_;
  assign new_n10234_ = ~new_n10232_ & ~new_n10233_;
  assign new_n10235_ = ~new_n3616_ & ~new_n10234_;
  assign new_n10236_ = ~new_n10230_ & ~new_n10235_;
  assign new_n10237_ = ~new_n10231_ & ~new_n10236_;
  assign new_n10238_ = new_n10226_ & new_n10237_;
  assign new_n10239_ = ~new_n10226_ & ~new_n10237_;
  assign new_n10240_ = ~new_n10238_ & ~new_n10239_;
  assign new_n10241_ = ~new_n10222_ & ~new_n10240_;
  assign new_n10242_ = ~new_n3674_ & ~new_n9141_;
  assign new_n10243_ = new_n3674_ & new_n9141_;
  assign new_n10244_ = ~new_n10242_ & ~new_n10243_;
  assign new_n10245_ = ~new_n3667_ & ~new_n10244_;
  assign new_n10246_ = ~new_n3719_ & ~new_n9148_;
  assign new_n10247_ = new_n3719_ & new_n9148_;
  assign new_n10248_ = ~new_n10246_ & ~new_n10247_;
  assign new_n10249_ = ~new_n3712_ & ~new_n10248_;
  assign new_n10250_ = ~new_n10245_ & new_n10249_;
  assign new_n10251_ = new_n10245_ & ~new_n10249_;
  assign new_n10252_ = ~new_n10250_ & ~new_n10251_;
  assign new_n10253_ = ~new_n3767_ & ~new_n9158_;
  assign new_n10254_ = new_n3767_ & new_n9158_;
  assign new_n10255_ = ~new_n10253_ & ~new_n10254_;
  assign new_n10256_ = ~new_n3760_ & ~new_n10255_;
  assign new_n10257_ = ~new_n3812_ & ~new_n9165_;
  assign new_n10258_ = new_n3812_ & new_n9165_;
  assign new_n10259_ = ~new_n10257_ & ~new_n10258_;
  assign new_n10260_ = ~new_n3805_ & ~new_n10259_;
  assign new_n10261_ = new_n10252_ & ~new_n10260_;
  assign new_n10262_ = ~new_n3858_ & ~new_n9173_;
  assign new_n10263_ = new_n3858_ & new_n9173_;
  assign new_n10264_ = ~new_n10262_ & ~new_n10263_;
  assign new_n10265_ = ~new_n3851_ & ~new_n10264_;
  assign new_n10266_ = ~new_n10260_ & ~new_n10265_;
  assign new_n10267_ = ~new_n10261_ & ~new_n10266_;
  assign new_n10268_ = new_n10256_ & new_n10267_;
  assign new_n10269_ = ~new_n10256_ & ~new_n10267_;
  assign new_n10270_ = ~new_n10268_ & ~new_n10269_;
  assign new_n10271_ = ~new_n10252_ & ~new_n10270_;
  assign new_n10272_ = ~new_n10241_ & new_n10271_;
  assign new_n10273_ = new_n10241_ & ~new_n10271_;
  assign new_n10274_ = ~new_n10272_ & ~new_n10273_;
  assign new_n10275_ = ~new_n3912_ & ~new_n9189_;
  assign new_n10276_ = new_n3912_ & new_n9189_;
  assign new_n10277_ = ~new_n10275_ & ~new_n10276_;
  assign new_n10278_ = ~new_n3905_ & ~new_n10277_;
  assign new_n10279_ = ~new_n3957_ & ~new_n9196_;
  assign new_n10280_ = new_n3957_ & new_n9196_;
  assign new_n10281_ = ~new_n10279_ & ~new_n10280_;
  assign new_n10282_ = ~new_n3950_ & ~new_n10281_;
  assign new_n10283_ = ~new_n10278_ & new_n10282_;
  assign new_n10284_ = new_n10278_ & ~new_n10282_;
  assign new_n10285_ = ~new_n10283_ & ~new_n10284_;
  assign new_n10286_ = ~new_n4005_ & ~new_n9206_;
  assign new_n10287_ = new_n4005_ & new_n9206_;
  assign new_n10288_ = ~new_n10286_ & ~new_n10287_;
  assign new_n10289_ = ~new_n3998_ & ~new_n10288_;
  assign new_n10290_ = ~new_n4050_ & ~new_n9213_;
  assign new_n10291_ = new_n4050_ & new_n9213_;
  assign new_n10292_ = ~new_n10290_ & ~new_n10291_;
  assign new_n10293_ = ~new_n4043_ & ~new_n10292_;
  assign new_n10294_ = new_n10285_ & ~new_n10293_;
  assign new_n10295_ = ~new_n4096_ & ~new_n9221_;
  assign new_n10296_ = new_n4096_ & new_n9221_;
  assign new_n10297_ = ~new_n10295_ & ~new_n10296_;
  assign new_n10298_ = ~new_n4089_ & ~new_n10297_;
  assign new_n10299_ = ~new_n10293_ & ~new_n10298_;
  assign new_n10300_ = ~new_n10294_ & ~new_n10299_;
  assign new_n10301_ = new_n10289_ & new_n10300_;
  assign new_n10302_ = ~new_n10289_ & ~new_n10300_;
  assign new_n10303_ = ~new_n10301_ & ~new_n10302_;
  assign new_n10304_ = ~new_n10285_ & ~new_n10303_;
  assign new_n10305_ = ~new_n4147_ & ~new_n9234_;
  assign new_n10306_ = new_n4147_ & new_n9234_;
  assign new_n10307_ = ~new_n10305_ & ~new_n10306_;
  assign new_n10308_ = ~new_n4140_ & ~new_n10307_;
  assign new_n10309_ = ~new_n4192_ & ~new_n9241_;
  assign new_n10310_ = new_n4192_ & new_n9241_;
  assign new_n10311_ = ~new_n10309_ & ~new_n10310_;
  assign new_n10312_ = ~new_n4185_ & ~new_n10311_;
  assign new_n10313_ = ~new_n10308_ & new_n10312_;
  assign new_n10314_ = new_n10308_ & ~new_n10312_;
  assign new_n10315_ = ~new_n10313_ & ~new_n10314_;
  assign new_n10316_ = ~new_n4240_ & ~new_n9251_;
  assign new_n10317_ = new_n4240_ & new_n9251_;
  assign new_n10318_ = ~new_n10316_ & ~new_n10317_;
  assign new_n10319_ = ~new_n4233_ & ~new_n10318_;
  assign new_n10320_ = ~new_n4285_ & ~new_n9258_;
  assign new_n10321_ = new_n4285_ & new_n9258_;
  assign new_n10322_ = ~new_n10320_ & ~new_n10321_;
  assign new_n10323_ = ~new_n4278_ & ~new_n10322_;
  assign new_n10324_ = new_n10315_ & ~new_n10323_;
  assign new_n10325_ = ~new_n4331_ & ~new_n9266_;
  assign new_n10326_ = new_n4331_ & new_n9266_;
  assign new_n10327_ = ~new_n10325_ & ~new_n10326_;
  assign new_n10328_ = ~new_n4324_ & ~new_n10327_;
  assign new_n10329_ = ~new_n10323_ & ~new_n10328_;
  assign new_n10330_ = ~new_n10324_ & ~new_n10329_;
  assign new_n10331_ = new_n10319_ & new_n10330_;
  assign new_n10332_ = ~new_n10319_ & ~new_n10330_;
  assign new_n10333_ = ~new_n10331_ & ~new_n10332_;
  assign new_n10334_ = ~new_n10315_ & ~new_n10333_;
  assign new_n10335_ = new_n10274_ & ~new_n10334_;
  assign new_n10336_ = ~new_n4383_ & ~new_n9280_;
  assign new_n10337_ = new_n4383_ & new_n9280_;
  assign new_n10338_ = ~new_n10336_ & ~new_n10337_;
  assign new_n10339_ = ~new_n4376_ & ~new_n10338_;
  assign new_n10340_ = ~new_n4428_ & ~new_n9287_;
  assign new_n10341_ = new_n4428_ & new_n9287_;
  assign new_n10342_ = ~new_n10340_ & ~new_n10341_;
  assign new_n10343_ = ~new_n4421_ & ~new_n10342_;
  assign new_n10344_ = ~new_n10339_ & new_n10343_;
  assign new_n10345_ = new_n10339_ & ~new_n10343_;
  assign new_n10346_ = ~new_n10344_ & ~new_n10345_;
  assign new_n10347_ = ~new_n4476_ & ~new_n9297_;
  assign new_n10348_ = new_n4476_ & new_n9297_;
  assign new_n10349_ = ~new_n10347_ & ~new_n10348_;
  assign new_n10350_ = ~new_n4469_ & ~new_n10349_;
  assign new_n10351_ = ~new_n4521_ & ~new_n9304_;
  assign new_n10352_ = new_n4521_ & new_n9304_;
  assign new_n10353_ = ~new_n10351_ & ~new_n10352_;
  assign new_n10354_ = ~new_n4514_ & ~new_n10353_;
  assign new_n10355_ = new_n10346_ & ~new_n10354_;
  assign new_n10356_ = ~new_n4567_ & ~new_n9312_;
  assign new_n10357_ = new_n4567_ & new_n9312_;
  assign new_n10358_ = ~new_n10356_ & ~new_n10357_;
  assign new_n10359_ = ~new_n4560_ & ~new_n10358_;
  assign new_n10360_ = ~new_n10354_ & ~new_n10359_;
  assign new_n10361_ = ~new_n10355_ & ~new_n10360_;
  assign new_n10362_ = new_n10350_ & new_n10361_;
  assign new_n10363_ = ~new_n10350_ & ~new_n10361_;
  assign new_n10364_ = ~new_n10362_ & ~new_n10363_;
  assign new_n10365_ = ~new_n10346_ & ~new_n10364_;
  assign new_n10366_ = ~new_n10334_ & ~new_n10365_;
  assign new_n10367_ = ~new_n10335_ & ~new_n10366_;
  assign new_n10368_ = new_n10304_ & new_n10367_;
  assign new_n10369_ = ~new_n10304_ & ~new_n10367_;
  assign new_n10370_ = ~new_n10368_ & ~new_n10369_;
  assign A6181 = ~new_n10274_ & ~new_n10370_;
  assign new_n10372_ = ~new_n10271_ & ~new_n10368_;
  assign A6180 = ~new_n10274_ & ~new_n10372_;
  assign new_n10374_ = new_n10271_ & new_n10304_;
  assign new_n10375_ = ~new_n10274_ & ~new_n10374_;
  assign new_n10376_ = new_n10274_ & ~new_n10375_;
  assign new_n10377_ = new_n10274_ & new_n10374_;
  assign new_n10378_ = new_n10376_ & ~new_n10377_;
  assign new_n10379_ = new_n10304_ & ~new_n10378_;
  assign A6179 = new_n10367_ | new_n10379_;
  assign new_n10381_ = new_n10334_ & new_n10365_;
  assign new_n10382_ = ~new_n10366_ & ~new_n10381_;
  assign new_n10383_ = ~new_n10274_ & ~new_n10334_;
  assign new_n10384_ = new_n10274_ & new_n10334_;
  assign new_n10385_ = ~new_n10383_ & ~new_n10384_;
  assign new_n10386_ = new_n10382_ & ~new_n10385_;
  assign A6178 = new_n10379_ | new_n10386_;
  assign new_n10388_ = new_n10304_ & ~new_n10386_;
  assign new_n10389_ = ~new_n10304_ & new_n10386_;
  assign new_n10390_ = ~new_n10388_ & ~new_n10389_;
  assign A6177 = ~new_n10274_ & ~new_n10390_;
  assign new_n10392_ = ~new_n4640_ & ~new_n9351_;
  assign new_n10393_ = new_n4640_ & new_n9351_;
  assign new_n10394_ = ~new_n10392_ & ~new_n10393_;
  assign new_n10395_ = ~new_n4633_ & ~new_n10394_;
  assign new_n10396_ = ~new_n4685_ & ~new_n9358_;
  assign new_n10397_ = new_n4685_ & new_n9358_;
  assign new_n10398_ = ~new_n10396_ & ~new_n10397_;
  assign new_n10399_ = ~new_n4678_ & ~new_n10398_;
  assign new_n10400_ = ~new_n10395_ & new_n10399_;
  assign new_n10401_ = new_n10395_ & ~new_n10399_;
  assign new_n10402_ = ~new_n10400_ & ~new_n10401_;
  assign new_n10403_ = ~new_n4733_ & ~new_n9368_;
  assign new_n10404_ = new_n4733_ & new_n9368_;
  assign new_n10405_ = ~new_n10403_ & ~new_n10404_;
  assign new_n10406_ = ~new_n4726_ & ~new_n10405_;
  assign new_n10407_ = ~new_n4778_ & ~new_n9375_;
  assign new_n10408_ = new_n4778_ & new_n9375_;
  assign new_n10409_ = ~new_n10407_ & ~new_n10408_;
  assign new_n10410_ = ~new_n4771_ & ~new_n10409_;
  assign new_n10411_ = new_n10402_ & ~new_n10410_;
  assign new_n10412_ = ~new_n4824_ & ~new_n9383_;
  assign new_n10413_ = new_n4824_ & new_n9383_;
  assign new_n10414_ = ~new_n10412_ & ~new_n10413_;
  assign new_n10415_ = ~new_n4817_ & ~new_n10414_;
  assign new_n10416_ = ~new_n10410_ & ~new_n10415_;
  assign new_n10417_ = ~new_n10411_ & ~new_n10416_;
  assign new_n10418_ = new_n10406_ & new_n10417_;
  assign new_n10419_ = ~new_n10406_ & ~new_n10417_;
  assign new_n10420_ = ~new_n10418_ & ~new_n10419_;
  assign new_n10421_ = ~new_n10402_ & ~new_n10420_;
  assign new_n10422_ = ~new_n4875_ & ~new_n9396_;
  assign new_n10423_ = new_n4875_ & new_n9396_;
  assign new_n10424_ = ~new_n10422_ & ~new_n10423_;
  assign new_n10425_ = ~new_n4868_ & ~new_n10424_;
  assign new_n10426_ = ~new_n4920_ & ~new_n9403_;
  assign new_n10427_ = new_n4920_ & new_n9403_;
  assign new_n10428_ = ~new_n10426_ & ~new_n10427_;
  assign new_n10429_ = ~new_n4913_ & ~new_n10428_;
  assign new_n10430_ = ~new_n10425_ & new_n10429_;
  assign new_n10431_ = new_n10425_ & ~new_n10429_;
  assign new_n10432_ = ~new_n10430_ & ~new_n10431_;
  assign new_n10433_ = ~new_n4968_ & ~new_n9413_;
  assign new_n10434_ = new_n4968_ & new_n9413_;
  assign new_n10435_ = ~new_n10433_ & ~new_n10434_;
  assign new_n10436_ = ~new_n4961_ & ~new_n10435_;
  assign new_n10437_ = ~new_n5013_ & ~new_n9420_;
  assign new_n10438_ = new_n5013_ & new_n9420_;
  assign new_n10439_ = ~new_n10437_ & ~new_n10438_;
  assign new_n10440_ = ~new_n5006_ & ~new_n10439_;
  assign new_n10441_ = new_n10432_ & ~new_n10440_;
  assign new_n10442_ = ~new_n5059_ & ~new_n9428_;
  assign new_n10443_ = new_n5059_ & new_n9428_;
  assign new_n10444_ = ~new_n10442_ & ~new_n10443_;
  assign new_n10445_ = ~new_n5052_ & ~new_n10444_;
  assign new_n10446_ = ~new_n10440_ & ~new_n10445_;
  assign new_n10447_ = ~new_n10441_ & ~new_n10446_;
  assign new_n10448_ = new_n10436_ & new_n10447_;
  assign new_n10449_ = ~new_n10436_ & ~new_n10447_;
  assign new_n10450_ = ~new_n10448_ & ~new_n10449_;
  assign new_n10451_ = ~new_n10432_ & ~new_n10450_;
  assign new_n10452_ = ~new_n10421_ & new_n10451_;
  assign new_n10453_ = new_n10421_ & ~new_n10451_;
  assign new_n10454_ = ~new_n10452_ & ~new_n10453_;
  assign new_n10455_ = ~new_n5113_ & ~new_n9444_;
  assign new_n10456_ = new_n5113_ & new_n9444_;
  assign new_n10457_ = ~new_n10455_ & ~new_n10456_;
  assign new_n10458_ = ~new_n5106_ & ~new_n10457_;
  assign new_n10459_ = ~new_n5158_ & ~new_n9451_;
  assign new_n10460_ = new_n5158_ & new_n9451_;
  assign new_n10461_ = ~new_n10459_ & ~new_n10460_;
  assign new_n10462_ = ~new_n5151_ & ~new_n10461_;
  assign new_n10463_ = ~new_n10458_ & new_n10462_;
  assign new_n10464_ = new_n10458_ & ~new_n10462_;
  assign new_n10465_ = ~new_n10463_ & ~new_n10464_;
  assign new_n10466_ = ~new_n5206_ & ~new_n9461_;
  assign new_n10467_ = new_n5206_ & new_n9461_;
  assign new_n10468_ = ~new_n10466_ & ~new_n10467_;
  assign new_n10469_ = ~new_n5199_ & ~new_n10468_;
  assign new_n10470_ = ~new_n5251_ & ~new_n9468_;
  assign new_n10471_ = new_n5251_ & new_n9468_;
  assign new_n10472_ = ~new_n10470_ & ~new_n10471_;
  assign new_n10473_ = ~new_n5244_ & ~new_n10472_;
  assign new_n10474_ = new_n10465_ & ~new_n10473_;
  assign new_n10475_ = ~new_n5297_ & ~new_n9476_;
  assign new_n10476_ = new_n5297_ & new_n9476_;
  assign new_n10477_ = ~new_n10475_ & ~new_n10476_;
  assign new_n10478_ = ~new_n5290_ & ~new_n10477_;
  assign new_n10479_ = ~new_n10473_ & ~new_n10478_;
  assign new_n10480_ = ~new_n10474_ & ~new_n10479_;
  assign new_n10481_ = new_n10469_ & new_n10480_;
  assign new_n10482_ = ~new_n10469_ & ~new_n10480_;
  assign new_n10483_ = ~new_n10481_ & ~new_n10482_;
  assign new_n10484_ = ~new_n10465_ & ~new_n10483_;
  assign new_n10485_ = ~new_n5348_ & ~new_n9489_;
  assign new_n10486_ = new_n5348_ & new_n9489_;
  assign new_n10487_ = ~new_n10485_ & ~new_n10486_;
  assign new_n10488_ = ~new_n5341_ & ~new_n10487_;
  assign new_n10489_ = ~new_n5393_ & ~new_n9496_;
  assign new_n10490_ = new_n5393_ & new_n9496_;
  assign new_n10491_ = ~new_n10489_ & ~new_n10490_;
  assign new_n10492_ = ~new_n5386_ & ~new_n10491_;
  assign new_n10493_ = ~new_n10488_ & new_n10492_;
  assign new_n10494_ = new_n10488_ & ~new_n10492_;
  assign new_n10495_ = ~new_n10493_ & ~new_n10494_;
  assign new_n10496_ = ~new_n5441_ & ~new_n9506_;
  assign new_n10497_ = new_n5441_ & new_n9506_;
  assign new_n10498_ = ~new_n10496_ & ~new_n10497_;
  assign new_n10499_ = ~new_n5434_ & ~new_n10498_;
  assign new_n10500_ = ~new_n5486_ & ~new_n9513_;
  assign new_n10501_ = new_n5486_ & new_n9513_;
  assign new_n10502_ = ~new_n10500_ & ~new_n10501_;
  assign new_n10503_ = ~new_n5479_ & ~new_n10502_;
  assign new_n10504_ = new_n10495_ & ~new_n10503_;
  assign new_n10505_ = ~new_n5532_ & ~new_n9521_;
  assign new_n10506_ = new_n5532_ & new_n9521_;
  assign new_n10507_ = ~new_n10505_ & ~new_n10506_;
  assign new_n10508_ = ~new_n5525_ & ~new_n10507_;
  assign new_n10509_ = ~new_n10503_ & ~new_n10508_;
  assign new_n10510_ = ~new_n10504_ & ~new_n10509_;
  assign new_n10511_ = new_n10499_ & new_n10510_;
  assign new_n10512_ = ~new_n10499_ & ~new_n10510_;
  assign new_n10513_ = ~new_n10511_ & ~new_n10512_;
  assign new_n10514_ = ~new_n10495_ & ~new_n10513_;
  assign new_n10515_ = new_n10454_ & ~new_n10514_;
  assign new_n10516_ = ~new_n5584_ & ~new_n9535_;
  assign new_n10517_ = new_n5584_ & new_n9535_;
  assign new_n10518_ = ~new_n10516_ & ~new_n10517_;
  assign new_n10519_ = ~new_n5577_ & ~new_n10518_;
  assign new_n10520_ = ~new_n5629_ & ~new_n9542_;
  assign new_n10521_ = new_n5629_ & new_n9542_;
  assign new_n10522_ = ~new_n10520_ & ~new_n10521_;
  assign new_n10523_ = ~new_n5622_ & ~new_n10522_;
  assign new_n10524_ = ~new_n10519_ & new_n10523_;
  assign new_n10525_ = new_n10519_ & ~new_n10523_;
  assign new_n10526_ = ~new_n10524_ & ~new_n10525_;
  assign new_n10527_ = ~new_n5677_ & ~new_n9552_;
  assign new_n10528_ = new_n5677_ & new_n9552_;
  assign new_n10529_ = ~new_n10527_ & ~new_n10528_;
  assign new_n10530_ = ~new_n5670_ & ~new_n10529_;
  assign new_n10531_ = ~new_n5722_ & ~new_n9559_;
  assign new_n10532_ = new_n5722_ & new_n9559_;
  assign new_n10533_ = ~new_n10531_ & ~new_n10532_;
  assign new_n10534_ = ~new_n5715_ & ~new_n10533_;
  assign new_n10535_ = new_n10526_ & ~new_n10534_;
  assign new_n10536_ = ~new_n5768_ & ~new_n9567_;
  assign new_n10537_ = new_n5768_ & new_n9567_;
  assign new_n10538_ = ~new_n10536_ & ~new_n10537_;
  assign new_n10539_ = ~new_n5761_ & ~new_n10538_;
  assign new_n10540_ = ~new_n10534_ & ~new_n10539_;
  assign new_n10541_ = ~new_n10535_ & ~new_n10540_;
  assign new_n10542_ = new_n10530_ & new_n10541_;
  assign new_n10543_ = ~new_n10530_ & ~new_n10541_;
  assign new_n10544_ = ~new_n10542_ & ~new_n10543_;
  assign new_n10545_ = ~new_n10526_ & ~new_n10544_;
  assign new_n10546_ = ~new_n10514_ & ~new_n10545_;
  assign new_n10547_ = ~new_n10515_ & ~new_n10546_;
  assign new_n10548_ = new_n10484_ & new_n10547_;
  assign new_n10549_ = ~new_n10484_ & ~new_n10547_;
  assign new_n10550_ = ~new_n10548_ & ~new_n10549_;
  assign A6148 = ~new_n10454_ & ~new_n10550_;
  assign new_n10552_ = ~new_n10451_ & ~new_n10548_;
  assign A6147 = ~new_n10454_ & ~new_n10552_;
  assign new_n10554_ = new_n10451_ & new_n10484_;
  assign new_n10555_ = ~new_n10454_ & ~new_n10554_;
  assign new_n10556_ = new_n10454_ & ~new_n10555_;
  assign new_n10557_ = new_n10454_ & new_n10554_;
  assign new_n10558_ = new_n10556_ & ~new_n10557_;
  assign new_n10559_ = new_n10484_ & ~new_n10558_;
  assign A6146 = new_n10547_ | new_n10559_;
  assign new_n10561_ = new_n10514_ & new_n10545_;
  assign new_n10562_ = ~new_n10546_ & ~new_n10561_;
  assign new_n10563_ = ~new_n10454_ & ~new_n10514_;
  assign new_n10564_ = new_n10454_ & new_n10514_;
  assign new_n10565_ = ~new_n10563_ & ~new_n10564_;
  assign new_n10566_ = new_n10562_ & ~new_n10565_;
  assign A6145 = new_n10559_ | new_n10566_;
  assign new_n10568_ = new_n10484_ & ~new_n10566_;
  assign new_n10569_ = ~new_n10484_ & new_n10566_;
  assign new_n10570_ = ~new_n10568_ & ~new_n10569_;
  assign A6144 = ~new_n10454_ & ~new_n10570_;
  assign new_n10572_ = new_n5869_ & ~new_n9609_;
  assign new_n10573_ = ~new_n5869_ & new_n9609_;
  assign new_n10574_ = ~new_n10572_ & ~new_n10573_;
  assign new_n10575_ = ~new_n5865_ & ~new_n10574_;
  assign new_n10576_ = ~new_n5850_ & ~new_n8331_;
  assign new_n10577_ = ~new_n9601_ & ~new_n10576_;
  assign new_n10578_ = ~new_n5842_ & ~new_n10577_;
  assign new_n10579_ = new_n10575_ & new_n10578_;
  assign new_n10580_ = ~new_n10575_ & ~new_n10578_;
  assign new_n10581_ = ~new_n10579_ & ~new_n10580_;
  assign new_n10582_ = new_n5963_ & ~new_n9634_;
  assign new_n10583_ = ~new_n5963_ & new_n9634_;
  assign new_n10584_ = ~new_n10582_ & ~new_n10583_;
  assign new_n10585_ = ~new_n5959_ & ~new_n10584_;
  assign new_n10586_ = new_n5932_ & ~new_n9626_;
  assign new_n10587_ = ~new_n5932_ & new_n9626_;
  assign new_n10588_ = ~new_n10586_ & ~new_n10587_;
  assign new_n10589_ = ~new_n5928_ & ~new_n10588_;
  assign new_n10590_ = ~new_n10585_ & new_n10589_;
  assign new_n10591_ = new_n10585_ & ~new_n10589_;
  assign new_n10592_ = ~new_n10590_ & ~new_n10591_;
  assign new_n10593_ = ~new_n10575_ & ~new_n10592_;
  assign new_n10594_ = new_n10575_ & new_n10592_;
  assign new_n10595_ = ~new_n10593_ & ~new_n10594_;
  assign new_n10596_ = new_n10581_ & ~new_n10595_;
  assign new_n10597_ = new_n5902_ & ~new_n9619_;
  assign new_n10598_ = ~new_n5902_ & new_n9619_;
  assign new_n10599_ = ~new_n10597_ & ~new_n10598_;
  assign new_n10600_ = ~new_n5898_ & ~new_n10599_;
  assign new_n10601_ = ~new_n10596_ & new_n10600_;
  assign new_n10602_ = new_n10596_ & ~new_n10600_;
  assign new_n10603_ = ~new_n10601_ & ~new_n10602_;
  assign new_n10604_ = ~new_n10592_ & ~new_n10603_;
  assign new_n10605_ = new_n5999_ & ~new_n9647_;
  assign new_n10606_ = ~new_n5999_ & new_n9647_;
  assign new_n10607_ = ~new_n10605_ & ~new_n10606_;
  assign new_n10608_ = ~new_n5995_ & ~new_n10607_;
  assign new_n10609_ = new_n6029_ & ~new_n9654_;
  assign new_n10610_ = ~new_n6029_ & new_n9654_;
  assign new_n10611_ = ~new_n10609_ & ~new_n10610_;
  assign new_n10612_ = ~new_n6025_ & ~new_n10611_;
  assign new_n10613_ = ~new_n10608_ & new_n10612_;
  assign new_n10614_ = new_n10608_ & ~new_n10612_;
  assign new_n10615_ = ~new_n10613_ & ~new_n10614_;
  assign new_n10616_ = new_n6062_ & ~new_n9664_;
  assign new_n10617_ = ~new_n6062_ & new_n9664_;
  assign new_n10618_ = ~new_n10616_ & ~new_n10617_;
  assign new_n10619_ = ~new_n6058_ & ~new_n10618_;
  assign new_n10620_ = new_n6092_ & ~new_n9671_;
  assign new_n10621_ = ~new_n6092_ & new_n9671_;
  assign new_n10622_ = ~new_n10620_ & ~new_n10621_;
  assign new_n10623_ = ~new_n6088_ & ~new_n10622_;
  assign new_n10624_ = new_n10615_ & ~new_n10623_;
  assign new_n10625_ = new_n6123_ & ~new_n9679_;
  assign new_n10626_ = ~new_n6123_ & new_n9679_;
  assign new_n10627_ = ~new_n10625_ & ~new_n10626_;
  assign new_n10628_ = ~new_n6119_ & ~new_n10627_;
  assign new_n10629_ = ~new_n10623_ & ~new_n10628_;
  assign new_n10630_ = ~new_n10624_ & ~new_n10629_;
  assign new_n10631_ = new_n10619_ & new_n10630_;
  assign new_n10632_ = ~new_n10619_ & ~new_n10630_;
  assign new_n10633_ = ~new_n10631_ & ~new_n10632_;
  assign new_n10634_ = ~new_n10615_ & ~new_n10633_;
  assign new_n10635_ = ~new_n10604_ & new_n10634_;
  assign new_n10636_ = new_n10604_ & ~new_n10634_;
  assign new_n10637_ = ~new_n10635_ & ~new_n10636_;
  assign new_n10638_ = new_n6162_ & ~new_n9695_;
  assign new_n10639_ = ~new_n6162_ & new_n9695_;
  assign new_n10640_ = ~new_n10638_ & ~new_n10639_;
  assign new_n10641_ = ~new_n6158_ & ~new_n10640_;
  assign new_n10642_ = new_n6192_ & ~new_n9702_;
  assign new_n10643_ = ~new_n6192_ & new_n9702_;
  assign new_n10644_ = ~new_n10642_ & ~new_n10643_;
  assign new_n10645_ = ~new_n6188_ & ~new_n10644_;
  assign new_n10646_ = ~new_n10641_ & new_n10645_;
  assign new_n10647_ = new_n10641_ & ~new_n10645_;
  assign new_n10648_ = ~new_n10646_ & ~new_n10647_;
  assign new_n10649_ = new_n6225_ & ~new_n9712_;
  assign new_n10650_ = ~new_n6225_ & new_n9712_;
  assign new_n10651_ = ~new_n10649_ & ~new_n10650_;
  assign new_n10652_ = ~new_n6221_ & ~new_n10651_;
  assign new_n10653_ = new_n6255_ & ~new_n9719_;
  assign new_n10654_ = ~new_n6255_ & new_n9719_;
  assign new_n10655_ = ~new_n10653_ & ~new_n10654_;
  assign new_n10656_ = ~new_n6251_ & ~new_n10655_;
  assign new_n10657_ = new_n10648_ & ~new_n10656_;
  assign new_n10658_ = new_n6286_ & ~new_n9727_;
  assign new_n10659_ = ~new_n6286_ & new_n9727_;
  assign new_n10660_ = ~new_n10658_ & ~new_n10659_;
  assign new_n10661_ = ~new_n6282_ & ~new_n10660_;
  assign new_n10662_ = ~new_n10656_ & ~new_n10661_;
  assign new_n10663_ = ~new_n10657_ & ~new_n10662_;
  assign new_n10664_ = new_n10652_ & new_n10663_;
  assign new_n10665_ = ~new_n10652_ & ~new_n10663_;
  assign new_n10666_ = ~new_n10664_ & ~new_n10665_;
  assign new_n10667_ = ~new_n10648_ & ~new_n10666_;
  assign new_n10668_ = new_n6322_ & ~new_n9740_;
  assign new_n10669_ = ~new_n6322_ & new_n9740_;
  assign new_n10670_ = ~new_n10668_ & ~new_n10669_;
  assign new_n10671_ = ~new_n6318_ & ~new_n10670_;
  assign new_n10672_ = new_n6352_ & ~new_n9747_;
  assign new_n10673_ = ~new_n6352_ & new_n9747_;
  assign new_n10674_ = ~new_n10672_ & ~new_n10673_;
  assign new_n10675_ = ~new_n6348_ & ~new_n10674_;
  assign new_n10676_ = ~new_n10671_ & new_n10675_;
  assign new_n10677_ = new_n10671_ & ~new_n10675_;
  assign new_n10678_ = ~new_n10676_ & ~new_n10677_;
  assign new_n10679_ = new_n6385_ & ~new_n9757_;
  assign new_n10680_ = ~new_n6385_ & new_n9757_;
  assign new_n10681_ = ~new_n10679_ & ~new_n10680_;
  assign new_n10682_ = ~new_n6381_ & ~new_n10681_;
  assign new_n10683_ = new_n6415_ & ~new_n9764_;
  assign new_n10684_ = ~new_n6415_ & new_n9764_;
  assign new_n10685_ = ~new_n10683_ & ~new_n10684_;
  assign new_n10686_ = ~new_n6411_ & ~new_n10685_;
  assign new_n10687_ = new_n10678_ & ~new_n10686_;
  assign new_n10688_ = new_n6446_ & ~new_n9772_;
  assign new_n10689_ = ~new_n6446_ & new_n9772_;
  assign new_n10690_ = ~new_n10688_ & ~new_n10689_;
  assign new_n10691_ = ~new_n6442_ & ~new_n10690_;
  assign new_n10692_ = ~new_n10686_ & ~new_n10691_;
  assign new_n10693_ = ~new_n10687_ & ~new_n10692_;
  assign new_n10694_ = new_n10682_ & new_n10693_;
  assign new_n10695_ = ~new_n10682_ & ~new_n10693_;
  assign new_n10696_ = ~new_n10694_ & ~new_n10695_;
  assign new_n10697_ = ~new_n10678_ & ~new_n10696_;
  assign new_n10698_ = new_n10637_ & ~new_n10697_;
  assign new_n10699_ = new_n6483_ & ~new_n9786_;
  assign new_n10700_ = ~new_n6483_ & new_n9786_;
  assign new_n10701_ = ~new_n10699_ & ~new_n10700_;
  assign new_n10702_ = ~new_n6479_ & ~new_n10701_;
  assign new_n10703_ = new_n6513_ & ~new_n9793_;
  assign new_n10704_ = ~new_n6513_ & new_n9793_;
  assign new_n10705_ = ~new_n10703_ & ~new_n10704_;
  assign new_n10706_ = ~new_n6509_ & ~new_n10705_;
  assign new_n10707_ = ~new_n10702_ & new_n10706_;
  assign new_n10708_ = new_n10702_ & ~new_n10706_;
  assign new_n10709_ = ~new_n10707_ & ~new_n10708_;
  assign new_n10710_ = new_n6546_ & ~new_n9803_;
  assign new_n10711_ = ~new_n6546_ & new_n9803_;
  assign new_n10712_ = ~new_n10710_ & ~new_n10711_;
  assign new_n10713_ = ~new_n6542_ & ~new_n10712_;
  assign new_n10714_ = new_n6576_ & ~new_n9810_;
  assign new_n10715_ = ~new_n6576_ & new_n9810_;
  assign new_n10716_ = ~new_n10714_ & ~new_n10715_;
  assign new_n10717_ = ~new_n6572_ & ~new_n10716_;
  assign new_n10718_ = new_n10709_ & ~new_n10717_;
  assign new_n10719_ = new_n6607_ & ~new_n9818_;
  assign new_n10720_ = ~new_n6607_ & new_n9818_;
  assign new_n10721_ = ~new_n10719_ & ~new_n10720_;
  assign new_n10722_ = ~new_n6603_ & ~new_n10721_;
  assign new_n10723_ = ~new_n10717_ & ~new_n10722_;
  assign new_n10724_ = ~new_n10718_ & ~new_n10723_;
  assign new_n10725_ = new_n10713_ & new_n10724_;
  assign new_n10726_ = ~new_n10713_ & ~new_n10724_;
  assign new_n10727_ = ~new_n10725_ & ~new_n10726_;
  assign new_n10728_ = ~new_n10709_ & ~new_n10727_;
  assign new_n10729_ = ~new_n10697_ & ~new_n10728_;
  assign new_n10730_ = ~new_n10698_ & ~new_n10729_;
  assign new_n10731_ = new_n10667_ & new_n10730_;
  assign new_n10732_ = ~new_n10667_ & ~new_n10730_;
  assign new_n10733_ = ~new_n10731_ & ~new_n10732_;
  assign A6115 = ~new_n10637_ & ~new_n10733_;
  assign new_n10735_ = ~new_n10634_ & ~new_n10731_;
  assign A6114 = ~new_n10637_ & ~new_n10735_;
  assign new_n10737_ = new_n10634_ & new_n10667_;
  assign new_n10738_ = ~new_n10637_ & ~new_n10737_;
  assign new_n10739_ = new_n10637_ & ~new_n10738_;
  assign new_n10740_ = new_n10637_ & new_n10737_;
  assign new_n10741_ = new_n10739_ & ~new_n10740_;
  assign new_n10742_ = new_n10667_ & ~new_n10741_;
  assign A6113 = new_n10730_ | new_n10742_;
  assign new_n10744_ = new_n10697_ & new_n10728_;
  assign new_n10745_ = ~new_n10729_ & ~new_n10744_;
  assign new_n10746_ = ~new_n10637_ & ~new_n10697_;
  assign new_n10747_ = new_n10637_ & new_n10697_;
  assign new_n10748_ = ~new_n10746_ & ~new_n10747_;
  assign new_n10749_ = new_n10745_ & ~new_n10748_;
  assign A6112 = new_n10742_ | new_n10749_;
  assign new_n10751_ = new_n10667_ & ~new_n10749_;
  assign new_n10752_ = ~new_n10667_ & new_n10749_;
  assign new_n10753_ = ~new_n10751_ & ~new_n10752_;
  assign A6111 = ~new_n10637_ & ~new_n10753_;
  assign new_n10755_ = ~new_n1374_ & ~new_n1561_;
  assign new_n10756_ = ~new_n1377_ & ~new_n10755_;
  assign new_n10757_ = ~new_n1684_ & ~new_n1871_;
  assign new_n10758_ = ~new_n1687_ & ~new_n10757_;
  assign new_n10759_ = ~new_n10756_ & new_n10758_;
  assign new_n10760_ = new_n10756_ & ~new_n10758_;
  assign new_n10761_ = ~new_n10759_ & ~new_n10760_;
  assign new_n10762_ = ~new_n1997_ & ~new_n2184_;
  assign new_n10763_ = ~new_n2000_ & ~new_n10762_;
  assign new_n10764_ = ~new_n2307_ & ~new_n2494_;
  assign new_n10765_ = ~new_n2310_ & ~new_n10764_;
  assign new_n10766_ = new_n10761_ & ~new_n10765_;
  assign new_n10767_ = ~new_n2618_ & ~new_n2805_;
  assign new_n10768_ = ~new_n2621_ & ~new_n10767_;
  assign new_n10769_ = ~new_n10765_ & ~new_n10768_;
  assign new_n10770_ = ~new_n10766_ & ~new_n10769_;
  assign new_n10771_ = new_n10763_ & new_n10770_;
  assign new_n10772_ = ~new_n10763_ & ~new_n10770_;
  assign new_n10773_ = ~new_n10771_ & ~new_n10772_;
  assign A6082 = ~new_n10761_ & ~new_n10773_;
  assign new_n10775_ = ~new_n10758_ & ~new_n10771_;
  assign A6081 = ~new_n10761_ & ~new_n10775_;
  assign new_n10777_ = new_n10758_ & new_n10763_;
  assign new_n10778_ = ~new_n10761_ & ~new_n10777_;
  assign new_n10779_ = new_n10761_ & ~new_n10778_;
  assign new_n10780_ = new_n10761_ & new_n10777_;
  assign new_n10781_ = new_n10779_ & ~new_n10780_;
  assign new_n10782_ = new_n10763_ & ~new_n10781_;
  assign A6080 = new_n10770_ | new_n10782_;
  assign new_n10784_ = new_n10765_ & new_n10768_;
  assign new_n10785_ = ~new_n10769_ & ~new_n10784_;
  assign new_n10786_ = ~new_n10761_ & ~new_n10765_;
  assign new_n10787_ = new_n10761_ & new_n10765_;
  assign new_n10788_ = ~new_n10786_ & ~new_n10787_;
  assign new_n10789_ = new_n10785_ & ~new_n10788_;
  assign A6079 = new_n10782_ | new_n10789_;
  assign new_n10791_ = new_n10763_ & ~new_n10789_;
  assign new_n10792_ = ~new_n10763_ & new_n10789_;
  assign new_n10793_ = ~new_n10791_ & ~new_n10792_;
  assign A6078 = ~new_n10761_ & ~new_n10793_;
  assign new_n10795_ = ~new_n2879_ & ~new_n2946_;
  assign new_n10796_ = ~new_n2882_ & ~new_n10795_;
  assign new_n10797_ = ~new_n2989_ & ~new_n3056_;
  assign new_n10798_ = ~new_n2992_ & ~new_n10797_;
  assign new_n10799_ = ~new_n10796_ & new_n10798_;
  assign new_n10800_ = new_n10796_ & ~new_n10798_;
  assign new_n10801_ = ~new_n10799_ & ~new_n10800_;
  assign new_n10802_ = ~new_n3102_ & ~new_n3169_;
  assign new_n10803_ = ~new_n3105_ & ~new_n10802_;
  assign new_n10804_ = ~new_n3212_ & ~new_n3279_;
  assign new_n10805_ = ~new_n3215_ & ~new_n10804_;
  assign new_n10806_ = new_n10801_ & ~new_n10805_;
  assign new_n10807_ = ~new_n3323_ & ~new_n3390_;
  assign new_n10808_ = ~new_n3326_ & ~new_n10807_;
  assign new_n10809_ = ~new_n10805_ & ~new_n10808_;
  assign new_n10810_ = ~new_n10806_ & ~new_n10809_;
  assign new_n10811_ = new_n10803_ & new_n10810_;
  assign new_n10812_ = ~new_n10803_ & ~new_n10810_;
  assign new_n10813_ = ~new_n10811_ & ~new_n10812_;
  assign A6049 = ~new_n10801_ & ~new_n10813_;
  assign new_n10815_ = ~new_n10798_ & ~new_n10811_;
  assign A6048 = ~new_n10801_ & ~new_n10815_;
  assign new_n10817_ = new_n10798_ & new_n10803_;
  assign new_n10818_ = ~new_n10801_ & ~new_n10817_;
  assign new_n10819_ = new_n10801_ & ~new_n10818_;
  assign new_n10820_ = new_n10801_ & new_n10817_;
  assign new_n10821_ = new_n10819_ & ~new_n10820_;
  assign new_n10822_ = new_n10803_ & ~new_n10821_;
  assign A6047 = new_n10810_ | new_n10822_;
  assign new_n10824_ = new_n10805_ & new_n10808_;
  assign new_n10825_ = ~new_n10809_ & ~new_n10824_;
  assign new_n10826_ = ~new_n10801_ & ~new_n10805_;
  assign new_n10827_ = new_n10801_ & new_n10805_;
  assign new_n10828_ = ~new_n10826_ & ~new_n10827_;
  assign new_n10829_ = new_n10825_ & ~new_n10828_;
  assign A6046 = new_n10822_ | new_n10829_;
  assign new_n10831_ = new_n10803_ & ~new_n10829_;
  assign new_n10832_ = ~new_n10803_ & new_n10829_;
  assign new_n10833_ = ~new_n10831_ & ~new_n10832_;
  assign A6045 = ~new_n10801_ & ~new_n10833_;
  assign new_n10835_ = ~new_n3505_ & ~new_n3647_;
  assign new_n10836_ = ~new_n3508_ & ~new_n10835_;
  assign new_n10837_ = ~new_n3740_ & ~new_n3882_;
  assign new_n10838_ = ~new_n3743_ & ~new_n10837_;
  assign new_n10839_ = ~new_n10836_ & new_n10838_;
  assign new_n10840_ = new_n10836_ & ~new_n10838_;
  assign new_n10841_ = ~new_n10839_ & ~new_n10840_;
  assign new_n10842_ = ~new_n3978_ & ~new_n4120_;
  assign new_n10843_ = ~new_n3981_ & ~new_n10842_;
  assign new_n10844_ = ~new_n4213_ & ~new_n4355_;
  assign new_n10845_ = ~new_n4216_ & ~new_n10844_;
  assign new_n10846_ = new_n10841_ & ~new_n10845_;
  assign new_n10847_ = ~new_n4449_ & ~new_n4591_;
  assign new_n10848_ = ~new_n4452_ & ~new_n10847_;
  assign new_n10849_ = ~new_n10845_ & ~new_n10848_;
  assign new_n10850_ = ~new_n10846_ & ~new_n10849_;
  assign new_n10851_ = new_n10843_ & new_n10850_;
  assign new_n10852_ = ~new_n10843_ & ~new_n10850_;
  assign new_n10853_ = ~new_n10851_ & ~new_n10852_;
  assign A6016 = ~new_n10841_ & ~new_n10853_;
  assign new_n10855_ = ~new_n10838_ & ~new_n10851_;
  assign A6015 = ~new_n10841_ & ~new_n10855_;
  assign new_n10857_ = new_n10838_ & new_n10843_;
  assign new_n10858_ = ~new_n10841_ & ~new_n10857_;
  assign new_n10859_ = new_n10841_ & ~new_n10858_;
  assign new_n10860_ = new_n10841_ & new_n10857_;
  assign new_n10861_ = new_n10859_ & ~new_n10860_;
  assign new_n10862_ = new_n10843_ & ~new_n10861_;
  assign A6014 = new_n10850_ | new_n10862_;
  assign new_n10864_ = new_n10845_ & new_n10848_;
  assign new_n10865_ = ~new_n10849_ & ~new_n10864_;
  assign new_n10866_ = ~new_n10841_ & ~new_n10845_;
  assign new_n10867_ = new_n10841_ & new_n10845_;
  assign new_n10868_ = ~new_n10866_ & ~new_n10867_;
  assign new_n10869_ = new_n10865_ & ~new_n10868_;
  assign A6013 = new_n10862_ | new_n10869_;
  assign new_n10871_ = new_n10843_ & ~new_n10869_;
  assign new_n10872_ = ~new_n10843_ & new_n10869_;
  assign new_n10873_ = ~new_n10871_ & ~new_n10872_;
  assign A6012 = ~new_n10841_ & ~new_n10873_;
  assign new_n10875_ = ~new_n4706_ & ~new_n4848_;
  assign new_n10876_ = ~new_n4709_ & ~new_n10875_;
  assign new_n10877_ = ~new_n4941_ & ~new_n5083_;
  assign new_n10878_ = ~new_n4944_ & ~new_n10877_;
  assign new_n10879_ = ~new_n10876_ & new_n10878_;
  assign new_n10880_ = new_n10876_ & ~new_n10878_;
  assign new_n10881_ = ~new_n10879_ & ~new_n10880_;
  assign new_n10882_ = ~new_n5179_ & ~new_n5321_;
  assign new_n10883_ = ~new_n5182_ & ~new_n10882_;
  assign new_n10884_ = ~new_n5414_ & ~new_n5556_;
  assign new_n10885_ = ~new_n5417_ & ~new_n10884_;
  assign new_n10886_ = new_n10881_ & ~new_n10885_;
  assign new_n10887_ = ~new_n5650_ & ~new_n5792_;
  assign new_n10888_ = ~new_n5653_ & ~new_n10887_;
  assign new_n10889_ = ~new_n10885_ & ~new_n10888_;
  assign new_n10890_ = ~new_n10886_ & ~new_n10889_;
  assign new_n10891_ = new_n10883_ & new_n10890_;
  assign new_n10892_ = ~new_n10883_ & ~new_n10890_;
  assign new_n10893_ = ~new_n10891_ & ~new_n10892_;
  assign A5983 = ~new_n10881_ & ~new_n10893_;
  assign new_n10895_ = ~new_n10878_ & ~new_n10891_;
  assign A5982 = ~new_n10881_ & ~new_n10895_;
  assign new_n10897_ = new_n10878_ & new_n10883_;
  assign new_n10898_ = ~new_n10881_ & ~new_n10897_;
  assign new_n10899_ = new_n10881_ & ~new_n10898_;
  assign new_n10900_ = new_n10881_ & new_n10897_;
  assign new_n10901_ = new_n10899_ & ~new_n10900_;
  assign new_n10902_ = new_n10883_ & ~new_n10901_;
  assign A5981 = new_n10890_ | new_n10902_;
  assign new_n10904_ = new_n10885_ & new_n10888_;
  assign new_n10905_ = ~new_n10889_ & ~new_n10904_;
  assign new_n10906_ = ~new_n10881_ & ~new_n10885_;
  assign new_n10907_ = new_n10881_ & new_n10885_;
  assign new_n10908_ = ~new_n10906_ & ~new_n10907_;
  assign new_n10909_ = new_n10905_ & ~new_n10908_;
  assign A5980 = new_n10902_ | new_n10909_;
  assign new_n10911_ = new_n10883_ & ~new_n10909_;
  assign new_n10912_ = ~new_n10883_ & new_n10909_;
  assign new_n10913_ = ~new_n10911_ & ~new_n10912_;
  assign A5979 = ~new_n10881_ & ~new_n10913_;
  assign new_n10915_ = ~new_n5884_ & ~new_n5981_;
  assign new_n10916_ = ~new_n5887_ & ~new_n10915_;
  assign new_n10917_ = ~new_n6044_ & ~new_n6141_;
  assign new_n10918_ = ~new_n6047_ & ~new_n10917_;
  assign new_n10919_ = ~new_n10916_ & new_n10918_;
  assign new_n10920_ = new_n10916_ & ~new_n10918_;
  assign new_n10921_ = ~new_n10919_ & ~new_n10920_;
  assign new_n10922_ = ~new_n6207_ & ~new_n6304_;
  assign new_n10923_ = ~new_n6210_ & ~new_n10922_;
  assign new_n10924_ = ~new_n6367_ & ~new_n6464_;
  assign new_n10925_ = ~new_n6370_ & ~new_n10924_;
  assign new_n10926_ = new_n10921_ & ~new_n10925_;
  assign new_n10927_ = ~new_n6528_ & ~new_n6625_;
  assign new_n10928_ = ~new_n6531_ & ~new_n10927_;
  assign new_n10929_ = ~new_n10925_ & ~new_n10928_;
  assign new_n10930_ = ~new_n10926_ & ~new_n10929_;
  assign new_n10931_ = new_n10923_ & new_n10930_;
  assign new_n10932_ = ~new_n10923_ & ~new_n10930_;
  assign new_n10933_ = ~new_n10931_ & ~new_n10932_;
  assign A5950 = ~new_n10921_ & ~new_n10933_;
  assign new_n10935_ = ~new_n10918_ & ~new_n10931_;
  assign A5949 = ~new_n10921_ & ~new_n10935_;
  assign new_n10937_ = new_n10918_ & new_n10923_;
  assign new_n10938_ = ~new_n10921_ & ~new_n10937_;
  assign new_n10939_ = new_n10921_ & ~new_n10938_;
  assign new_n10940_ = new_n10921_ & new_n10937_;
  assign new_n10941_ = new_n10939_ & ~new_n10940_;
  assign new_n10942_ = new_n10923_ & ~new_n10941_;
  assign A5948 = new_n10930_ | new_n10942_;
  assign new_n10944_ = new_n10925_ & new_n10928_;
  assign new_n10945_ = ~new_n10929_ & ~new_n10944_;
  assign new_n10946_ = ~new_n10921_ & ~new_n10925_;
  assign new_n10947_ = new_n10921_ & new_n10925_;
  assign new_n10948_ = ~new_n10946_ & ~new_n10947_;
  assign new_n10949_ = new_n10945_ & ~new_n10948_;
  assign A5947 = new_n10942_ | new_n10949_;
  assign new_n10951_ = new_n10923_ & ~new_n10949_;
  assign new_n10952_ = ~new_n10923_ & new_n10949_;
  assign new_n10953_ = ~new_n10951_ & ~new_n10952_;
  assign A5946 = ~new_n10921_ & ~new_n10953_;
  assign new_n10955_ = ~new_n6658_ & ~new_n6671_;
  assign new_n10956_ = ~new_n6661_ & ~new_n10955_;
  assign new_n10957_ = ~new_n6678_ & ~new_n6691_;
  assign new_n10958_ = ~new_n6681_ & ~new_n10957_;
  assign new_n10959_ = ~new_n10956_ & new_n10958_;
  assign new_n10960_ = new_n10956_ & ~new_n10958_;
  assign new_n10961_ = ~new_n10959_ & ~new_n10960_;
  assign new_n10962_ = ~new_n6701_ & ~new_n6714_;
  assign new_n10963_ = ~new_n6704_ & ~new_n10962_;
  assign new_n10964_ = ~new_n6721_ & ~new_n6734_;
  assign new_n10965_ = ~new_n6724_ & ~new_n10964_;
  assign new_n10966_ = new_n10961_ & ~new_n10965_;
  assign new_n10967_ = ~new_n6742_ & ~new_n6755_;
  assign new_n10968_ = ~new_n6745_ & ~new_n10967_;
  assign new_n10969_ = ~new_n10965_ & ~new_n10968_;
  assign new_n10970_ = ~new_n10966_ & ~new_n10969_;
  assign new_n10971_ = new_n10963_ & new_n10970_;
  assign new_n10972_ = ~new_n10963_ & ~new_n10970_;
  assign new_n10973_ = ~new_n10971_ & ~new_n10972_;
  assign A5917 = ~new_n10961_ & ~new_n10973_;
  assign new_n10975_ = ~new_n10958_ & ~new_n10971_;
  assign A5916 = ~new_n10961_ & ~new_n10975_;
  assign new_n10977_ = new_n10958_ & new_n10963_;
  assign new_n10978_ = ~new_n10961_ & ~new_n10977_;
  assign new_n10979_ = new_n10961_ & ~new_n10978_;
  assign new_n10980_ = new_n10961_ & new_n10977_;
  assign new_n10981_ = new_n10979_ & ~new_n10980_;
  assign new_n10982_ = new_n10963_ & ~new_n10981_;
  assign A5915 = new_n10970_ | new_n10982_;
  assign new_n10984_ = new_n10965_ & new_n10968_;
  assign new_n10985_ = ~new_n10969_ & ~new_n10984_;
  assign new_n10986_ = ~new_n10961_ & ~new_n10965_;
  assign new_n10987_ = new_n10961_ & new_n10965_;
  assign new_n10988_ = ~new_n10986_ & ~new_n10987_;
  assign new_n10989_ = new_n10985_ & ~new_n10988_;
  assign A5914 = new_n10982_ | new_n10989_;
  assign new_n10991_ = new_n10963_ & ~new_n10989_;
  assign new_n10992_ = ~new_n10963_ & new_n10989_;
  assign new_n10993_ = ~new_n10991_ & ~new_n10992_;
  assign A5913 = ~new_n10961_ & ~new_n10993_;
  assign new_n10995_ = ~new_n6788_ & ~new_n6801_;
  assign new_n10996_ = ~new_n6791_ & ~new_n10995_;
  assign new_n10997_ = ~new_n6808_ & ~new_n6821_;
  assign new_n10998_ = ~new_n6811_ & ~new_n10997_;
  assign new_n10999_ = ~new_n10996_ & new_n10998_;
  assign new_n11000_ = new_n10996_ & ~new_n10998_;
  assign new_n11001_ = ~new_n10999_ & ~new_n11000_;
  assign new_n11002_ = ~new_n6831_ & ~new_n6844_;
  assign new_n11003_ = ~new_n6834_ & ~new_n11002_;
  assign new_n11004_ = ~new_n6851_ & ~new_n6864_;
  assign new_n11005_ = ~new_n6854_ & ~new_n11004_;
  assign new_n11006_ = new_n11001_ & ~new_n11005_;
  assign new_n11007_ = ~new_n6872_ & ~new_n6885_;
  assign new_n11008_ = ~new_n6875_ & ~new_n11007_;
  assign new_n11009_ = ~new_n11005_ & ~new_n11008_;
  assign new_n11010_ = ~new_n11006_ & ~new_n11009_;
  assign new_n11011_ = new_n11003_ & new_n11010_;
  assign new_n11012_ = ~new_n11003_ & ~new_n11010_;
  assign new_n11013_ = ~new_n11011_ & ~new_n11012_;
  assign A5884 = ~new_n11001_ & ~new_n11013_;
  assign new_n11015_ = ~new_n10998_ & ~new_n11011_;
  assign A5883 = ~new_n11001_ & ~new_n11015_;
  assign new_n11017_ = new_n10998_ & new_n11003_;
  assign new_n11018_ = ~new_n11001_ & ~new_n11017_;
  assign new_n11019_ = new_n11001_ & ~new_n11018_;
  assign new_n11020_ = new_n11001_ & new_n11017_;
  assign new_n11021_ = new_n11019_ & ~new_n11020_;
  assign new_n11022_ = new_n11003_ & ~new_n11021_;
  assign A5882 = new_n11010_ | new_n11022_;
  assign new_n11024_ = new_n11005_ & new_n11008_;
  assign new_n11025_ = ~new_n11009_ & ~new_n11024_;
  assign new_n11026_ = ~new_n11001_ & ~new_n11005_;
  assign new_n11027_ = new_n11001_ & new_n11005_;
  assign new_n11028_ = ~new_n11026_ & ~new_n11027_;
  assign new_n11029_ = new_n11025_ & ~new_n11028_;
  assign A5881 = new_n11022_ | new_n11029_;
  assign new_n11031_ = new_n11003_ & ~new_n11029_;
  assign new_n11032_ = ~new_n11003_ & new_n11029_;
  assign new_n11033_ = ~new_n11031_ & ~new_n11032_;
  assign A5880 = ~new_n11001_ & ~new_n11033_;
  assign new_n11035_ = ~new_n6918_ & ~new_n6931_;
  assign new_n11036_ = ~new_n6921_ & ~new_n11035_;
  assign new_n11037_ = ~new_n6938_ & ~new_n6951_;
  assign new_n11038_ = ~new_n6941_ & ~new_n11037_;
  assign new_n11039_ = ~new_n11036_ & new_n11038_;
  assign new_n11040_ = new_n11036_ & ~new_n11038_;
  assign new_n11041_ = ~new_n11039_ & ~new_n11040_;
  assign new_n11042_ = ~new_n6961_ & ~new_n6974_;
  assign new_n11043_ = ~new_n6964_ & ~new_n11042_;
  assign new_n11044_ = ~new_n6981_ & ~new_n6994_;
  assign new_n11045_ = ~new_n6984_ & ~new_n11044_;
  assign new_n11046_ = new_n11041_ & ~new_n11045_;
  assign new_n11047_ = ~new_n7002_ & ~new_n7015_;
  assign new_n11048_ = ~new_n7005_ & ~new_n11047_;
  assign new_n11049_ = ~new_n11045_ & ~new_n11048_;
  assign new_n11050_ = ~new_n11046_ & ~new_n11049_;
  assign new_n11051_ = new_n11043_ & new_n11050_;
  assign new_n11052_ = ~new_n11043_ & ~new_n11050_;
  assign new_n11053_ = ~new_n11051_ & ~new_n11052_;
  assign A5851 = ~new_n11041_ & ~new_n11053_;
  assign new_n11055_ = ~new_n11038_ & ~new_n11051_;
  assign A5850 = ~new_n11041_ & ~new_n11055_;
  assign new_n11057_ = new_n11038_ & new_n11043_;
  assign new_n11058_ = ~new_n11041_ & ~new_n11057_;
  assign new_n11059_ = new_n11041_ & ~new_n11058_;
  assign new_n11060_ = new_n11041_ & new_n11057_;
  assign new_n11061_ = new_n11059_ & ~new_n11060_;
  assign new_n11062_ = new_n11043_ & ~new_n11061_;
  assign A5849 = new_n11050_ | new_n11062_;
  assign new_n11064_ = new_n11045_ & new_n11048_;
  assign new_n11065_ = ~new_n11049_ & ~new_n11064_;
  assign new_n11066_ = ~new_n11041_ & ~new_n11045_;
  assign new_n11067_ = new_n11041_ & new_n11045_;
  assign new_n11068_ = ~new_n11066_ & ~new_n11067_;
  assign new_n11069_ = new_n11065_ & ~new_n11068_;
  assign A5848 = new_n11062_ | new_n11069_;
  assign new_n11071_ = new_n11043_ & ~new_n11069_;
  assign new_n11072_ = ~new_n11043_ & new_n11069_;
  assign new_n11073_ = ~new_n11071_ & ~new_n11072_;
  assign A5847 = ~new_n11041_ & ~new_n11073_;
  assign new_n11075_ = ~new_n7048_ & ~new_n7061_;
  assign new_n11076_ = ~new_n7051_ & ~new_n11075_;
  assign new_n11077_ = ~new_n7068_ & ~new_n7081_;
  assign new_n11078_ = ~new_n7071_ & ~new_n11077_;
  assign new_n11079_ = ~new_n11076_ & new_n11078_;
  assign new_n11080_ = new_n11076_ & ~new_n11078_;
  assign new_n11081_ = ~new_n11079_ & ~new_n11080_;
  assign new_n11082_ = ~new_n7091_ & ~new_n7104_;
  assign new_n11083_ = ~new_n7094_ & ~new_n11082_;
  assign new_n11084_ = ~new_n7111_ & ~new_n7124_;
  assign new_n11085_ = ~new_n7114_ & ~new_n11084_;
  assign new_n11086_ = new_n11081_ & ~new_n11085_;
  assign new_n11087_ = ~new_n7132_ & ~new_n7145_;
  assign new_n11088_ = ~new_n7135_ & ~new_n11087_;
  assign new_n11089_ = ~new_n11085_ & ~new_n11088_;
  assign new_n11090_ = ~new_n11086_ & ~new_n11089_;
  assign new_n11091_ = new_n11083_ & new_n11090_;
  assign new_n11092_ = ~new_n11083_ & ~new_n11090_;
  assign new_n11093_ = ~new_n11091_ & ~new_n11092_;
  assign A5818 = ~new_n11081_ & ~new_n11093_;
  assign new_n11095_ = ~new_n11078_ & ~new_n11091_;
  assign A5817 = ~new_n11081_ & ~new_n11095_;
  assign new_n11097_ = new_n11078_ & new_n11083_;
  assign new_n11098_ = ~new_n11081_ & ~new_n11097_;
  assign new_n11099_ = new_n11081_ & ~new_n11098_;
  assign new_n11100_ = new_n11081_ & new_n11097_;
  assign new_n11101_ = new_n11099_ & ~new_n11100_;
  assign new_n11102_ = new_n11083_ & ~new_n11101_;
  assign A5816 = new_n11090_ | new_n11102_;
  assign new_n11104_ = new_n11085_ & new_n11088_;
  assign new_n11105_ = ~new_n11089_ & ~new_n11104_;
  assign new_n11106_ = ~new_n11081_ & ~new_n11085_;
  assign new_n11107_ = new_n11081_ & new_n11085_;
  assign new_n11108_ = ~new_n11106_ & ~new_n11107_;
  assign new_n11109_ = new_n11105_ & ~new_n11108_;
  assign A5815 = new_n11102_ | new_n11109_;
  assign new_n11111_ = new_n11083_ & ~new_n11109_;
  assign new_n11112_ = ~new_n11083_ & new_n11109_;
  assign new_n11113_ = ~new_n11111_ & ~new_n11112_;
  assign A5814 = ~new_n11081_ & ~new_n11113_;
  assign new_n11115_ = ~new_n7183_ & ~new_n7196_;
  assign new_n11116_ = ~new_n7186_ & ~new_n11115_;
  assign new_n11117_ = ~new_n7203_ & ~new_n7216_;
  assign new_n11118_ = ~new_n7206_ & ~new_n11117_;
  assign new_n11119_ = ~new_n11116_ & new_n11118_;
  assign new_n11120_ = new_n11116_ & ~new_n11118_;
  assign new_n11121_ = ~new_n11119_ & ~new_n11120_;
  assign new_n11122_ = ~new_n7226_ & ~new_n7239_;
  assign new_n11123_ = ~new_n7229_ & ~new_n11122_;
  assign new_n11124_ = ~new_n7246_ & ~new_n7259_;
  assign new_n11125_ = ~new_n7249_ & ~new_n11124_;
  assign new_n11126_ = new_n11121_ & ~new_n11125_;
  assign new_n11127_ = ~new_n7267_ & ~new_n7280_;
  assign new_n11128_ = ~new_n7270_ & ~new_n11127_;
  assign new_n11129_ = ~new_n11125_ & ~new_n11128_;
  assign new_n11130_ = ~new_n11126_ & ~new_n11129_;
  assign new_n11131_ = new_n11123_ & new_n11130_;
  assign new_n11132_ = ~new_n11123_ & ~new_n11130_;
  assign new_n11133_ = ~new_n11131_ & ~new_n11132_;
  assign A5785 = ~new_n11121_ & ~new_n11133_;
  assign new_n11135_ = ~new_n11118_ & ~new_n11131_;
  assign A5784 = ~new_n11121_ & ~new_n11135_;
  assign new_n11137_ = new_n11118_ & new_n11123_;
  assign new_n11138_ = ~new_n11121_ & ~new_n11137_;
  assign new_n11139_ = new_n11121_ & ~new_n11138_;
  assign new_n11140_ = new_n11121_ & new_n11137_;
  assign new_n11141_ = new_n11139_ & ~new_n11140_;
  assign new_n11142_ = new_n11123_ & ~new_n11141_;
  assign A5783 = new_n11130_ | new_n11142_;
  assign new_n11144_ = new_n11125_ & new_n11128_;
  assign new_n11145_ = ~new_n11129_ & ~new_n11144_;
  assign new_n11146_ = ~new_n11121_ & ~new_n11125_;
  assign new_n11147_ = new_n11121_ & new_n11125_;
  assign new_n11148_ = ~new_n11146_ & ~new_n11147_;
  assign new_n11149_ = new_n11145_ & ~new_n11148_;
  assign A5782 = new_n11142_ | new_n11149_;
  assign new_n11151_ = new_n11123_ & ~new_n11149_;
  assign new_n11152_ = ~new_n11123_ & new_n11149_;
  assign new_n11153_ = ~new_n11151_ & ~new_n11152_;
  assign A5781 = ~new_n11121_ & ~new_n11153_;
  assign new_n11155_ = new_n7323_ & ~new_n7351_;
  assign new_n11156_ = ~new_n7326_ & ~new_n11155_;
  assign new_n11157_ = new_n7368_ & ~new_n7396_;
  assign new_n11158_ = ~new_n7371_ & ~new_n11157_;
  assign new_n11159_ = ~new_n11156_ & new_n11158_;
  assign new_n11160_ = new_n11156_ & ~new_n11158_;
  assign new_n11161_ = ~new_n11159_ & ~new_n11160_;
  assign new_n11162_ = new_n7416_ & ~new_n7444_;
  assign new_n11163_ = ~new_n7419_ & ~new_n11162_;
  assign new_n11164_ = new_n7461_ & ~new_n7489_;
  assign new_n11165_ = ~new_n7464_ & ~new_n11164_;
  assign new_n11166_ = new_n11161_ & ~new_n11165_;
  assign new_n11167_ = new_n7507_ & ~new_n7535_;
  assign new_n11168_ = ~new_n7510_ & ~new_n11167_;
  assign new_n11169_ = ~new_n11165_ & ~new_n11168_;
  assign new_n11170_ = ~new_n11166_ & ~new_n11169_;
  assign new_n11171_ = new_n11163_ & new_n11170_;
  assign new_n11172_ = ~new_n11163_ & ~new_n11170_;
  assign new_n11173_ = ~new_n11171_ & ~new_n11172_;
  assign A5752 = ~new_n11161_ & ~new_n11173_;
  assign new_n11175_ = ~new_n11158_ & ~new_n11171_;
  assign A5751 = ~new_n11161_ & ~new_n11175_;
  assign new_n11177_ = new_n11158_ & new_n11163_;
  assign new_n11178_ = ~new_n11161_ & ~new_n11177_;
  assign new_n11179_ = new_n11161_ & ~new_n11178_;
  assign new_n11180_ = new_n11161_ & new_n11177_;
  assign new_n11181_ = new_n11179_ & ~new_n11180_;
  assign new_n11182_ = new_n11163_ & ~new_n11181_;
  assign A5750 = new_n11170_ | new_n11182_;
  assign new_n11184_ = new_n11165_ & new_n11168_;
  assign new_n11185_ = ~new_n11169_ & ~new_n11184_;
  assign new_n11186_ = ~new_n11161_ & ~new_n11165_;
  assign new_n11187_ = new_n11161_ & new_n11165_;
  assign new_n11188_ = ~new_n11186_ & ~new_n11187_;
  assign new_n11189_ = new_n11185_ & ~new_n11188_;
  assign A5749 = new_n11182_ | new_n11189_;
  assign new_n11191_ = new_n11163_ & ~new_n11189_;
  assign new_n11192_ = ~new_n11163_ & new_n11189_;
  assign new_n11193_ = ~new_n11191_ & ~new_n11192_;
  assign A5748 = ~new_n11161_ & ~new_n11193_;
  assign new_n11195_ = new_n7578_ & ~new_n7606_;
  assign new_n11196_ = ~new_n7581_ & ~new_n11195_;
  assign new_n11197_ = new_n7623_ & ~new_n7651_;
  assign new_n11198_ = ~new_n7626_ & ~new_n11197_;
  assign new_n11199_ = ~new_n11196_ & new_n11198_;
  assign new_n11200_ = new_n11196_ & ~new_n11198_;
  assign new_n11201_ = ~new_n11199_ & ~new_n11200_;
  assign new_n11202_ = new_n7671_ & ~new_n7699_;
  assign new_n11203_ = ~new_n7674_ & ~new_n11202_;
  assign new_n11204_ = new_n7716_ & ~new_n7744_;
  assign new_n11205_ = ~new_n7719_ & ~new_n11204_;
  assign new_n11206_ = new_n11201_ & ~new_n11205_;
  assign new_n11207_ = new_n7762_ & ~new_n7790_;
  assign new_n11208_ = ~new_n7765_ & ~new_n11207_;
  assign new_n11209_ = ~new_n11205_ & ~new_n11208_;
  assign new_n11210_ = ~new_n11206_ & ~new_n11209_;
  assign new_n11211_ = new_n11203_ & new_n11210_;
  assign new_n11212_ = ~new_n11203_ & ~new_n11210_;
  assign new_n11213_ = ~new_n11211_ & ~new_n11212_;
  assign A5719 = ~new_n11201_ & ~new_n11213_;
  assign new_n11215_ = ~new_n11198_ & ~new_n11211_;
  assign A5718 = ~new_n11201_ & ~new_n11215_;
  assign new_n11217_ = new_n11198_ & new_n11203_;
  assign new_n11218_ = ~new_n11201_ & ~new_n11217_;
  assign new_n11219_ = new_n11201_ & ~new_n11218_;
  assign new_n11220_ = new_n11201_ & new_n11217_;
  assign new_n11221_ = new_n11219_ & ~new_n11220_;
  assign new_n11222_ = new_n11203_ & ~new_n11221_;
  assign A5717 = new_n11210_ | new_n11222_;
  assign new_n11224_ = new_n11205_ & new_n11208_;
  assign new_n11225_ = ~new_n11209_ & ~new_n11224_;
  assign new_n11226_ = ~new_n11201_ & ~new_n11205_;
  assign new_n11227_ = new_n11201_ & new_n11205_;
  assign new_n11228_ = ~new_n11226_ & ~new_n11227_;
  assign new_n11229_ = new_n11225_ & ~new_n11228_;
  assign A5716 = new_n11222_ | new_n11229_;
  assign new_n11231_ = new_n11203_ & ~new_n11229_;
  assign new_n11232_ = ~new_n11203_ & new_n11229_;
  assign new_n11233_ = ~new_n11231_ & ~new_n11232_;
  assign A5715 = ~new_n11201_ & ~new_n11233_;
  assign new_n11235_ = new_n7833_ & ~new_n7861_;
  assign new_n11236_ = ~new_n7836_ & ~new_n11235_;
  assign new_n11237_ = new_n7878_ & ~new_n7906_;
  assign new_n11238_ = ~new_n7881_ & ~new_n11237_;
  assign new_n11239_ = ~new_n11236_ & new_n11238_;
  assign new_n11240_ = new_n11236_ & ~new_n11238_;
  assign new_n11241_ = ~new_n11239_ & ~new_n11240_;
  assign new_n11242_ = new_n7926_ & ~new_n7954_;
  assign new_n11243_ = ~new_n7929_ & ~new_n11242_;
  assign new_n11244_ = new_n7971_ & ~new_n7999_;
  assign new_n11245_ = ~new_n7974_ & ~new_n11244_;
  assign new_n11246_ = new_n11241_ & ~new_n11245_;
  assign new_n11247_ = new_n8017_ & ~new_n8045_;
  assign new_n11248_ = ~new_n8020_ & ~new_n11247_;
  assign new_n11249_ = ~new_n11245_ & ~new_n11248_;
  assign new_n11250_ = ~new_n11246_ & ~new_n11249_;
  assign new_n11251_ = new_n11243_ & new_n11250_;
  assign new_n11252_ = ~new_n11243_ & ~new_n11250_;
  assign new_n11253_ = ~new_n11251_ & ~new_n11252_;
  assign A5686 = ~new_n11241_ & ~new_n11253_;
  assign new_n11255_ = ~new_n11238_ & ~new_n11251_;
  assign A5685 = ~new_n11241_ & ~new_n11255_;
  assign new_n11257_ = new_n11238_ & new_n11243_;
  assign new_n11258_ = ~new_n11241_ & ~new_n11257_;
  assign new_n11259_ = new_n11241_ & ~new_n11258_;
  assign new_n11260_ = new_n11241_ & new_n11257_;
  assign new_n11261_ = new_n11259_ & ~new_n11260_;
  assign new_n11262_ = new_n11243_ & ~new_n11261_;
  assign A5684 = new_n11250_ | new_n11262_;
  assign new_n11264_ = new_n11245_ & new_n11248_;
  assign new_n11265_ = ~new_n11249_ & ~new_n11264_;
  assign new_n11266_ = ~new_n11241_ & ~new_n11245_;
  assign new_n11267_ = new_n11241_ & new_n11245_;
  assign new_n11268_ = ~new_n11266_ & ~new_n11267_;
  assign new_n11269_ = new_n11265_ & ~new_n11268_;
  assign A5683 = new_n11262_ | new_n11269_;
  assign new_n11271_ = new_n11243_ & ~new_n11269_;
  assign new_n11272_ = ~new_n11243_ & new_n11269_;
  assign new_n11273_ = ~new_n11271_ & ~new_n11272_;
  assign A5682 = ~new_n11241_ & ~new_n11273_;
  assign new_n11275_ = new_n8088_ & ~new_n8116_;
  assign new_n11276_ = ~new_n8091_ & ~new_n11275_;
  assign new_n11277_ = new_n8133_ & ~new_n8161_;
  assign new_n11278_ = ~new_n8136_ & ~new_n11277_;
  assign new_n11279_ = ~new_n11276_ & new_n11278_;
  assign new_n11280_ = new_n11276_ & ~new_n11278_;
  assign new_n11281_ = ~new_n11279_ & ~new_n11280_;
  assign new_n11282_ = new_n8181_ & ~new_n8209_;
  assign new_n11283_ = ~new_n8184_ & ~new_n11282_;
  assign new_n11284_ = new_n8226_ & ~new_n8254_;
  assign new_n11285_ = ~new_n8229_ & ~new_n11284_;
  assign new_n11286_ = new_n11281_ & ~new_n11285_;
  assign new_n11287_ = new_n8272_ & ~new_n8300_;
  assign new_n11288_ = ~new_n8275_ & ~new_n11287_;
  assign new_n11289_ = ~new_n11285_ & ~new_n11288_;
  assign new_n11290_ = ~new_n11286_ & ~new_n11289_;
  assign new_n11291_ = new_n11283_ & new_n11290_;
  assign new_n11292_ = ~new_n11283_ & ~new_n11290_;
  assign new_n11293_ = ~new_n11291_ & ~new_n11292_;
  assign A5653 = ~new_n11281_ & ~new_n11293_;
  assign new_n11295_ = ~new_n11278_ & ~new_n11291_;
  assign A5652 = ~new_n11281_ & ~new_n11295_;
  assign new_n11297_ = new_n11278_ & new_n11283_;
  assign new_n11298_ = ~new_n11281_ & ~new_n11297_;
  assign new_n11299_ = new_n11281_ & ~new_n11298_;
  assign new_n11300_ = new_n11281_ & new_n11297_;
  assign new_n11301_ = new_n11299_ & ~new_n11300_;
  assign new_n11302_ = new_n11283_ & ~new_n11301_;
  assign A5651 = new_n11290_ | new_n11302_;
  assign new_n11304_ = new_n11285_ & new_n11288_;
  assign new_n11305_ = ~new_n11289_ & ~new_n11304_;
  assign new_n11306_ = ~new_n11281_ & ~new_n11285_;
  assign new_n11307_ = new_n11281_ & new_n11285_;
  assign new_n11308_ = ~new_n11306_ & ~new_n11307_;
  assign new_n11309_ = new_n11305_ & ~new_n11308_;
  assign A5650 = new_n11302_ | new_n11309_;
  assign new_n11311_ = new_n11283_ & ~new_n11309_;
  assign new_n11312_ = ~new_n11283_ & new_n11309_;
  assign new_n11313_ = ~new_n11311_ & ~new_n11312_;
  assign A5649 = ~new_n11281_ & ~new_n11313_;
  assign new_n11315_ = new_n8339_ & ~new_n8367_;
  assign new_n11316_ = ~new_n8342_ & ~new_n11315_;
  assign new_n11317_ = new_n8384_ & ~new_n8412_;
  assign new_n11318_ = ~new_n8387_ & ~new_n11317_;
  assign new_n11319_ = ~new_n11316_ & new_n11318_;
  assign new_n11320_ = new_n11316_ & ~new_n11318_;
  assign new_n11321_ = ~new_n11319_ & ~new_n11320_;
  assign new_n11322_ = new_n8432_ & ~new_n8460_;
  assign new_n11323_ = ~new_n8435_ & ~new_n11322_;
  assign new_n11324_ = new_n8477_ & ~new_n8505_;
  assign new_n11325_ = ~new_n8480_ & ~new_n11324_;
  assign new_n11326_ = new_n11321_ & ~new_n11325_;
  assign new_n11327_ = new_n8523_ & ~new_n8551_;
  assign new_n11328_ = ~new_n8526_ & ~new_n11327_;
  assign new_n11329_ = ~new_n11325_ & ~new_n11328_;
  assign new_n11330_ = ~new_n11326_ & ~new_n11329_;
  assign new_n11331_ = new_n11323_ & new_n11330_;
  assign new_n11332_ = ~new_n11323_ & ~new_n11330_;
  assign new_n11333_ = ~new_n11331_ & ~new_n11332_;
  assign A5620 = ~new_n11321_ & ~new_n11333_;
  assign new_n11335_ = ~new_n11318_ & ~new_n11331_;
  assign A5619 = ~new_n11321_ & ~new_n11335_;
  assign new_n11337_ = new_n11318_ & new_n11323_;
  assign new_n11338_ = ~new_n11321_ & ~new_n11337_;
  assign new_n11339_ = new_n11321_ & ~new_n11338_;
  assign new_n11340_ = new_n11321_ & new_n11337_;
  assign new_n11341_ = new_n11339_ & ~new_n11340_;
  assign new_n11342_ = new_n11323_ & ~new_n11341_;
  assign A5618 = new_n11330_ | new_n11342_;
  assign new_n11344_ = new_n11325_ & new_n11328_;
  assign new_n11345_ = ~new_n11329_ & ~new_n11344_;
  assign new_n11346_ = ~new_n11321_ & ~new_n11325_;
  assign new_n11347_ = new_n11321_ & new_n11325_;
  assign new_n11348_ = ~new_n11346_ & ~new_n11347_;
  assign new_n11349_ = new_n11345_ & ~new_n11348_;
  assign A5617 = new_n11342_ | new_n11349_;
  assign new_n11351_ = new_n11323_ & ~new_n11349_;
  assign new_n11352_ = ~new_n11323_ & new_n11349_;
  assign new_n11353_ = ~new_n11351_ & ~new_n11352_;
  assign A5616 = ~new_n11321_ & ~new_n11353_;
  assign new_n11355_ = new_n8594_ & ~new_n8622_;
  assign new_n11356_ = ~new_n8597_ & ~new_n11355_;
  assign new_n11357_ = new_n8639_ & ~new_n8667_;
  assign new_n11358_ = ~new_n8642_ & ~new_n11357_;
  assign new_n11359_ = ~new_n11356_ & new_n11358_;
  assign new_n11360_ = new_n11356_ & ~new_n11358_;
  assign new_n11361_ = ~new_n11359_ & ~new_n11360_;
  assign new_n11362_ = new_n8687_ & ~new_n8715_;
  assign new_n11363_ = ~new_n8690_ & ~new_n11362_;
  assign new_n11364_ = new_n8732_ & ~new_n8760_;
  assign new_n11365_ = ~new_n8735_ & ~new_n11364_;
  assign new_n11366_ = new_n11361_ & ~new_n11365_;
  assign new_n11367_ = new_n8778_ & ~new_n8806_;
  assign new_n11368_ = ~new_n8781_ & ~new_n11367_;
  assign new_n11369_ = ~new_n11365_ & ~new_n11368_;
  assign new_n11370_ = ~new_n11366_ & ~new_n11369_;
  assign new_n11371_ = new_n11363_ & new_n11370_;
  assign new_n11372_ = ~new_n11363_ & ~new_n11370_;
  assign new_n11373_ = ~new_n11371_ & ~new_n11372_;
  assign A5587 = ~new_n11361_ & ~new_n11373_;
  assign new_n11375_ = ~new_n11358_ & ~new_n11371_;
  assign A5586 = ~new_n11361_ & ~new_n11375_;
  assign new_n11377_ = new_n11358_ & new_n11363_;
  assign new_n11378_ = ~new_n11361_ & ~new_n11377_;
  assign new_n11379_ = new_n11361_ & ~new_n11378_;
  assign new_n11380_ = new_n11361_ & new_n11377_;
  assign new_n11381_ = new_n11379_ & ~new_n11380_;
  assign new_n11382_ = new_n11363_ & ~new_n11381_;
  assign A5585 = new_n11370_ | new_n11382_;
  assign new_n11384_ = new_n11365_ & new_n11368_;
  assign new_n11385_ = ~new_n11369_ & ~new_n11384_;
  assign new_n11386_ = ~new_n11361_ & ~new_n11365_;
  assign new_n11387_ = new_n11361_ & new_n11365_;
  assign new_n11388_ = ~new_n11386_ & ~new_n11387_;
  assign new_n11389_ = new_n11385_ & ~new_n11388_;
  assign A5584 = new_n11382_ | new_n11389_;
  assign new_n11391_ = new_n11363_ & ~new_n11389_;
  assign new_n11392_ = ~new_n11363_ & new_n11389_;
  assign new_n11393_ = ~new_n11391_ & ~new_n11392_;
  assign A5583 = ~new_n11361_ & ~new_n11393_;
  assign new_n11395_ = new_n8849_ & ~new_n8877_;
  assign new_n11396_ = ~new_n8852_ & ~new_n11395_;
  assign new_n11397_ = new_n8894_ & ~new_n8922_;
  assign new_n11398_ = ~new_n8897_ & ~new_n11397_;
  assign new_n11399_ = ~new_n11396_ & new_n11398_;
  assign new_n11400_ = new_n11396_ & ~new_n11398_;
  assign new_n11401_ = ~new_n11399_ & ~new_n11400_;
  assign new_n11402_ = new_n8942_ & ~new_n8970_;
  assign new_n11403_ = ~new_n8945_ & ~new_n11402_;
  assign new_n11404_ = new_n8987_ & ~new_n9015_;
  assign new_n11405_ = ~new_n8990_ & ~new_n11404_;
  assign new_n11406_ = new_n11401_ & ~new_n11405_;
  assign new_n11407_ = new_n9033_ & ~new_n9061_;
  assign new_n11408_ = ~new_n9036_ & ~new_n11407_;
  assign new_n11409_ = ~new_n11405_ & ~new_n11408_;
  assign new_n11410_ = ~new_n11406_ & ~new_n11409_;
  assign new_n11411_ = new_n11403_ & new_n11410_;
  assign new_n11412_ = ~new_n11403_ & ~new_n11410_;
  assign new_n11413_ = ~new_n11411_ & ~new_n11412_;
  assign A5554 = ~new_n11401_ & ~new_n11413_;
  assign new_n11415_ = ~new_n11398_ & ~new_n11411_;
  assign A5553 = ~new_n11401_ & ~new_n11415_;
  assign new_n11417_ = new_n11398_ & new_n11403_;
  assign new_n11418_ = ~new_n11401_ & ~new_n11417_;
  assign new_n11419_ = new_n11401_ & ~new_n11418_;
  assign new_n11420_ = new_n11401_ & new_n11417_;
  assign new_n11421_ = new_n11419_ & ~new_n11420_;
  assign new_n11422_ = new_n11403_ & ~new_n11421_;
  assign A5552 = new_n11410_ | new_n11422_;
  assign new_n11424_ = new_n11405_ & new_n11408_;
  assign new_n11425_ = ~new_n11409_ & ~new_n11424_;
  assign new_n11426_ = ~new_n11401_ & ~new_n11405_;
  assign new_n11427_ = new_n11401_ & new_n11405_;
  assign new_n11428_ = ~new_n11426_ & ~new_n11427_;
  assign new_n11429_ = new_n11425_ & ~new_n11428_;
  assign A5551 = new_n11422_ | new_n11429_;
  assign new_n11431_ = new_n11403_ & ~new_n11429_;
  assign new_n11432_ = ~new_n11403_ & new_n11429_;
  assign new_n11433_ = ~new_n11431_ & ~new_n11432_;
  assign A5550 = ~new_n11401_ & ~new_n11433_;
  assign new_n11435_ = new_n9104_ & ~new_n9132_;
  assign new_n11436_ = ~new_n9107_ & ~new_n11435_;
  assign new_n11437_ = new_n9149_ & ~new_n9177_;
  assign new_n11438_ = ~new_n9152_ & ~new_n11437_;
  assign new_n11439_ = ~new_n11436_ & new_n11438_;
  assign new_n11440_ = new_n11436_ & ~new_n11438_;
  assign new_n11441_ = ~new_n11439_ & ~new_n11440_;
  assign new_n11442_ = new_n9197_ & ~new_n9225_;
  assign new_n11443_ = ~new_n9200_ & ~new_n11442_;
  assign new_n11444_ = new_n9242_ & ~new_n9270_;
  assign new_n11445_ = ~new_n9245_ & ~new_n11444_;
  assign new_n11446_ = new_n11441_ & ~new_n11445_;
  assign new_n11447_ = new_n9288_ & ~new_n9316_;
  assign new_n11448_ = ~new_n9291_ & ~new_n11447_;
  assign new_n11449_ = ~new_n11445_ & ~new_n11448_;
  assign new_n11450_ = ~new_n11446_ & ~new_n11449_;
  assign new_n11451_ = new_n11443_ & new_n11450_;
  assign new_n11452_ = ~new_n11443_ & ~new_n11450_;
  assign new_n11453_ = ~new_n11451_ & ~new_n11452_;
  assign A5521 = ~new_n11441_ & ~new_n11453_;
  assign new_n11455_ = ~new_n11438_ & ~new_n11451_;
  assign A5520 = ~new_n11441_ & ~new_n11455_;
  assign new_n11457_ = new_n11438_ & new_n11443_;
  assign new_n11458_ = ~new_n11441_ & ~new_n11457_;
  assign new_n11459_ = new_n11441_ & ~new_n11458_;
  assign new_n11460_ = new_n11441_ & new_n11457_;
  assign new_n11461_ = new_n11459_ & ~new_n11460_;
  assign new_n11462_ = new_n11443_ & ~new_n11461_;
  assign A5519 = new_n11450_ | new_n11462_;
  assign new_n11464_ = new_n11445_ & new_n11448_;
  assign new_n11465_ = ~new_n11449_ & ~new_n11464_;
  assign new_n11466_ = ~new_n11441_ & ~new_n11445_;
  assign new_n11467_ = new_n11441_ & new_n11445_;
  assign new_n11468_ = ~new_n11466_ & ~new_n11467_;
  assign new_n11469_ = new_n11465_ & ~new_n11468_;
  assign A5518 = new_n11462_ | new_n11469_;
  assign new_n11471_ = new_n11443_ & ~new_n11469_;
  assign new_n11472_ = ~new_n11443_ & new_n11469_;
  assign new_n11473_ = ~new_n11471_ & ~new_n11472_;
  assign A5517 = ~new_n11441_ & ~new_n11473_;
  assign new_n11475_ = new_n9359_ & ~new_n9387_;
  assign new_n11476_ = ~new_n9362_ & ~new_n11475_;
  assign new_n11477_ = new_n9404_ & ~new_n9432_;
  assign new_n11478_ = ~new_n9407_ & ~new_n11477_;
  assign new_n11479_ = ~new_n11476_ & new_n11478_;
  assign new_n11480_ = new_n11476_ & ~new_n11478_;
  assign new_n11481_ = ~new_n11479_ & ~new_n11480_;
  assign new_n11482_ = new_n9452_ & ~new_n9480_;
  assign new_n11483_ = ~new_n9455_ & ~new_n11482_;
  assign new_n11484_ = new_n9497_ & ~new_n9525_;
  assign new_n11485_ = ~new_n9500_ & ~new_n11484_;
  assign new_n11486_ = new_n11481_ & ~new_n11485_;
  assign new_n11487_ = new_n9543_ & ~new_n9571_;
  assign new_n11488_ = ~new_n9546_ & ~new_n11487_;
  assign new_n11489_ = ~new_n11485_ & ~new_n11488_;
  assign new_n11490_ = ~new_n11486_ & ~new_n11489_;
  assign new_n11491_ = new_n11483_ & new_n11490_;
  assign new_n11492_ = ~new_n11483_ & ~new_n11490_;
  assign new_n11493_ = ~new_n11491_ & ~new_n11492_;
  assign A5488 = ~new_n11481_ & ~new_n11493_;
  assign new_n11495_ = ~new_n11478_ & ~new_n11491_;
  assign A5487 = ~new_n11481_ & ~new_n11495_;
  assign new_n11497_ = new_n11478_ & new_n11483_;
  assign new_n11498_ = ~new_n11481_ & ~new_n11497_;
  assign new_n11499_ = new_n11481_ & ~new_n11498_;
  assign new_n11500_ = new_n11481_ & new_n11497_;
  assign new_n11501_ = new_n11499_ & ~new_n11500_;
  assign new_n11502_ = new_n11483_ & ~new_n11501_;
  assign A5486 = new_n11490_ | new_n11502_;
  assign new_n11504_ = new_n11485_ & new_n11488_;
  assign new_n11505_ = ~new_n11489_ & ~new_n11504_;
  assign new_n11506_ = ~new_n11481_ & ~new_n11485_;
  assign new_n11507_ = new_n11481_ & new_n11485_;
  assign new_n11508_ = ~new_n11506_ & ~new_n11507_;
  assign new_n11509_ = new_n11505_ & ~new_n11508_;
  assign A5485 = new_n11502_ | new_n11509_;
  assign new_n11511_ = new_n11483_ & ~new_n11509_;
  assign new_n11512_ = ~new_n11483_ & new_n11509_;
  assign new_n11513_ = ~new_n11511_ & ~new_n11512_;
  assign A5484 = ~new_n11481_ & ~new_n11513_;
  assign new_n11515_ = new_n9610_ & ~new_n9638_;
  assign new_n11516_ = ~new_n9613_ & ~new_n11515_;
  assign new_n11517_ = new_n9655_ & ~new_n9683_;
  assign new_n11518_ = ~new_n9658_ & ~new_n11517_;
  assign new_n11519_ = ~new_n11516_ & new_n11518_;
  assign new_n11520_ = new_n11516_ & ~new_n11518_;
  assign new_n11521_ = ~new_n11519_ & ~new_n11520_;
  assign new_n11522_ = new_n9703_ & ~new_n9731_;
  assign new_n11523_ = ~new_n9706_ & ~new_n11522_;
  assign new_n11524_ = new_n9748_ & ~new_n9776_;
  assign new_n11525_ = ~new_n9751_ & ~new_n11524_;
  assign new_n11526_ = new_n11521_ & ~new_n11525_;
  assign new_n11527_ = new_n9794_ & ~new_n9822_;
  assign new_n11528_ = ~new_n9797_ & ~new_n11527_;
  assign new_n11529_ = ~new_n11525_ & ~new_n11528_;
  assign new_n11530_ = ~new_n11526_ & ~new_n11529_;
  assign new_n11531_ = new_n11523_ & new_n11530_;
  assign new_n11532_ = ~new_n11523_ & ~new_n11530_;
  assign new_n11533_ = ~new_n11531_ & ~new_n11532_;
  assign A5455 = ~new_n11521_ & ~new_n11533_;
  assign new_n11535_ = ~new_n11518_ & ~new_n11531_;
  assign A5454 = ~new_n11521_ & ~new_n11535_;
  assign new_n11537_ = new_n11518_ & new_n11523_;
  assign new_n11538_ = ~new_n11521_ & ~new_n11537_;
  assign new_n11539_ = new_n11521_ & ~new_n11538_;
  assign new_n11540_ = new_n11521_ & new_n11537_;
  assign new_n11541_ = new_n11539_ & ~new_n11540_;
  assign new_n11542_ = new_n11523_ & ~new_n11541_;
  assign A5453 = new_n11530_ | new_n11542_;
  assign new_n11544_ = new_n11525_ & new_n11528_;
  assign new_n11545_ = ~new_n11529_ & ~new_n11544_;
  assign new_n11546_ = ~new_n11521_ & ~new_n11525_;
  assign new_n11547_ = new_n11521_ & new_n11525_;
  assign new_n11548_ = ~new_n11546_ & ~new_n11547_;
  assign new_n11549_ = new_n11545_ & ~new_n11548_;
  assign A5452 = new_n11542_ | new_n11549_;
  assign new_n11551_ = new_n11523_ & ~new_n11549_;
  assign new_n11552_ = ~new_n11523_ & new_n11549_;
  assign new_n11553_ = ~new_n11551_ & ~new_n11552_;
  assign A5451 = ~new_n11521_ & ~new_n11553_;
  assign new_n11555_ = ~new_n9859_ & ~new_n9878_;
  assign new_n11556_ = ~new_n9862_ & ~new_n11555_;
  assign new_n11557_ = ~new_n9889_ & ~new_n9908_;
  assign new_n11558_ = ~new_n9892_ & ~new_n11557_;
  assign new_n11559_ = ~new_n11556_ & new_n11558_;
  assign new_n11560_ = new_n11556_ & ~new_n11558_;
  assign new_n11561_ = ~new_n11559_ & ~new_n11560_;
  assign new_n11562_ = ~new_n9922_ & ~new_n9941_;
  assign new_n11563_ = ~new_n9925_ & ~new_n11562_;
  assign new_n11564_ = ~new_n9952_ & ~new_n9971_;
  assign new_n11565_ = ~new_n9955_ & ~new_n11564_;
  assign new_n11566_ = new_n11561_ & ~new_n11565_;
  assign new_n11567_ = ~new_n9983_ & ~new_n10002_;
  assign new_n11568_ = ~new_n9986_ & ~new_n11567_;
  assign new_n11569_ = ~new_n11565_ & ~new_n11568_;
  assign new_n11570_ = ~new_n11566_ & ~new_n11569_;
  assign new_n11571_ = new_n11563_ & new_n11570_;
  assign new_n11572_ = ~new_n11563_ & ~new_n11570_;
  assign new_n11573_ = ~new_n11571_ & ~new_n11572_;
  assign A5422 = ~new_n11561_ & ~new_n11573_;
  assign new_n11575_ = ~new_n11558_ & ~new_n11571_;
  assign A5421 = ~new_n11561_ & ~new_n11575_;
  assign new_n11577_ = new_n11558_ & new_n11563_;
  assign new_n11578_ = ~new_n11561_ & ~new_n11577_;
  assign new_n11579_ = new_n11561_ & ~new_n11578_;
  assign new_n11580_ = new_n11561_ & new_n11577_;
  assign new_n11581_ = new_n11579_ & ~new_n11580_;
  assign new_n11582_ = new_n11563_ & ~new_n11581_;
  assign A5420 = new_n11570_ | new_n11582_;
  assign new_n11584_ = new_n11565_ & new_n11568_;
  assign new_n11585_ = ~new_n11569_ & ~new_n11584_;
  assign new_n11586_ = ~new_n11561_ & ~new_n11565_;
  assign new_n11587_ = new_n11561_ & new_n11565_;
  assign new_n11588_ = ~new_n11586_ & ~new_n11587_;
  assign new_n11589_ = new_n11585_ & ~new_n11588_;
  assign A5419 = new_n11582_ | new_n11589_;
  assign new_n11591_ = new_n11563_ & ~new_n11589_;
  assign new_n11592_ = ~new_n11563_ & new_n11589_;
  assign new_n11593_ = ~new_n11591_ & ~new_n11592_;
  assign A5418 = ~new_n11561_ & ~new_n11593_;
  assign new_n11595_ = ~new_n10039_ & ~new_n10058_;
  assign new_n11596_ = ~new_n10042_ & ~new_n11595_;
  assign new_n11597_ = ~new_n10069_ & ~new_n10088_;
  assign new_n11598_ = ~new_n10072_ & ~new_n11597_;
  assign new_n11599_ = ~new_n11596_ & new_n11598_;
  assign new_n11600_ = new_n11596_ & ~new_n11598_;
  assign new_n11601_ = ~new_n11599_ & ~new_n11600_;
  assign new_n11602_ = ~new_n10102_ & ~new_n10121_;
  assign new_n11603_ = ~new_n10105_ & ~new_n11602_;
  assign new_n11604_ = ~new_n10132_ & ~new_n10151_;
  assign new_n11605_ = ~new_n10135_ & ~new_n11604_;
  assign new_n11606_ = new_n11601_ & ~new_n11605_;
  assign new_n11607_ = ~new_n10163_ & ~new_n10182_;
  assign new_n11608_ = ~new_n10166_ & ~new_n11607_;
  assign new_n11609_ = ~new_n11605_ & ~new_n11608_;
  assign new_n11610_ = ~new_n11606_ & ~new_n11609_;
  assign new_n11611_ = new_n11603_ & new_n11610_;
  assign new_n11612_ = ~new_n11603_ & ~new_n11610_;
  assign new_n11613_ = ~new_n11611_ & ~new_n11612_;
  assign A5389 = ~new_n11601_ & ~new_n11613_;
  assign new_n11615_ = ~new_n11598_ & ~new_n11611_;
  assign A5388 = ~new_n11601_ & ~new_n11615_;
  assign new_n11617_ = new_n11598_ & new_n11603_;
  assign new_n11618_ = ~new_n11601_ & ~new_n11617_;
  assign new_n11619_ = new_n11601_ & ~new_n11618_;
  assign new_n11620_ = new_n11601_ & new_n11617_;
  assign new_n11621_ = new_n11619_ & ~new_n11620_;
  assign new_n11622_ = new_n11603_ & ~new_n11621_;
  assign A5387 = new_n11610_ | new_n11622_;
  assign new_n11624_ = new_n11605_ & new_n11608_;
  assign new_n11625_ = ~new_n11609_ & ~new_n11624_;
  assign new_n11626_ = ~new_n11601_ & ~new_n11605_;
  assign new_n11627_ = new_n11601_ & new_n11605_;
  assign new_n11628_ = ~new_n11626_ & ~new_n11627_;
  assign new_n11629_ = new_n11625_ & ~new_n11628_;
  assign A5386 = new_n11622_ | new_n11629_;
  assign new_n11631_ = new_n11603_ & ~new_n11629_;
  assign new_n11632_ = ~new_n11603_ & new_n11629_;
  assign new_n11633_ = ~new_n11631_ & ~new_n11632_;
  assign A5385 = ~new_n11601_ & ~new_n11633_;
  assign new_n11635_ = ~new_n10219_ & ~new_n10238_;
  assign new_n11636_ = ~new_n10222_ & ~new_n11635_;
  assign new_n11637_ = ~new_n10249_ & ~new_n10268_;
  assign new_n11638_ = ~new_n10252_ & ~new_n11637_;
  assign new_n11639_ = ~new_n11636_ & new_n11638_;
  assign new_n11640_ = new_n11636_ & ~new_n11638_;
  assign new_n11641_ = ~new_n11639_ & ~new_n11640_;
  assign new_n11642_ = ~new_n10282_ & ~new_n10301_;
  assign new_n11643_ = ~new_n10285_ & ~new_n11642_;
  assign new_n11644_ = ~new_n10312_ & ~new_n10331_;
  assign new_n11645_ = ~new_n10315_ & ~new_n11644_;
  assign new_n11646_ = new_n11641_ & ~new_n11645_;
  assign new_n11647_ = ~new_n10343_ & ~new_n10362_;
  assign new_n11648_ = ~new_n10346_ & ~new_n11647_;
  assign new_n11649_ = ~new_n11645_ & ~new_n11648_;
  assign new_n11650_ = ~new_n11646_ & ~new_n11649_;
  assign new_n11651_ = new_n11643_ & new_n11650_;
  assign new_n11652_ = ~new_n11643_ & ~new_n11650_;
  assign new_n11653_ = ~new_n11651_ & ~new_n11652_;
  assign A5356 = ~new_n11641_ & ~new_n11653_;
  assign new_n11655_ = ~new_n11638_ & ~new_n11651_;
  assign A5355 = ~new_n11641_ & ~new_n11655_;
  assign new_n11657_ = new_n11638_ & new_n11643_;
  assign new_n11658_ = ~new_n11641_ & ~new_n11657_;
  assign new_n11659_ = new_n11641_ & ~new_n11658_;
  assign new_n11660_ = new_n11641_ & new_n11657_;
  assign new_n11661_ = new_n11659_ & ~new_n11660_;
  assign new_n11662_ = new_n11643_ & ~new_n11661_;
  assign A5354 = new_n11650_ | new_n11662_;
  assign new_n11664_ = new_n11645_ & new_n11648_;
  assign new_n11665_ = ~new_n11649_ & ~new_n11664_;
  assign new_n11666_ = ~new_n11641_ & ~new_n11645_;
  assign new_n11667_ = new_n11641_ & new_n11645_;
  assign new_n11668_ = ~new_n11666_ & ~new_n11667_;
  assign new_n11669_ = new_n11665_ & ~new_n11668_;
  assign A5353 = new_n11662_ | new_n11669_;
  assign new_n11671_ = new_n11643_ & ~new_n11669_;
  assign new_n11672_ = ~new_n11643_ & new_n11669_;
  assign new_n11673_ = ~new_n11671_ & ~new_n11672_;
  assign A5352 = ~new_n11641_ & ~new_n11673_;
  assign new_n11675_ = ~new_n10399_ & ~new_n10418_;
  assign new_n11676_ = ~new_n10402_ & ~new_n11675_;
  assign new_n11677_ = ~new_n10429_ & ~new_n10448_;
  assign new_n11678_ = ~new_n10432_ & ~new_n11677_;
  assign new_n11679_ = ~new_n11676_ & new_n11678_;
  assign new_n11680_ = new_n11676_ & ~new_n11678_;
  assign new_n11681_ = ~new_n11679_ & ~new_n11680_;
  assign new_n11682_ = ~new_n10462_ & ~new_n10481_;
  assign new_n11683_ = ~new_n10465_ & ~new_n11682_;
  assign new_n11684_ = ~new_n10492_ & ~new_n10511_;
  assign new_n11685_ = ~new_n10495_ & ~new_n11684_;
  assign new_n11686_ = new_n11681_ & ~new_n11685_;
  assign new_n11687_ = ~new_n10523_ & ~new_n10542_;
  assign new_n11688_ = ~new_n10526_ & ~new_n11687_;
  assign new_n11689_ = ~new_n11685_ & ~new_n11688_;
  assign new_n11690_ = ~new_n11686_ & ~new_n11689_;
  assign new_n11691_ = new_n11683_ & new_n11690_;
  assign new_n11692_ = ~new_n11683_ & ~new_n11690_;
  assign new_n11693_ = ~new_n11691_ & ~new_n11692_;
  assign A5323 = ~new_n11681_ & ~new_n11693_;
  assign new_n11695_ = ~new_n11678_ & ~new_n11691_;
  assign A5322 = ~new_n11681_ & ~new_n11695_;
  assign new_n11697_ = new_n11678_ & new_n11683_;
  assign new_n11698_ = ~new_n11681_ & ~new_n11697_;
  assign new_n11699_ = new_n11681_ & ~new_n11698_;
  assign new_n11700_ = new_n11681_ & new_n11697_;
  assign new_n11701_ = new_n11699_ & ~new_n11700_;
  assign new_n11702_ = new_n11683_ & ~new_n11701_;
  assign A5321 = new_n11690_ | new_n11702_;
  assign new_n11704_ = new_n11685_ & new_n11688_;
  assign new_n11705_ = ~new_n11689_ & ~new_n11704_;
  assign new_n11706_ = ~new_n11681_ & ~new_n11685_;
  assign new_n11707_ = new_n11681_ & new_n11685_;
  assign new_n11708_ = ~new_n11706_ & ~new_n11707_;
  assign new_n11709_ = new_n11705_ & ~new_n11708_;
  assign A5320 = new_n11702_ | new_n11709_;
  assign new_n11711_ = new_n11683_ & ~new_n11709_;
  assign new_n11712_ = ~new_n11683_ & new_n11709_;
  assign new_n11713_ = ~new_n11711_ & ~new_n11712_;
  assign A5319 = ~new_n11681_ & ~new_n11713_;
  assign new_n11715_ = new_n10589_ & new_n10600_;
  assign new_n11716_ = ~new_n10592_ & ~new_n11715_;
  assign new_n11717_ = new_n10592_ & ~new_n11716_;
  assign new_n11718_ = new_n10592_ & new_n11715_;
  assign new_n11719_ = new_n11717_ & ~new_n11718_;
  assign new_n11720_ = new_n10600_ & ~new_n11719_;
  assign new_n11721_ = ~new_n10596_ & ~new_n11720_;
  assign new_n11722_ = ~new_n10612_ & ~new_n10631_;
  assign new_n11723_ = ~new_n10615_ & ~new_n11722_;
  assign new_n11724_ = new_n11721_ & new_n11723_;
  assign new_n11725_ = ~new_n11721_ & ~new_n11723_;
  assign new_n11726_ = ~new_n11724_ & ~new_n11725_;
  assign new_n11727_ = ~new_n10645_ & ~new_n10664_;
  assign new_n11728_ = ~new_n10648_ & ~new_n11727_;
  assign new_n11729_ = ~new_n10675_ & ~new_n10694_;
  assign new_n11730_ = ~new_n10678_ & ~new_n11729_;
  assign new_n11731_ = new_n11726_ & ~new_n11730_;
  assign new_n11732_ = ~new_n10706_ & ~new_n10725_;
  assign new_n11733_ = ~new_n10709_ & ~new_n11732_;
  assign new_n11734_ = ~new_n11730_ & ~new_n11733_;
  assign new_n11735_ = ~new_n11731_ & ~new_n11734_;
  assign new_n11736_ = new_n11728_ & new_n11735_;
  assign new_n11737_ = ~new_n11728_ & ~new_n11735_;
  assign new_n11738_ = ~new_n11736_ & ~new_n11737_;
  assign A5290 = ~new_n11726_ & ~new_n11738_;
  assign new_n11740_ = ~new_n11723_ & ~new_n11736_;
  assign A5289 = ~new_n11726_ & ~new_n11740_;
  assign new_n11742_ = new_n11723_ & new_n11728_;
  assign new_n11743_ = ~new_n11726_ & ~new_n11742_;
  assign new_n11744_ = new_n11726_ & ~new_n11743_;
  assign new_n11745_ = new_n11726_ & new_n11742_;
  assign new_n11746_ = new_n11744_ & ~new_n11745_;
  assign new_n11747_ = new_n11728_ & ~new_n11746_;
  assign A5288 = new_n11735_ | new_n11747_;
  assign new_n11749_ = new_n11730_ & new_n11733_;
  assign new_n11750_ = ~new_n11734_ & ~new_n11749_;
  assign new_n11751_ = ~new_n11726_ & ~new_n11730_;
  assign new_n11752_ = new_n11726_ & new_n11730_;
  assign new_n11753_ = ~new_n11751_ & ~new_n11752_;
  assign new_n11754_ = new_n11750_ & ~new_n11753_;
  assign A5287 = new_n11747_ | new_n11754_;
  assign new_n11756_ = new_n11728_ & ~new_n11754_;
  assign new_n11757_ = ~new_n11728_ & new_n11754_;
  assign new_n11758_ = ~new_n11756_ & ~new_n11757_;
  assign A5286 = ~new_n11726_ & ~new_n11758_;
  assign new_n11760_ = new_n1374_ & new_n1437_;
  assign new_n11761_ = ~new_n1377_ & ~new_n11760_;
  assign new_n11762_ = new_n1377_ & ~new_n11761_;
  assign new_n11763_ = new_n1377_ & new_n11760_;
  assign new_n11764_ = new_n11762_ & ~new_n11763_;
  assign new_n11765_ = new_n1437_ & ~new_n11764_;
  assign new_n11766_ = ~new_n1560_ & ~new_n11765_;
  assign new_n11767_ = new_n1684_ & new_n1747_;
  assign new_n11768_ = ~new_n1687_ & ~new_n11767_;
  assign new_n11769_ = new_n1687_ & ~new_n11768_;
  assign new_n11770_ = new_n1687_ & new_n11767_;
  assign new_n11771_ = new_n11769_ & ~new_n11770_;
  assign new_n11772_ = new_n1747_ & ~new_n11771_;
  assign new_n11773_ = ~new_n1870_ & ~new_n11772_;
  assign new_n11774_ = new_n11766_ & ~new_n11773_;
  assign new_n11775_ = ~new_n11766_ & new_n11773_;
  assign new_n11776_ = ~new_n11774_ & ~new_n11775_;
  assign new_n11777_ = new_n1997_ & new_n2060_;
  assign new_n11778_ = ~new_n2000_ & ~new_n11777_;
  assign new_n11779_ = new_n2000_ & ~new_n11778_;
  assign new_n11780_ = new_n2000_ & new_n11777_;
  assign new_n11781_ = new_n11779_ & ~new_n11780_;
  assign new_n11782_ = new_n2060_ & ~new_n11781_;
  assign new_n11783_ = ~new_n2183_ & ~new_n11782_;
  assign new_n11784_ = new_n2307_ & new_n2370_;
  assign new_n11785_ = ~new_n2310_ & ~new_n11784_;
  assign new_n11786_ = new_n2310_ & ~new_n11785_;
  assign new_n11787_ = new_n2310_ & new_n11784_;
  assign new_n11788_ = new_n11786_ & ~new_n11787_;
  assign new_n11789_ = new_n2370_ & ~new_n11788_;
  assign new_n11790_ = ~new_n2493_ & ~new_n11789_;
  assign new_n11791_ = new_n11776_ & new_n11790_;
  assign new_n11792_ = new_n2618_ & new_n2681_;
  assign new_n11793_ = ~new_n2621_ & ~new_n11792_;
  assign new_n11794_ = new_n2621_ & ~new_n11793_;
  assign new_n11795_ = new_n2621_ & new_n11792_;
  assign new_n11796_ = new_n11794_ & ~new_n11795_;
  assign new_n11797_ = new_n2681_ & ~new_n11796_;
  assign new_n11798_ = ~new_n2804_ & ~new_n11797_;
  assign new_n11799_ = new_n11790_ & new_n11798_;
  assign new_n11800_ = ~new_n11791_ & ~new_n11799_;
  assign new_n11801_ = ~new_n11783_ & new_n11800_;
  assign new_n11802_ = new_n11783_ & ~new_n11800_;
  assign new_n11803_ = ~new_n11801_ & ~new_n11802_;
  assign A5257 = ~new_n11776_ & ~new_n11803_;
  assign new_n11805_ = new_n11773_ & ~new_n11801_;
  assign A5256 = ~new_n11776_ & ~new_n11805_;
  assign new_n11807_ = ~new_n11773_ & ~new_n11783_;
  assign new_n11808_ = ~new_n11776_ & ~new_n11807_;
  assign new_n11809_ = new_n11776_ & ~new_n11808_;
  assign new_n11810_ = new_n11776_ & new_n11807_;
  assign new_n11811_ = new_n11809_ & ~new_n11810_;
  assign new_n11812_ = ~new_n11783_ & ~new_n11811_;
  assign A5255 = new_n11800_ | new_n11812_;
  assign new_n11814_ = ~new_n11790_ & ~new_n11798_;
  assign new_n11815_ = ~new_n11799_ & ~new_n11814_;
  assign new_n11816_ = ~new_n11776_ & new_n11790_;
  assign new_n11817_ = new_n11776_ & ~new_n11790_;
  assign new_n11818_ = ~new_n11816_ & ~new_n11817_;
  assign new_n11819_ = new_n11815_ & ~new_n11818_;
  assign A5254 = new_n11812_ | new_n11819_;
  assign new_n11821_ = ~new_n11783_ & ~new_n11819_;
  assign new_n11822_ = new_n11783_ & new_n11819_;
  assign new_n11823_ = ~new_n11821_ & ~new_n11822_;
  assign A5253 = ~new_n11776_ & ~new_n11823_;
  assign new_n11825_ = new_n2879_ & new_n2902_;
  assign new_n11826_ = ~new_n2882_ & ~new_n11825_;
  assign new_n11827_ = new_n2882_ & ~new_n11826_;
  assign new_n11828_ = new_n2882_ & new_n11825_;
  assign new_n11829_ = new_n11827_ & ~new_n11828_;
  assign new_n11830_ = new_n2902_ & ~new_n11829_;
  assign new_n11831_ = ~new_n2945_ & ~new_n11830_;
  assign new_n11832_ = new_n2989_ & new_n3012_;
  assign new_n11833_ = ~new_n2992_ & ~new_n11832_;
  assign new_n11834_ = new_n2992_ & ~new_n11833_;
  assign new_n11835_ = new_n2992_ & new_n11832_;
  assign new_n11836_ = new_n11834_ & ~new_n11835_;
  assign new_n11837_ = new_n3012_ & ~new_n11836_;
  assign new_n11838_ = ~new_n3055_ & ~new_n11837_;
  assign new_n11839_ = new_n11831_ & ~new_n11838_;
  assign new_n11840_ = ~new_n11831_ & new_n11838_;
  assign new_n11841_ = ~new_n11839_ & ~new_n11840_;
  assign new_n11842_ = new_n3102_ & new_n3125_;
  assign new_n11843_ = ~new_n3105_ & ~new_n11842_;
  assign new_n11844_ = new_n3105_ & ~new_n11843_;
  assign new_n11845_ = new_n3105_ & new_n11842_;
  assign new_n11846_ = new_n11844_ & ~new_n11845_;
  assign new_n11847_ = new_n3125_ & ~new_n11846_;
  assign new_n11848_ = ~new_n3168_ & ~new_n11847_;
  assign new_n11849_ = new_n3212_ & new_n3235_;
  assign new_n11850_ = ~new_n3215_ & ~new_n11849_;
  assign new_n11851_ = new_n3215_ & ~new_n11850_;
  assign new_n11852_ = new_n3215_ & new_n11849_;
  assign new_n11853_ = new_n11851_ & ~new_n11852_;
  assign new_n11854_ = new_n3235_ & ~new_n11853_;
  assign new_n11855_ = ~new_n3278_ & ~new_n11854_;
  assign new_n11856_ = new_n11841_ & new_n11855_;
  assign new_n11857_ = new_n3323_ & new_n3346_;
  assign new_n11858_ = ~new_n3326_ & ~new_n11857_;
  assign new_n11859_ = new_n3326_ & ~new_n11858_;
  assign new_n11860_ = new_n3326_ & new_n11857_;
  assign new_n11861_ = new_n11859_ & ~new_n11860_;
  assign new_n11862_ = new_n3346_ & ~new_n11861_;
  assign new_n11863_ = ~new_n3389_ & ~new_n11862_;
  assign new_n11864_ = new_n11855_ & new_n11863_;
  assign new_n11865_ = ~new_n11856_ & ~new_n11864_;
  assign new_n11866_ = ~new_n11848_ & new_n11865_;
  assign new_n11867_ = new_n11848_ & ~new_n11865_;
  assign new_n11868_ = ~new_n11866_ & ~new_n11867_;
  assign A5224 = ~new_n11841_ & ~new_n11868_;
  assign new_n11870_ = new_n11838_ & ~new_n11866_;
  assign A5223 = ~new_n11841_ & ~new_n11870_;
  assign new_n11872_ = ~new_n11838_ & ~new_n11848_;
  assign new_n11873_ = ~new_n11841_ & ~new_n11872_;
  assign new_n11874_ = new_n11841_ & ~new_n11873_;
  assign new_n11875_ = new_n11841_ & new_n11872_;
  assign new_n11876_ = new_n11874_ & ~new_n11875_;
  assign new_n11877_ = ~new_n11848_ & ~new_n11876_;
  assign A5222 = new_n11865_ | new_n11877_;
  assign new_n11879_ = ~new_n11855_ & ~new_n11863_;
  assign new_n11880_ = ~new_n11864_ & ~new_n11879_;
  assign new_n11881_ = ~new_n11841_ & new_n11855_;
  assign new_n11882_ = new_n11841_ & ~new_n11855_;
  assign new_n11883_ = ~new_n11881_ & ~new_n11882_;
  assign new_n11884_ = new_n11880_ & ~new_n11883_;
  assign A5221 = new_n11877_ | new_n11884_;
  assign new_n11886_ = ~new_n11848_ & ~new_n11884_;
  assign new_n11887_ = new_n11848_ & new_n11884_;
  assign new_n11888_ = ~new_n11886_ & ~new_n11887_;
  assign A5220 = ~new_n11841_ & ~new_n11888_;
  assign new_n11890_ = new_n3505_ & new_n3553_;
  assign new_n11891_ = ~new_n3508_ & ~new_n11890_;
  assign new_n11892_ = new_n3508_ & ~new_n11891_;
  assign new_n11893_ = new_n3508_ & new_n11890_;
  assign new_n11894_ = new_n11892_ & ~new_n11893_;
  assign new_n11895_ = new_n3553_ & ~new_n11894_;
  assign new_n11896_ = ~new_n3646_ & ~new_n11895_;
  assign new_n11897_ = new_n3740_ & new_n3788_;
  assign new_n11898_ = ~new_n3743_ & ~new_n11897_;
  assign new_n11899_ = new_n3743_ & ~new_n11898_;
  assign new_n11900_ = new_n3743_ & new_n11897_;
  assign new_n11901_ = new_n11899_ & ~new_n11900_;
  assign new_n11902_ = new_n3788_ & ~new_n11901_;
  assign new_n11903_ = ~new_n3881_ & ~new_n11902_;
  assign new_n11904_ = new_n11896_ & ~new_n11903_;
  assign new_n11905_ = ~new_n11896_ & new_n11903_;
  assign new_n11906_ = ~new_n11904_ & ~new_n11905_;
  assign new_n11907_ = new_n3978_ & new_n4026_;
  assign new_n11908_ = ~new_n3981_ & ~new_n11907_;
  assign new_n11909_ = new_n3981_ & ~new_n11908_;
  assign new_n11910_ = new_n3981_ & new_n11907_;
  assign new_n11911_ = new_n11909_ & ~new_n11910_;
  assign new_n11912_ = new_n4026_ & ~new_n11911_;
  assign new_n11913_ = ~new_n4119_ & ~new_n11912_;
  assign new_n11914_ = new_n4213_ & new_n4261_;
  assign new_n11915_ = ~new_n4216_ & ~new_n11914_;
  assign new_n11916_ = new_n4216_ & ~new_n11915_;
  assign new_n11917_ = new_n4216_ & new_n11914_;
  assign new_n11918_ = new_n11916_ & ~new_n11917_;
  assign new_n11919_ = new_n4261_ & ~new_n11918_;
  assign new_n11920_ = ~new_n4354_ & ~new_n11919_;
  assign new_n11921_ = new_n11906_ & new_n11920_;
  assign new_n11922_ = new_n4449_ & new_n4497_;
  assign new_n11923_ = ~new_n4452_ & ~new_n11922_;
  assign new_n11924_ = new_n4452_ & ~new_n11923_;
  assign new_n11925_ = new_n4452_ & new_n11922_;
  assign new_n11926_ = new_n11924_ & ~new_n11925_;
  assign new_n11927_ = new_n4497_ & ~new_n11926_;
  assign new_n11928_ = ~new_n4590_ & ~new_n11927_;
  assign new_n11929_ = new_n11920_ & new_n11928_;
  assign new_n11930_ = ~new_n11921_ & ~new_n11929_;
  assign new_n11931_ = ~new_n11913_ & new_n11930_;
  assign new_n11932_ = new_n11913_ & ~new_n11930_;
  assign new_n11933_ = ~new_n11931_ & ~new_n11932_;
  assign A5191 = ~new_n11906_ & ~new_n11933_;
  assign new_n11935_ = new_n11903_ & ~new_n11931_;
  assign A5190 = ~new_n11906_ & ~new_n11935_;
  assign new_n11937_ = ~new_n11903_ & ~new_n11913_;
  assign new_n11938_ = ~new_n11906_ & ~new_n11937_;
  assign new_n11939_ = new_n11906_ & ~new_n11938_;
  assign new_n11940_ = new_n11906_ & new_n11937_;
  assign new_n11941_ = new_n11939_ & ~new_n11940_;
  assign new_n11942_ = ~new_n11913_ & ~new_n11941_;
  assign A5189 = new_n11930_ | new_n11942_;
  assign new_n11944_ = ~new_n11920_ & ~new_n11928_;
  assign new_n11945_ = ~new_n11929_ & ~new_n11944_;
  assign new_n11946_ = ~new_n11906_ & new_n11920_;
  assign new_n11947_ = new_n11906_ & ~new_n11920_;
  assign new_n11948_ = ~new_n11946_ & ~new_n11947_;
  assign new_n11949_ = new_n11945_ & ~new_n11948_;
  assign A5188 = new_n11942_ | new_n11949_;
  assign new_n11951_ = ~new_n11913_ & ~new_n11949_;
  assign new_n11952_ = new_n11913_ & new_n11949_;
  assign new_n11953_ = ~new_n11951_ & ~new_n11952_;
  assign A5187 = ~new_n11906_ & ~new_n11953_;
  assign new_n11955_ = new_n4706_ & new_n4754_;
  assign new_n11956_ = ~new_n4709_ & ~new_n11955_;
  assign new_n11957_ = new_n4709_ & ~new_n11956_;
  assign new_n11958_ = new_n4709_ & new_n11955_;
  assign new_n11959_ = new_n11957_ & ~new_n11958_;
  assign new_n11960_ = new_n4754_ & ~new_n11959_;
  assign new_n11961_ = ~new_n4847_ & ~new_n11960_;
  assign new_n11962_ = new_n4941_ & new_n4989_;
  assign new_n11963_ = ~new_n4944_ & ~new_n11962_;
  assign new_n11964_ = new_n4944_ & ~new_n11963_;
  assign new_n11965_ = new_n4944_ & new_n11962_;
  assign new_n11966_ = new_n11964_ & ~new_n11965_;
  assign new_n11967_ = new_n4989_ & ~new_n11966_;
  assign new_n11968_ = ~new_n5082_ & ~new_n11967_;
  assign new_n11969_ = new_n11961_ & ~new_n11968_;
  assign new_n11970_ = ~new_n11961_ & new_n11968_;
  assign new_n11971_ = ~new_n11969_ & ~new_n11970_;
  assign new_n11972_ = new_n5179_ & new_n5227_;
  assign new_n11973_ = ~new_n5182_ & ~new_n11972_;
  assign new_n11974_ = new_n5182_ & ~new_n11973_;
  assign new_n11975_ = new_n5182_ & new_n11972_;
  assign new_n11976_ = new_n11974_ & ~new_n11975_;
  assign new_n11977_ = new_n5227_ & ~new_n11976_;
  assign new_n11978_ = ~new_n5320_ & ~new_n11977_;
  assign new_n11979_ = new_n5414_ & new_n5462_;
  assign new_n11980_ = ~new_n5417_ & ~new_n11979_;
  assign new_n11981_ = new_n5417_ & ~new_n11980_;
  assign new_n11982_ = new_n5417_ & new_n11979_;
  assign new_n11983_ = new_n11981_ & ~new_n11982_;
  assign new_n11984_ = new_n5462_ & ~new_n11983_;
  assign new_n11985_ = ~new_n5555_ & ~new_n11984_;
  assign new_n11986_ = new_n11971_ & new_n11985_;
  assign new_n11987_ = new_n5650_ & new_n5698_;
  assign new_n11988_ = ~new_n5653_ & ~new_n11987_;
  assign new_n11989_ = new_n5653_ & ~new_n11988_;
  assign new_n11990_ = new_n5653_ & new_n11987_;
  assign new_n11991_ = new_n11989_ & ~new_n11990_;
  assign new_n11992_ = new_n5698_ & ~new_n11991_;
  assign new_n11993_ = ~new_n5791_ & ~new_n11992_;
  assign new_n11994_ = new_n11985_ & new_n11993_;
  assign new_n11995_ = ~new_n11986_ & ~new_n11994_;
  assign new_n11996_ = ~new_n11978_ & new_n11995_;
  assign new_n11997_ = new_n11978_ & ~new_n11995_;
  assign new_n11998_ = ~new_n11996_ & ~new_n11997_;
  assign A5158 = ~new_n11971_ & ~new_n11998_;
  assign new_n12000_ = new_n11968_ & ~new_n11996_;
  assign A5157 = ~new_n11971_ & ~new_n12000_;
  assign new_n12002_ = ~new_n11968_ & ~new_n11978_;
  assign new_n12003_ = ~new_n11971_ & ~new_n12002_;
  assign new_n12004_ = new_n11971_ & ~new_n12003_;
  assign new_n12005_ = new_n11971_ & new_n12002_;
  assign new_n12006_ = new_n12004_ & ~new_n12005_;
  assign new_n12007_ = ~new_n11978_ & ~new_n12006_;
  assign A5156 = new_n11995_ | new_n12007_;
  assign new_n12009_ = ~new_n11985_ & ~new_n11993_;
  assign new_n12010_ = ~new_n11994_ & ~new_n12009_;
  assign new_n12011_ = ~new_n11971_ & new_n11985_;
  assign new_n12012_ = new_n11971_ & ~new_n11985_;
  assign new_n12013_ = ~new_n12011_ & ~new_n12012_;
  assign new_n12014_ = new_n12010_ & ~new_n12013_;
  assign A5155 = new_n12007_ | new_n12014_;
  assign new_n12016_ = ~new_n11978_ & ~new_n12014_;
  assign new_n12017_ = new_n11978_ & new_n12014_;
  assign new_n12018_ = ~new_n12016_ & ~new_n12017_;
  assign A5154 = ~new_n11971_ & ~new_n12018_;
  assign new_n12020_ = new_n5884_ & new_n5917_;
  assign new_n12021_ = ~new_n5887_ & ~new_n12020_;
  assign new_n12022_ = new_n5887_ & ~new_n12021_;
  assign new_n12023_ = new_n5887_ & new_n12020_;
  assign new_n12024_ = new_n12022_ & ~new_n12023_;
  assign new_n12025_ = new_n5917_ & ~new_n12024_;
  assign new_n12026_ = ~new_n5980_ & ~new_n12025_;
  assign new_n12027_ = new_n6044_ & new_n6077_;
  assign new_n12028_ = ~new_n6047_ & ~new_n12027_;
  assign new_n12029_ = new_n6047_ & ~new_n12028_;
  assign new_n12030_ = new_n6047_ & new_n12027_;
  assign new_n12031_ = new_n12029_ & ~new_n12030_;
  assign new_n12032_ = new_n6077_ & ~new_n12031_;
  assign new_n12033_ = ~new_n6140_ & ~new_n12032_;
  assign new_n12034_ = new_n12026_ & ~new_n12033_;
  assign new_n12035_ = ~new_n12026_ & new_n12033_;
  assign new_n12036_ = ~new_n12034_ & ~new_n12035_;
  assign new_n12037_ = new_n6207_ & new_n6240_;
  assign new_n12038_ = ~new_n6210_ & ~new_n12037_;
  assign new_n12039_ = new_n6210_ & ~new_n12038_;
  assign new_n12040_ = new_n6210_ & new_n12037_;
  assign new_n12041_ = new_n12039_ & ~new_n12040_;
  assign new_n12042_ = new_n6240_ & ~new_n12041_;
  assign new_n12043_ = ~new_n6303_ & ~new_n12042_;
  assign new_n12044_ = new_n6367_ & new_n6400_;
  assign new_n12045_ = ~new_n6370_ & ~new_n12044_;
  assign new_n12046_ = new_n6370_ & ~new_n12045_;
  assign new_n12047_ = new_n6370_ & new_n12044_;
  assign new_n12048_ = new_n12046_ & ~new_n12047_;
  assign new_n12049_ = new_n6400_ & ~new_n12048_;
  assign new_n12050_ = ~new_n6463_ & ~new_n12049_;
  assign new_n12051_ = new_n12036_ & new_n12050_;
  assign new_n12052_ = new_n6528_ & new_n6561_;
  assign new_n12053_ = ~new_n6531_ & ~new_n12052_;
  assign new_n12054_ = new_n6531_ & ~new_n12053_;
  assign new_n12055_ = new_n6531_ & new_n12052_;
  assign new_n12056_ = new_n12054_ & ~new_n12055_;
  assign new_n12057_ = new_n6561_ & ~new_n12056_;
  assign new_n12058_ = ~new_n6624_ & ~new_n12057_;
  assign new_n12059_ = new_n12050_ & new_n12058_;
  assign new_n12060_ = ~new_n12051_ & ~new_n12059_;
  assign new_n12061_ = ~new_n12043_ & new_n12060_;
  assign new_n12062_ = new_n12043_ & ~new_n12060_;
  assign new_n12063_ = ~new_n12061_ & ~new_n12062_;
  assign A5125 = ~new_n12036_ & ~new_n12063_;
  assign new_n12065_ = new_n12033_ & ~new_n12061_;
  assign A5124 = ~new_n12036_ & ~new_n12065_;
  assign new_n12067_ = ~new_n12033_ & ~new_n12043_;
  assign new_n12068_ = ~new_n12036_ & ~new_n12067_;
  assign new_n12069_ = new_n12036_ & ~new_n12068_;
  assign new_n12070_ = new_n12036_ & new_n12067_;
  assign new_n12071_ = new_n12069_ & ~new_n12070_;
  assign new_n12072_ = ~new_n12043_ & ~new_n12071_;
  assign A5123 = new_n12060_ | new_n12072_;
  assign new_n12074_ = ~new_n12050_ & ~new_n12058_;
  assign new_n12075_ = ~new_n12059_ & ~new_n12074_;
  assign new_n12076_ = ~new_n12036_ & new_n12050_;
  assign new_n12077_ = new_n12036_ & ~new_n12050_;
  assign new_n12078_ = ~new_n12076_ & ~new_n12077_;
  assign new_n12079_ = new_n12075_ & ~new_n12078_;
  assign A5122 = new_n12072_ | new_n12079_;
  assign new_n12081_ = ~new_n12043_ & ~new_n12079_;
  assign new_n12082_ = new_n12043_ & new_n12079_;
  assign new_n12083_ = ~new_n12081_ & ~new_n12082_;
  assign A5121 = ~new_n12036_ & ~new_n12083_;
  assign new_n12085_ = new_n6658_ & new_n6663_;
  assign new_n12086_ = ~new_n6661_ & ~new_n12085_;
  assign new_n12087_ = new_n6661_ & ~new_n12086_;
  assign new_n12088_ = new_n6661_ & new_n12085_;
  assign new_n12089_ = new_n12087_ & ~new_n12088_;
  assign new_n12090_ = new_n6663_ & ~new_n12089_;
  assign new_n12091_ = ~new_n6670_ & ~new_n12090_;
  assign new_n12092_ = new_n6678_ & new_n6683_;
  assign new_n12093_ = ~new_n6681_ & ~new_n12092_;
  assign new_n12094_ = new_n6681_ & ~new_n12093_;
  assign new_n12095_ = new_n6681_ & new_n12092_;
  assign new_n12096_ = new_n12094_ & ~new_n12095_;
  assign new_n12097_ = new_n6683_ & ~new_n12096_;
  assign new_n12098_ = ~new_n6690_ & ~new_n12097_;
  assign new_n12099_ = new_n12091_ & ~new_n12098_;
  assign new_n12100_ = ~new_n12091_ & new_n12098_;
  assign new_n12101_ = ~new_n12099_ & ~new_n12100_;
  assign new_n12102_ = new_n6701_ & new_n6706_;
  assign new_n12103_ = ~new_n6704_ & ~new_n12102_;
  assign new_n12104_ = new_n6704_ & ~new_n12103_;
  assign new_n12105_ = new_n6704_ & new_n12102_;
  assign new_n12106_ = new_n12104_ & ~new_n12105_;
  assign new_n12107_ = new_n6706_ & ~new_n12106_;
  assign new_n12108_ = ~new_n6713_ & ~new_n12107_;
  assign new_n12109_ = new_n6721_ & new_n6726_;
  assign new_n12110_ = ~new_n6724_ & ~new_n12109_;
  assign new_n12111_ = new_n6724_ & ~new_n12110_;
  assign new_n12112_ = new_n6724_ & new_n12109_;
  assign new_n12113_ = new_n12111_ & ~new_n12112_;
  assign new_n12114_ = new_n6726_ & ~new_n12113_;
  assign new_n12115_ = ~new_n6733_ & ~new_n12114_;
  assign new_n12116_ = new_n12101_ & new_n12115_;
  assign new_n12117_ = new_n6742_ & new_n6747_;
  assign new_n12118_ = ~new_n6745_ & ~new_n12117_;
  assign new_n12119_ = new_n6745_ & ~new_n12118_;
  assign new_n12120_ = new_n6745_ & new_n12117_;
  assign new_n12121_ = new_n12119_ & ~new_n12120_;
  assign new_n12122_ = new_n6747_ & ~new_n12121_;
  assign new_n12123_ = ~new_n6754_ & ~new_n12122_;
  assign new_n12124_ = new_n12115_ & new_n12123_;
  assign new_n12125_ = ~new_n12116_ & ~new_n12124_;
  assign new_n12126_ = ~new_n12108_ & new_n12125_;
  assign new_n12127_ = new_n12108_ & ~new_n12125_;
  assign new_n12128_ = ~new_n12126_ & ~new_n12127_;
  assign A5092 = ~new_n12101_ & ~new_n12128_;
  assign new_n12130_ = new_n12098_ & ~new_n12126_;
  assign A5091 = ~new_n12101_ & ~new_n12130_;
  assign new_n12132_ = ~new_n12098_ & ~new_n12108_;
  assign new_n12133_ = ~new_n12101_ & ~new_n12132_;
  assign new_n12134_ = new_n12101_ & ~new_n12133_;
  assign new_n12135_ = new_n12101_ & new_n12132_;
  assign new_n12136_ = new_n12134_ & ~new_n12135_;
  assign new_n12137_ = ~new_n12108_ & ~new_n12136_;
  assign A5090 = new_n12125_ | new_n12137_;
  assign new_n12139_ = ~new_n12115_ & ~new_n12123_;
  assign new_n12140_ = ~new_n12124_ & ~new_n12139_;
  assign new_n12141_ = ~new_n12101_ & new_n12115_;
  assign new_n12142_ = new_n12101_ & ~new_n12115_;
  assign new_n12143_ = ~new_n12141_ & ~new_n12142_;
  assign new_n12144_ = new_n12140_ & ~new_n12143_;
  assign A5089 = new_n12137_ | new_n12144_;
  assign new_n12146_ = ~new_n12108_ & ~new_n12144_;
  assign new_n12147_ = new_n12108_ & new_n12144_;
  assign new_n12148_ = ~new_n12146_ & ~new_n12147_;
  assign A5088 = ~new_n12101_ & ~new_n12148_;
  assign new_n12150_ = new_n6788_ & new_n6793_;
  assign new_n12151_ = ~new_n6791_ & ~new_n12150_;
  assign new_n12152_ = new_n6791_ & ~new_n12151_;
  assign new_n12153_ = new_n6791_ & new_n12150_;
  assign new_n12154_ = new_n12152_ & ~new_n12153_;
  assign new_n12155_ = new_n6793_ & ~new_n12154_;
  assign new_n12156_ = ~new_n6800_ & ~new_n12155_;
  assign new_n12157_ = new_n6808_ & new_n6813_;
  assign new_n12158_ = ~new_n6811_ & ~new_n12157_;
  assign new_n12159_ = new_n6811_ & ~new_n12158_;
  assign new_n12160_ = new_n6811_ & new_n12157_;
  assign new_n12161_ = new_n12159_ & ~new_n12160_;
  assign new_n12162_ = new_n6813_ & ~new_n12161_;
  assign new_n12163_ = ~new_n6820_ & ~new_n12162_;
  assign new_n12164_ = new_n12156_ & ~new_n12163_;
  assign new_n12165_ = ~new_n12156_ & new_n12163_;
  assign new_n12166_ = ~new_n12164_ & ~new_n12165_;
  assign new_n12167_ = new_n6831_ & new_n6836_;
  assign new_n12168_ = ~new_n6834_ & ~new_n12167_;
  assign new_n12169_ = new_n6834_ & ~new_n12168_;
  assign new_n12170_ = new_n6834_ & new_n12167_;
  assign new_n12171_ = new_n12169_ & ~new_n12170_;
  assign new_n12172_ = new_n6836_ & ~new_n12171_;
  assign new_n12173_ = ~new_n6843_ & ~new_n12172_;
  assign new_n12174_ = new_n6851_ & new_n6856_;
  assign new_n12175_ = ~new_n6854_ & ~new_n12174_;
  assign new_n12176_ = new_n6854_ & ~new_n12175_;
  assign new_n12177_ = new_n6854_ & new_n12174_;
  assign new_n12178_ = new_n12176_ & ~new_n12177_;
  assign new_n12179_ = new_n6856_ & ~new_n12178_;
  assign new_n12180_ = ~new_n6863_ & ~new_n12179_;
  assign new_n12181_ = new_n12166_ & new_n12180_;
  assign new_n12182_ = new_n6872_ & new_n6877_;
  assign new_n12183_ = ~new_n6875_ & ~new_n12182_;
  assign new_n12184_ = new_n6875_ & ~new_n12183_;
  assign new_n12185_ = new_n6875_ & new_n12182_;
  assign new_n12186_ = new_n12184_ & ~new_n12185_;
  assign new_n12187_ = new_n6877_ & ~new_n12186_;
  assign new_n12188_ = ~new_n6884_ & ~new_n12187_;
  assign new_n12189_ = new_n12180_ & new_n12188_;
  assign new_n12190_ = ~new_n12181_ & ~new_n12189_;
  assign new_n12191_ = ~new_n12173_ & new_n12190_;
  assign new_n12192_ = new_n12173_ & ~new_n12190_;
  assign new_n12193_ = ~new_n12191_ & ~new_n12192_;
  assign A5059 = ~new_n12166_ & ~new_n12193_;
  assign new_n12195_ = new_n12163_ & ~new_n12191_;
  assign A5058 = ~new_n12166_ & ~new_n12195_;
  assign new_n12197_ = ~new_n12163_ & ~new_n12173_;
  assign new_n12198_ = ~new_n12166_ & ~new_n12197_;
  assign new_n12199_ = new_n12166_ & ~new_n12198_;
  assign new_n12200_ = new_n12166_ & new_n12197_;
  assign new_n12201_ = new_n12199_ & ~new_n12200_;
  assign new_n12202_ = ~new_n12173_ & ~new_n12201_;
  assign A5057 = new_n12190_ | new_n12202_;
  assign new_n12204_ = ~new_n12180_ & ~new_n12188_;
  assign new_n12205_ = ~new_n12189_ & ~new_n12204_;
  assign new_n12206_ = ~new_n12166_ & new_n12180_;
  assign new_n12207_ = new_n12166_ & ~new_n12180_;
  assign new_n12208_ = ~new_n12206_ & ~new_n12207_;
  assign new_n12209_ = new_n12205_ & ~new_n12208_;
  assign A5056 = new_n12202_ | new_n12209_;
  assign new_n12211_ = ~new_n12173_ & ~new_n12209_;
  assign new_n12212_ = new_n12173_ & new_n12209_;
  assign new_n12213_ = ~new_n12211_ & ~new_n12212_;
  assign A5055 = ~new_n12166_ & ~new_n12213_;
  assign new_n12215_ = new_n6918_ & new_n6923_;
  assign new_n12216_ = ~new_n6921_ & ~new_n12215_;
  assign new_n12217_ = new_n6921_ & ~new_n12216_;
  assign new_n12218_ = new_n6921_ & new_n12215_;
  assign new_n12219_ = new_n12217_ & ~new_n12218_;
  assign new_n12220_ = new_n6923_ & ~new_n12219_;
  assign new_n12221_ = ~new_n6930_ & ~new_n12220_;
  assign new_n12222_ = new_n6938_ & new_n6943_;
  assign new_n12223_ = ~new_n6941_ & ~new_n12222_;
  assign new_n12224_ = new_n6941_ & ~new_n12223_;
  assign new_n12225_ = new_n6941_ & new_n12222_;
  assign new_n12226_ = new_n12224_ & ~new_n12225_;
  assign new_n12227_ = new_n6943_ & ~new_n12226_;
  assign new_n12228_ = ~new_n6950_ & ~new_n12227_;
  assign new_n12229_ = new_n12221_ & ~new_n12228_;
  assign new_n12230_ = ~new_n12221_ & new_n12228_;
  assign new_n12231_ = ~new_n12229_ & ~new_n12230_;
  assign new_n12232_ = new_n6961_ & new_n6966_;
  assign new_n12233_ = ~new_n6964_ & ~new_n12232_;
  assign new_n12234_ = new_n6964_ & ~new_n12233_;
  assign new_n12235_ = new_n6964_ & new_n12232_;
  assign new_n12236_ = new_n12234_ & ~new_n12235_;
  assign new_n12237_ = new_n6966_ & ~new_n12236_;
  assign new_n12238_ = ~new_n6973_ & ~new_n12237_;
  assign new_n12239_ = new_n6981_ & new_n6986_;
  assign new_n12240_ = ~new_n6984_ & ~new_n12239_;
  assign new_n12241_ = new_n6984_ & ~new_n12240_;
  assign new_n12242_ = new_n6984_ & new_n12239_;
  assign new_n12243_ = new_n12241_ & ~new_n12242_;
  assign new_n12244_ = new_n6986_ & ~new_n12243_;
  assign new_n12245_ = ~new_n6993_ & ~new_n12244_;
  assign new_n12246_ = new_n12231_ & new_n12245_;
  assign new_n12247_ = new_n7002_ & new_n7007_;
  assign new_n12248_ = ~new_n7005_ & ~new_n12247_;
  assign new_n12249_ = new_n7005_ & ~new_n12248_;
  assign new_n12250_ = new_n7005_ & new_n12247_;
  assign new_n12251_ = new_n12249_ & ~new_n12250_;
  assign new_n12252_ = new_n7007_ & ~new_n12251_;
  assign new_n12253_ = ~new_n7014_ & ~new_n12252_;
  assign new_n12254_ = new_n12245_ & new_n12253_;
  assign new_n12255_ = ~new_n12246_ & ~new_n12254_;
  assign new_n12256_ = ~new_n12238_ & new_n12255_;
  assign new_n12257_ = new_n12238_ & ~new_n12255_;
  assign new_n12258_ = ~new_n12256_ & ~new_n12257_;
  assign A5026 = ~new_n12231_ & ~new_n12258_;
  assign new_n12260_ = new_n12228_ & ~new_n12256_;
  assign A5025 = ~new_n12231_ & ~new_n12260_;
  assign new_n12262_ = ~new_n12228_ & ~new_n12238_;
  assign new_n12263_ = ~new_n12231_ & ~new_n12262_;
  assign new_n12264_ = new_n12231_ & ~new_n12263_;
  assign new_n12265_ = new_n12231_ & new_n12262_;
  assign new_n12266_ = new_n12264_ & ~new_n12265_;
  assign new_n12267_ = ~new_n12238_ & ~new_n12266_;
  assign A5024 = new_n12255_ | new_n12267_;
  assign new_n12269_ = ~new_n12245_ & ~new_n12253_;
  assign new_n12270_ = ~new_n12254_ & ~new_n12269_;
  assign new_n12271_ = ~new_n12231_ & new_n12245_;
  assign new_n12272_ = new_n12231_ & ~new_n12245_;
  assign new_n12273_ = ~new_n12271_ & ~new_n12272_;
  assign new_n12274_ = new_n12270_ & ~new_n12273_;
  assign A5023 = new_n12267_ | new_n12274_;
  assign new_n12276_ = ~new_n12238_ & ~new_n12274_;
  assign new_n12277_ = new_n12238_ & new_n12274_;
  assign new_n12278_ = ~new_n12276_ & ~new_n12277_;
  assign A5022 = ~new_n12231_ & ~new_n12278_;
  assign new_n12280_ = new_n7048_ & new_n7053_;
  assign new_n12281_ = ~new_n7051_ & ~new_n12280_;
  assign new_n12282_ = new_n7051_ & ~new_n12281_;
  assign new_n12283_ = new_n7051_ & new_n12280_;
  assign new_n12284_ = new_n12282_ & ~new_n12283_;
  assign new_n12285_ = new_n7053_ & ~new_n12284_;
  assign new_n12286_ = ~new_n7060_ & ~new_n12285_;
  assign new_n12287_ = new_n7068_ & new_n7073_;
  assign new_n12288_ = ~new_n7071_ & ~new_n12287_;
  assign new_n12289_ = new_n7071_ & ~new_n12288_;
  assign new_n12290_ = new_n7071_ & new_n12287_;
  assign new_n12291_ = new_n12289_ & ~new_n12290_;
  assign new_n12292_ = new_n7073_ & ~new_n12291_;
  assign new_n12293_ = ~new_n7080_ & ~new_n12292_;
  assign new_n12294_ = new_n12286_ & ~new_n12293_;
  assign new_n12295_ = ~new_n12286_ & new_n12293_;
  assign new_n12296_ = ~new_n12294_ & ~new_n12295_;
  assign new_n12297_ = new_n7091_ & new_n7096_;
  assign new_n12298_ = ~new_n7094_ & ~new_n12297_;
  assign new_n12299_ = new_n7094_ & ~new_n12298_;
  assign new_n12300_ = new_n7094_ & new_n12297_;
  assign new_n12301_ = new_n12299_ & ~new_n12300_;
  assign new_n12302_ = new_n7096_ & ~new_n12301_;
  assign new_n12303_ = ~new_n7103_ & ~new_n12302_;
  assign new_n12304_ = new_n7111_ & new_n7116_;
  assign new_n12305_ = ~new_n7114_ & ~new_n12304_;
  assign new_n12306_ = new_n7114_ & ~new_n12305_;
  assign new_n12307_ = new_n7114_ & new_n12304_;
  assign new_n12308_ = new_n12306_ & ~new_n12307_;
  assign new_n12309_ = new_n7116_ & ~new_n12308_;
  assign new_n12310_ = ~new_n7123_ & ~new_n12309_;
  assign new_n12311_ = new_n12296_ & new_n12310_;
  assign new_n12312_ = new_n7132_ & new_n7137_;
  assign new_n12313_ = ~new_n7135_ & ~new_n12312_;
  assign new_n12314_ = new_n7135_ & ~new_n12313_;
  assign new_n12315_ = new_n7135_ & new_n12312_;
  assign new_n12316_ = new_n12314_ & ~new_n12315_;
  assign new_n12317_ = new_n7137_ & ~new_n12316_;
  assign new_n12318_ = ~new_n7144_ & ~new_n12317_;
  assign new_n12319_ = new_n12310_ & new_n12318_;
  assign new_n12320_ = ~new_n12311_ & ~new_n12319_;
  assign new_n12321_ = ~new_n12303_ & new_n12320_;
  assign new_n12322_ = new_n12303_ & ~new_n12320_;
  assign new_n12323_ = ~new_n12321_ & ~new_n12322_;
  assign A4993 = ~new_n12296_ & ~new_n12323_;
  assign new_n12325_ = new_n12293_ & ~new_n12321_;
  assign A4992 = ~new_n12296_ & ~new_n12325_;
  assign new_n12327_ = ~new_n12293_ & ~new_n12303_;
  assign new_n12328_ = ~new_n12296_ & ~new_n12327_;
  assign new_n12329_ = new_n12296_ & ~new_n12328_;
  assign new_n12330_ = new_n12296_ & new_n12327_;
  assign new_n12331_ = new_n12329_ & ~new_n12330_;
  assign new_n12332_ = ~new_n12303_ & ~new_n12331_;
  assign A4991 = new_n12320_ | new_n12332_;
  assign new_n12334_ = ~new_n12310_ & ~new_n12318_;
  assign new_n12335_ = ~new_n12319_ & ~new_n12334_;
  assign new_n12336_ = ~new_n12296_ & new_n12310_;
  assign new_n12337_ = new_n12296_ & ~new_n12310_;
  assign new_n12338_ = ~new_n12336_ & ~new_n12337_;
  assign new_n12339_ = new_n12335_ & ~new_n12338_;
  assign A4990 = new_n12332_ | new_n12339_;
  assign new_n12341_ = ~new_n12303_ & ~new_n12339_;
  assign new_n12342_ = new_n12303_ & new_n12339_;
  assign new_n12343_ = ~new_n12341_ & ~new_n12342_;
  assign A4989 = ~new_n12296_ & ~new_n12343_;
  assign new_n12345_ = new_n7183_ & new_n7188_;
  assign new_n12346_ = ~new_n7186_ & ~new_n12345_;
  assign new_n12347_ = new_n7186_ & ~new_n12346_;
  assign new_n12348_ = new_n7186_ & new_n12345_;
  assign new_n12349_ = new_n12347_ & ~new_n12348_;
  assign new_n12350_ = new_n7188_ & ~new_n12349_;
  assign new_n12351_ = ~new_n7195_ & ~new_n12350_;
  assign new_n12352_ = new_n7203_ & new_n7208_;
  assign new_n12353_ = ~new_n7206_ & ~new_n12352_;
  assign new_n12354_ = new_n7206_ & ~new_n12353_;
  assign new_n12355_ = new_n7206_ & new_n12352_;
  assign new_n12356_ = new_n12354_ & ~new_n12355_;
  assign new_n12357_ = new_n7208_ & ~new_n12356_;
  assign new_n12358_ = ~new_n7215_ & ~new_n12357_;
  assign new_n12359_ = new_n12351_ & ~new_n12358_;
  assign new_n12360_ = ~new_n12351_ & new_n12358_;
  assign new_n12361_ = ~new_n12359_ & ~new_n12360_;
  assign new_n12362_ = new_n7226_ & new_n7231_;
  assign new_n12363_ = ~new_n7229_ & ~new_n12362_;
  assign new_n12364_ = new_n7229_ & ~new_n12363_;
  assign new_n12365_ = new_n7229_ & new_n12362_;
  assign new_n12366_ = new_n12364_ & ~new_n12365_;
  assign new_n12367_ = new_n7231_ & ~new_n12366_;
  assign new_n12368_ = ~new_n7238_ & ~new_n12367_;
  assign new_n12369_ = new_n7246_ & new_n7251_;
  assign new_n12370_ = ~new_n7249_ & ~new_n12369_;
  assign new_n12371_ = new_n7249_ & ~new_n12370_;
  assign new_n12372_ = new_n7249_ & new_n12369_;
  assign new_n12373_ = new_n12371_ & ~new_n12372_;
  assign new_n12374_ = new_n7251_ & ~new_n12373_;
  assign new_n12375_ = ~new_n7258_ & ~new_n12374_;
  assign new_n12376_ = new_n12361_ & new_n12375_;
  assign new_n12377_ = new_n7267_ & new_n7272_;
  assign new_n12378_ = ~new_n7270_ & ~new_n12377_;
  assign new_n12379_ = new_n7270_ & ~new_n12378_;
  assign new_n12380_ = new_n7270_ & new_n12377_;
  assign new_n12381_ = new_n12379_ & ~new_n12380_;
  assign new_n12382_ = new_n7272_ & ~new_n12381_;
  assign new_n12383_ = ~new_n7279_ & ~new_n12382_;
  assign new_n12384_ = new_n12375_ & new_n12383_;
  assign new_n12385_ = ~new_n12376_ & ~new_n12384_;
  assign new_n12386_ = ~new_n12368_ & new_n12385_;
  assign new_n12387_ = new_n12368_ & ~new_n12385_;
  assign new_n12388_ = ~new_n12386_ & ~new_n12387_;
  assign A4960 = ~new_n12361_ & ~new_n12388_;
  assign new_n12390_ = new_n12358_ & ~new_n12386_;
  assign A4959 = ~new_n12361_ & ~new_n12390_;
  assign new_n12392_ = ~new_n12358_ & ~new_n12368_;
  assign new_n12393_ = ~new_n12361_ & ~new_n12392_;
  assign new_n12394_ = new_n12361_ & ~new_n12393_;
  assign new_n12395_ = new_n12361_ & new_n12392_;
  assign new_n12396_ = new_n12394_ & ~new_n12395_;
  assign new_n12397_ = ~new_n12368_ & ~new_n12396_;
  assign A4958 = new_n12385_ | new_n12397_;
  assign new_n12399_ = ~new_n12375_ & ~new_n12383_;
  assign new_n12400_ = ~new_n12384_ & ~new_n12399_;
  assign new_n12401_ = ~new_n12361_ & new_n12375_;
  assign new_n12402_ = new_n12361_ & ~new_n12375_;
  assign new_n12403_ = ~new_n12401_ & ~new_n12402_;
  assign new_n12404_ = new_n12400_ & ~new_n12403_;
  assign A4957 = new_n12397_ | new_n12404_;
  assign new_n12406_ = ~new_n12368_ & ~new_n12404_;
  assign new_n12407_ = new_n12368_ & new_n12404_;
  assign new_n12408_ = ~new_n12406_ & ~new_n12407_;
  assign A4956 = ~new_n12361_ & ~new_n12408_;
  assign new_n12410_ = ~new_n7323_ & ~new_n7333_;
  assign new_n12411_ = ~new_n7326_ & ~new_n12410_;
  assign new_n12412_ = new_n7326_ & ~new_n12411_;
  assign new_n12413_ = new_n7326_ & new_n12410_;
  assign new_n12414_ = new_n12412_ & ~new_n12413_;
  assign new_n12415_ = ~new_n7333_ & ~new_n12414_;
  assign new_n12416_ = ~new_n7350_ & ~new_n12415_;
  assign new_n12417_ = ~new_n7368_ & ~new_n7378_;
  assign new_n12418_ = ~new_n7371_ & ~new_n12417_;
  assign new_n12419_ = new_n7371_ & ~new_n12418_;
  assign new_n12420_ = new_n7371_ & new_n12417_;
  assign new_n12421_ = new_n12419_ & ~new_n12420_;
  assign new_n12422_ = ~new_n7378_ & ~new_n12421_;
  assign new_n12423_ = ~new_n7395_ & ~new_n12422_;
  assign new_n12424_ = new_n12416_ & ~new_n12423_;
  assign new_n12425_ = ~new_n12416_ & new_n12423_;
  assign new_n12426_ = ~new_n12424_ & ~new_n12425_;
  assign new_n12427_ = ~new_n7416_ & ~new_n7426_;
  assign new_n12428_ = ~new_n7419_ & ~new_n12427_;
  assign new_n12429_ = new_n7419_ & ~new_n12428_;
  assign new_n12430_ = new_n7419_ & new_n12427_;
  assign new_n12431_ = new_n12429_ & ~new_n12430_;
  assign new_n12432_ = ~new_n7426_ & ~new_n12431_;
  assign new_n12433_ = ~new_n7443_ & ~new_n12432_;
  assign new_n12434_ = ~new_n7461_ & ~new_n7471_;
  assign new_n12435_ = ~new_n7464_ & ~new_n12434_;
  assign new_n12436_ = new_n7464_ & ~new_n12435_;
  assign new_n12437_ = new_n7464_ & new_n12434_;
  assign new_n12438_ = new_n12436_ & ~new_n12437_;
  assign new_n12439_ = ~new_n7471_ & ~new_n12438_;
  assign new_n12440_ = ~new_n7488_ & ~new_n12439_;
  assign new_n12441_ = new_n12426_ & new_n12440_;
  assign new_n12442_ = ~new_n7507_ & ~new_n7517_;
  assign new_n12443_ = ~new_n7510_ & ~new_n12442_;
  assign new_n12444_ = new_n7510_ & ~new_n12443_;
  assign new_n12445_ = new_n7510_ & new_n12442_;
  assign new_n12446_ = new_n12444_ & ~new_n12445_;
  assign new_n12447_ = ~new_n7517_ & ~new_n12446_;
  assign new_n12448_ = ~new_n7534_ & ~new_n12447_;
  assign new_n12449_ = new_n12440_ & new_n12448_;
  assign new_n12450_ = ~new_n12441_ & ~new_n12449_;
  assign new_n12451_ = ~new_n12433_ & new_n12450_;
  assign new_n12452_ = new_n12433_ & ~new_n12450_;
  assign new_n12453_ = ~new_n12451_ & ~new_n12452_;
  assign A4927 = ~new_n12426_ & ~new_n12453_;
  assign new_n12455_ = new_n12423_ & ~new_n12451_;
  assign A4926 = ~new_n12426_ & ~new_n12455_;
  assign new_n12457_ = ~new_n12423_ & ~new_n12433_;
  assign new_n12458_ = ~new_n12426_ & ~new_n12457_;
  assign new_n12459_ = new_n12426_ & ~new_n12458_;
  assign new_n12460_ = new_n12426_ & new_n12457_;
  assign new_n12461_ = new_n12459_ & ~new_n12460_;
  assign new_n12462_ = ~new_n12433_ & ~new_n12461_;
  assign A4925 = new_n12450_ | new_n12462_;
  assign new_n12464_ = ~new_n12440_ & ~new_n12448_;
  assign new_n12465_ = ~new_n12449_ & ~new_n12464_;
  assign new_n12466_ = ~new_n12426_ & new_n12440_;
  assign new_n12467_ = new_n12426_ & ~new_n12440_;
  assign new_n12468_ = ~new_n12466_ & ~new_n12467_;
  assign new_n12469_ = new_n12465_ & ~new_n12468_;
  assign A4924 = new_n12462_ | new_n12469_;
  assign new_n12471_ = ~new_n12433_ & ~new_n12469_;
  assign new_n12472_ = new_n12433_ & new_n12469_;
  assign new_n12473_ = ~new_n12471_ & ~new_n12472_;
  assign A4923 = ~new_n12426_ & ~new_n12473_;
  assign new_n12475_ = ~new_n7578_ & ~new_n7588_;
  assign new_n12476_ = ~new_n7581_ & ~new_n12475_;
  assign new_n12477_ = new_n7581_ & ~new_n12476_;
  assign new_n12478_ = new_n7581_ & new_n12475_;
  assign new_n12479_ = new_n12477_ & ~new_n12478_;
  assign new_n12480_ = ~new_n7588_ & ~new_n12479_;
  assign new_n12481_ = ~new_n7605_ & ~new_n12480_;
  assign new_n12482_ = ~new_n7623_ & ~new_n7633_;
  assign new_n12483_ = ~new_n7626_ & ~new_n12482_;
  assign new_n12484_ = new_n7626_ & ~new_n12483_;
  assign new_n12485_ = new_n7626_ & new_n12482_;
  assign new_n12486_ = new_n12484_ & ~new_n12485_;
  assign new_n12487_ = ~new_n7633_ & ~new_n12486_;
  assign new_n12488_ = ~new_n7650_ & ~new_n12487_;
  assign new_n12489_ = new_n12481_ & ~new_n12488_;
  assign new_n12490_ = ~new_n12481_ & new_n12488_;
  assign new_n12491_ = ~new_n12489_ & ~new_n12490_;
  assign new_n12492_ = ~new_n7671_ & ~new_n7681_;
  assign new_n12493_ = ~new_n7674_ & ~new_n12492_;
  assign new_n12494_ = new_n7674_ & ~new_n12493_;
  assign new_n12495_ = new_n7674_ & new_n12492_;
  assign new_n12496_ = new_n12494_ & ~new_n12495_;
  assign new_n12497_ = ~new_n7681_ & ~new_n12496_;
  assign new_n12498_ = ~new_n7698_ & ~new_n12497_;
  assign new_n12499_ = ~new_n7716_ & ~new_n7726_;
  assign new_n12500_ = ~new_n7719_ & ~new_n12499_;
  assign new_n12501_ = new_n7719_ & ~new_n12500_;
  assign new_n12502_ = new_n7719_ & new_n12499_;
  assign new_n12503_ = new_n12501_ & ~new_n12502_;
  assign new_n12504_ = ~new_n7726_ & ~new_n12503_;
  assign new_n12505_ = ~new_n7743_ & ~new_n12504_;
  assign new_n12506_ = new_n12491_ & new_n12505_;
  assign new_n12507_ = ~new_n7762_ & ~new_n7772_;
  assign new_n12508_ = ~new_n7765_ & ~new_n12507_;
  assign new_n12509_ = new_n7765_ & ~new_n12508_;
  assign new_n12510_ = new_n7765_ & new_n12507_;
  assign new_n12511_ = new_n12509_ & ~new_n12510_;
  assign new_n12512_ = ~new_n7772_ & ~new_n12511_;
  assign new_n12513_ = ~new_n7789_ & ~new_n12512_;
  assign new_n12514_ = new_n12505_ & new_n12513_;
  assign new_n12515_ = ~new_n12506_ & ~new_n12514_;
  assign new_n12516_ = ~new_n12498_ & new_n12515_;
  assign new_n12517_ = new_n12498_ & ~new_n12515_;
  assign new_n12518_ = ~new_n12516_ & ~new_n12517_;
  assign A4894 = ~new_n12491_ & ~new_n12518_;
  assign new_n12520_ = new_n12488_ & ~new_n12516_;
  assign A4893 = ~new_n12491_ & ~new_n12520_;
  assign new_n12522_ = ~new_n12488_ & ~new_n12498_;
  assign new_n12523_ = ~new_n12491_ & ~new_n12522_;
  assign new_n12524_ = new_n12491_ & ~new_n12523_;
  assign new_n12525_ = new_n12491_ & new_n12522_;
  assign new_n12526_ = new_n12524_ & ~new_n12525_;
  assign new_n12527_ = ~new_n12498_ & ~new_n12526_;
  assign A4892 = new_n12515_ | new_n12527_;
  assign new_n12529_ = ~new_n12505_ & ~new_n12513_;
  assign new_n12530_ = ~new_n12514_ & ~new_n12529_;
  assign new_n12531_ = ~new_n12491_ & new_n12505_;
  assign new_n12532_ = new_n12491_ & ~new_n12505_;
  assign new_n12533_ = ~new_n12531_ & ~new_n12532_;
  assign new_n12534_ = new_n12530_ & ~new_n12533_;
  assign A4891 = new_n12527_ | new_n12534_;
  assign new_n12536_ = ~new_n12498_ & ~new_n12534_;
  assign new_n12537_ = new_n12498_ & new_n12534_;
  assign new_n12538_ = ~new_n12536_ & ~new_n12537_;
  assign A4890 = ~new_n12491_ & ~new_n12538_;
  assign new_n12540_ = ~new_n7833_ & ~new_n7843_;
  assign new_n12541_ = ~new_n7836_ & ~new_n12540_;
  assign new_n12542_ = new_n7836_ & ~new_n12541_;
  assign new_n12543_ = new_n7836_ & new_n12540_;
  assign new_n12544_ = new_n12542_ & ~new_n12543_;
  assign new_n12545_ = ~new_n7843_ & ~new_n12544_;
  assign new_n12546_ = ~new_n7860_ & ~new_n12545_;
  assign new_n12547_ = ~new_n7878_ & ~new_n7888_;
  assign new_n12548_ = ~new_n7881_ & ~new_n12547_;
  assign new_n12549_ = new_n7881_ & ~new_n12548_;
  assign new_n12550_ = new_n7881_ & new_n12547_;
  assign new_n12551_ = new_n12549_ & ~new_n12550_;
  assign new_n12552_ = ~new_n7888_ & ~new_n12551_;
  assign new_n12553_ = ~new_n7905_ & ~new_n12552_;
  assign new_n12554_ = new_n12546_ & ~new_n12553_;
  assign new_n12555_ = ~new_n12546_ & new_n12553_;
  assign new_n12556_ = ~new_n12554_ & ~new_n12555_;
  assign new_n12557_ = ~new_n7926_ & ~new_n7936_;
  assign new_n12558_ = ~new_n7929_ & ~new_n12557_;
  assign new_n12559_ = new_n7929_ & ~new_n12558_;
  assign new_n12560_ = new_n7929_ & new_n12557_;
  assign new_n12561_ = new_n12559_ & ~new_n12560_;
  assign new_n12562_ = ~new_n7936_ & ~new_n12561_;
  assign new_n12563_ = ~new_n7953_ & ~new_n12562_;
  assign new_n12564_ = ~new_n7971_ & ~new_n7981_;
  assign new_n12565_ = ~new_n7974_ & ~new_n12564_;
  assign new_n12566_ = new_n7974_ & ~new_n12565_;
  assign new_n12567_ = new_n7974_ & new_n12564_;
  assign new_n12568_ = new_n12566_ & ~new_n12567_;
  assign new_n12569_ = ~new_n7981_ & ~new_n12568_;
  assign new_n12570_ = ~new_n7998_ & ~new_n12569_;
  assign new_n12571_ = new_n12556_ & new_n12570_;
  assign new_n12572_ = ~new_n8017_ & ~new_n8027_;
  assign new_n12573_ = ~new_n8020_ & ~new_n12572_;
  assign new_n12574_ = new_n8020_ & ~new_n12573_;
  assign new_n12575_ = new_n8020_ & new_n12572_;
  assign new_n12576_ = new_n12574_ & ~new_n12575_;
  assign new_n12577_ = ~new_n8027_ & ~new_n12576_;
  assign new_n12578_ = ~new_n8044_ & ~new_n12577_;
  assign new_n12579_ = new_n12570_ & new_n12578_;
  assign new_n12580_ = ~new_n12571_ & ~new_n12579_;
  assign new_n12581_ = ~new_n12563_ & new_n12580_;
  assign new_n12582_ = new_n12563_ & ~new_n12580_;
  assign new_n12583_ = ~new_n12581_ & ~new_n12582_;
  assign A4861 = ~new_n12556_ & ~new_n12583_;
  assign new_n12585_ = new_n12553_ & ~new_n12581_;
  assign A4860 = ~new_n12556_ & ~new_n12585_;
  assign new_n12587_ = ~new_n12553_ & ~new_n12563_;
  assign new_n12588_ = ~new_n12556_ & ~new_n12587_;
  assign new_n12589_ = new_n12556_ & ~new_n12588_;
  assign new_n12590_ = new_n12556_ & new_n12587_;
  assign new_n12591_ = new_n12589_ & ~new_n12590_;
  assign new_n12592_ = ~new_n12563_ & ~new_n12591_;
  assign A4859 = new_n12580_ | new_n12592_;
  assign new_n12594_ = ~new_n12570_ & ~new_n12578_;
  assign new_n12595_ = ~new_n12579_ & ~new_n12594_;
  assign new_n12596_ = ~new_n12556_ & new_n12570_;
  assign new_n12597_ = new_n12556_ & ~new_n12570_;
  assign new_n12598_ = ~new_n12596_ & ~new_n12597_;
  assign new_n12599_ = new_n12595_ & ~new_n12598_;
  assign A4858 = new_n12592_ | new_n12599_;
  assign new_n12601_ = ~new_n12563_ & ~new_n12599_;
  assign new_n12602_ = new_n12563_ & new_n12599_;
  assign new_n12603_ = ~new_n12601_ & ~new_n12602_;
  assign A4857 = ~new_n12556_ & ~new_n12603_;
  assign new_n12605_ = ~new_n8088_ & ~new_n8098_;
  assign new_n12606_ = ~new_n8091_ & ~new_n12605_;
  assign new_n12607_ = new_n8091_ & ~new_n12606_;
  assign new_n12608_ = new_n8091_ & new_n12605_;
  assign new_n12609_ = new_n12607_ & ~new_n12608_;
  assign new_n12610_ = ~new_n8098_ & ~new_n12609_;
  assign new_n12611_ = ~new_n8115_ & ~new_n12610_;
  assign new_n12612_ = ~new_n8133_ & ~new_n8143_;
  assign new_n12613_ = ~new_n8136_ & ~new_n12612_;
  assign new_n12614_ = new_n8136_ & ~new_n12613_;
  assign new_n12615_ = new_n8136_ & new_n12612_;
  assign new_n12616_ = new_n12614_ & ~new_n12615_;
  assign new_n12617_ = ~new_n8143_ & ~new_n12616_;
  assign new_n12618_ = ~new_n8160_ & ~new_n12617_;
  assign new_n12619_ = new_n12611_ & ~new_n12618_;
  assign new_n12620_ = ~new_n12611_ & new_n12618_;
  assign new_n12621_ = ~new_n12619_ & ~new_n12620_;
  assign new_n12622_ = ~new_n8181_ & ~new_n8191_;
  assign new_n12623_ = ~new_n8184_ & ~new_n12622_;
  assign new_n12624_ = new_n8184_ & ~new_n12623_;
  assign new_n12625_ = new_n8184_ & new_n12622_;
  assign new_n12626_ = new_n12624_ & ~new_n12625_;
  assign new_n12627_ = ~new_n8191_ & ~new_n12626_;
  assign new_n12628_ = ~new_n8208_ & ~new_n12627_;
  assign new_n12629_ = ~new_n8226_ & ~new_n8236_;
  assign new_n12630_ = ~new_n8229_ & ~new_n12629_;
  assign new_n12631_ = new_n8229_ & ~new_n12630_;
  assign new_n12632_ = new_n8229_ & new_n12629_;
  assign new_n12633_ = new_n12631_ & ~new_n12632_;
  assign new_n12634_ = ~new_n8236_ & ~new_n12633_;
  assign new_n12635_ = ~new_n8253_ & ~new_n12634_;
  assign new_n12636_ = new_n12621_ & new_n12635_;
  assign new_n12637_ = ~new_n8272_ & ~new_n8282_;
  assign new_n12638_ = ~new_n8275_ & ~new_n12637_;
  assign new_n12639_ = new_n8275_ & ~new_n12638_;
  assign new_n12640_ = new_n8275_ & new_n12637_;
  assign new_n12641_ = new_n12639_ & ~new_n12640_;
  assign new_n12642_ = ~new_n8282_ & ~new_n12641_;
  assign new_n12643_ = ~new_n8299_ & ~new_n12642_;
  assign new_n12644_ = new_n12635_ & new_n12643_;
  assign new_n12645_ = ~new_n12636_ & ~new_n12644_;
  assign new_n12646_ = ~new_n12628_ & new_n12645_;
  assign new_n12647_ = new_n12628_ & ~new_n12645_;
  assign new_n12648_ = ~new_n12646_ & ~new_n12647_;
  assign A4828 = ~new_n12621_ & ~new_n12648_;
  assign new_n12650_ = new_n12618_ & ~new_n12646_;
  assign A4827 = ~new_n12621_ & ~new_n12650_;
  assign new_n12652_ = ~new_n12618_ & ~new_n12628_;
  assign new_n12653_ = ~new_n12621_ & ~new_n12652_;
  assign new_n12654_ = new_n12621_ & ~new_n12653_;
  assign new_n12655_ = new_n12621_ & new_n12652_;
  assign new_n12656_ = new_n12654_ & ~new_n12655_;
  assign new_n12657_ = ~new_n12628_ & ~new_n12656_;
  assign A4826 = new_n12645_ | new_n12657_;
  assign new_n12659_ = ~new_n12635_ & ~new_n12643_;
  assign new_n12660_ = ~new_n12644_ & ~new_n12659_;
  assign new_n12661_ = ~new_n12621_ & new_n12635_;
  assign new_n12662_ = new_n12621_ & ~new_n12635_;
  assign new_n12663_ = ~new_n12661_ & ~new_n12662_;
  assign new_n12664_ = new_n12660_ & ~new_n12663_;
  assign A4825 = new_n12657_ | new_n12664_;
  assign new_n12666_ = ~new_n12628_ & ~new_n12664_;
  assign new_n12667_ = new_n12628_ & new_n12664_;
  assign new_n12668_ = ~new_n12666_ & ~new_n12667_;
  assign A4824 = ~new_n12621_ & ~new_n12668_;
  assign new_n12670_ = ~new_n8339_ & ~new_n8349_;
  assign new_n12671_ = ~new_n8342_ & ~new_n12670_;
  assign new_n12672_ = new_n8342_ & ~new_n12671_;
  assign new_n12673_ = new_n8342_ & new_n12670_;
  assign new_n12674_ = new_n12672_ & ~new_n12673_;
  assign new_n12675_ = ~new_n8349_ & ~new_n12674_;
  assign new_n12676_ = ~new_n8366_ & ~new_n12675_;
  assign new_n12677_ = ~new_n8384_ & ~new_n8394_;
  assign new_n12678_ = ~new_n8387_ & ~new_n12677_;
  assign new_n12679_ = new_n8387_ & ~new_n12678_;
  assign new_n12680_ = new_n8387_ & new_n12677_;
  assign new_n12681_ = new_n12679_ & ~new_n12680_;
  assign new_n12682_ = ~new_n8394_ & ~new_n12681_;
  assign new_n12683_ = ~new_n8411_ & ~new_n12682_;
  assign new_n12684_ = new_n12676_ & ~new_n12683_;
  assign new_n12685_ = ~new_n12676_ & new_n12683_;
  assign new_n12686_ = ~new_n12684_ & ~new_n12685_;
  assign new_n12687_ = ~new_n8432_ & ~new_n8442_;
  assign new_n12688_ = ~new_n8435_ & ~new_n12687_;
  assign new_n12689_ = new_n8435_ & ~new_n12688_;
  assign new_n12690_ = new_n8435_ & new_n12687_;
  assign new_n12691_ = new_n12689_ & ~new_n12690_;
  assign new_n12692_ = ~new_n8442_ & ~new_n12691_;
  assign new_n12693_ = ~new_n8459_ & ~new_n12692_;
  assign new_n12694_ = ~new_n8477_ & ~new_n8487_;
  assign new_n12695_ = ~new_n8480_ & ~new_n12694_;
  assign new_n12696_ = new_n8480_ & ~new_n12695_;
  assign new_n12697_ = new_n8480_ & new_n12694_;
  assign new_n12698_ = new_n12696_ & ~new_n12697_;
  assign new_n12699_ = ~new_n8487_ & ~new_n12698_;
  assign new_n12700_ = ~new_n8504_ & ~new_n12699_;
  assign new_n12701_ = new_n12686_ & new_n12700_;
  assign new_n12702_ = ~new_n8523_ & ~new_n8533_;
  assign new_n12703_ = ~new_n8526_ & ~new_n12702_;
  assign new_n12704_ = new_n8526_ & ~new_n12703_;
  assign new_n12705_ = new_n8526_ & new_n12702_;
  assign new_n12706_ = new_n12704_ & ~new_n12705_;
  assign new_n12707_ = ~new_n8533_ & ~new_n12706_;
  assign new_n12708_ = ~new_n8550_ & ~new_n12707_;
  assign new_n12709_ = new_n12700_ & new_n12708_;
  assign new_n12710_ = ~new_n12701_ & ~new_n12709_;
  assign new_n12711_ = ~new_n12693_ & new_n12710_;
  assign new_n12712_ = new_n12693_ & ~new_n12710_;
  assign new_n12713_ = ~new_n12711_ & ~new_n12712_;
  assign A4795 = ~new_n12686_ & ~new_n12713_;
  assign new_n12715_ = new_n12683_ & ~new_n12711_;
  assign A4794 = ~new_n12686_ & ~new_n12715_;
  assign new_n12717_ = ~new_n12683_ & ~new_n12693_;
  assign new_n12718_ = ~new_n12686_ & ~new_n12717_;
  assign new_n12719_ = new_n12686_ & ~new_n12718_;
  assign new_n12720_ = new_n12686_ & new_n12717_;
  assign new_n12721_ = new_n12719_ & ~new_n12720_;
  assign new_n12722_ = ~new_n12693_ & ~new_n12721_;
  assign A4793 = new_n12710_ | new_n12722_;
  assign new_n12724_ = ~new_n12700_ & ~new_n12708_;
  assign new_n12725_ = ~new_n12709_ & ~new_n12724_;
  assign new_n12726_ = ~new_n12686_ & new_n12700_;
  assign new_n12727_ = new_n12686_ & ~new_n12700_;
  assign new_n12728_ = ~new_n12726_ & ~new_n12727_;
  assign new_n12729_ = new_n12725_ & ~new_n12728_;
  assign A4792 = new_n12722_ | new_n12729_;
  assign new_n12731_ = ~new_n12693_ & ~new_n12729_;
  assign new_n12732_ = new_n12693_ & new_n12729_;
  assign new_n12733_ = ~new_n12731_ & ~new_n12732_;
  assign A4791 = ~new_n12686_ & ~new_n12733_;
  assign new_n12735_ = ~new_n8594_ & ~new_n8604_;
  assign new_n12736_ = ~new_n8597_ & ~new_n12735_;
  assign new_n12737_ = new_n8597_ & ~new_n12736_;
  assign new_n12738_ = new_n8597_ & new_n12735_;
  assign new_n12739_ = new_n12737_ & ~new_n12738_;
  assign new_n12740_ = ~new_n8604_ & ~new_n12739_;
  assign new_n12741_ = ~new_n8621_ & ~new_n12740_;
  assign new_n12742_ = ~new_n8639_ & ~new_n8649_;
  assign new_n12743_ = ~new_n8642_ & ~new_n12742_;
  assign new_n12744_ = new_n8642_ & ~new_n12743_;
  assign new_n12745_ = new_n8642_ & new_n12742_;
  assign new_n12746_ = new_n12744_ & ~new_n12745_;
  assign new_n12747_ = ~new_n8649_ & ~new_n12746_;
  assign new_n12748_ = ~new_n8666_ & ~new_n12747_;
  assign new_n12749_ = new_n12741_ & ~new_n12748_;
  assign new_n12750_ = ~new_n12741_ & new_n12748_;
  assign new_n12751_ = ~new_n12749_ & ~new_n12750_;
  assign new_n12752_ = ~new_n8687_ & ~new_n8697_;
  assign new_n12753_ = ~new_n8690_ & ~new_n12752_;
  assign new_n12754_ = new_n8690_ & ~new_n12753_;
  assign new_n12755_ = new_n8690_ & new_n12752_;
  assign new_n12756_ = new_n12754_ & ~new_n12755_;
  assign new_n12757_ = ~new_n8697_ & ~new_n12756_;
  assign new_n12758_ = ~new_n8714_ & ~new_n12757_;
  assign new_n12759_ = ~new_n8732_ & ~new_n8742_;
  assign new_n12760_ = ~new_n8735_ & ~new_n12759_;
  assign new_n12761_ = new_n8735_ & ~new_n12760_;
  assign new_n12762_ = new_n8735_ & new_n12759_;
  assign new_n12763_ = new_n12761_ & ~new_n12762_;
  assign new_n12764_ = ~new_n8742_ & ~new_n12763_;
  assign new_n12765_ = ~new_n8759_ & ~new_n12764_;
  assign new_n12766_ = new_n12751_ & new_n12765_;
  assign new_n12767_ = ~new_n8778_ & ~new_n8788_;
  assign new_n12768_ = ~new_n8781_ & ~new_n12767_;
  assign new_n12769_ = new_n8781_ & ~new_n12768_;
  assign new_n12770_ = new_n8781_ & new_n12767_;
  assign new_n12771_ = new_n12769_ & ~new_n12770_;
  assign new_n12772_ = ~new_n8788_ & ~new_n12771_;
  assign new_n12773_ = ~new_n8805_ & ~new_n12772_;
  assign new_n12774_ = new_n12765_ & new_n12773_;
  assign new_n12775_ = ~new_n12766_ & ~new_n12774_;
  assign new_n12776_ = ~new_n12758_ & new_n12775_;
  assign new_n12777_ = new_n12758_ & ~new_n12775_;
  assign new_n12778_ = ~new_n12776_ & ~new_n12777_;
  assign A4762 = ~new_n12751_ & ~new_n12778_;
  assign new_n12780_ = new_n12748_ & ~new_n12776_;
  assign A4761 = ~new_n12751_ & ~new_n12780_;
  assign new_n12782_ = ~new_n12748_ & ~new_n12758_;
  assign new_n12783_ = ~new_n12751_ & ~new_n12782_;
  assign new_n12784_ = new_n12751_ & ~new_n12783_;
  assign new_n12785_ = new_n12751_ & new_n12782_;
  assign new_n12786_ = new_n12784_ & ~new_n12785_;
  assign new_n12787_ = ~new_n12758_ & ~new_n12786_;
  assign A4760 = new_n12775_ | new_n12787_;
  assign new_n12789_ = ~new_n12765_ & ~new_n12773_;
  assign new_n12790_ = ~new_n12774_ & ~new_n12789_;
  assign new_n12791_ = ~new_n12751_ & new_n12765_;
  assign new_n12792_ = new_n12751_ & ~new_n12765_;
  assign new_n12793_ = ~new_n12791_ & ~new_n12792_;
  assign new_n12794_ = new_n12790_ & ~new_n12793_;
  assign A4759 = new_n12787_ | new_n12794_;
  assign new_n12796_ = ~new_n12758_ & ~new_n12794_;
  assign new_n12797_ = new_n12758_ & new_n12794_;
  assign new_n12798_ = ~new_n12796_ & ~new_n12797_;
  assign A4758 = ~new_n12751_ & ~new_n12798_;
  assign new_n12800_ = ~new_n8849_ & ~new_n8859_;
  assign new_n12801_ = ~new_n8852_ & ~new_n12800_;
  assign new_n12802_ = new_n8852_ & ~new_n12801_;
  assign new_n12803_ = new_n8852_ & new_n12800_;
  assign new_n12804_ = new_n12802_ & ~new_n12803_;
  assign new_n12805_ = ~new_n8859_ & ~new_n12804_;
  assign new_n12806_ = ~new_n8876_ & ~new_n12805_;
  assign new_n12807_ = ~new_n8894_ & ~new_n8904_;
  assign new_n12808_ = ~new_n8897_ & ~new_n12807_;
  assign new_n12809_ = new_n8897_ & ~new_n12808_;
  assign new_n12810_ = new_n8897_ & new_n12807_;
  assign new_n12811_ = new_n12809_ & ~new_n12810_;
  assign new_n12812_ = ~new_n8904_ & ~new_n12811_;
  assign new_n12813_ = ~new_n8921_ & ~new_n12812_;
  assign new_n12814_ = new_n12806_ & ~new_n12813_;
  assign new_n12815_ = ~new_n12806_ & new_n12813_;
  assign new_n12816_ = ~new_n12814_ & ~new_n12815_;
  assign new_n12817_ = ~new_n8942_ & ~new_n8952_;
  assign new_n12818_ = ~new_n8945_ & ~new_n12817_;
  assign new_n12819_ = new_n8945_ & ~new_n12818_;
  assign new_n12820_ = new_n8945_ & new_n12817_;
  assign new_n12821_ = new_n12819_ & ~new_n12820_;
  assign new_n12822_ = ~new_n8952_ & ~new_n12821_;
  assign new_n12823_ = ~new_n8969_ & ~new_n12822_;
  assign new_n12824_ = ~new_n8987_ & ~new_n8997_;
  assign new_n12825_ = ~new_n8990_ & ~new_n12824_;
  assign new_n12826_ = new_n8990_ & ~new_n12825_;
  assign new_n12827_ = new_n8990_ & new_n12824_;
  assign new_n12828_ = new_n12826_ & ~new_n12827_;
  assign new_n12829_ = ~new_n8997_ & ~new_n12828_;
  assign new_n12830_ = ~new_n9014_ & ~new_n12829_;
  assign new_n12831_ = new_n12816_ & new_n12830_;
  assign new_n12832_ = ~new_n9033_ & ~new_n9043_;
  assign new_n12833_ = ~new_n9036_ & ~new_n12832_;
  assign new_n12834_ = new_n9036_ & ~new_n12833_;
  assign new_n12835_ = new_n9036_ & new_n12832_;
  assign new_n12836_ = new_n12834_ & ~new_n12835_;
  assign new_n12837_ = ~new_n9043_ & ~new_n12836_;
  assign new_n12838_ = ~new_n9060_ & ~new_n12837_;
  assign new_n12839_ = new_n12830_ & new_n12838_;
  assign new_n12840_ = ~new_n12831_ & ~new_n12839_;
  assign new_n12841_ = ~new_n12823_ & new_n12840_;
  assign new_n12842_ = new_n12823_ & ~new_n12840_;
  assign new_n12843_ = ~new_n12841_ & ~new_n12842_;
  assign A4729 = ~new_n12816_ & ~new_n12843_;
  assign new_n12845_ = new_n12813_ & ~new_n12841_;
  assign A4728 = ~new_n12816_ & ~new_n12845_;
  assign new_n12847_ = ~new_n12813_ & ~new_n12823_;
  assign new_n12848_ = ~new_n12816_ & ~new_n12847_;
  assign new_n12849_ = new_n12816_ & ~new_n12848_;
  assign new_n12850_ = new_n12816_ & new_n12847_;
  assign new_n12851_ = new_n12849_ & ~new_n12850_;
  assign new_n12852_ = ~new_n12823_ & ~new_n12851_;
  assign A4727 = new_n12840_ | new_n12852_;
  assign new_n12854_ = ~new_n12830_ & ~new_n12838_;
  assign new_n12855_ = ~new_n12839_ & ~new_n12854_;
  assign new_n12856_ = ~new_n12816_ & new_n12830_;
  assign new_n12857_ = new_n12816_ & ~new_n12830_;
  assign new_n12858_ = ~new_n12856_ & ~new_n12857_;
  assign new_n12859_ = new_n12855_ & ~new_n12858_;
  assign A4726 = new_n12852_ | new_n12859_;
  assign new_n12861_ = ~new_n12823_ & ~new_n12859_;
  assign new_n12862_ = new_n12823_ & new_n12859_;
  assign new_n12863_ = ~new_n12861_ & ~new_n12862_;
  assign A4725 = ~new_n12816_ & ~new_n12863_;
  assign new_n12865_ = ~new_n9104_ & ~new_n9114_;
  assign new_n12866_ = ~new_n9107_ & ~new_n12865_;
  assign new_n12867_ = new_n9107_ & ~new_n12866_;
  assign new_n12868_ = new_n9107_ & new_n12865_;
  assign new_n12869_ = new_n12867_ & ~new_n12868_;
  assign new_n12870_ = ~new_n9114_ & ~new_n12869_;
  assign new_n12871_ = ~new_n9131_ & ~new_n12870_;
  assign new_n12872_ = ~new_n9149_ & ~new_n9159_;
  assign new_n12873_ = ~new_n9152_ & ~new_n12872_;
  assign new_n12874_ = new_n9152_ & ~new_n12873_;
  assign new_n12875_ = new_n9152_ & new_n12872_;
  assign new_n12876_ = new_n12874_ & ~new_n12875_;
  assign new_n12877_ = ~new_n9159_ & ~new_n12876_;
  assign new_n12878_ = ~new_n9176_ & ~new_n12877_;
  assign new_n12879_ = new_n12871_ & ~new_n12878_;
  assign new_n12880_ = ~new_n12871_ & new_n12878_;
  assign new_n12881_ = ~new_n12879_ & ~new_n12880_;
  assign new_n12882_ = ~new_n9197_ & ~new_n9207_;
  assign new_n12883_ = ~new_n9200_ & ~new_n12882_;
  assign new_n12884_ = new_n9200_ & ~new_n12883_;
  assign new_n12885_ = new_n9200_ & new_n12882_;
  assign new_n12886_ = new_n12884_ & ~new_n12885_;
  assign new_n12887_ = ~new_n9207_ & ~new_n12886_;
  assign new_n12888_ = ~new_n9224_ & ~new_n12887_;
  assign new_n12889_ = ~new_n9242_ & ~new_n9252_;
  assign new_n12890_ = ~new_n9245_ & ~new_n12889_;
  assign new_n12891_ = new_n9245_ & ~new_n12890_;
  assign new_n12892_ = new_n9245_ & new_n12889_;
  assign new_n12893_ = new_n12891_ & ~new_n12892_;
  assign new_n12894_ = ~new_n9252_ & ~new_n12893_;
  assign new_n12895_ = ~new_n9269_ & ~new_n12894_;
  assign new_n12896_ = new_n12881_ & new_n12895_;
  assign new_n12897_ = ~new_n9288_ & ~new_n9298_;
  assign new_n12898_ = ~new_n9291_ & ~new_n12897_;
  assign new_n12899_ = new_n9291_ & ~new_n12898_;
  assign new_n12900_ = new_n9291_ & new_n12897_;
  assign new_n12901_ = new_n12899_ & ~new_n12900_;
  assign new_n12902_ = ~new_n9298_ & ~new_n12901_;
  assign new_n12903_ = ~new_n9315_ & ~new_n12902_;
  assign new_n12904_ = new_n12895_ & new_n12903_;
  assign new_n12905_ = ~new_n12896_ & ~new_n12904_;
  assign new_n12906_ = ~new_n12888_ & new_n12905_;
  assign new_n12907_ = new_n12888_ & ~new_n12905_;
  assign new_n12908_ = ~new_n12906_ & ~new_n12907_;
  assign A4696 = ~new_n12881_ & ~new_n12908_;
  assign new_n12910_ = new_n12878_ & ~new_n12906_;
  assign A4695 = ~new_n12881_ & ~new_n12910_;
  assign new_n12912_ = ~new_n12878_ & ~new_n12888_;
  assign new_n12913_ = ~new_n12881_ & ~new_n12912_;
  assign new_n12914_ = new_n12881_ & ~new_n12913_;
  assign new_n12915_ = new_n12881_ & new_n12912_;
  assign new_n12916_ = new_n12914_ & ~new_n12915_;
  assign new_n12917_ = ~new_n12888_ & ~new_n12916_;
  assign A4694 = new_n12905_ | new_n12917_;
  assign new_n12919_ = ~new_n12895_ & ~new_n12903_;
  assign new_n12920_ = ~new_n12904_ & ~new_n12919_;
  assign new_n12921_ = ~new_n12881_ & new_n12895_;
  assign new_n12922_ = new_n12881_ & ~new_n12895_;
  assign new_n12923_ = ~new_n12921_ & ~new_n12922_;
  assign new_n12924_ = new_n12920_ & ~new_n12923_;
  assign A4693 = new_n12917_ | new_n12924_;
  assign new_n12926_ = ~new_n12888_ & ~new_n12924_;
  assign new_n12927_ = new_n12888_ & new_n12924_;
  assign new_n12928_ = ~new_n12926_ & ~new_n12927_;
  assign A4692 = ~new_n12881_ & ~new_n12928_;
  assign new_n12930_ = ~new_n9359_ & ~new_n9369_;
  assign new_n12931_ = ~new_n9362_ & ~new_n12930_;
  assign new_n12932_ = new_n9362_ & ~new_n12931_;
  assign new_n12933_ = new_n9362_ & new_n12930_;
  assign new_n12934_ = new_n12932_ & ~new_n12933_;
  assign new_n12935_ = ~new_n9369_ & ~new_n12934_;
  assign new_n12936_ = ~new_n9386_ & ~new_n12935_;
  assign new_n12937_ = ~new_n9404_ & ~new_n9414_;
  assign new_n12938_ = ~new_n9407_ & ~new_n12937_;
  assign new_n12939_ = new_n9407_ & ~new_n12938_;
  assign new_n12940_ = new_n9407_ & new_n12937_;
  assign new_n12941_ = new_n12939_ & ~new_n12940_;
  assign new_n12942_ = ~new_n9414_ & ~new_n12941_;
  assign new_n12943_ = ~new_n9431_ & ~new_n12942_;
  assign new_n12944_ = new_n12936_ & ~new_n12943_;
  assign new_n12945_ = ~new_n12936_ & new_n12943_;
  assign new_n12946_ = ~new_n12944_ & ~new_n12945_;
  assign new_n12947_ = ~new_n9452_ & ~new_n9462_;
  assign new_n12948_ = ~new_n9455_ & ~new_n12947_;
  assign new_n12949_ = new_n9455_ & ~new_n12948_;
  assign new_n12950_ = new_n9455_ & new_n12947_;
  assign new_n12951_ = new_n12949_ & ~new_n12950_;
  assign new_n12952_ = ~new_n9462_ & ~new_n12951_;
  assign new_n12953_ = ~new_n9479_ & ~new_n12952_;
  assign new_n12954_ = ~new_n9497_ & ~new_n9507_;
  assign new_n12955_ = ~new_n9500_ & ~new_n12954_;
  assign new_n12956_ = new_n9500_ & ~new_n12955_;
  assign new_n12957_ = new_n9500_ & new_n12954_;
  assign new_n12958_ = new_n12956_ & ~new_n12957_;
  assign new_n12959_ = ~new_n9507_ & ~new_n12958_;
  assign new_n12960_ = ~new_n9524_ & ~new_n12959_;
  assign new_n12961_ = new_n12946_ & new_n12960_;
  assign new_n12962_ = ~new_n9543_ & ~new_n9553_;
  assign new_n12963_ = ~new_n9546_ & ~new_n12962_;
  assign new_n12964_ = new_n9546_ & ~new_n12963_;
  assign new_n12965_ = new_n9546_ & new_n12962_;
  assign new_n12966_ = new_n12964_ & ~new_n12965_;
  assign new_n12967_ = ~new_n9553_ & ~new_n12966_;
  assign new_n12968_ = ~new_n9570_ & ~new_n12967_;
  assign new_n12969_ = new_n12960_ & new_n12968_;
  assign new_n12970_ = ~new_n12961_ & ~new_n12969_;
  assign new_n12971_ = ~new_n12953_ & new_n12970_;
  assign new_n12972_ = new_n12953_ & ~new_n12970_;
  assign new_n12973_ = ~new_n12971_ & ~new_n12972_;
  assign A4663 = ~new_n12946_ & ~new_n12973_;
  assign new_n12975_ = new_n12943_ & ~new_n12971_;
  assign A4662 = ~new_n12946_ & ~new_n12975_;
  assign new_n12977_ = ~new_n12943_ & ~new_n12953_;
  assign new_n12978_ = ~new_n12946_ & ~new_n12977_;
  assign new_n12979_ = new_n12946_ & ~new_n12978_;
  assign new_n12980_ = new_n12946_ & new_n12977_;
  assign new_n12981_ = new_n12979_ & ~new_n12980_;
  assign new_n12982_ = ~new_n12953_ & ~new_n12981_;
  assign A4661 = new_n12970_ | new_n12982_;
  assign new_n12984_ = ~new_n12960_ & ~new_n12968_;
  assign new_n12985_ = ~new_n12969_ & ~new_n12984_;
  assign new_n12986_ = ~new_n12946_ & new_n12960_;
  assign new_n12987_ = new_n12946_ & ~new_n12960_;
  assign new_n12988_ = ~new_n12986_ & ~new_n12987_;
  assign new_n12989_ = new_n12985_ & ~new_n12988_;
  assign A4660 = new_n12982_ | new_n12989_;
  assign new_n12991_ = ~new_n12953_ & ~new_n12989_;
  assign new_n12992_ = new_n12953_ & new_n12989_;
  assign new_n12993_ = ~new_n12991_ & ~new_n12992_;
  assign A4659 = ~new_n12946_ & ~new_n12993_;
  assign new_n12995_ = ~new_n9610_ & ~new_n9620_;
  assign new_n12996_ = ~new_n9613_ & ~new_n12995_;
  assign new_n12997_ = new_n9613_ & ~new_n12996_;
  assign new_n12998_ = new_n9613_ & new_n12995_;
  assign new_n12999_ = new_n12997_ & ~new_n12998_;
  assign new_n13000_ = ~new_n9620_ & ~new_n12999_;
  assign new_n13001_ = ~new_n9637_ & ~new_n13000_;
  assign new_n13002_ = ~new_n9655_ & ~new_n9665_;
  assign new_n13003_ = ~new_n9658_ & ~new_n13002_;
  assign new_n13004_ = new_n9658_ & ~new_n13003_;
  assign new_n13005_ = new_n9658_ & new_n13002_;
  assign new_n13006_ = new_n13004_ & ~new_n13005_;
  assign new_n13007_ = ~new_n9665_ & ~new_n13006_;
  assign new_n13008_ = ~new_n9682_ & ~new_n13007_;
  assign new_n13009_ = new_n13001_ & ~new_n13008_;
  assign new_n13010_ = ~new_n13001_ & new_n13008_;
  assign new_n13011_ = ~new_n13009_ & ~new_n13010_;
  assign new_n13012_ = ~new_n9703_ & ~new_n9713_;
  assign new_n13013_ = ~new_n9706_ & ~new_n13012_;
  assign new_n13014_ = new_n9706_ & ~new_n13013_;
  assign new_n13015_ = new_n9706_ & new_n13012_;
  assign new_n13016_ = new_n13014_ & ~new_n13015_;
  assign new_n13017_ = ~new_n9713_ & ~new_n13016_;
  assign new_n13018_ = ~new_n9730_ & ~new_n13017_;
  assign new_n13019_ = ~new_n9748_ & ~new_n9758_;
  assign new_n13020_ = ~new_n9751_ & ~new_n13019_;
  assign new_n13021_ = new_n9751_ & ~new_n13020_;
  assign new_n13022_ = new_n9751_ & new_n13019_;
  assign new_n13023_ = new_n13021_ & ~new_n13022_;
  assign new_n13024_ = ~new_n9758_ & ~new_n13023_;
  assign new_n13025_ = ~new_n9775_ & ~new_n13024_;
  assign new_n13026_ = new_n13011_ & new_n13025_;
  assign new_n13027_ = ~new_n9794_ & ~new_n9804_;
  assign new_n13028_ = ~new_n9797_ & ~new_n13027_;
  assign new_n13029_ = new_n9797_ & ~new_n13028_;
  assign new_n13030_ = new_n9797_ & new_n13027_;
  assign new_n13031_ = new_n13029_ & ~new_n13030_;
  assign new_n13032_ = ~new_n9804_ & ~new_n13031_;
  assign new_n13033_ = ~new_n9821_ & ~new_n13032_;
  assign new_n13034_ = new_n13025_ & new_n13033_;
  assign new_n13035_ = ~new_n13026_ & ~new_n13034_;
  assign new_n13036_ = ~new_n13018_ & new_n13035_;
  assign new_n13037_ = new_n13018_ & ~new_n13035_;
  assign new_n13038_ = ~new_n13036_ & ~new_n13037_;
  assign A4630 = ~new_n13011_ & ~new_n13038_;
  assign new_n13040_ = new_n13008_ & ~new_n13036_;
  assign A4629 = ~new_n13011_ & ~new_n13040_;
  assign new_n13042_ = ~new_n13008_ & ~new_n13018_;
  assign new_n13043_ = ~new_n13011_ & ~new_n13042_;
  assign new_n13044_ = new_n13011_ & ~new_n13043_;
  assign new_n13045_ = new_n13011_ & new_n13042_;
  assign new_n13046_ = new_n13044_ & ~new_n13045_;
  assign new_n13047_ = ~new_n13018_ & ~new_n13046_;
  assign A4628 = new_n13035_ | new_n13047_;
  assign new_n13049_ = ~new_n13025_ & ~new_n13033_;
  assign new_n13050_ = ~new_n13034_ & ~new_n13049_;
  assign new_n13051_ = ~new_n13011_ & new_n13025_;
  assign new_n13052_ = new_n13011_ & ~new_n13025_;
  assign new_n13053_ = ~new_n13051_ & ~new_n13052_;
  assign new_n13054_ = new_n13050_ & ~new_n13053_;
  assign A4627 = new_n13047_ | new_n13054_;
  assign new_n13056_ = ~new_n13018_ & ~new_n13054_;
  assign new_n13057_ = new_n13018_ & new_n13054_;
  assign new_n13058_ = ~new_n13056_ & ~new_n13057_;
  assign A4626 = ~new_n13011_ & ~new_n13058_;
  assign new_n13060_ = new_n9859_ & new_n9866_;
  assign new_n13061_ = ~new_n9862_ & ~new_n13060_;
  assign new_n13062_ = new_n9862_ & ~new_n13061_;
  assign new_n13063_ = new_n9862_ & new_n13060_;
  assign new_n13064_ = new_n13062_ & ~new_n13063_;
  assign new_n13065_ = new_n9866_ & ~new_n13064_;
  assign new_n13066_ = ~new_n9877_ & ~new_n13065_;
  assign new_n13067_ = new_n9889_ & new_n9896_;
  assign new_n13068_ = ~new_n9892_ & ~new_n13067_;
  assign new_n13069_ = new_n9892_ & ~new_n13068_;
  assign new_n13070_ = new_n9892_ & new_n13067_;
  assign new_n13071_ = new_n13069_ & ~new_n13070_;
  assign new_n13072_ = new_n9896_ & ~new_n13071_;
  assign new_n13073_ = ~new_n9907_ & ~new_n13072_;
  assign new_n13074_ = new_n13066_ & ~new_n13073_;
  assign new_n13075_ = ~new_n13066_ & new_n13073_;
  assign new_n13076_ = ~new_n13074_ & ~new_n13075_;
  assign new_n13077_ = new_n9922_ & new_n9929_;
  assign new_n13078_ = ~new_n9925_ & ~new_n13077_;
  assign new_n13079_ = new_n9925_ & ~new_n13078_;
  assign new_n13080_ = new_n9925_ & new_n13077_;
  assign new_n13081_ = new_n13079_ & ~new_n13080_;
  assign new_n13082_ = new_n9929_ & ~new_n13081_;
  assign new_n13083_ = ~new_n9940_ & ~new_n13082_;
  assign new_n13084_ = new_n9952_ & new_n9959_;
  assign new_n13085_ = ~new_n9955_ & ~new_n13084_;
  assign new_n13086_ = new_n9955_ & ~new_n13085_;
  assign new_n13087_ = new_n9955_ & new_n13084_;
  assign new_n13088_ = new_n13086_ & ~new_n13087_;
  assign new_n13089_ = new_n9959_ & ~new_n13088_;
  assign new_n13090_ = ~new_n9970_ & ~new_n13089_;
  assign new_n13091_ = new_n13076_ & new_n13090_;
  assign new_n13092_ = new_n9983_ & new_n9990_;
  assign new_n13093_ = ~new_n9986_ & ~new_n13092_;
  assign new_n13094_ = new_n9986_ & ~new_n13093_;
  assign new_n13095_ = new_n9986_ & new_n13092_;
  assign new_n13096_ = new_n13094_ & ~new_n13095_;
  assign new_n13097_ = new_n9990_ & ~new_n13096_;
  assign new_n13098_ = ~new_n10001_ & ~new_n13097_;
  assign new_n13099_ = new_n13090_ & new_n13098_;
  assign new_n13100_ = ~new_n13091_ & ~new_n13099_;
  assign new_n13101_ = ~new_n13083_ & new_n13100_;
  assign new_n13102_ = new_n13083_ & ~new_n13100_;
  assign new_n13103_ = ~new_n13101_ & ~new_n13102_;
  assign A4597 = ~new_n13076_ & ~new_n13103_;
  assign new_n13105_ = new_n13073_ & ~new_n13101_;
  assign A4596 = ~new_n13076_ & ~new_n13105_;
  assign new_n13107_ = ~new_n13073_ & ~new_n13083_;
  assign new_n13108_ = ~new_n13076_ & ~new_n13107_;
  assign new_n13109_ = new_n13076_ & ~new_n13108_;
  assign new_n13110_ = new_n13076_ & new_n13107_;
  assign new_n13111_ = new_n13109_ & ~new_n13110_;
  assign new_n13112_ = ~new_n13083_ & ~new_n13111_;
  assign A4595 = new_n13100_ | new_n13112_;
  assign new_n13114_ = ~new_n13090_ & ~new_n13098_;
  assign new_n13115_ = ~new_n13099_ & ~new_n13114_;
  assign new_n13116_ = ~new_n13076_ & new_n13090_;
  assign new_n13117_ = new_n13076_ & ~new_n13090_;
  assign new_n13118_ = ~new_n13116_ & ~new_n13117_;
  assign new_n13119_ = new_n13115_ & ~new_n13118_;
  assign A4594 = new_n13112_ | new_n13119_;
  assign new_n13121_ = ~new_n13083_ & ~new_n13119_;
  assign new_n13122_ = new_n13083_ & new_n13119_;
  assign new_n13123_ = ~new_n13121_ & ~new_n13122_;
  assign A4593 = ~new_n13076_ & ~new_n13123_;
  assign new_n13125_ = new_n10039_ & new_n10046_;
  assign new_n13126_ = ~new_n10042_ & ~new_n13125_;
  assign new_n13127_ = new_n10042_ & ~new_n13126_;
  assign new_n13128_ = new_n10042_ & new_n13125_;
  assign new_n13129_ = new_n13127_ & ~new_n13128_;
  assign new_n13130_ = new_n10046_ & ~new_n13129_;
  assign new_n13131_ = ~new_n10057_ & ~new_n13130_;
  assign new_n13132_ = new_n10069_ & new_n10076_;
  assign new_n13133_ = ~new_n10072_ & ~new_n13132_;
  assign new_n13134_ = new_n10072_ & ~new_n13133_;
  assign new_n13135_ = new_n10072_ & new_n13132_;
  assign new_n13136_ = new_n13134_ & ~new_n13135_;
  assign new_n13137_ = new_n10076_ & ~new_n13136_;
  assign new_n13138_ = ~new_n10087_ & ~new_n13137_;
  assign new_n13139_ = new_n13131_ & ~new_n13138_;
  assign new_n13140_ = ~new_n13131_ & new_n13138_;
  assign new_n13141_ = ~new_n13139_ & ~new_n13140_;
  assign new_n13142_ = new_n10102_ & new_n10109_;
  assign new_n13143_ = ~new_n10105_ & ~new_n13142_;
  assign new_n13144_ = new_n10105_ & ~new_n13143_;
  assign new_n13145_ = new_n10105_ & new_n13142_;
  assign new_n13146_ = new_n13144_ & ~new_n13145_;
  assign new_n13147_ = new_n10109_ & ~new_n13146_;
  assign new_n13148_ = ~new_n10120_ & ~new_n13147_;
  assign new_n13149_ = new_n10132_ & new_n10139_;
  assign new_n13150_ = ~new_n10135_ & ~new_n13149_;
  assign new_n13151_ = new_n10135_ & ~new_n13150_;
  assign new_n13152_ = new_n10135_ & new_n13149_;
  assign new_n13153_ = new_n13151_ & ~new_n13152_;
  assign new_n13154_ = new_n10139_ & ~new_n13153_;
  assign new_n13155_ = ~new_n10150_ & ~new_n13154_;
  assign new_n13156_ = new_n13141_ & new_n13155_;
  assign new_n13157_ = new_n10163_ & new_n10170_;
  assign new_n13158_ = ~new_n10166_ & ~new_n13157_;
  assign new_n13159_ = new_n10166_ & ~new_n13158_;
  assign new_n13160_ = new_n10166_ & new_n13157_;
  assign new_n13161_ = new_n13159_ & ~new_n13160_;
  assign new_n13162_ = new_n10170_ & ~new_n13161_;
  assign new_n13163_ = ~new_n10181_ & ~new_n13162_;
  assign new_n13164_ = new_n13155_ & new_n13163_;
  assign new_n13165_ = ~new_n13156_ & ~new_n13164_;
  assign new_n13166_ = ~new_n13148_ & new_n13165_;
  assign new_n13167_ = new_n13148_ & ~new_n13165_;
  assign new_n13168_ = ~new_n13166_ & ~new_n13167_;
  assign A4564 = ~new_n13141_ & ~new_n13168_;
  assign new_n13170_ = new_n13138_ & ~new_n13166_;
  assign A4563 = ~new_n13141_ & ~new_n13170_;
  assign new_n13172_ = ~new_n13138_ & ~new_n13148_;
  assign new_n13173_ = ~new_n13141_ & ~new_n13172_;
  assign new_n13174_ = new_n13141_ & ~new_n13173_;
  assign new_n13175_ = new_n13141_ & new_n13172_;
  assign new_n13176_ = new_n13174_ & ~new_n13175_;
  assign new_n13177_ = ~new_n13148_ & ~new_n13176_;
  assign A4562 = new_n13165_ | new_n13177_;
  assign new_n13179_ = ~new_n13155_ & ~new_n13163_;
  assign new_n13180_ = ~new_n13164_ & ~new_n13179_;
  assign new_n13181_ = ~new_n13141_ & new_n13155_;
  assign new_n13182_ = new_n13141_ & ~new_n13155_;
  assign new_n13183_ = ~new_n13181_ & ~new_n13182_;
  assign new_n13184_ = new_n13180_ & ~new_n13183_;
  assign A4561 = new_n13177_ | new_n13184_;
  assign new_n13186_ = ~new_n13148_ & ~new_n13184_;
  assign new_n13187_ = new_n13148_ & new_n13184_;
  assign new_n13188_ = ~new_n13186_ & ~new_n13187_;
  assign A4560 = ~new_n13141_ & ~new_n13188_;
  assign new_n13190_ = new_n10219_ & new_n10226_;
  assign new_n13191_ = ~new_n10222_ & ~new_n13190_;
  assign new_n13192_ = new_n10222_ & ~new_n13191_;
  assign new_n13193_ = new_n10222_ & new_n13190_;
  assign new_n13194_ = new_n13192_ & ~new_n13193_;
  assign new_n13195_ = new_n10226_ & ~new_n13194_;
  assign new_n13196_ = ~new_n10237_ & ~new_n13195_;
  assign new_n13197_ = new_n10249_ & new_n10256_;
  assign new_n13198_ = ~new_n10252_ & ~new_n13197_;
  assign new_n13199_ = new_n10252_ & ~new_n13198_;
  assign new_n13200_ = new_n10252_ & new_n13197_;
  assign new_n13201_ = new_n13199_ & ~new_n13200_;
  assign new_n13202_ = new_n10256_ & ~new_n13201_;
  assign new_n13203_ = ~new_n10267_ & ~new_n13202_;
  assign new_n13204_ = new_n13196_ & ~new_n13203_;
  assign new_n13205_ = ~new_n13196_ & new_n13203_;
  assign new_n13206_ = ~new_n13204_ & ~new_n13205_;
  assign new_n13207_ = new_n10282_ & new_n10289_;
  assign new_n13208_ = ~new_n10285_ & ~new_n13207_;
  assign new_n13209_ = new_n10285_ & ~new_n13208_;
  assign new_n13210_ = new_n10285_ & new_n13207_;
  assign new_n13211_ = new_n13209_ & ~new_n13210_;
  assign new_n13212_ = new_n10289_ & ~new_n13211_;
  assign new_n13213_ = ~new_n10300_ & ~new_n13212_;
  assign new_n13214_ = new_n10312_ & new_n10319_;
  assign new_n13215_ = ~new_n10315_ & ~new_n13214_;
  assign new_n13216_ = new_n10315_ & ~new_n13215_;
  assign new_n13217_ = new_n10315_ & new_n13214_;
  assign new_n13218_ = new_n13216_ & ~new_n13217_;
  assign new_n13219_ = new_n10319_ & ~new_n13218_;
  assign new_n13220_ = ~new_n10330_ & ~new_n13219_;
  assign new_n13221_ = new_n13206_ & new_n13220_;
  assign new_n13222_ = new_n10343_ & new_n10350_;
  assign new_n13223_ = ~new_n10346_ & ~new_n13222_;
  assign new_n13224_ = new_n10346_ & ~new_n13223_;
  assign new_n13225_ = new_n10346_ & new_n13222_;
  assign new_n13226_ = new_n13224_ & ~new_n13225_;
  assign new_n13227_ = new_n10350_ & ~new_n13226_;
  assign new_n13228_ = ~new_n10361_ & ~new_n13227_;
  assign new_n13229_ = new_n13220_ & new_n13228_;
  assign new_n13230_ = ~new_n13221_ & ~new_n13229_;
  assign new_n13231_ = ~new_n13213_ & new_n13230_;
  assign new_n13232_ = new_n13213_ & ~new_n13230_;
  assign new_n13233_ = ~new_n13231_ & ~new_n13232_;
  assign A4531 = ~new_n13206_ & ~new_n13233_;
  assign new_n13235_ = new_n13203_ & ~new_n13231_;
  assign A4530 = ~new_n13206_ & ~new_n13235_;
  assign new_n13237_ = ~new_n13203_ & ~new_n13213_;
  assign new_n13238_ = ~new_n13206_ & ~new_n13237_;
  assign new_n13239_ = new_n13206_ & ~new_n13238_;
  assign new_n13240_ = new_n13206_ & new_n13237_;
  assign new_n13241_ = new_n13239_ & ~new_n13240_;
  assign new_n13242_ = ~new_n13213_ & ~new_n13241_;
  assign A4529 = new_n13230_ | new_n13242_;
  assign new_n13244_ = ~new_n13220_ & ~new_n13228_;
  assign new_n13245_ = ~new_n13229_ & ~new_n13244_;
  assign new_n13246_ = ~new_n13206_ & new_n13220_;
  assign new_n13247_ = new_n13206_ & ~new_n13220_;
  assign new_n13248_ = ~new_n13246_ & ~new_n13247_;
  assign new_n13249_ = new_n13245_ & ~new_n13248_;
  assign A4528 = new_n13242_ | new_n13249_;
  assign new_n13251_ = ~new_n13213_ & ~new_n13249_;
  assign new_n13252_ = new_n13213_ & new_n13249_;
  assign new_n13253_ = ~new_n13251_ & ~new_n13252_;
  assign A4527 = ~new_n13206_ & ~new_n13253_;
  assign new_n13255_ = new_n10399_ & new_n10406_;
  assign new_n13256_ = ~new_n10402_ & ~new_n13255_;
  assign new_n13257_ = new_n10402_ & ~new_n13256_;
  assign new_n13258_ = new_n10402_ & new_n13255_;
  assign new_n13259_ = new_n13257_ & ~new_n13258_;
  assign new_n13260_ = new_n10406_ & ~new_n13259_;
  assign new_n13261_ = ~new_n10417_ & ~new_n13260_;
  assign new_n13262_ = new_n10429_ & new_n10436_;
  assign new_n13263_ = ~new_n10432_ & ~new_n13262_;
  assign new_n13264_ = new_n10432_ & ~new_n13263_;
  assign new_n13265_ = new_n10432_ & new_n13262_;
  assign new_n13266_ = new_n13264_ & ~new_n13265_;
  assign new_n13267_ = new_n10436_ & ~new_n13266_;
  assign new_n13268_ = ~new_n10447_ & ~new_n13267_;
  assign new_n13269_ = new_n13261_ & ~new_n13268_;
  assign new_n13270_ = ~new_n13261_ & new_n13268_;
  assign new_n13271_ = ~new_n13269_ & ~new_n13270_;
  assign new_n13272_ = new_n10462_ & new_n10469_;
  assign new_n13273_ = ~new_n10465_ & ~new_n13272_;
  assign new_n13274_ = new_n10465_ & ~new_n13273_;
  assign new_n13275_ = new_n10465_ & new_n13272_;
  assign new_n13276_ = new_n13274_ & ~new_n13275_;
  assign new_n13277_ = new_n10469_ & ~new_n13276_;
  assign new_n13278_ = ~new_n10480_ & ~new_n13277_;
  assign new_n13279_ = new_n10492_ & new_n10499_;
  assign new_n13280_ = ~new_n10495_ & ~new_n13279_;
  assign new_n13281_ = new_n10495_ & ~new_n13280_;
  assign new_n13282_ = new_n10495_ & new_n13279_;
  assign new_n13283_ = new_n13281_ & ~new_n13282_;
  assign new_n13284_ = new_n10499_ & ~new_n13283_;
  assign new_n13285_ = ~new_n10510_ & ~new_n13284_;
  assign new_n13286_ = new_n13271_ & new_n13285_;
  assign new_n13287_ = new_n10523_ & new_n10530_;
  assign new_n13288_ = ~new_n10526_ & ~new_n13287_;
  assign new_n13289_ = new_n10526_ & ~new_n13288_;
  assign new_n13290_ = new_n10526_ & new_n13287_;
  assign new_n13291_ = new_n13289_ & ~new_n13290_;
  assign new_n13292_ = new_n10530_ & ~new_n13291_;
  assign new_n13293_ = ~new_n10541_ & ~new_n13292_;
  assign new_n13294_ = new_n13285_ & new_n13293_;
  assign new_n13295_ = ~new_n13286_ & ~new_n13294_;
  assign new_n13296_ = ~new_n13278_ & new_n13295_;
  assign new_n13297_ = new_n13278_ & ~new_n13295_;
  assign new_n13298_ = ~new_n13296_ & ~new_n13297_;
  assign A4498 = ~new_n13271_ & ~new_n13298_;
  assign new_n13300_ = new_n13268_ & ~new_n13296_;
  assign A4497 = ~new_n13271_ & ~new_n13300_;
  assign new_n13302_ = ~new_n13268_ & ~new_n13278_;
  assign new_n13303_ = ~new_n13271_ & ~new_n13302_;
  assign new_n13304_ = new_n13271_ & ~new_n13303_;
  assign new_n13305_ = new_n13271_ & new_n13302_;
  assign new_n13306_ = new_n13304_ & ~new_n13305_;
  assign new_n13307_ = ~new_n13278_ & ~new_n13306_;
  assign A4496 = new_n13295_ | new_n13307_;
  assign new_n13309_ = ~new_n13285_ & ~new_n13293_;
  assign new_n13310_ = ~new_n13294_ & ~new_n13309_;
  assign new_n13311_ = ~new_n13271_ & new_n13285_;
  assign new_n13312_ = new_n13271_ & ~new_n13285_;
  assign new_n13313_ = ~new_n13311_ & ~new_n13312_;
  assign new_n13314_ = new_n13310_ & ~new_n13313_;
  assign A4495 = new_n13307_ | new_n13314_;
  assign new_n13316_ = ~new_n13278_ & ~new_n13314_;
  assign new_n13317_ = new_n13278_ & new_n13314_;
  assign new_n13318_ = ~new_n13316_ & ~new_n13317_;
  assign A4494 = ~new_n13271_ & ~new_n13318_;
  assign new_n13320_ = ~new_n10575_ & new_n10592_;
  assign new_n13321_ = ~new_n10580_ & ~new_n13320_;
  assign new_n13322_ = ~new_n11720_ & ~new_n13321_;
  assign new_n13323_ = new_n10612_ & new_n10619_;
  assign new_n13324_ = ~new_n10615_ & ~new_n13323_;
  assign new_n13325_ = new_n10615_ & ~new_n13324_;
  assign new_n13326_ = new_n10615_ & new_n13323_;
  assign new_n13327_ = new_n13325_ & ~new_n13326_;
  assign new_n13328_ = new_n10619_ & ~new_n13327_;
  assign new_n13329_ = ~new_n10630_ & ~new_n13328_;
  assign new_n13330_ = new_n13322_ & ~new_n13329_;
  assign new_n13331_ = ~new_n13322_ & new_n13329_;
  assign new_n13332_ = ~new_n13330_ & ~new_n13331_;
  assign new_n13333_ = new_n10645_ & new_n10652_;
  assign new_n13334_ = ~new_n10648_ & ~new_n13333_;
  assign new_n13335_ = new_n10648_ & ~new_n13334_;
  assign new_n13336_ = new_n10648_ & new_n13333_;
  assign new_n13337_ = new_n13335_ & ~new_n13336_;
  assign new_n13338_ = new_n10652_ & ~new_n13337_;
  assign new_n13339_ = ~new_n10663_ & ~new_n13338_;
  assign new_n13340_ = new_n10675_ & new_n10682_;
  assign new_n13341_ = ~new_n10678_ & ~new_n13340_;
  assign new_n13342_ = new_n10678_ & ~new_n13341_;
  assign new_n13343_ = new_n10678_ & new_n13340_;
  assign new_n13344_ = new_n13342_ & ~new_n13343_;
  assign new_n13345_ = new_n10682_ & ~new_n13344_;
  assign new_n13346_ = ~new_n10693_ & ~new_n13345_;
  assign new_n13347_ = new_n13332_ & new_n13346_;
  assign new_n13348_ = new_n10706_ & new_n10713_;
  assign new_n13349_ = ~new_n10709_ & ~new_n13348_;
  assign new_n13350_ = new_n10709_ & ~new_n13349_;
  assign new_n13351_ = new_n10709_ & new_n13348_;
  assign new_n13352_ = new_n13350_ & ~new_n13351_;
  assign new_n13353_ = new_n10713_ & ~new_n13352_;
  assign new_n13354_ = ~new_n10724_ & ~new_n13353_;
  assign new_n13355_ = new_n13346_ & new_n13354_;
  assign new_n13356_ = ~new_n13347_ & ~new_n13355_;
  assign new_n13357_ = ~new_n13339_ & new_n13356_;
  assign new_n13358_ = new_n13339_ & ~new_n13356_;
  assign new_n13359_ = ~new_n13357_ & ~new_n13358_;
  assign A4465 = ~new_n13332_ & ~new_n13359_;
  assign new_n13361_ = new_n13329_ & ~new_n13357_;
  assign A4464 = ~new_n13332_ & ~new_n13361_;
  assign new_n13363_ = ~new_n13329_ & ~new_n13339_;
  assign new_n13364_ = ~new_n13332_ & ~new_n13363_;
  assign new_n13365_ = new_n13332_ & ~new_n13364_;
  assign new_n13366_ = new_n13332_ & new_n13363_;
  assign new_n13367_ = new_n13365_ & ~new_n13366_;
  assign new_n13368_ = ~new_n13339_ & ~new_n13367_;
  assign A4463 = new_n13356_ | new_n13368_;
  assign new_n13370_ = ~new_n13346_ & ~new_n13354_;
  assign new_n13371_ = ~new_n13355_ & ~new_n13370_;
  assign new_n13372_ = ~new_n13332_ & new_n13346_;
  assign new_n13373_ = new_n13332_ & ~new_n13346_;
  assign new_n13374_ = ~new_n13372_ & ~new_n13373_;
  assign new_n13375_ = new_n13371_ & ~new_n13374_;
  assign A4462 = new_n13368_ | new_n13375_;
  assign new_n13377_ = ~new_n13339_ & ~new_n13375_;
  assign new_n13378_ = new_n13339_ & new_n13375_;
  assign new_n13379_ = ~new_n13377_ & ~new_n13378_;
  assign A4461 = ~new_n13332_ & ~new_n13379_;
  assign new_n13381_ = new_n1497_ & new_n1558_;
  assign new_n13382_ = ~new_n1559_ & ~new_n13381_;
  assign new_n13383_ = ~new_n1377_ & ~new_n1497_;
  assign new_n13384_ = new_n1377_ & new_n1497_;
  assign new_n13385_ = ~new_n13383_ & ~new_n13384_;
  assign new_n13386_ = new_n13382_ & ~new_n13385_;
  assign new_n13387_ = ~new_n11765_ & ~new_n13386_;
  assign new_n13388_ = new_n1807_ & new_n1868_;
  assign new_n13389_ = ~new_n1869_ & ~new_n13388_;
  assign new_n13390_ = ~new_n1687_ & ~new_n1807_;
  assign new_n13391_ = new_n1687_ & new_n1807_;
  assign new_n13392_ = ~new_n13390_ & ~new_n13391_;
  assign new_n13393_ = new_n13389_ & ~new_n13392_;
  assign new_n13394_ = ~new_n11772_ & ~new_n13393_;
  assign new_n13395_ = new_n13387_ & ~new_n13394_;
  assign new_n13396_ = ~new_n13387_ & new_n13394_;
  assign new_n13397_ = ~new_n13395_ & ~new_n13396_;
  assign new_n13398_ = new_n2120_ & new_n2181_;
  assign new_n13399_ = ~new_n2182_ & ~new_n13398_;
  assign new_n13400_ = ~new_n2000_ & ~new_n2120_;
  assign new_n13401_ = new_n2000_ & new_n2120_;
  assign new_n13402_ = ~new_n13400_ & ~new_n13401_;
  assign new_n13403_ = new_n13399_ & ~new_n13402_;
  assign new_n13404_ = ~new_n11782_ & ~new_n13403_;
  assign new_n13405_ = new_n2430_ & new_n2491_;
  assign new_n13406_ = ~new_n2492_ & ~new_n13405_;
  assign new_n13407_ = ~new_n2310_ & ~new_n2430_;
  assign new_n13408_ = new_n2310_ & new_n2430_;
  assign new_n13409_ = ~new_n13407_ & ~new_n13408_;
  assign new_n13410_ = new_n13406_ & ~new_n13409_;
  assign new_n13411_ = ~new_n11789_ & ~new_n13410_;
  assign new_n13412_ = new_n13397_ & new_n13411_;
  assign new_n13413_ = new_n2741_ & new_n2802_;
  assign new_n13414_ = ~new_n2803_ & ~new_n13413_;
  assign new_n13415_ = ~new_n2621_ & ~new_n2741_;
  assign new_n13416_ = new_n2621_ & new_n2741_;
  assign new_n13417_ = ~new_n13415_ & ~new_n13416_;
  assign new_n13418_ = new_n13414_ & ~new_n13417_;
  assign new_n13419_ = ~new_n11797_ & ~new_n13418_;
  assign new_n13420_ = new_n13411_ & new_n13419_;
  assign new_n13421_ = ~new_n13412_ & ~new_n13420_;
  assign new_n13422_ = ~new_n13404_ & new_n13421_;
  assign new_n13423_ = new_n13404_ & ~new_n13421_;
  assign new_n13424_ = ~new_n13422_ & ~new_n13423_;
  assign A4432 = ~new_n13397_ & ~new_n13424_;
  assign new_n13426_ = new_n13394_ & ~new_n13422_;
  assign A4431 = ~new_n13397_ & ~new_n13426_;
  assign new_n13428_ = ~new_n13394_ & ~new_n13404_;
  assign new_n13429_ = ~new_n13397_ & ~new_n13428_;
  assign new_n13430_ = new_n13397_ & ~new_n13429_;
  assign new_n13431_ = new_n13397_ & new_n13428_;
  assign new_n13432_ = new_n13430_ & ~new_n13431_;
  assign new_n13433_ = ~new_n13404_ & ~new_n13432_;
  assign A4430 = new_n13421_ | new_n13433_;
  assign new_n13435_ = ~new_n13411_ & ~new_n13419_;
  assign new_n13436_ = ~new_n13420_ & ~new_n13435_;
  assign new_n13437_ = ~new_n13397_ & new_n13411_;
  assign new_n13438_ = new_n13397_ & ~new_n13411_;
  assign new_n13439_ = ~new_n13437_ & ~new_n13438_;
  assign new_n13440_ = new_n13436_ & ~new_n13439_;
  assign A4429 = new_n13433_ | new_n13440_;
  assign new_n13442_ = ~new_n13404_ & ~new_n13440_;
  assign new_n13443_ = new_n13404_ & new_n13440_;
  assign new_n13444_ = ~new_n13442_ & ~new_n13443_;
  assign A4428 = ~new_n13397_ & ~new_n13444_;
  assign new_n13446_ = new_n2922_ & new_n2943_;
  assign new_n13447_ = ~new_n2944_ & ~new_n13446_;
  assign new_n13448_ = ~new_n2882_ & ~new_n2922_;
  assign new_n13449_ = new_n2882_ & new_n2922_;
  assign new_n13450_ = ~new_n13448_ & ~new_n13449_;
  assign new_n13451_ = new_n13447_ & ~new_n13450_;
  assign new_n13452_ = ~new_n11830_ & ~new_n13451_;
  assign new_n13453_ = new_n3032_ & new_n3053_;
  assign new_n13454_ = ~new_n3054_ & ~new_n13453_;
  assign new_n13455_ = ~new_n2992_ & ~new_n3032_;
  assign new_n13456_ = new_n2992_ & new_n3032_;
  assign new_n13457_ = ~new_n13455_ & ~new_n13456_;
  assign new_n13458_ = new_n13454_ & ~new_n13457_;
  assign new_n13459_ = ~new_n11837_ & ~new_n13458_;
  assign new_n13460_ = new_n13452_ & ~new_n13459_;
  assign new_n13461_ = ~new_n13452_ & new_n13459_;
  assign new_n13462_ = ~new_n13460_ & ~new_n13461_;
  assign new_n13463_ = new_n3145_ & new_n3166_;
  assign new_n13464_ = ~new_n3167_ & ~new_n13463_;
  assign new_n13465_ = ~new_n3105_ & ~new_n3145_;
  assign new_n13466_ = new_n3105_ & new_n3145_;
  assign new_n13467_ = ~new_n13465_ & ~new_n13466_;
  assign new_n13468_ = new_n13464_ & ~new_n13467_;
  assign new_n13469_ = ~new_n11847_ & ~new_n13468_;
  assign new_n13470_ = new_n3255_ & new_n3276_;
  assign new_n13471_ = ~new_n3277_ & ~new_n13470_;
  assign new_n13472_ = ~new_n3215_ & ~new_n3255_;
  assign new_n13473_ = new_n3215_ & new_n3255_;
  assign new_n13474_ = ~new_n13472_ & ~new_n13473_;
  assign new_n13475_ = new_n13471_ & ~new_n13474_;
  assign new_n13476_ = ~new_n11854_ & ~new_n13475_;
  assign new_n13477_ = new_n13462_ & new_n13476_;
  assign new_n13478_ = new_n3366_ & new_n3387_;
  assign new_n13479_ = ~new_n3388_ & ~new_n13478_;
  assign new_n13480_ = ~new_n3326_ & ~new_n3366_;
  assign new_n13481_ = new_n3326_ & new_n3366_;
  assign new_n13482_ = ~new_n13480_ & ~new_n13481_;
  assign new_n13483_ = new_n13479_ & ~new_n13482_;
  assign new_n13484_ = ~new_n11862_ & ~new_n13483_;
  assign new_n13485_ = new_n13476_ & new_n13484_;
  assign new_n13486_ = ~new_n13477_ & ~new_n13485_;
  assign new_n13487_ = ~new_n13469_ & new_n13486_;
  assign new_n13488_ = new_n13469_ & ~new_n13486_;
  assign new_n13489_ = ~new_n13487_ & ~new_n13488_;
  assign A4399 = ~new_n13462_ & ~new_n13489_;
  assign new_n13491_ = new_n13459_ & ~new_n13487_;
  assign A4398 = ~new_n13462_ & ~new_n13491_;
  assign new_n13493_ = ~new_n13459_ & ~new_n13469_;
  assign new_n13494_ = ~new_n13462_ & ~new_n13493_;
  assign new_n13495_ = new_n13462_ & ~new_n13494_;
  assign new_n13496_ = new_n13462_ & new_n13493_;
  assign new_n13497_ = new_n13495_ & ~new_n13496_;
  assign new_n13498_ = ~new_n13469_ & ~new_n13497_;
  assign A4397 = new_n13486_ | new_n13498_;
  assign new_n13500_ = ~new_n13476_ & ~new_n13484_;
  assign new_n13501_ = ~new_n13485_ & ~new_n13500_;
  assign new_n13502_ = ~new_n13462_ & new_n13476_;
  assign new_n13503_ = new_n13462_ & ~new_n13476_;
  assign new_n13504_ = ~new_n13502_ & ~new_n13503_;
  assign new_n13505_ = new_n13501_ & ~new_n13504_;
  assign A4396 = new_n13498_ | new_n13505_;
  assign new_n13507_ = ~new_n13469_ & ~new_n13505_;
  assign new_n13508_ = new_n13469_ & new_n13505_;
  assign new_n13509_ = ~new_n13507_ & ~new_n13508_;
  assign A4395 = ~new_n13462_ & ~new_n13509_;
  assign new_n13511_ = new_n3598_ & new_n3644_;
  assign new_n13512_ = ~new_n3645_ & ~new_n13511_;
  assign new_n13513_ = ~new_n3508_ & ~new_n3598_;
  assign new_n13514_ = new_n3508_ & new_n3598_;
  assign new_n13515_ = ~new_n13513_ & ~new_n13514_;
  assign new_n13516_ = new_n13512_ & ~new_n13515_;
  assign new_n13517_ = ~new_n11895_ & ~new_n13516_;
  assign new_n13518_ = new_n3833_ & new_n3879_;
  assign new_n13519_ = ~new_n3880_ & ~new_n13518_;
  assign new_n13520_ = ~new_n3743_ & ~new_n3833_;
  assign new_n13521_ = new_n3743_ & new_n3833_;
  assign new_n13522_ = ~new_n13520_ & ~new_n13521_;
  assign new_n13523_ = new_n13519_ & ~new_n13522_;
  assign new_n13524_ = ~new_n11902_ & ~new_n13523_;
  assign new_n13525_ = new_n13517_ & ~new_n13524_;
  assign new_n13526_ = ~new_n13517_ & new_n13524_;
  assign new_n13527_ = ~new_n13525_ & ~new_n13526_;
  assign new_n13528_ = new_n4071_ & new_n4117_;
  assign new_n13529_ = ~new_n4118_ & ~new_n13528_;
  assign new_n13530_ = ~new_n3981_ & ~new_n4071_;
  assign new_n13531_ = new_n3981_ & new_n4071_;
  assign new_n13532_ = ~new_n13530_ & ~new_n13531_;
  assign new_n13533_ = new_n13529_ & ~new_n13532_;
  assign new_n13534_ = ~new_n11912_ & ~new_n13533_;
  assign new_n13535_ = new_n4306_ & new_n4352_;
  assign new_n13536_ = ~new_n4353_ & ~new_n13535_;
  assign new_n13537_ = ~new_n4216_ & ~new_n4306_;
  assign new_n13538_ = new_n4216_ & new_n4306_;
  assign new_n13539_ = ~new_n13537_ & ~new_n13538_;
  assign new_n13540_ = new_n13536_ & ~new_n13539_;
  assign new_n13541_ = ~new_n11919_ & ~new_n13540_;
  assign new_n13542_ = new_n13527_ & new_n13541_;
  assign new_n13543_ = new_n4542_ & new_n4588_;
  assign new_n13544_ = ~new_n4589_ & ~new_n13543_;
  assign new_n13545_ = ~new_n4452_ & ~new_n4542_;
  assign new_n13546_ = new_n4452_ & new_n4542_;
  assign new_n13547_ = ~new_n13545_ & ~new_n13546_;
  assign new_n13548_ = new_n13544_ & ~new_n13547_;
  assign new_n13549_ = ~new_n11927_ & ~new_n13548_;
  assign new_n13550_ = new_n13541_ & new_n13549_;
  assign new_n13551_ = ~new_n13542_ & ~new_n13550_;
  assign new_n13552_ = ~new_n13534_ & new_n13551_;
  assign new_n13553_ = new_n13534_ & ~new_n13551_;
  assign new_n13554_ = ~new_n13552_ & ~new_n13553_;
  assign A4366 = ~new_n13527_ & ~new_n13554_;
  assign new_n13556_ = new_n13524_ & ~new_n13552_;
  assign A4365 = ~new_n13527_ & ~new_n13556_;
  assign new_n13558_ = ~new_n13524_ & ~new_n13534_;
  assign new_n13559_ = ~new_n13527_ & ~new_n13558_;
  assign new_n13560_ = new_n13527_ & ~new_n13559_;
  assign new_n13561_ = new_n13527_ & new_n13558_;
  assign new_n13562_ = new_n13560_ & ~new_n13561_;
  assign new_n13563_ = ~new_n13534_ & ~new_n13562_;
  assign A4364 = new_n13551_ | new_n13563_;
  assign new_n13565_ = ~new_n13541_ & ~new_n13549_;
  assign new_n13566_ = ~new_n13550_ & ~new_n13565_;
  assign new_n13567_ = ~new_n13527_ & new_n13541_;
  assign new_n13568_ = new_n13527_ & ~new_n13541_;
  assign new_n13569_ = ~new_n13567_ & ~new_n13568_;
  assign new_n13570_ = new_n13566_ & ~new_n13569_;
  assign A4363 = new_n13563_ | new_n13570_;
  assign new_n13572_ = ~new_n13534_ & ~new_n13570_;
  assign new_n13573_ = new_n13534_ & new_n13570_;
  assign new_n13574_ = ~new_n13572_ & ~new_n13573_;
  assign A4362 = ~new_n13527_ & ~new_n13574_;
  assign new_n13576_ = new_n4799_ & new_n4845_;
  assign new_n13577_ = ~new_n4846_ & ~new_n13576_;
  assign new_n13578_ = ~new_n4709_ & ~new_n4799_;
  assign new_n13579_ = new_n4709_ & new_n4799_;
  assign new_n13580_ = ~new_n13578_ & ~new_n13579_;
  assign new_n13581_ = new_n13577_ & ~new_n13580_;
  assign new_n13582_ = ~new_n11960_ & ~new_n13581_;
  assign new_n13583_ = new_n5034_ & new_n5080_;
  assign new_n13584_ = ~new_n5081_ & ~new_n13583_;
  assign new_n13585_ = ~new_n4944_ & ~new_n5034_;
  assign new_n13586_ = new_n4944_ & new_n5034_;
  assign new_n13587_ = ~new_n13585_ & ~new_n13586_;
  assign new_n13588_ = new_n13584_ & ~new_n13587_;
  assign new_n13589_ = ~new_n11967_ & ~new_n13588_;
  assign new_n13590_ = new_n13582_ & ~new_n13589_;
  assign new_n13591_ = ~new_n13582_ & new_n13589_;
  assign new_n13592_ = ~new_n13590_ & ~new_n13591_;
  assign new_n13593_ = new_n5272_ & new_n5318_;
  assign new_n13594_ = ~new_n5319_ & ~new_n13593_;
  assign new_n13595_ = ~new_n5182_ & ~new_n5272_;
  assign new_n13596_ = new_n5182_ & new_n5272_;
  assign new_n13597_ = ~new_n13595_ & ~new_n13596_;
  assign new_n13598_ = new_n13594_ & ~new_n13597_;
  assign new_n13599_ = ~new_n11977_ & ~new_n13598_;
  assign new_n13600_ = new_n5507_ & new_n5553_;
  assign new_n13601_ = ~new_n5554_ & ~new_n13600_;
  assign new_n13602_ = ~new_n5417_ & ~new_n5507_;
  assign new_n13603_ = new_n5417_ & new_n5507_;
  assign new_n13604_ = ~new_n13602_ & ~new_n13603_;
  assign new_n13605_ = new_n13601_ & ~new_n13604_;
  assign new_n13606_ = ~new_n11984_ & ~new_n13605_;
  assign new_n13607_ = new_n13592_ & new_n13606_;
  assign new_n13608_ = new_n5743_ & new_n5789_;
  assign new_n13609_ = ~new_n5790_ & ~new_n13608_;
  assign new_n13610_ = ~new_n5653_ & ~new_n5743_;
  assign new_n13611_ = new_n5653_ & new_n5743_;
  assign new_n13612_ = ~new_n13610_ & ~new_n13611_;
  assign new_n13613_ = new_n13609_ & ~new_n13612_;
  assign new_n13614_ = ~new_n11992_ & ~new_n13613_;
  assign new_n13615_ = new_n13606_ & new_n13614_;
  assign new_n13616_ = ~new_n13607_ & ~new_n13615_;
  assign new_n13617_ = ~new_n13599_ & new_n13616_;
  assign new_n13618_ = new_n13599_ & ~new_n13616_;
  assign new_n13619_ = ~new_n13617_ & ~new_n13618_;
  assign A4333 = ~new_n13592_ & ~new_n13619_;
  assign new_n13621_ = new_n13589_ & ~new_n13617_;
  assign A4332 = ~new_n13592_ & ~new_n13621_;
  assign new_n13623_ = ~new_n13589_ & ~new_n13599_;
  assign new_n13624_ = ~new_n13592_ & ~new_n13623_;
  assign new_n13625_ = new_n13592_ & ~new_n13624_;
  assign new_n13626_ = new_n13592_ & new_n13623_;
  assign new_n13627_ = new_n13625_ & ~new_n13626_;
  assign new_n13628_ = ~new_n13599_ & ~new_n13627_;
  assign A4331 = new_n13616_ | new_n13628_;
  assign new_n13630_ = ~new_n13606_ & ~new_n13614_;
  assign new_n13631_ = ~new_n13615_ & ~new_n13630_;
  assign new_n13632_ = ~new_n13592_ & new_n13606_;
  assign new_n13633_ = new_n13592_ & ~new_n13606_;
  assign new_n13634_ = ~new_n13632_ & ~new_n13633_;
  assign new_n13635_ = new_n13631_ & ~new_n13634_;
  assign A4330 = new_n13628_ | new_n13635_;
  assign new_n13637_ = ~new_n13599_ & ~new_n13635_;
  assign new_n13638_ = new_n13599_ & new_n13635_;
  assign new_n13639_ = ~new_n13637_ & ~new_n13638_;
  assign A4329 = ~new_n13592_ & ~new_n13639_;
  assign new_n13641_ = new_n5947_ & new_n5978_;
  assign new_n13642_ = ~new_n5979_ & ~new_n13641_;
  assign new_n13643_ = ~new_n5887_ & ~new_n5947_;
  assign new_n13644_ = new_n5887_ & new_n5947_;
  assign new_n13645_ = ~new_n13643_ & ~new_n13644_;
  assign new_n13646_ = new_n13642_ & ~new_n13645_;
  assign new_n13647_ = ~new_n12025_ & ~new_n13646_;
  assign new_n13648_ = new_n6107_ & new_n6138_;
  assign new_n13649_ = ~new_n6139_ & ~new_n13648_;
  assign new_n13650_ = ~new_n6047_ & ~new_n6107_;
  assign new_n13651_ = new_n6047_ & new_n6107_;
  assign new_n13652_ = ~new_n13650_ & ~new_n13651_;
  assign new_n13653_ = new_n13649_ & ~new_n13652_;
  assign new_n13654_ = ~new_n12032_ & ~new_n13653_;
  assign new_n13655_ = new_n13647_ & ~new_n13654_;
  assign new_n13656_ = ~new_n13647_ & new_n13654_;
  assign new_n13657_ = ~new_n13655_ & ~new_n13656_;
  assign new_n13658_ = new_n6270_ & new_n6301_;
  assign new_n13659_ = ~new_n6302_ & ~new_n13658_;
  assign new_n13660_ = ~new_n6210_ & ~new_n6270_;
  assign new_n13661_ = new_n6210_ & new_n6270_;
  assign new_n13662_ = ~new_n13660_ & ~new_n13661_;
  assign new_n13663_ = new_n13659_ & ~new_n13662_;
  assign new_n13664_ = ~new_n12042_ & ~new_n13663_;
  assign new_n13665_ = new_n6430_ & new_n6461_;
  assign new_n13666_ = ~new_n6462_ & ~new_n13665_;
  assign new_n13667_ = ~new_n6370_ & ~new_n6430_;
  assign new_n13668_ = new_n6370_ & new_n6430_;
  assign new_n13669_ = ~new_n13667_ & ~new_n13668_;
  assign new_n13670_ = new_n13666_ & ~new_n13669_;
  assign new_n13671_ = ~new_n12049_ & ~new_n13670_;
  assign new_n13672_ = new_n13657_ & new_n13671_;
  assign new_n13673_ = new_n6591_ & new_n6622_;
  assign new_n13674_ = ~new_n6623_ & ~new_n13673_;
  assign new_n13675_ = ~new_n6531_ & ~new_n6591_;
  assign new_n13676_ = new_n6531_ & new_n6591_;
  assign new_n13677_ = ~new_n13675_ & ~new_n13676_;
  assign new_n13678_ = new_n13674_ & ~new_n13677_;
  assign new_n13679_ = ~new_n12057_ & ~new_n13678_;
  assign new_n13680_ = new_n13671_ & new_n13679_;
  assign new_n13681_ = ~new_n13672_ & ~new_n13680_;
  assign new_n13682_ = ~new_n13664_ & new_n13681_;
  assign new_n13683_ = new_n13664_ & ~new_n13681_;
  assign new_n13684_ = ~new_n13682_ & ~new_n13683_;
  assign A4300 = ~new_n13657_ & ~new_n13684_;
  assign new_n13686_ = new_n13654_ & ~new_n13682_;
  assign A4299 = ~new_n13657_ & ~new_n13686_;
  assign new_n13688_ = ~new_n13654_ & ~new_n13664_;
  assign new_n13689_ = ~new_n13657_ & ~new_n13688_;
  assign new_n13690_ = new_n13657_ & ~new_n13689_;
  assign new_n13691_ = new_n13657_ & new_n13688_;
  assign new_n13692_ = new_n13690_ & ~new_n13691_;
  assign new_n13693_ = ~new_n13664_ & ~new_n13692_;
  assign A4298 = new_n13681_ | new_n13693_;
  assign new_n13695_ = ~new_n13671_ & ~new_n13679_;
  assign new_n13696_ = ~new_n13680_ & ~new_n13695_;
  assign new_n13697_ = ~new_n13657_ & new_n13671_;
  assign new_n13698_ = new_n13657_ & ~new_n13671_;
  assign new_n13699_ = ~new_n13697_ & ~new_n13698_;
  assign new_n13700_ = new_n13696_ & ~new_n13699_;
  assign A4297 = new_n13693_ | new_n13700_;
  assign new_n13702_ = ~new_n13664_ & ~new_n13700_;
  assign new_n13703_ = new_n13664_ & new_n13700_;
  assign new_n13704_ = ~new_n13702_ & ~new_n13703_;
  assign A4296 = ~new_n13657_ & ~new_n13704_;
  assign new_n13706_ = new_n6665_ & new_n6668_;
  assign new_n13707_ = ~new_n6669_ & ~new_n13706_;
  assign new_n13708_ = ~new_n6661_ & ~new_n6665_;
  assign new_n13709_ = new_n6661_ & new_n6665_;
  assign new_n13710_ = ~new_n13708_ & ~new_n13709_;
  assign new_n13711_ = new_n13707_ & ~new_n13710_;
  assign new_n13712_ = ~new_n12090_ & ~new_n13711_;
  assign new_n13713_ = new_n6685_ & new_n6688_;
  assign new_n13714_ = ~new_n6689_ & ~new_n13713_;
  assign new_n13715_ = ~new_n6681_ & ~new_n6685_;
  assign new_n13716_ = new_n6681_ & new_n6685_;
  assign new_n13717_ = ~new_n13715_ & ~new_n13716_;
  assign new_n13718_ = new_n13714_ & ~new_n13717_;
  assign new_n13719_ = ~new_n12097_ & ~new_n13718_;
  assign new_n13720_ = new_n13712_ & ~new_n13719_;
  assign new_n13721_ = ~new_n13712_ & new_n13719_;
  assign new_n13722_ = ~new_n13720_ & ~new_n13721_;
  assign new_n13723_ = new_n6708_ & new_n6711_;
  assign new_n13724_ = ~new_n6712_ & ~new_n13723_;
  assign new_n13725_ = ~new_n6704_ & ~new_n6708_;
  assign new_n13726_ = new_n6704_ & new_n6708_;
  assign new_n13727_ = ~new_n13725_ & ~new_n13726_;
  assign new_n13728_ = new_n13724_ & ~new_n13727_;
  assign new_n13729_ = ~new_n12107_ & ~new_n13728_;
  assign new_n13730_ = new_n6728_ & new_n6731_;
  assign new_n13731_ = ~new_n6732_ & ~new_n13730_;
  assign new_n13732_ = ~new_n6724_ & ~new_n6728_;
  assign new_n13733_ = new_n6724_ & new_n6728_;
  assign new_n13734_ = ~new_n13732_ & ~new_n13733_;
  assign new_n13735_ = new_n13731_ & ~new_n13734_;
  assign new_n13736_ = ~new_n12114_ & ~new_n13735_;
  assign new_n13737_ = new_n13722_ & new_n13736_;
  assign new_n13738_ = new_n6749_ & new_n6752_;
  assign new_n13739_ = ~new_n6753_ & ~new_n13738_;
  assign new_n13740_ = ~new_n6745_ & ~new_n6749_;
  assign new_n13741_ = new_n6745_ & new_n6749_;
  assign new_n13742_ = ~new_n13740_ & ~new_n13741_;
  assign new_n13743_ = new_n13739_ & ~new_n13742_;
  assign new_n13744_ = ~new_n12122_ & ~new_n13743_;
  assign new_n13745_ = new_n13736_ & new_n13744_;
  assign new_n13746_ = ~new_n13737_ & ~new_n13745_;
  assign new_n13747_ = ~new_n13729_ & new_n13746_;
  assign new_n13748_ = new_n13729_ & ~new_n13746_;
  assign new_n13749_ = ~new_n13747_ & ~new_n13748_;
  assign A4267 = ~new_n13722_ & ~new_n13749_;
  assign new_n13751_ = new_n13719_ & ~new_n13747_;
  assign A4266 = ~new_n13722_ & ~new_n13751_;
  assign new_n13753_ = ~new_n13719_ & ~new_n13729_;
  assign new_n13754_ = ~new_n13722_ & ~new_n13753_;
  assign new_n13755_ = new_n13722_ & ~new_n13754_;
  assign new_n13756_ = new_n13722_ & new_n13753_;
  assign new_n13757_ = new_n13755_ & ~new_n13756_;
  assign new_n13758_ = ~new_n13729_ & ~new_n13757_;
  assign A4265 = new_n13746_ | new_n13758_;
  assign new_n13760_ = ~new_n13736_ & ~new_n13744_;
  assign new_n13761_ = ~new_n13745_ & ~new_n13760_;
  assign new_n13762_ = ~new_n13722_ & new_n13736_;
  assign new_n13763_ = new_n13722_ & ~new_n13736_;
  assign new_n13764_ = ~new_n13762_ & ~new_n13763_;
  assign new_n13765_ = new_n13761_ & ~new_n13764_;
  assign A4264 = new_n13758_ | new_n13765_;
  assign new_n13767_ = ~new_n13729_ & ~new_n13765_;
  assign new_n13768_ = new_n13729_ & new_n13765_;
  assign new_n13769_ = ~new_n13767_ & ~new_n13768_;
  assign A4263 = ~new_n13722_ & ~new_n13769_;
  assign new_n13771_ = new_n6795_ & new_n6798_;
  assign new_n13772_ = ~new_n6799_ & ~new_n13771_;
  assign new_n13773_ = ~new_n6791_ & ~new_n6795_;
  assign new_n13774_ = new_n6791_ & new_n6795_;
  assign new_n13775_ = ~new_n13773_ & ~new_n13774_;
  assign new_n13776_ = new_n13772_ & ~new_n13775_;
  assign new_n13777_ = ~new_n12155_ & ~new_n13776_;
  assign new_n13778_ = new_n6815_ & new_n6818_;
  assign new_n13779_ = ~new_n6819_ & ~new_n13778_;
  assign new_n13780_ = ~new_n6811_ & ~new_n6815_;
  assign new_n13781_ = new_n6811_ & new_n6815_;
  assign new_n13782_ = ~new_n13780_ & ~new_n13781_;
  assign new_n13783_ = new_n13779_ & ~new_n13782_;
  assign new_n13784_ = ~new_n12162_ & ~new_n13783_;
  assign new_n13785_ = new_n13777_ & ~new_n13784_;
  assign new_n13786_ = ~new_n13777_ & new_n13784_;
  assign new_n13787_ = ~new_n13785_ & ~new_n13786_;
  assign new_n13788_ = new_n6838_ & new_n6841_;
  assign new_n13789_ = ~new_n6842_ & ~new_n13788_;
  assign new_n13790_ = ~new_n6834_ & ~new_n6838_;
  assign new_n13791_ = new_n6834_ & new_n6838_;
  assign new_n13792_ = ~new_n13790_ & ~new_n13791_;
  assign new_n13793_ = new_n13789_ & ~new_n13792_;
  assign new_n13794_ = ~new_n12172_ & ~new_n13793_;
  assign new_n13795_ = new_n6858_ & new_n6861_;
  assign new_n13796_ = ~new_n6862_ & ~new_n13795_;
  assign new_n13797_ = ~new_n6854_ & ~new_n6858_;
  assign new_n13798_ = new_n6854_ & new_n6858_;
  assign new_n13799_ = ~new_n13797_ & ~new_n13798_;
  assign new_n13800_ = new_n13796_ & ~new_n13799_;
  assign new_n13801_ = ~new_n12179_ & ~new_n13800_;
  assign new_n13802_ = new_n13787_ & new_n13801_;
  assign new_n13803_ = new_n6879_ & new_n6882_;
  assign new_n13804_ = ~new_n6883_ & ~new_n13803_;
  assign new_n13805_ = ~new_n6875_ & ~new_n6879_;
  assign new_n13806_ = new_n6875_ & new_n6879_;
  assign new_n13807_ = ~new_n13805_ & ~new_n13806_;
  assign new_n13808_ = new_n13804_ & ~new_n13807_;
  assign new_n13809_ = ~new_n12187_ & ~new_n13808_;
  assign new_n13810_ = new_n13801_ & new_n13809_;
  assign new_n13811_ = ~new_n13802_ & ~new_n13810_;
  assign new_n13812_ = ~new_n13794_ & new_n13811_;
  assign new_n13813_ = new_n13794_ & ~new_n13811_;
  assign new_n13814_ = ~new_n13812_ & ~new_n13813_;
  assign A4234 = ~new_n13787_ & ~new_n13814_;
  assign new_n13816_ = new_n13784_ & ~new_n13812_;
  assign A4233 = ~new_n13787_ & ~new_n13816_;
  assign new_n13818_ = ~new_n13784_ & ~new_n13794_;
  assign new_n13819_ = ~new_n13787_ & ~new_n13818_;
  assign new_n13820_ = new_n13787_ & ~new_n13819_;
  assign new_n13821_ = new_n13787_ & new_n13818_;
  assign new_n13822_ = new_n13820_ & ~new_n13821_;
  assign new_n13823_ = ~new_n13794_ & ~new_n13822_;
  assign A4232 = new_n13811_ | new_n13823_;
  assign new_n13825_ = ~new_n13801_ & ~new_n13809_;
  assign new_n13826_ = ~new_n13810_ & ~new_n13825_;
  assign new_n13827_ = ~new_n13787_ & new_n13801_;
  assign new_n13828_ = new_n13787_ & ~new_n13801_;
  assign new_n13829_ = ~new_n13827_ & ~new_n13828_;
  assign new_n13830_ = new_n13826_ & ~new_n13829_;
  assign A4231 = new_n13823_ | new_n13830_;
  assign new_n13832_ = ~new_n13794_ & ~new_n13830_;
  assign new_n13833_ = new_n13794_ & new_n13830_;
  assign new_n13834_ = ~new_n13832_ & ~new_n13833_;
  assign A4230 = ~new_n13787_ & ~new_n13834_;
  assign new_n13836_ = new_n6925_ & new_n6928_;
  assign new_n13837_ = ~new_n6929_ & ~new_n13836_;
  assign new_n13838_ = ~new_n6921_ & ~new_n6925_;
  assign new_n13839_ = new_n6921_ & new_n6925_;
  assign new_n13840_ = ~new_n13838_ & ~new_n13839_;
  assign new_n13841_ = new_n13837_ & ~new_n13840_;
  assign new_n13842_ = ~new_n12220_ & ~new_n13841_;
  assign new_n13843_ = new_n6945_ & new_n6948_;
  assign new_n13844_ = ~new_n6949_ & ~new_n13843_;
  assign new_n13845_ = ~new_n6941_ & ~new_n6945_;
  assign new_n13846_ = new_n6941_ & new_n6945_;
  assign new_n13847_ = ~new_n13845_ & ~new_n13846_;
  assign new_n13848_ = new_n13844_ & ~new_n13847_;
  assign new_n13849_ = ~new_n12227_ & ~new_n13848_;
  assign new_n13850_ = new_n13842_ & ~new_n13849_;
  assign new_n13851_ = ~new_n13842_ & new_n13849_;
  assign new_n13852_ = ~new_n13850_ & ~new_n13851_;
  assign new_n13853_ = new_n6968_ & new_n6971_;
  assign new_n13854_ = ~new_n6972_ & ~new_n13853_;
  assign new_n13855_ = ~new_n6964_ & ~new_n6968_;
  assign new_n13856_ = new_n6964_ & new_n6968_;
  assign new_n13857_ = ~new_n13855_ & ~new_n13856_;
  assign new_n13858_ = new_n13854_ & ~new_n13857_;
  assign new_n13859_ = ~new_n12237_ & ~new_n13858_;
  assign new_n13860_ = new_n6988_ & new_n6991_;
  assign new_n13861_ = ~new_n6992_ & ~new_n13860_;
  assign new_n13862_ = ~new_n6984_ & ~new_n6988_;
  assign new_n13863_ = new_n6984_ & new_n6988_;
  assign new_n13864_ = ~new_n13862_ & ~new_n13863_;
  assign new_n13865_ = new_n13861_ & ~new_n13864_;
  assign new_n13866_ = ~new_n12244_ & ~new_n13865_;
  assign new_n13867_ = new_n13852_ & new_n13866_;
  assign new_n13868_ = new_n7009_ & new_n7012_;
  assign new_n13869_ = ~new_n7013_ & ~new_n13868_;
  assign new_n13870_ = ~new_n7005_ & ~new_n7009_;
  assign new_n13871_ = new_n7005_ & new_n7009_;
  assign new_n13872_ = ~new_n13870_ & ~new_n13871_;
  assign new_n13873_ = new_n13869_ & ~new_n13872_;
  assign new_n13874_ = ~new_n12252_ & ~new_n13873_;
  assign new_n13875_ = new_n13866_ & new_n13874_;
  assign new_n13876_ = ~new_n13867_ & ~new_n13875_;
  assign new_n13877_ = ~new_n13859_ & new_n13876_;
  assign new_n13878_ = new_n13859_ & ~new_n13876_;
  assign new_n13879_ = ~new_n13877_ & ~new_n13878_;
  assign A4201 = ~new_n13852_ & ~new_n13879_;
  assign new_n13881_ = new_n13849_ & ~new_n13877_;
  assign A4200 = ~new_n13852_ & ~new_n13881_;
  assign new_n13883_ = ~new_n13849_ & ~new_n13859_;
  assign new_n13884_ = ~new_n13852_ & ~new_n13883_;
  assign new_n13885_ = new_n13852_ & ~new_n13884_;
  assign new_n13886_ = new_n13852_ & new_n13883_;
  assign new_n13887_ = new_n13885_ & ~new_n13886_;
  assign new_n13888_ = ~new_n13859_ & ~new_n13887_;
  assign A4199 = new_n13876_ | new_n13888_;
  assign new_n13890_ = ~new_n13866_ & ~new_n13874_;
  assign new_n13891_ = ~new_n13875_ & ~new_n13890_;
  assign new_n13892_ = ~new_n13852_ & new_n13866_;
  assign new_n13893_ = new_n13852_ & ~new_n13866_;
  assign new_n13894_ = ~new_n13892_ & ~new_n13893_;
  assign new_n13895_ = new_n13891_ & ~new_n13894_;
  assign A4198 = new_n13888_ | new_n13895_;
  assign new_n13897_ = ~new_n13859_ & ~new_n13895_;
  assign new_n13898_ = new_n13859_ & new_n13895_;
  assign new_n13899_ = ~new_n13897_ & ~new_n13898_;
  assign A4197 = ~new_n13852_ & ~new_n13899_;
  assign new_n13901_ = new_n7055_ & new_n7058_;
  assign new_n13902_ = ~new_n7059_ & ~new_n13901_;
  assign new_n13903_ = ~new_n7051_ & ~new_n7055_;
  assign new_n13904_ = new_n7051_ & new_n7055_;
  assign new_n13905_ = ~new_n13903_ & ~new_n13904_;
  assign new_n13906_ = new_n13902_ & ~new_n13905_;
  assign new_n13907_ = ~new_n12285_ & ~new_n13906_;
  assign new_n13908_ = new_n7075_ & new_n7078_;
  assign new_n13909_ = ~new_n7079_ & ~new_n13908_;
  assign new_n13910_ = ~new_n7071_ & ~new_n7075_;
  assign new_n13911_ = new_n7071_ & new_n7075_;
  assign new_n13912_ = ~new_n13910_ & ~new_n13911_;
  assign new_n13913_ = new_n13909_ & ~new_n13912_;
  assign new_n13914_ = ~new_n12292_ & ~new_n13913_;
  assign new_n13915_ = new_n13907_ & ~new_n13914_;
  assign new_n13916_ = ~new_n13907_ & new_n13914_;
  assign new_n13917_ = ~new_n13915_ & ~new_n13916_;
  assign new_n13918_ = new_n7098_ & new_n7101_;
  assign new_n13919_ = ~new_n7102_ & ~new_n13918_;
  assign new_n13920_ = ~new_n7094_ & ~new_n7098_;
  assign new_n13921_ = new_n7094_ & new_n7098_;
  assign new_n13922_ = ~new_n13920_ & ~new_n13921_;
  assign new_n13923_ = new_n13919_ & ~new_n13922_;
  assign new_n13924_ = ~new_n12302_ & ~new_n13923_;
  assign new_n13925_ = new_n7118_ & new_n7121_;
  assign new_n13926_ = ~new_n7122_ & ~new_n13925_;
  assign new_n13927_ = ~new_n7114_ & ~new_n7118_;
  assign new_n13928_ = new_n7114_ & new_n7118_;
  assign new_n13929_ = ~new_n13927_ & ~new_n13928_;
  assign new_n13930_ = new_n13926_ & ~new_n13929_;
  assign new_n13931_ = ~new_n12309_ & ~new_n13930_;
  assign new_n13932_ = new_n13917_ & new_n13931_;
  assign new_n13933_ = new_n7139_ & new_n7142_;
  assign new_n13934_ = ~new_n7143_ & ~new_n13933_;
  assign new_n13935_ = ~new_n7135_ & ~new_n7139_;
  assign new_n13936_ = new_n7135_ & new_n7139_;
  assign new_n13937_ = ~new_n13935_ & ~new_n13936_;
  assign new_n13938_ = new_n13934_ & ~new_n13937_;
  assign new_n13939_ = ~new_n12317_ & ~new_n13938_;
  assign new_n13940_ = new_n13931_ & new_n13939_;
  assign new_n13941_ = ~new_n13932_ & ~new_n13940_;
  assign new_n13942_ = ~new_n13924_ & new_n13941_;
  assign new_n13943_ = new_n13924_ & ~new_n13941_;
  assign new_n13944_ = ~new_n13942_ & ~new_n13943_;
  assign A4168 = ~new_n13917_ & ~new_n13944_;
  assign new_n13946_ = new_n13914_ & ~new_n13942_;
  assign A4167 = ~new_n13917_ & ~new_n13946_;
  assign new_n13948_ = ~new_n13914_ & ~new_n13924_;
  assign new_n13949_ = ~new_n13917_ & ~new_n13948_;
  assign new_n13950_ = new_n13917_ & ~new_n13949_;
  assign new_n13951_ = new_n13917_ & new_n13948_;
  assign new_n13952_ = new_n13950_ & ~new_n13951_;
  assign new_n13953_ = ~new_n13924_ & ~new_n13952_;
  assign A4166 = new_n13941_ | new_n13953_;
  assign new_n13955_ = ~new_n13931_ & ~new_n13939_;
  assign new_n13956_ = ~new_n13940_ & ~new_n13955_;
  assign new_n13957_ = ~new_n13917_ & new_n13931_;
  assign new_n13958_ = new_n13917_ & ~new_n13931_;
  assign new_n13959_ = ~new_n13957_ & ~new_n13958_;
  assign new_n13960_ = new_n13956_ & ~new_n13959_;
  assign A4165 = new_n13953_ | new_n13960_;
  assign new_n13962_ = ~new_n13924_ & ~new_n13960_;
  assign new_n13963_ = new_n13924_ & new_n13960_;
  assign new_n13964_ = ~new_n13962_ & ~new_n13963_;
  assign A4164 = ~new_n13917_ & ~new_n13964_;
  assign new_n13966_ = new_n7190_ & new_n7193_;
  assign new_n13967_ = ~new_n7194_ & ~new_n13966_;
  assign new_n13968_ = ~new_n7186_ & ~new_n7190_;
  assign new_n13969_ = new_n7186_ & new_n7190_;
  assign new_n13970_ = ~new_n13968_ & ~new_n13969_;
  assign new_n13971_ = new_n13967_ & ~new_n13970_;
  assign new_n13972_ = ~new_n12350_ & ~new_n13971_;
  assign new_n13973_ = new_n7210_ & new_n7213_;
  assign new_n13974_ = ~new_n7214_ & ~new_n13973_;
  assign new_n13975_ = ~new_n7206_ & ~new_n7210_;
  assign new_n13976_ = new_n7206_ & new_n7210_;
  assign new_n13977_ = ~new_n13975_ & ~new_n13976_;
  assign new_n13978_ = new_n13974_ & ~new_n13977_;
  assign new_n13979_ = ~new_n12357_ & ~new_n13978_;
  assign new_n13980_ = new_n13972_ & ~new_n13979_;
  assign new_n13981_ = ~new_n13972_ & new_n13979_;
  assign new_n13982_ = ~new_n13980_ & ~new_n13981_;
  assign new_n13983_ = new_n7233_ & new_n7236_;
  assign new_n13984_ = ~new_n7237_ & ~new_n13983_;
  assign new_n13985_ = ~new_n7229_ & ~new_n7233_;
  assign new_n13986_ = new_n7229_ & new_n7233_;
  assign new_n13987_ = ~new_n13985_ & ~new_n13986_;
  assign new_n13988_ = new_n13984_ & ~new_n13987_;
  assign new_n13989_ = ~new_n12367_ & ~new_n13988_;
  assign new_n13990_ = new_n7253_ & new_n7256_;
  assign new_n13991_ = ~new_n7257_ & ~new_n13990_;
  assign new_n13992_ = ~new_n7249_ & ~new_n7253_;
  assign new_n13993_ = new_n7249_ & new_n7253_;
  assign new_n13994_ = ~new_n13992_ & ~new_n13993_;
  assign new_n13995_ = new_n13991_ & ~new_n13994_;
  assign new_n13996_ = ~new_n12374_ & ~new_n13995_;
  assign new_n13997_ = new_n13982_ & new_n13996_;
  assign new_n13998_ = new_n7274_ & new_n7277_;
  assign new_n13999_ = ~new_n7278_ & ~new_n13998_;
  assign new_n14000_ = ~new_n7270_ & ~new_n7274_;
  assign new_n14001_ = new_n7270_ & new_n7274_;
  assign new_n14002_ = ~new_n14000_ & ~new_n14001_;
  assign new_n14003_ = new_n13999_ & ~new_n14002_;
  assign new_n14004_ = ~new_n12382_ & ~new_n14003_;
  assign new_n14005_ = new_n13996_ & new_n14004_;
  assign new_n14006_ = ~new_n13997_ & ~new_n14005_;
  assign new_n14007_ = ~new_n13989_ & new_n14006_;
  assign new_n14008_ = new_n13989_ & ~new_n14006_;
  assign new_n14009_ = ~new_n14007_ & ~new_n14008_;
  assign A4135 = ~new_n13982_ & ~new_n14009_;
  assign new_n14011_ = new_n13979_ & ~new_n14007_;
  assign A4134 = ~new_n13982_ & ~new_n14011_;
  assign new_n14013_ = ~new_n13979_ & ~new_n13989_;
  assign new_n14014_ = ~new_n13982_ & ~new_n14013_;
  assign new_n14015_ = new_n13982_ & ~new_n14014_;
  assign new_n14016_ = new_n13982_ & new_n14013_;
  assign new_n14017_ = new_n14015_ & ~new_n14016_;
  assign new_n14018_ = ~new_n13989_ & ~new_n14017_;
  assign A4133 = new_n14006_ | new_n14018_;
  assign new_n14020_ = ~new_n13996_ & ~new_n14004_;
  assign new_n14021_ = ~new_n14005_ & ~new_n14020_;
  assign new_n14022_ = ~new_n13982_ & new_n13996_;
  assign new_n14023_ = new_n13982_ & ~new_n13996_;
  assign new_n14024_ = ~new_n14022_ & ~new_n14023_;
  assign new_n14025_ = new_n14021_ & ~new_n14024_;
  assign A4132 = new_n14018_ | new_n14025_;
  assign new_n14027_ = ~new_n13989_ & ~new_n14025_;
  assign new_n14028_ = new_n13989_ & new_n14025_;
  assign new_n14029_ = ~new_n14027_ & ~new_n14028_;
  assign A4131 = ~new_n13982_ & ~new_n14029_;
  assign new_n14031_ = ~new_n7340_ & ~new_n7348_;
  assign new_n14032_ = ~new_n7349_ & ~new_n14031_;
  assign new_n14033_ = ~new_n7326_ & new_n7340_;
  assign new_n14034_ = new_n7326_ & ~new_n7340_;
  assign new_n14035_ = ~new_n14033_ & ~new_n14034_;
  assign new_n14036_ = new_n14032_ & ~new_n14035_;
  assign new_n14037_ = ~new_n12415_ & ~new_n14036_;
  assign new_n14038_ = ~new_n7385_ & ~new_n7393_;
  assign new_n14039_ = ~new_n7394_ & ~new_n14038_;
  assign new_n14040_ = ~new_n7371_ & new_n7385_;
  assign new_n14041_ = new_n7371_ & ~new_n7385_;
  assign new_n14042_ = ~new_n14040_ & ~new_n14041_;
  assign new_n14043_ = new_n14039_ & ~new_n14042_;
  assign new_n14044_ = ~new_n12422_ & ~new_n14043_;
  assign new_n14045_ = new_n14037_ & ~new_n14044_;
  assign new_n14046_ = ~new_n14037_ & new_n14044_;
  assign new_n14047_ = ~new_n14045_ & ~new_n14046_;
  assign new_n14048_ = ~new_n7433_ & ~new_n7441_;
  assign new_n14049_ = ~new_n7442_ & ~new_n14048_;
  assign new_n14050_ = ~new_n7419_ & new_n7433_;
  assign new_n14051_ = new_n7419_ & ~new_n7433_;
  assign new_n14052_ = ~new_n14050_ & ~new_n14051_;
  assign new_n14053_ = new_n14049_ & ~new_n14052_;
  assign new_n14054_ = ~new_n12432_ & ~new_n14053_;
  assign new_n14055_ = ~new_n7478_ & ~new_n7486_;
  assign new_n14056_ = ~new_n7487_ & ~new_n14055_;
  assign new_n14057_ = ~new_n7464_ & new_n7478_;
  assign new_n14058_ = new_n7464_ & ~new_n7478_;
  assign new_n14059_ = ~new_n14057_ & ~new_n14058_;
  assign new_n14060_ = new_n14056_ & ~new_n14059_;
  assign new_n14061_ = ~new_n12439_ & ~new_n14060_;
  assign new_n14062_ = new_n14047_ & new_n14061_;
  assign new_n14063_ = ~new_n7524_ & ~new_n7532_;
  assign new_n14064_ = ~new_n7533_ & ~new_n14063_;
  assign new_n14065_ = ~new_n7510_ & new_n7524_;
  assign new_n14066_ = new_n7510_ & ~new_n7524_;
  assign new_n14067_ = ~new_n14065_ & ~new_n14066_;
  assign new_n14068_ = new_n14064_ & ~new_n14067_;
  assign new_n14069_ = ~new_n12447_ & ~new_n14068_;
  assign new_n14070_ = new_n14061_ & new_n14069_;
  assign new_n14071_ = ~new_n14062_ & ~new_n14070_;
  assign new_n14072_ = ~new_n14054_ & new_n14071_;
  assign new_n14073_ = new_n14054_ & ~new_n14071_;
  assign new_n14074_ = ~new_n14072_ & ~new_n14073_;
  assign A4102 = ~new_n14047_ & ~new_n14074_;
  assign new_n14076_ = new_n14044_ & ~new_n14072_;
  assign A4101 = ~new_n14047_ & ~new_n14076_;
  assign new_n14078_ = ~new_n14044_ & ~new_n14054_;
  assign new_n14079_ = ~new_n14047_ & ~new_n14078_;
  assign new_n14080_ = new_n14047_ & ~new_n14079_;
  assign new_n14081_ = new_n14047_ & new_n14078_;
  assign new_n14082_ = new_n14080_ & ~new_n14081_;
  assign new_n14083_ = ~new_n14054_ & ~new_n14082_;
  assign A4100 = new_n14071_ | new_n14083_;
  assign new_n14085_ = ~new_n14061_ & ~new_n14069_;
  assign new_n14086_ = ~new_n14070_ & ~new_n14085_;
  assign new_n14087_ = ~new_n14047_ & new_n14061_;
  assign new_n14088_ = new_n14047_ & ~new_n14061_;
  assign new_n14089_ = ~new_n14087_ & ~new_n14088_;
  assign new_n14090_ = new_n14086_ & ~new_n14089_;
  assign A4099 = new_n14083_ | new_n14090_;
  assign new_n14092_ = ~new_n14054_ & ~new_n14090_;
  assign new_n14093_ = new_n14054_ & new_n14090_;
  assign new_n14094_ = ~new_n14092_ & ~new_n14093_;
  assign A4098 = ~new_n14047_ & ~new_n14094_;
  assign new_n14096_ = ~new_n7595_ & ~new_n7603_;
  assign new_n14097_ = ~new_n7604_ & ~new_n14096_;
  assign new_n14098_ = ~new_n7581_ & new_n7595_;
  assign new_n14099_ = new_n7581_ & ~new_n7595_;
  assign new_n14100_ = ~new_n14098_ & ~new_n14099_;
  assign new_n14101_ = new_n14097_ & ~new_n14100_;
  assign new_n14102_ = ~new_n12480_ & ~new_n14101_;
  assign new_n14103_ = ~new_n7640_ & ~new_n7648_;
  assign new_n14104_ = ~new_n7649_ & ~new_n14103_;
  assign new_n14105_ = ~new_n7626_ & new_n7640_;
  assign new_n14106_ = new_n7626_ & ~new_n7640_;
  assign new_n14107_ = ~new_n14105_ & ~new_n14106_;
  assign new_n14108_ = new_n14104_ & ~new_n14107_;
  assign new_n14109_ = ~new_n12487_ & ~new_n14108_;
  assign new_n14110_ = new_n14102_ & ~new_n14109_;
  assign new_n14111_ = ~new_n14102_ & new_n14109_;
  assign new_n14112_ = ~new_n14110_ & ~new_n14111_;
  assign new_n14113_ = ~new_n7688_ & ~new_n7696_;
  assign new_n14114_ = ~new_n7697_ & ~new_n14113_;
  assign new_n14115_ = ~new_n7674_ & new_n7688_;
  assign new_n14116_ = new_n7674_ & ~new_n7688_;
  assign new_n14117_ = ~new_n14115_ & ~new_n14116_;
  assign new_n14118_ = new_n14114_ & ~new_n14117_;
  assign new_n14119_ = ~new_n12497_ & ~new_n14118_;
  assign new_n14120_ = ~new_n7733_ & ~new_n7741_;
  assign new_n14121_ = ~new_n7742_ & ~new_n14120_;
  assign new_n14122_ = ~new_n7719_ & new_n7733_;
  assign new_n14123_ = new_n7719_ & ~new_n7733_;
  assign new_n14124_ = ~new_n14122_ & ~new_n14123_;
  assign new_n14125_ = new_n14121_ & ~new_n14124_;
  assign new_n14126_ = ~new_n12504_ & ~new_n14125_;
  assign new_n14127_ = new_n14112_ & new_n14126_;
  assign new_n14128_ = ~new_n7779_ & ~new_n7787_;
  assign new_n14129_ = ~new_n7788_ & ~new_n14128_;
  assign new_n14130_ = ~new_n7765_ & new_n7779_;
  assign new_n14131_ = new_n7765_ & ~new_n7779_;
  assign new_n14132_ = ~new_n14130_ & ~new_n14131_;
  assign new_n14133_ = new_n14129_ & ~new_n14132_;
  assign new_n14134_ = ~new_n12512_ & ~new_n14133_;
  assign new_n14135_ = new_n14126_ & new_n14134_;
  assign new_n14136_ = ~new_n14127_ & ~new_n14135_;
  assign new_n14137_ = ~new_n14119_ & new_n14136_;
  assign new_n14138_ = new_n14119_ & ~new_n14136_;
  assign new_n14139_ = ~new_n14137_ & ~new_n14138_;
  assign A4069 = ~new_n14112_ & ~new_n14139_;
  assign new_n14141_ = new_n14109_ & ~new_n14137_;
  assign A4068 = ~new_n14112_ & ~new_n14141_;
  assign new_n14143_ = ~new_n14109_ & ~new_n14119_;
  assign new_n14144_ = ~new_n14112_ & ~new_n14143_;
  assign new_n14145_ = new_n14112_ & ~new_n14144_;
  assign new_n14146_ = new_n14112_ & new_n14143_;
  assign new_n14147_ = new_n14145_ & ~new_n14146_;
  assign new_n14148_ = ~new_n14119_ & ~new_n14147_;
  assign A4067 = new_n14136_ | new_n14148_;
  assign new_n14150_ = ~new_n14126_ & ~new_n14134_;
  assign new_n14151_ = ~new_n14135_ & ~new_n14150_;
  assign new_n14152_ = ~new_n14112_ & new_n14126_;
  assign new_n14153_ = new_n14112_ & ~new_n14126_;
  assign new_n14154_ = ~new_n14152_ & ~new_n14153_;
  assign new_n14155_ = new_n14151_ & ~new_n14154_;
  assign A4066 = new_n14148_ | new_n14155_;
  assign new_n14157_ = ~new_n14119_ & ~new_n14155_;
  assign new_n14158_ = new_n14119_ & new_n14155_;
  assign new_n14159_ = ~new_n14157_ & ~new_n14158_;
  assign A4065 = ~new_n14112_ & ~new_n14159_;
  assign new_n14161_ = ~new_n7850_ & ~new_n7858_;
  assign new_n14162_ = ~new_n7859_ & ~new_n14161_;
  assign new_n14163_ = ~new_n7836_ & new_n7850_;
  assign new_n14164_ = new_n7836_ & ~new_n7850_;
  assign new_n14165_ = ~new_n14163_ & ~new_n14164_;
  assign new_n14166_ = new_n14162_ & ~new_n14165_;
  assign new_n14167_ = ~new_n12545_ & ~new_n14166_;
  assign new_n14168_ = ~new_n7895_ & ~new_n7903_;
  assign new_n14169_ = ~new_n7904_ & ~new_n14168_;
  assign new_n14170_ = ~new_n7881_ & new_n7895_;
  assign new_n14171_ = new_n7881_ & ~new_n7895_;
  assign new_n14172_ = ~new_n14170_ & ~new_n14171_;
  assign new_n14173_ = new_n14169_ & ~new_n14172_;
  assign new_n14174_ = ~new_n12552_ & ~new_n14173_;
  assign new_n14175_ = new_n14167_ & ~new_n14174_;
  assign new_n14176_ = ~new_n14167_ & new_n14174_;
  assign new_n14177_ = ~new_n14175_ & ~new_n14176_;
  assign new_n14178_ = ~new_n7943_ & ~new_n7951_;
  assign new_n14179_ = ~new_n7952_ & ~new_n14178_;
  assign new_n14180_ = ~new_n7929_ & new_n7943_;
  assign new_n14181_ = new_n7929_ & ~new_n7943_;
  assign new_n14182_ = ~new_n14180_ & ~new_n14181_;
  assign new_n14183_ = new_n14179_ & ~new_n14182_;
  assign new_n14184_ = ~new_n12562_ & ~new_n14183_;
  assign new_n14185_ = ~new_n7988_ & ~new_n7996_;
  assign new_n14186_ = ~new_n7997_ & ~new_n14185_;
  assign new_n14187_ = ~new_n7974_ & new_n7988_;
  assign new_n14188_ = new_n7974_ & ~new_n7988_;
  assign new_n14189_ = ~new_n14187_ & ~new_n14188_;
  assign new_n14190_ = new_n14186_ & ~new_n14189_;
  assign new_n14191_ = ~new_n12569_ & ~new_n14190_;
  assign new_n14192_ = new_n14177_ & new_n14191_;
  assign new_n14193_ = ~new_n8034_ & ~new_n8042_;
  assign new_n14194_ = ~new_n8043_ & ~new_n14193_;
  assign new_n14195_ = ~new_n8020_ & new_n8034_;
  assign new_n14196_ = new_n8020_ & ~new_n8034_;
  assign new_n14197_ = ~new_n14195_ & ~new_n14196_;
  assign new_n14198_ = new_n14194_ & ~new_n14197_;
  assign new_n14199_ = ~new_n12577_ & ~new_n14198_;
  assign new_n14200_ = new_n14191_ & new_n14199_;
  assign new_n14201_ = ~new_n14192_ & ~new_n14200_;
  assign new_n14202_ = ~new_n14184_ & new_n14201_;
  assign new_n14203_ = new_n14184_ & ~new_n14201_;
  assign new_n14204_ = ~new_n14202_ & ~new_n14203_;
  assign A4036 = ~new_n14177_ & ~new_n14204_;
  assign new_n14206_ = new_n14174_ & ~new_n14202_;
  assign A4035 = ~new_n14177_ & ~new_n14206_;
  assign new_n14208_ = ~new_n14174_ & ~new_n14184_;
  assign new_n14209_ = ~new_n14177_ & ~new_n14208_;
  assign new_n14210_ = new_n14177_ & ~new_n14209_;
  assign new_n14211_ = new_n14177_ & new_n14208_;
  assign new_n14212_ = new_n14210_ & ~new_n14211_;
  assign new_n14213_ = ~new_n14184_ & ~new_n14212_;
  assign A4034 = new_n14201_ | new_n14213_;
  assign new_n14215_ = ~new_n14191_ & ~new_n14199_;
  assign new_n14216_ = ~new_n14200_ & ~new_n14215_;
  assign new_n14217_ = ~new_n14177_ & new_n14191_;
  assign new_n14218_ = new_n14177_ & ~new_n14191_;
  assign new_n14219_ = ~new_n14217_ & ~new_n14218_;
  assign new_n14220_ = new_n14216_ & ~new_n14219_;
  assign A4033 = new_n14213_ | new_n14220_;
  assign new_n14222_ = ~new_n14184_ & ~new_n14220_;
  assign new_n14223_ = new_n14184_ & new_n14220_;
  assign new_n14224_ = ~new_n14222_ & ~new_n14223_;
  assign A4032 = ~new_n14177_ & ~new_n14224_;
  assign new_n14226_ = ~new_n8105_ & ~new_n8113_;
  assign new_n14227_ = ~new_n8114_ & ~new_n14226_;
  assign new_n14228_ = ~new_n8091_ & new_n8105_;
  assign new_n14229_ = new_n8091_ & ~new_n8105_;
  assign new_n14230_ = ~new_n14228_ & ~new_n14229_;
  assign new_n14231_ = new_n14227_ & ~new_n14230_;
  assign new_n14232_ = ~new_n12610_ & ~new_n14231_;
  assign new_n14233_ = ~new_n8150_ & ~new_n8158_;
  assign new_n14234_ = ~new_n8159_ & ~new_n14233_;
  assign new_n14235_ = ~new_n8136_ & new_n8150_;
  assign new_n14236_ = new_n8136_ & ~new_n8150_;
  assign new_n14237_ = ~new_n14235_ & ~new_n14236_;
  assign new_n14238_ = new_n14234_ & ~new_n14237_;
  assign new_n14239_ = ~new_n12617_ & ~new_n14238_;
  assign new_n14240_ = new_n14232_ & ~new_n14239_;
  assign new_n14241_ = ~new_n14232_ & new_n14239_;
  assign new_n14242_ = ~new_n14240_ & ~new_n14241_;
  assign new_n14243_ = ~new_n8198_ & ~new_n8206_;
  assign new_n14244_ = ~new_n8207_ & ~new_n14243_;
  assign new_n14245_ = ~new_n8184_ & new_n8198_;
  assign new_n14246_ = new_n8184_ & ~new_n8198_;
  assign new_n14247_ = ~new_n14245_ & ~new_n14246_;
  assign new_n14248_ = new_n14244_ & ~new_n14247_;
  assign new_n14249_ = ~new_n12627_ & ~new_n14248_;
  assign new_n14250_ = ~new_n8243_ & ~new_n8251_;
  assign new_n14251_ = ~new_n8252_ & ~new_n14250_;
  assign new_n14252_ = ~new_n8229_ & new_n8243_;
  assign new_n14253_ = new_n8229_ & ~new_n8243_;
  assign new_n14254_ = ~new_n14252_ & ~new_n14253_;
  assign new_n14255_ = new_n14251_ & ~new_n14254_;
  assign new_n14256_ = ~new_n12634_ & ~new_n14255_;
  assign new_n14257_ = new_n14242_ & new_n14256_;
  assign new_n14258_ = ~new_n8289_ & ~new_n8297_;
  assign new_n14259_ = ~new_n8298_ & ~new_n14258_;
  assign new_n14260_ = ~new_n8275_ & new_n8289_;
  assign new_n14261_ = new_n8275_ & ~new_n8289_;
  assign new_n14262_ = ~new_n14260_ & ~new_n14261_;
  assign new_n14263_ = new_n14259_ & ~new_n14262_;
  assign new_n14264_ = ~new_n12642_ & ~new_n14263_;
  assign new_n14265_ = new_n14256_ & new_n14264_;
  assign new_n14266_ = ~new_n14257_ & ~new_n14265_;
  assign new_n14267_ = ~new_n14249_ & new_n14266_;
  assign new_n14268_ = new_n14249_ & ~new_n14266_;
  assign new_n14269_ = ~new_n14267_ & ~new_n14268_;
  assign A4003 = ~new_n14242_ & ~new_n14269_;
  assign new_n14271_ = new_n14239_ & ~new_n14267_;
  assign A4002 = ~new_n14242_ & ~new_n14271_;
  assign new_n14273_ = ~new_n14239_ & ~new_n14249_;
  assign new_n14274_ = ~new_n14242_ & ~new_n14273_;
  assign new_n14275_ = new_n14242_ & ~new_n14274_;
  assign new_n14276_ = new_n14242_ & new_n14273_;
  assign new_n14277_ = new_n14275_ & ~new_n14276_;
  assign new_n14278_ = ~new_n14249_ & ~new_n14277_;
  assign A4001 = new_n14266_ | new_n14278_;
  assign new_n14280_ = ~new_n14256_ & ~new_n14264_;
  assign new_n14281_ = ~new_n14265_ & ~new_n14280_;
  assign new_n14282_ = ~new_n14242_ & new_n14256_;
  assign new_n14283_ = new_n14242_ & ~new_n14256_;
  assign new_n14284_ = ~new_n14282_ & ~new_n14283_;
  assign new_n14285_ = new_n14281_ & ~new_n14284_;
  assign A4000 = new_n14278_ | new_n14285_;
  assign new_n14287_ = ~new_n14249_ & ~new_n14285_;
  assign new_n14288_ = new_n14249_ & new_n14285_;
  assign new_n14289_ = ~new_n14287_ & ~new_n14288_;
  assign A3999 = ~new_n14242_ & ~new_n14289_;
  assign new_n14291_ = ~new_n8356_ & ~new_n8364_;
  assign new_n14292_ = ~new_n8365_ & ~new_n14291_;
  assign new_n14293_ = ~new_n8342_ & new_n8356_;
  assign new_n14294_ = new_n8342_ & ~new_n8356_;
  assign new_n14295_ = ~new_n14293_ & ~new_n14294_;
  assign new_n14296_ = new_n14292_ & ~new_n14295_;
  assign new_n14297_ = ~new_n12675_ & ~new_n14296_;
  assign new_n14298_ = ~new_n8401_ & ~new_n8409_;
  assign new_n14299_ = ~new_n8410_ & ~new_n14298_;
  assign new_n14300_ = ~new_n8387_ & new_n8401_;
  assign new_n14301_ = new_n8387_ & ~new_n8401_;
  assign new_n14302_ = ~new_n14300_ & ~new_n14301_;
  assign new_n14303_ = new_n14299_ & ~new_n14302_;
  assign new_n14304_ = ~new_n12682_ & ~new_n14303_;
  assign new_n14305_ = new_n14297_ & ~new_n14304_;
  assign new_n14306_ = ~new_n14297_ & new_n14304_;
  assign new_n14307_ = ~new_n14305_ & ~new_n14306_;
  assign new_n14308_ = ~new_n8449_ & ~new_n8457_;
  assign new_n14309_ = ~new_n8458_ & ~new_n14308_;
  assign new_n14310_ = ~new_n8435_ & new_n8449_;
  assign new_n14311_ = new_n8435_ & ~new_n8449_;
  assign new_n14312_ = ~new_n14310_ & ~new_n14311_;
  assign new_n14313_ = new_n14309_ & ~new_n14312_;
  assign new_n14314_ = ~new_n12692_ & ~new_n14313_;
  assign new_n14315_ = ~new_n8494_ & ~new_n8502_;
  assign new_n14316_ = ~new_n8503_ & ~new_n14315_;
  assign new_n14317_ = ~new_n8480_ & new_n8494_;
  assign new_n14318_ = new_n8480_ & ~new_n8494_;
  assign new_n14319_ = ~new_n14317_ & ~new_n14318_;
  assign new_n14320_ = new_n14316_ & ~new_n14319_;
  assign new_n14321_ = ~new_n12699_ & ~new_n14320_;
  assign new_n14322_ = new_n14307_ & new_n14321_;
  assign new_n14323_ = ~new_n8540_ & ~new_n8548_;
  assign new_n14324_ = ~new_n8549_ & ~new_n14323_;
  assign new_n14325_ = ~new_n8526_ & new_n8540_;
  assign new_n14326_ = new_n8526_ & ~new_n8540_;
  assign new_n14327_ = ~new_n14325_ & ~new_n14326_;
  assign new_n14328_ = new_n14324_ & ~new_n14327_;
  assign new_n14329_ = ~new_n12707_ & ~new_n14328_;
  assign new_n14330_ = new_n14321_ & new_n14329_;
  assign new_n14331_ = ~new_n14322_ & ~new_n14330_;
  assign new_n14332_ = ~new_n14314_ & new_n14331_;
  assign new_n14333_ = new_n14314_ & ~new_n14331_;
  assign new_n14334_ = ~new_n14332_ & ~new_n14333_;
  assign A3970 = ~new_n14307_ & ~new_n14334_;
  assign new_n14336_ = new_n14304_ & ~new_n14332_;
  assign A3969 = ~new_n14307_ & ~new_n14336_;
  assign new_n14338_ = ~new_n14304_ & ~new_n14314_;
  assign new_n14339_ = ~new_n14307_ & ~new_n14338_;
  assign new_n14340_ = new_n14307_ & ~new_n14339_;
  assign new_n14341_ = new_n14307_ & new_n14338_;
  assign new_n14342_ = new_n14340_ & ~new_n14341_;
  assign new_n14343_ = ~new_n14314_ & ~new_n14342_;
  assign A3968 = new_n14331_ | new_n14343_;
  assign new_n14345_ = ~new_n14321_ & ~new_n14329_;
  assign new_n14346_ = ~new_n14330_ & ~new_n14345_;
  assign new_n14347_ = ~new_n14307_ & new_n14321_;
  assign new_n14348_ = new_n14307_ & ~new_n14321_;
  assign new_n14349_ = ~new_n14347_ & ~new_n14348_;
  assign new_n14350_ = new_n14346_ & ~new_n14349_;
  assign A3967 = new_n14343_ | new_n14350_;
  assign new_n14352_ = ~new_n14314_ & ~new_n14350_;
  assign new_n14353_ = new_n14314_ & new_n14350_;
  assign new_n14354_ = ~new_n14352_ & ~new_n14353_;
  assign A3966 = ~new_n14307_ & ~new_n14354_;
  assign new_n14356_ = ~new_n8611_ & ~new_n8619_;
  assign new_n14357_ = ~new_n8620_ & ~new_n14356_;
  assign new_n14358_ = ~new_n8597_ & new_n8611_;
  assign new_n14359_ = new_n8597_ & ~new_n8611_;
  assign new_n14360_ = ~new_n14358_ & ~new_n14359_;
  assign new_n14361_ = new_n14357_ & ~new_n14360_;
  assign new_n14362_ = ~new_n12740_ & ~new_n14361_;
  assign new_n14363_ = ~new_n8656_ & ~new_n8664_;
  assign new_n14364_ = ~new_n8665_ & ~new_n14363_;
  assign new_n14365_ = ~new_n8642_ & new_n8656_;
  assign new_n14366_ = new_n8642_ & ~new_n8656_;
  assign new_n14367_ = ~new_n14365_ & ~new_n14366_;
  assign new_n14368_ = new_n14364_ & ~new_n14367_;
  assign new_n14369_ = ~new_n12747_ & ~new_n14368_;
  assign new_n14370_ = new_n14362_ & ~new_n14369_;
  assign new_n14371_ = ~new_n14362_ & new_n14369_;
  assign new_n14372_ = ~new_n14370_ & ~new_n14371_;
  assign new_n14373_ = ~new_n8704_ & ~new_n8712_;
  assign new_n14374_ = ~new_n8713_ & ~new_n14373_;
  assign new_n14375_ = ~new_n8690_ & new_n8704_;
  assign new_n14376_ = new_n8690_ & ~new_n8704_;
  assign new_n14377_ = ~new_n14375_ & ~new_n14376_;
  assign new_n14378_ = new_n14374_ & ~new_n14377_;
  assign new_n14379_ = ~new_n12757_ & ~new_n14378_;
  assign new_n14380_ = ~new_n8749_ & ~new_n8757_;
  assign new_n14381_ = ~new_n8758_ & ~new_n14380_;
  assign new_n14382_ = ~new_n8735_ & new_n8749_;
  assign new_n14383_ = new_n8735_ & ~new_n8749_;
  assign new_n14384_ = ~new_n14382_ & ~new_n14383_;
  assign new_n14385_ = new_n14381_ & ~new_n14384_;
  assign new_n14386_ = ~new_n12764_ & ~new_n14385_;
  assign new_n14387_ = new_n14372_ & new_n14386_;
  assign new_n14388_ = ~new_n8795_ & ~new_n8803_;
  assign new_n14389_ = ~new_n8804_ & ~new_n14388_;
  assign new_n14390_ = ~new_n8781_ & new_n8795_;
  assign new_n14391_ = new_n8781_ & ~new_n8795_;
  assign new_n14392_ = ~new_n14390_ & ~new_n14391_;
  assign new_n14393_ = new_n14389_ & ~new_n14392_;
  assign new_n14394_ = ~new_n12772_ & ~new_n14393_;
  assign new_n14395_ = new_n14386_ & new_n14394_;
  assign new_n14396_ = ~new_n14387_ & ~new_n14395_;
  assign new_n14397_ = ~new_n14379_ & new_n14396_;
  assign new_n14398_ = new_n14379_ & ~new_n14396_;
  assign new_n14399_ = ~new_n14397_ & ~new_n14398_;
  assign A3937 = ~new_n14372_ & ~new_n14399_;
  assign new_n14401_ = new_n14369_ & ~new_n14397_;
  assign A3936 = ~new_n14372_ & ~new_n14401_;
  assign new_n14403_ = ~new_n14369_ & ~new_n14379_;
  assign new_n14404_ = ~new_n14372_ & ~new_n14403_;
  assign new_n14405_ = new_n14372_ & ~new_n14404_;
  assign new_n14406_ = new_n14372_ & new_n14403_;
  assign new_n14407_ = new_n14405_ & ~new_n14406_;
  assign new_n14408_ = ~new_n14379_ & ~new_n14407_;
  assign A3935 = new_n14396_ | new_n14408_;
  assign new_n14410_ = ~new_n14386_ & ~new_n14394_;
  assign new_n14411_ = ~new_n14395_ & ~new_n14410_;
  assign new_n14412_ = ~new_n14372_ & new_n14386_;
  assign new_n14413_ = new_n14372_ & ~new_n14386_;
  assign new_n14414_ = ~new_n14412_ & ~new_n14413_;
  assign new_n14415_ = new_n14411_ & ~new_n14414_;
  assign A3934 = new_n14408_ | new_n14415_;
  assign new_n14417_ = ~new_n14379_ & ~new_n14415_;
  assign new_n14418_ = new_n14379_ & new_n14415_;
  assign new_n14419_ = ~new_n14417_ & ~new_n14418_;
  assign A3933 = ~new_n14372_ & ~new_n14419_;
  assign new_n14421_ = ~new_n8866_ & ~new_n8874_;
  assign new_n14422_ = ~new_n8875_ & ~new_n14421_;
  assign new_n14423_ = ~new_n8852_ & new_n8866_;
  assign new_n14424_ = new_n8852_ & ~new_n8866_;
  assign new_n14425_ = ~new_n14423_ & ~new_n14424_;
  assign new_n14426_ = new_n14422_ & ~new_n14425_;
  assign new_n14427_ = ~new_n12805_ & ~new_n14426_;
  assign new_n14428_ = ~new_n8911_ & ~new_n8919_;
  assign new_n14429_ = ~new_n8920_ & ~new_n14428_;
  assign new_n14430_ = ~new_n8897_ & new_n8911_;
  assign new_n14431_ = new_n8897_ & ~new_n8911_;
  assign new_n14432_ = ~new_n14430_ & ~new_n14431_;
  assign new_n14433_ = new_n14429_ & ~new_n14432_;
  assign new_n14434_ = ~new_n12812_ & ~new_n14433_;
  assign new_n14435_ = new_n14427_ & ~new_n14434_;
  assign new_n14436_ = ~new_n14427_ & new_n14434_;
  assign new_n14437_ = ~new_n14435_ & ~new_n14436_;
  assign new_n14438_ = ~new_n8959_ & ~new_n8967_;
  assign new_n14439_ = ~new_n8968_ & ~new_n14438_;
  assign new_n14440_ = ~new_n8945_ & new_n8959_;
  assign new_n14441_ = new_n8945_ & ~new_n8959_;
  assign new_n14442_ = ~new_n14440_ & ~new_n14441_;
  assign new_n14443_ = new_n14439_ & ~new_n14442_;
  assign new_n14444_ = ~new_n12822_ & ~new_n14443_;
  assign new_n14445_ = ~new_n9004_ & ~new_n9012_;
  assign new_n14446_ = ~new_n9013_ & ~new_n14445_;
  assign new_n14447_ = ~new_n8990_ & new_n9004_;
  assign new_n14448_ = new_n8990_ & ~new_n9004_;
  assign new_n14449_ = ~new_n14447_ & ~new_n14448_;
  assign new_n14450_ = new_n14446_ & ~new_n14449_;
  assign new_n14451_ = ~new_n12829_ & ~new_n14450_;
  assign new_n14452_ = new_n14437_ & new_n14451_;
  assign new_n14453_ = ~new_n9050_ & ~new_n9058_;
  assign new_n14454_ = ~new_n9059_ & ~new_n14453_;
  assign new_n14455_ = ~new_n9036_ & new_n9050_;
  assign new_n14456_ = new_n9036_ & ~new_n9050_;
  assign new_n14457_ = ~new_n14455_ & ~new_n14456_;
  assign new_n14458_ = new_n14454_ & ~new_n14457_;
  assign new_n14459_ = ~new_n12837_ & ~new_n14458_;
  assign new_n14460_ = new_n14451_ & new_n14459_;
  assign new_n14461_ = ~new_n14452_ & ~new_n14460_;
  assign new_n14462_ = ~new_n14444_ & new_n14461_;
  assign new_n14463_ = new_n14444_ & ~new_n14461_;
  assign new_n14464_ = ~new_n14462_ & ~new_n14463_;
  assign A3904 = ~new_n14437_ & ~new_n14464_;
  assign new_n14466_ = new_n14434_ & ~new_n14462_;
  assign A3903 = ~new_n14437_ & ~new_n14466_;
  assign new_n14468_ = ~new_n14434_ & ~new_n14444_;
  assign new_n14469_ = ~new_n14437_ & ~new_n14468_;
  assign new_n14470_ = new_n14437_ & ~new_n14469_;
  assign new_n14471_ = new_n14437_ & new_n14468_;
  assign new_n14472_ = new_n14470_ & ~new_n14471_;
  assign new_n14473_ = ~new_n14444_ & ~new_n14472_;
  assign A3902 = new_n14461_ | new_n14473_;
  assign new_n14475_ = ~new_n14451_ & ~new_n14459_;
  assign new_n14476_ = ~new_n14460_ & ~new_n14475_;
  assign new_n14477_ = ~new_n14437_ & new_n14451_;
  assign new_n14478_ = new_n14437_ & ~new_n14451_;
  assign new_n14479_ = ~new_n14477_ & ~new_n14478_;
  assign new_n14480_ = new_n14476_ & ~new_n14479_;
  assign A3901 = new_n14473_ | new_n14480_;
  assign new_n14482_ = ~new_n14444_ & ~new_n14480_;
  assign new_n14483_ = new_n14444_ & new_n14480_;
  assign new_n14484_ = ~new_n14482_ & ~new_n14483_;
  assign A3900 = ~new_n14437_ & ~new_n14484_;
  assign new_n14486_ = ~new_n9121_ & ~new_n9129_;
  assign new_n14487_ = ~new_n9130_ & ~new_n14486_;
  assign new_n14488_ = ~new_n9107_ & new_n9121_;
  assign new_n14489_ = new_n9107_ & ~new_n9121_;
  assign new_n14490_ = ~new_n14488_ & ~new_n14489_;
  assign new_n14491_ = new_n14487_ & ~new_n14490_;
  assign new_n14492_ = ~new_n12870_ & ~new_n14491_;
  assign new_n14493_ = ~new_n9166_ & ~new_n9174_;
  assign new_n14494_ = ~new_n9175_ & ~new_n14493_;
  assign new_n14495_ = ~new_n9152_ & new_n9166_;
  assign new_n14496_ = new_n9152_ & ~new_n9166_;
  assign new_n14497_ = ~new_n14495_ & ~new_n14496_;
  assign new_n14498_ = new_n14494_ & ~new_n14497_;
  assign new_n14499_ = ~new_n12877_ & ~new_n14498_;
  assign new_n14500_ = new_n14492_ & ~new_n14499_;
  assign new_n14501_ = ~new_n14492_ & new_n14499_;
  assign new_n14502_ = ~new_n14500_ & ~new_n14501_;
  assign new_n14503_ = ~new_n9214_ & ~new_n9222_;
  assign new_n14504_ = ~new_n9223_ & ~new_n14503_;
  assign new_n14505_ = ~new_n9200_ & new_n9214_;
  assign new_n14506_ = new_n9200_ & ~new_n9214_;
  assign new_n14507_ = ~new_n14505_ & ~new_n14506_;
  assign new_n14508_ = new_n14504_ & ~new_n14507_;
  assign new_n14509_ = ~new_n12887_ & ~new_n14508_;
  assign new_n14510_ = ~new_n9259_ & ~new_n9267_;
  assign new_n14511_ = ~new_n9268_ & ~new_n14510_;
  assign new_n14512_ = ~new_n9245_ & new_n9259_;
  assign new_n14513_ = new_n9245_ & ~new_n9259_;
  assign new_n14514_ = ~new_n14512_ & ~new_n14513_;
  assign new_n14515_ = new_n14511_ & ~new_n14514_;
  assign new_n14516_ = ~new_n12894_ & ~new_n14515_;
  assign new_n14517_ = new_n14502_ & new_n14516_;
  assign new_n14518_ = ~new_n9305_ & ~new_n9313_;
  assign new_n14519_ = ~new_n9314_ & ~new_n14518_;
  assign new_n14520_ = ~new_n9291_ & new_n9305_;
  assign new_n14521_ = new_n9291_ & ~new_n9305_;
  assign new_n14522_ = ~new_n14520_ & ~new_n14521_;
  assign new_n14523_ = new_n14519_ & ~new_n14522_;
  assign new_n14524_ = ~new_n12902_ & ~new_n14523_;
  assign new_n14525_ = new_n14516_ & new_n14524_;
  assign new_n14526_ = ~new_n14517_ & ~new_n14525_;
  assign new_n14527_ = ~new_n14509_ & new_n14526_;
  assign new_n14528_ = new_n14509_ & ~new_n14526_;
  assign new_n14529_ = ~new_n14527_ & ~new_n14528_;
  assign A3871 = ~new_n14502_ & ~new_n14529_;
  assign new_n14531_ = new_n14499_ & ~new_n14527_;
  assign A3870 = ~new_n14502_ & ~new_n14531_;
  assign new_n14533_ = ~new_n14499_ & ~new_n14509_;
  assign new_n14534_ = ~new_n14502_ & ~new_n14533_;
  assign new_n14535_ = new_n14502_ & ~new_n14534_;
  assign new_n14536_ = new_n14502_ & new_n14533_;
  assign new_n14537_ = new_n14535_ & ~new_n14536_;
  assign new_n14538_ = ~new_n14509_ & ~new_n14537_;
  assign A3869 = new_n14526_ | new_n14538_;
  assign new_n14540_ = ~new_n14516_ & ~new_n14524_;
  assign new_n14541_ = ~new_n14525_ & ~new_n14540_;
  assign new_n14542_ = ~new_n14502_ & new_n14516_;
  assign new_n14543_ = new_n14502_ & ~new_n14516_;
  assign new_n14544_ = ~new_n14542_ & ~new_n14543_;
  assign new_n14545_ = new_n14541_ & ~new_n14544_;
  assign A3868 = new_n14538_ | new_n14545_;
  assign new_n14547_ = ~new_n14509_ & ~new_n14545_;
  assign new_n14548_ = new_n14509_ & new_n14545_;
  assign new_n14549_ = ~new_n14547_ & ~new_n14548_;
  assign A3867 = ~new_n14502_ & ~new_n14549_;
  assign new_n14551_ = ~new_n9376_ & ~new_n9384_;
  assign new_n14552_ = ~new_n9385_ & ~new_n14551_;
  assign new_n14553_ = ~new_n9362_ & new_n9376_;
  assign new_n14554_ = new_n9362_ & ~new_n9376_;
  assign new_n14555_ = ~new_n14553_ & ~new_n14554_;
  assign new_n14556_ = new_n14552_ & ~new_n14555_;
  assign new_n14557_ = ~new_n12935_ & ~new_n14556_;
  assign new_n14558_ = ~new_n9421_ & ~new_n9429_;
  assign new_n14559_ = ~new_n9430_ & ~new_n14558_;
  assign new_n14560_ = ~new_n9407_ & new_n9421_;
  assign new_n14561_ = new_n9407_ & ~new_n9421_;
  assign new_n14562_ = ~new_n14560_ & ~new_n14561_;
  assign new_n14563_ = new_n14559_ & ~new_n14562_;
  assign new_n14564_ = ~new_n12942_ & ~new_n14563_;
  assign new_n14565_ = new_n14557_ & ~new_n14564_;
  assign new_n14566_ = ~new_n14557_ & new_n14564_;
  assign new_n14567_ = ~new_n14565_ & ~new_n14566_;
  assign new_n14568_ = ~new_n9469_ & ~new_n9477_;
  assign new_n14569_ = ~new_n9478_ & ~new_n14568_;
  assign new_n14570_ = ~new_n9455_ & new_n9469_;
  assign new_n14571_ = new_n9455_ & ~new_n9469_;
  assign new_n14572_ = ~new_n14570_ & ~new_n14571_;
  assign new_n14573_ = new_n14569_ & ~new_n14572_;
  assign new_n14574_ = ~new_n12952_ & ~new_n14573_;
  assign new_n14575_ = ~new_n9514_ & ~new_n9522_;
  assign new_n14576_ = ~new_n9523_ & ~new_n14575_;
  assign new_n14577_ = ~new_n9500_ & new_n9514_;
  assign new_n14578_ = new_n9500_ & ~new_n9514_;
  assign new_n14579_ = ~new_n14577_ & ~new_n14578_;
  assign new_n14580_ = new_n14576_ & ~new_n14579_;
  assign new_n14581_ = ~new_n12959_ & ~new_n14580_;
  assign new_n14582_ = new_n14567_ & new_n14581_;
  assign new_n14583_ = ~new_n9560_ & ~new_n9568_;
  assign new_n14584_ = ~new_n9569_ & ~new_n14583_;
  assign new_n14585_ = ~new_n9546_ & new_n9560_;
  assign new_n14586_ = new_n9546_ & ~new_n9560_;
  assign new_n14587_ = ~new_n14585_ & ~new_n14586_;
  assign new_n14588_ = new_n14584_ & ~new_n14587_;
  assign new_n14589_ = ~new_n12967_ & ~new_n14588_;
  assign new_n14590_ = new_n14581_ & new_n14589_;
  assign new_n14591_ = ~new_n14582_ & ~new_n14590_;
  assign new_n14592_ = ~new_n14574_ & new_n14591_;
  assign new_n14593_ = new_n14574_ & ~new_n14591_;
  assign new_n14594_ = ~new_n14592_ & ~new_n14593_;
  assign A3838 = ~new_n14567_ & ~new_n14594_;
  assign new_n14596_ = new_n14564_ & ~new_n14592_;
  assign A3837 = ~new_n14567_ & ~new_n14596_;
  assign new_n14598_ = ~new_n14564_ & ~new_n14574_;
  assign new_n14599_ = ~new_n14567_ & ~new_n14598_;
  assign new_n14600_ = new_n14567_ & ~new_n14599_;
  assign new_n14601_ = new_n14567_ & new_n14598_;
  assign new_n14602_ = new_n14600_ & ~new_n14601_;
  assign new_n14603_ = ~new_n14574_ & ~new_n14602_;
  assign A3836 = new_n14591_ | new_n14603_;
  assign new_n14605_ = ~new_n14581_ & ~new_n14589_;
  assign new_n14606_ = ~new_n14590_ & ~new_n14605_;
  assign new_n14607_ = ~new_n14567_ & new_n14581_;
  assign new_n14608_ = new_n14567_ & ~new_n14581_;
  assign new_n14609_ = ~new_n14607_ & ~new_n14608_;
  assign new_n14610_ = new_n14606_ & ~new_n14609_;
  assign A3835 = new_n14603_ | new_n14610_;
  assign new_n14612_ = ~new_n14574_ & ~new_n14610_;
  assign new_n14613_ = new_n14574_ & new_n14610_;
  assign new_n14614_ = ~new_n14612_ & ~new_n14613_;
  assign A3834 = ~new_n14567_ & ~new_n14614_;
  assign new_n14616_ = ~new_n9627_ & ~new_n9635_;
  assign new_n14617_ = ~new_n9636_ & ~new_n14616_;
  assign new_n14618_ = ~new_n9613_ & new_n9627_;
  assign new_n14619_ = new_n9613_ & ~new_n9627_;
  assign new_n14620_ = ~new_n14618_ & ~new_n14619_;
  assign new_n14621_ = new_n14617_ & ~new_n14620_;
  assign new_n14622_ = ~new_n13000_ & ~new_n14621_;
  assign new_n14623_ = ~new_n9672_ & ~new_n9680_;
  assign new_n14624_ = ~new_n9681_ & ~new_n14623_;
  assign new_n14625_ = ~new_n9658_ & new_n9672_;
  assign new_n14626_ = new_n9658_ & ~new_n9672_;
  assign new_n14627_ = ~new_n14625_ & ~new_n14626_;
  assign new_n14628_ = new_n14624_ & ~new_n14627_;
  assign new_n14629_ = ~new_n13007_ & ~new_n14628_;
  assign new_n14630_ = new_n14622_ & ~new_n14629_;
  assign new_n14631_ = ~new_n14622_ & new_n14629_;
  assign new_n14632_ = ~new_n14630_ & ~new_n14631_;
  assign new_n14633_ = ~new_n9720_ & ~new_n9728_;
  assign new_n14634_ = ~new_n9729_ & ~new_n14633_;
  assign new_n14635_ = ~new_n9706_ & new_n9720_;
  assign new_n14636_ = new_n9706_ & ~new_n9720_;
  assign new_n14637_ = ~new_n14635_ & ~new_n14636_;
  assign new_n14638_ = new_n14634_ & ~new_n14637_;
  assign new_n14639_ = ~new_n13017_ & ~new_n14638_;
  assign new_n14640_ = ~new_n9765_ & ~new_n9773_;
  assign new_n14641_ = ~new_n9774_ & ~new_n14640_;
  assign new_n14642_ = ~new_n9751_ & new_n9765_;
  assign new_n14643_ = new_n9751_ & ~new_n9765_;
  assign new_n14644_ = ~new_n14642_ & ~new_n14643_;
  assign new_n14645_ = new_n14641_ & ~new_n14644_;
  assign new_n14646_ = ~new_n13024_ & ~new_n14645_;
  assign new_n14647_ = new_n14632_ & new_n14646_;
  assign new_n14648_ = ~new_n9811_ & ~new_n9819_;
  assign new_n14649_ = ~new_n9820_ & ~new_n14648_;
  assign new_n14650_ = ~new_n9797_ & new_n9811_;
  assign new_n14651_ = new_n9797_ & ~new_n9811_;
  assign new_n14652_ = ~new_n14650_ & ~new_n14651_;
  assign new_n14653_ = new_n14649_ & ~new_n14652_;
  assign new_n14654_ = ~new_n13032_ & ~new_n14653_;
  assign new_n14655_ = new_n14646_ & new_n14654_;
  assign new_n14656_ = ~new_n14647_ & ~new_n14655_;
  assign new_n14657_ = ~new_n14639_ & new_n14656_;
  assign new_n14658_ = new_n14639_ & ~new_n14656_;
  assign new_n14659_ = ~new_n14657_ & ~new_n14658_;
  assign A3805 = ~new_n14632_ & ~new_n14659_;
  assign new_n14661_ = new_n14629_ & ~new_n14657_;
  assign A3804 = ~new_n14632_ & ~new_n14661_;
  assign new_n14663_ = ~new_n14629_ & ~new_n14639_;
  assign new_n14664_ = ~new_n14632_ & ~new_n14663_;
  assign new_n14665_ = new_n14632_ & ~new_n14664_;
  assign new_n14666_ = new_n14632_ & new_n14663_;
  assign new_n14667_ = new_n14665_ & ~new_n14666_;
  assign new_n14668_ = ~new_n14639_ & ~new_n14667_;
  assign A3803 = new_n14656_ | new_n14668_;
  assign new_n14670_ = ~new_n14646_ & ~new_n14654_;
  assign new_n14671_ = ~new_n14655_ & ~new_n14670_;
  assign new_n14672_ = ~new_n14632_ & new_n14646_;
  assign new_n14673_ = new_n14632_ & ~new_n14646_;
  assign new_n14674_ = ~new_n14672_ & ~new_n14673_;
  assign new_n14675_ = new_n14671_ & ~new_n14674_;
  assign A3802 = new_n14668_ | new_n14675_;
  assign new_n14677_ = ~new_n14639_ & ~new_n14675_;
  assign new_n14678_ = new_n14639_ & new_n14675_;
  assign new_n14679_ = ~new_n14677_ & ~new_n14678_;
  assign A3801 = ~new_n14632_ & ~new_n14679_;
  assign new_n14681_ = new_n9870_ & new_n9875_;
  assign new_n14682_ = ~new_n9876_ & ~new_n14681_;
  assign new_n14683_ = ~new_n9862_ & ~new_n9870_;
  assign new_n14684_ = new_n9862_ & new_n9870_;
  assign new_n14685_ = ~new_n14683_ & ~new_n14684_;
  assign new_n14686_ = new_n14682_ & ~new_n14685_;
  assign new_n14687_ = ~new_n13065_ & ~new_n14686_;
  assign new_n14688_ = new_n9900_ & new_n9905_;
  assign new_n14689_ = ~new_n9906_ & ~new_n14688_;
  assign new_n14690_ = ~new_n9892_ & ~new_n9900_;
  assign new_n14691_ = new_n9892_ & new_n9900_;
  assign new_n14692_ = ~new_n14690_ & ~new_n14691_;
  assign new_n14693_ = new_n14689_ & ~new_n14692_;
  assign new_n14694_ = ~new_n13072_ & ~new_n14693_;
  assign new_n14695_ = new_n14687_ & ~new_n14694_;
  assign new_n14696_ = ~new_n14687_ & new_n14694_;
  assign new_n14697_ = ~new_n14695_ & ~new_n14696_;
  assign new_n14698_ = new_n9933_ & new_n9938_;
  assign new_n14699_ = ~new_n9939_ & ~new_n14698_;
  assign new_n14700_ = ~new_n9925_ & ~new_n9933_;
  assign new_n14701_ = new_n9925_ & new_n9933_;
  assign new_n14702_ = ~new_n14700_ & ~new_n14701_;
  assign new_n14703_ = new_n14699_ & ~new_n14702_;
  assign new_n14704_ = ~new_n13082_ & ~new_n14703_;
  assign new_n14705_ = new_n9963_ & new_n9968_;
  assign new_n14706_ = ~new_n9969_ & ~new_n14705_;
  assign new_n14707_ = ~new_n9955_ & ~new_n9963_;
  assign new_n14708_ = new_n9955_ & new_n9963_;
  assign new_n14709_ = ~new_n14707_ & ~new_n14708_;
  assign new_n14710_ = new_n14706_ & ~new_n14709_;
  assign new_n14711_ = ~new_n13089_ & ~new_n14710_;
  assign new_n14712_ = new_n14697_ & new_n14711_;
  assign new_n14713_ = new_n9994_ & new_n9999_;
  assign new_n14714_ = ~new_n10000_ & ~new_n14713_;
  assign new_n14715_ = ~new_n9986_ & ~new_n9994_;
  assign new_n14716_ = new_n9986_ & new_n9994_;
  assign new_n14717_ = ~new_n14715_ & ~new_n14716_;
  assign new_n14718_ = new_n14714_ & ~new_n14717_;
  assign new_n14719_ = ~new_n13097_ & ~new_n14718_;
  assign new_n14720_ = new_n14711_ & new_n14719_;
  assign new_n14721_ = ~new_n14712_ & ~new_n14720_;
  assign new_n14722_ = ~new_n14704_ & new_n14721_;
  assign new_n14723_ = new_n14704_ & ~new_n14721_;
  assign new_n14724_ = ~new_n14722_ & ~new_n14723_;
  assign A3772 = ~new_n14697_ & ~new_n14724_;
  assign new_n14726_ = new_n14694_ & ~new_n14722_;
  assign A3771 = ~new_n14697_ & ~new_n14726_;
  assign new_n14728_ = ~new_n14694_ & ~new_n14704_;
  assign new_n14729_ = ~new_n14697_ & ~new_n14728_;
  assign new_n14730_ = new_n14697_ & ~new_n14729_;
  assign new_n14731_ = new_n14697_ & new_n14728_;
  assign new_n14732_ = new_n14730_ & ~new_n14731_;
  assign new_n14733_ = ~new_n14704_ & ~new_n14732_;
  assign A3770 = new_n14721_ | new_n14733_;
  assign new_n14735_ = ~new_n14711_ & ~new_n14719_;
  assign new_n14736_ = ~new_n14720_ & ~new_n14735_;
  assign new_n14737_ = ~new_n14697_ & new_n14711_;
  assign new_n14738_ = new_n14697_ & ~new_n14711_;
  assign new_n14739_ = ~new_n14737_ & ~new_n14738_;
  assign new_n14740_ = new_n14736_ & ~new_n14739_;
  assign A3769 = new_n14733_ | new_n14740_;
  assign new_n14742_ = ~new_n14704_ & ~new_n14740_;
  assign new_n14743_ = new_n14704_ & new_n14740_;
  assign new_n14744_ = ~new_n14742_ & ~new_n14743_;
  assign A3768 = ~new_n14697_ & ~new_n14744_;
  assign new_n14746_ = new_n10050_ & new_n10055_;
  assign new_n14747_ = ~new_n10056_ & ~new_n14746_;
  assign new_n14748_ = ~new_n10042_ & ~new_n10050_;
  assign new_n14749_ = new_n10042_ & new_n10050_;
  assign new_n14750_ = ~new_n14748_ & ~new_n14749_;
  assign new_n14751_ = new_n14747_ & ~new_n14750_;
  assign new_n14752_ = ~new_n13130_ & ~new_n14751_;
  assign new_n14753_ = new_n10080_ & new_n10085_;
  assign new_n14754_ = ~new_n10086_ & ~new_n14753_;
  assign new_n14755_ = ~new_n10072_ & ~new_n10080_;
  assign new_n14756_ = new_n10072_ & new_n10080_;
  assign new_n14757_ = ~new_n14755_ & ~new_n14756_;
  assign new_n14758_ = new_n14754_ & ~new_n14757_;
  assign new_n14759_ = ~new_n13137_ & ~new_n14758_;
  assign new_n14760_ = new_n14752_ & ~new_n14759_;
  assign new_n14761_ = ~new_n14752_ & new_n14759_;
  assign new_n14762_ = ~new_n14760_ & ~new_n14761_;
  assign new_n14763_ = new_n10113_ & new_n10118_;
  assign new_n14764_ = ~new_n10119_ & ~new_n14763_;
  assign new_n14765_ = ~new_n10105_ & ~new_n10113_;
  assign new_n14766_ = new_n10105_ & new_n10113_;
  assign new_n14767_ = ~new_n14765_ & ~new_n14766_;
  assign new_n14768_ = new_n14764_ & ~new_n14767_;
  assign new_n14769_ = ~new_n13147_ & ~new_n14768_;
  assign new_n14770_ = new_n10143_ & new_n10148_;
  assign new_n14771_ = ~new_n10149_ & ~new_n14770_;
  assign new_n14772_ = ~new_n10135_ & ~new_n10143_;
  assign new_n14773_ = new_n10135_ & new_n10143_;
  assign new_n14774_ = ~new_n14772_ & ~new_n14773_;
  assign new_n14775_ = new_n14771_ & ~new_n14774_;
  assign new_n14776_ = ~new_n13154_ & ~new_n14775_;
  assign new_n14777_ = new_n14762_ & new_n14776_;
  assign new_n14778_ = new_n10174_ & new_n10179_;
  assign new_n14779_ = ~new_n10180_ & ~new_n14778_;
  assign new_n14780_ = ~new_n10166_ & ~new_n10174_;
  assign new_n14781_ = new_n10166_ & new_n10174_;
  assign new_n14782_ = ~new_n14780_ & ~new_n14781_;
  assign new_n14783_ = new_n14779_ & ~new_n14782_;
  assign new_n14784_ = ~new_n13162_ & ~new_n14783_;
  assign new_n14785_ = new_n14776_ & new_n14784_;
  assign new_n14786_ = ~new_n14777_ & ~new_n14785_;
  assign new_n14787_ = ~new_n14769_ & new_n14786_;
  assign new_n14788_ = new_n14769_ & ~new_n14786_;
  assign new_n14789_ = ~new_n14787_ & ~new_n14788_;
  assign A3739 = ~new_n14762_ & ~new_n14789_;
  assign new_n14791_ = new_n14759_ & ~new_n14787_;
  assign A3738 = ~new_n14762_ & ~new_n14791_;
  assign new_n14793_ = ~new_n14759_ & ~new_n14769_;
  assign new_n14794_ = ~new_n14762_ & ~new_n14793_;
  assign new_n14795_ = new_n14762_ & ~new_n14794_;
  assign new_n14796_ = new_n14762_ & new_n14793_;
  assign new_n14797_ = new_n14795_ & ~new_n14796_;
  assign new_n14798_ = ~new_n14769_ & ~new_n14797_;
  assign A3737 = new_n14786_ | new_n14798_;
  assign new_n14800_ = ~new_n14776_ & ~new_n14784_;
  assign new_n14801_ = ~new_n14785_ & ~new_n14800_;
  assign new_n14802_ = ~new_n14762_ & new_n14776_;
  assign new_n14803_ = new_n14762_ & ~new_n14776_;
  assign new_n14804_ = ~new_n14802_ & ~new_n14803_;
  assign new_n14805_ = new_n14801_ & ~new_n14804_;
  assign A3736 = new_n14798_ | new_n14805_;
  assign new_n14807_ = ~new_n14769_ & ~new_n14805_;
  assign new_n14808_ = new_n14769_ & new_n14805_;
  assign new_n14809_ = ~new_n14807_ & ~new_n14808_;
  assign A3735 = ~new_n14762_ & ~new_n14809_;
  assign new_n14811_ = new_n10230_ & new_n10235_;
  assign new_n14812_ = ~new_n10236_ & ~new_n14811_;
  assign new_n14813_ = ~new_n10222_ & ~new_n10230_;
  assign new_n14814_ = new_n10222_ & new_n10230_;
  assign new_n14815_ = ~new_n14813_ & ~new_n14814_;
  assign new_n14816_ = new_n14812_ & ~new_n14815_;
  assign new_n14817_ = ~new_n13195_ & ~new_n14816_;
  assign new_n14818_ = new_n10260_ & new_n10265_;
  assign new_n14819_ = ~new_n10266_ & ~new_n14818_;
  assign new_n14820_ = ~new_n10252_ & ~new_n10260_;
  assign new_n14821_ = new_n10252_ & new_n10260_;
  assign new_n14822_ = ~new_n14820_ & ~new_n14821_;
  assign new_n14823_ = new_n14819_ & ~new_n14822_;
  assign new_n14824_ = ~new_n13202_ & ~new_n14823_;
  assign new_n14825_ = new_n14817_ & ~new_n14824_;
  assign new_n14826_ = ~new_n14817_ & new_n14824_;
  assign new_n14827_ = ~new_n14825_ & ~new_n14826_;
  assign new_n14828_ = new_n10293_ & new_n10298_;
  assign new_n14829_ = ~new_n10299_ & ~new_n14828_;
  assign new_n14830_ = ~new_n10285_ & ~new_n10293_;
  assign new_n14831_ = new_n10285_ & new_n10293_;
  assign new_n14832_ = ~new_n14830_ & ~new_n14831_;
  assign new_n14833_ = new_n14829_ & ~new_n14832_;
  assign new_n14834_ = ~new_n13212_ & ~new_n14833_;
  assign new_n14835_ = new_n10323_ & new_n10328_;
  assign new_n14836_ = ~new_n10329_ & ~new_n14835_;
  assign new_n14837_ = ~new_n10315_ & ~new_n10323_;
  assign new_n14838_ = new_n10315_ & new_n10323_;
  assign new_n14839_ = ~new_n14837_ & ~new_n14838_;
  assign new_n14840_ = new_n14836_ & ~new_n14839_;
  assign new_n14841_ = ~new_n13219_ & ~new_n14840_;
  assign new_n14842_ = new_n14827_ & new_n14841_;
  assign new_n14843_ = new_n10354_ & new_n10359_;
  assign new_n14844_ = ~new_n10360_ & ~new_n14843_;
  assign new_n14845_ = ~new_n10346_ & ~new_n10354_;
  assign new_n14846_ = new_n10346_ & new_n10354_;
  assign new_n14847_ = ~new_n14845_ & ~new_n14846_;
  assign new_n14848_ = new_n14844_ & ~new_n14847_;
  assign new_n14849_ = ~new_n13227_ & ~new_n14848_;
  assign new_n14850_ = new_n14841_ & new_n14849_;
  assign new_n14851_ = ~new_n14842_ & ~new_n14850_;
  assign new_n14852_ = ~new_n14834_ & new_n14851_;
  assign new_n14853_ = new_n14834_ & ~new_n14851_;
  assign new_n14854_ = ~new_n14852_ & ~new_n14853_;
  assign A3706 = ~new_n14827_ & ~new_n14854_;
  assign new_n14856_ = new_n14824_ & ~new_n14852_;
  assign A3705 = ~new_n14827_ & ~new_n14856_;
  assign new_n14858_ = ~new_n14824_ & ~new_n14834_;
  assign new_n14859_ = ~new_n14827_ & ~new_n14858_;
  assign new_n14860_ = new_n14827_ & ~new_n14859_;
  assign new_n14861_ = new_n14827_ & new_n14858_;
  assign new_n14862_ = new_n14860_ & ~new_n14861_;
  assign new_n14863_ = ~new_n14834_ & ~new_n14862_;
  assign A3704 = new_n14851_ | new_n14863_;
  assign new_n14865_ = ~new_n14841_ & ~new_n14849_;
  assign new_n14866_ = ~new_n14850_ & ~new_n14865_;
  assign new_n14867_ = ~new_n14827_ & new_n14841_;
  assign new_n14868_ = new_n14827_ & ~new_n14841_;
  assign new_n14869_ = ~new_n14867_ & ~new_n14868_;
  assign new_n14870_ = new_n14866_ & ~new_n14869_;
  assign A3703 = new_n14863_ | new_n14870_;
  assign new_n14872_ = ~new_n14834_ & ~new_n14870_;
  assign new_n14873_ = new_n14834_ & new_n14870_;
  assign new_n14874_ = ~new_n14872_ & ~new_n14873_;
  assign A3702 = ~new_n14827_ & ~new_n14874_;
  assign new_n14876_ = new_n10410_ & new_n10415_;
  assign new_n14877_ = ~new_n10416_ & ~new_n14876_;
  assign new_n14878_ = ~new_n10402_ & ~new_n10410_;
  assign new_n14879_ = new_n10402_ & new_n10410_;
  assign new_n14880_ = ~new_n14878_ & ~new_n14879_;
  assign new_n14881_ = new_n14877_ & ~new_n14880_;
  assign new_n14882_ = ~new_n13260_ & ~new_n14881_;
  assign new_n14883_ = new_n10440_ & new_n10445_;
  assign new_n14884_ = ~new_n10446_ & ~new_n14883_;
  assign new_n14885_ = ~new_n10432_ & ~new_n10440_;
  assign new_n14886_ = new_n10432_ & new_n10440_;
  assign new_n14887_ = ~new_n14885_ & ~new_n14886_;
  assign new_n14888_ = new_n14884_ & ~new_n14887_;
  assign new_n14889_ = ~new_n13267_ & ~new_n14888_;
  assign new_n14890_ = new_n14882_ & ~new_n14889_;
  assign new_n14891_ = ~new_n14882_ & new_n14889_;
  assign new_n14892_ = ~new_n14890_ & ~new_n14891_;
  assign new_n14893_ = new_n10473_ & new_n10478_;
  assign new_n14894_ = ~new_n10479_ & ~new_n14893_;
  assign new_n14895_ = ~new_n10465_ & ~new_n10473_;
  assign new_n14896_ = new_n10465_ & new_n10473_;
  assign new_n14897_ = ~new_n14895_ & ~new_n14896_;
  assign new_n14898_ = new_n14894_ & ~new_n14897_;
  assign new_n14899_ = ~new_n13277_ & ~new_n14898_;
  assign new_n14900_ = new_n10503_ & new_n10508_;
  assign new_n14901_ = ~new_n10509_ & ~new_n14900_;
  assign new_n14902_ = ~new_n10495_ & ~new_n10503_;
  assign new_n14903_ = new_n10495_ & new_n10503_;
  assign new_n14904_ = ~new_n14902_ & ~new_n14903_;
  assign new_n14905_ = new_n14901_ & ~new_n14904_;
  assign new_n14906_ = ~new_n13284_ & ~new_n14905_;
  assign new_n14907_ = new_n14892_ & new_n14906_;
  assign new_n14908_ = new_n10534_ & new_n10539_;
  assign new_n14909_ = ~new_n10540_ & ~new_n14908_;
  assign new_n14910_ = ~new_n10526_ & ~new_n10534_;
  assign new_n14911_ = new_n10526_ & new_n10534_;
  assign new_n14912_ = ~new_n14910_ & ~new_n14911_;
  assign new_n14913_ = new_n14909_ & ~new_n14912_;
  assign new_n14914_ = ~new_n13292_ & ~new_n14913_;
  assign new_n14915_ = new_n14906_ & new_n14914_;
  assign new_n14916_ = ~new_n14907_ & ~new_n14915_;
  assign new_n14917_ = ~new_n14899_ & new_n14916_;
  assign new_n14918_ = new_n14899_ & ~new_n14916_;
  assign new_n14919_ = ~new_n14917_ & ~new_n14918_;
  assign A3673 = ~new_n14892_ & ~new_n14919_;
  assign new_n14921_ = new_n14889_ & ~new_n14917_;
  assign A3672 = ~new_n14892_ & ~new_n14921_;
  assign new_n14923_ = ~new_n14889_ & ~new_n14899_;
  assign new_n14924_ = ~new_n14892_ & ~new_n14923_;
  assign new_n14925_ = new_n14892_ & ~new_n14924_;
  assign new_n14926_ = new_n14892_ & new_n14923_;
  assign new_n14927_ = new_n14925_ & ~new_n14926_;
  assign new_n14928_ = ~new_n14899_ & ~new_n14927_;
  assign A3671 = new_n14916_ | new_n14928_;
  assign new_n14930_ = ~new_n14906_ & ~new_n14914_;
  assign new_n14931_ = ~new_n14915_ & ~new_n14930_;
  assign new_n14932_ = ~new_n14892_ & new_n14906_;
  assign new_n14933_ = new_n14892_ & ~new_n14906_;
  assign new_n14934_ = ~new_n14932_ & ~new_n14933_;
  assign new_n14935_ = new_n14931_ & ~new_n14934_;
  assign A3670 = new_n14928_ | new_n14935_;
  assign new_n14937_ = ~new_n14899_ & ~new_n14935_;
  assign new_n14938_ = new_n14899_ & new_n14935_;
  assign new_n14939_ = ~new_n14937_ & ~new_n14938_;
  assign A3669 = ~new_n14892_ & ~new_n14939_;
  assign new_n14941_ = new_n10600_ & new_n13321_;
  assign new_n14942_ = ~new_n10589_ & ~new_n14941_;
  assign new_n14943_ = ~new_n10592_ & ~new_n14942_;
  assign new_n14944_ = new_n10623_ & new_n10628_;
  assign new_n14945_ = ~new_n10629_ & ~new_n14944_;
  assign new_n14946_ = ~new_n10615_ & ~new_n10623_;
  assign new_n14947_ = new_n10615_ & new_n10623_;
  assign new_n14948_ = ~new_n14946_ & ~new_n14947_;
  assign new_n14949_ = new_n14945_ & ~new_n14948_;
  assign new_n14950_ = ~new_n13328_ & ~new_n14949_;
  assign new_n14951_ = ~new_n14943_ & ~new_n14950_;
  assign new_n14952_ = new_n14943_ & new_n14950_;
  assign new_n14953_ = ~new_n14951_ & ~new_n14952_;
  assign new_n14954_ = new_n10656_ & new_n10661_;
  assign new_n14955_ = ~new_n10662_ & ~new_n14954_;
  assign new_n14956_ = ~new_n10648_ & ~new_n10656_;
  assign new_n14957_ = new_n10648_ & new_n10656_;
  assign new_n14958_ = ~new_n14956_ & ~new_n14957_;
  assign new_n14959_ = new_n14955_ & ~new_n14958_;
  assign new_n14960_ = ~new_n13338_ & ~new_n14959_;
  assign new_n14961_ = new_n10686_ & new_n10691_;
  assign new_n14962_ = ~new_n10692_ & ~new_n14961_;
  assign new_n14963_ = ~new_n10678_ & ~new_n10686_;
  assign new_n14964_ = new_n10678_ & new_n10686_;
  assign new_n14965_ = ~new_n14963_ & ~new_n14964_;
  assign new_n14966_ = new_n14962_ & ~new_n14965_;
  assign new_n14967_ = ~new_n13345_ & ~new_n14966_;
  assign new_n14968_ = new_n14953_ & new_n14967_;
  assign new_n14969_ = new_n10717_ & new_n10722_;
  assign new_n14970_ = ~new_n10723_ & ~new_n14969_;
  assign new_n14971_ = ~new_n10709_ & ~new_n10717_;
  assign new_n14972_ = new_n10709_ & new_n10717_;
  assign new_n14973_ = ~new_n14971_ & ~new_n14972_;
  assign new_n14974_ = new_n14970_ & ~new_n14973_;
  assign new_n14975_ = ~new_n13353_ & ~new_n14974_;
  assign new_n14976_ = new_n14967_ & new_n14975_;
  assign new_n14977_ = ~new_n14968_ & ~new_n14976_;
  assign new_n14978_ = ~new_n14960_ & new_n14977_;
  assign new_n14979_ = new_n14960_ & ~new_n14977_;
  assign new_n14980_ = ~new_n14978_ & ~new_n14979_;
  assign A3640 = ~new_n14953_ & ~new_n14980_;
  assign new_n14982_ = new_n14950_ & ~new_n14978_;
  assign A3639 = ~new_n14953_ & ~new_n14982_;
  assign new_n14984_ = ~new_n14950_ & ~new_n14960_;
  assign new_n14985_ = ~new_n14953_ & ~new_n14984_;
  assign new_n14986_ = new_n14953_ & ~new_n14985_;
  assign new_n14987_ = new_n14953_ & new_n14984_;
  assign new_n14988_ = new_n14986_ & ~new_n14987_;
  assign new_n14989_ = ~new_n14960_ & ~new_n14988_;
  assign A3638 = new_n14977_ | new_n14989_;
  assign new_n14991_ = ~new_n14967_ & ~new_n14975_;
  assign new_n14992_ = ~new_n14976_ & ~new_n14991_;
  assign new_n14993_ = ~new_n14953_ & new_n14967_;
  assign new_n14994_ = new_n14953_ & ~new_n14967_;
  assign new_n14995_ = ~new_n14993_ & ~new_n14994_;
  assign new_n14996_ = new_n14992_ & ~new_n14995_;
  assign A3637 = new_n14989_ | new_n14996_;
  assign new_n14998_ = ~new_n14960_ & ~new_n14996_;
  assign new_n14999_ = new_n14960_ & new_n14996_;
  assign new_n15000_ = ~new_n14998_ & ~new_n14999_;
  assign A3636 = ~new_n14953_ & ~new_n15000_;
  assign new_n15002_ = new_n1437_ & ~new_n13386_;
  assign new_n15003_ = ~new_n1437_ & new_n13386_;
  assign new_n15004_ = ~new_n15002_ & ~new_n15003_;
  assign new_n15005_ = ~new_n1377_ & ~new_n15004_;
  assign new_n15006_ = new_n1747_ & ~new_n13393_;
  assign new_n15007_ = ~new_n1747_ & new_n13393_;
  assign new_n15008_ = ~new_n15006_ & ~new_n15007_;
  assign new_n15009_ = ~new_n1687_ & ~new_n15008_;
  assign new_n15010_ = ~new_n15005_ & new_n15009_;
  assign new_n15011_ = new_n15005_ & ~new_n15009_;
  assign new_n15012_ = ~new_n15010_ & ~new_n15011_;
  assign new_n15013_ = new_n2060_ & ~new_n13403_;
  assign new_n15014_ = ~new_n2060_ & new_n13403_;
  assign new_n15015_ = ~new_n15013_ & ~new_n15014_;
  assign new_n15016_ = ~new_n2000_ & ~new_n15015_;
  assign new_n15017_ = new_n2370_ & ~new_n13410_;
  assign new_n15018_ = ~new_n2370_ & new_n13410_;
  assign new_n15019_ = ~new_n15017_ & ~new_n15018_;
  assign new_n15020_ = ~new_n2310_ & ~new_n15019_;
  assign new_n15021_ = new_n15012_ & ~new_n15020_;
  assign new_n15022_ = new_n2681_ & ~new_n13418_;
  assign new_n15023_ = ~new_n2681_ & new_n13418_;
  assign new_n15024_ = ~new_n15022_ & ~new_n15023_;
  assign new_n15025_ = ~new_n2621_ & ~new_n15024_;
  assign new_n15026_ = ~new_n15020_ & ~new_n15025_;
  assign new_n15027_ = ~new_n15021_ & ~new_n15026_;
  assign new_n15028_ = new_n15016_ & new_n15027_;
  assign new_n15029_ = ~new_n15016_ & ~new_n15027_;
  assign new_n15030_ = ~new_n15028_ & ~new_n15029_;
  assign A3607 = ~new_n15012_ & ~new_n15030_;
  assign new_n15032_ = ~new_n15009_ & ~new_n15028_;
  assign A3606 = ~new_n15012_ & ~new_n15032_;
  assign new_n15034_ = new_n15009_ & new_n15016_;
  assign new_n15035_ = ~new_n15012_ & ~new_n15034_;
  assign new_n15036_ = new_n15012_ & ~new_n15035_;
  assign new_n15037_ = new_n15012_ & new_n15034_;
  assign new_n15038_ = new_n15036_ & ~new_n15037_;
  assign new_n15039_ = new_n15016_ & ~new_n15038_;
  assign A3605 = new_n15027_ | new_n15039_;
  assign new_n15041_ = new_n15020_ & new_n15025_;
  assign new_n15042_ = ~new_n15026_ & ~new_n15041_;
  assign new_n15043_ = ~new_n15012_ & ~new_n15020_;
  assign new_n15044_ = new_n15012_ & new_n15020_;
  assign new_n15045_ = ~new_n15043_ & ~new_n15044_;
  assign new_n15046_ = new_n15042_ & ~new_n15045_;
  assign A3604 = new_n15039_ | new_n15046_;
  assign new_n15048_ = new_n15016_ & ~new_n15046_;
  assign new_n15049_ = ~new_n15016_ & new_n15046_;
  assign new_n15050_ = ~new_n15048_ & ~new_n15049_;
  assign A3603 = ~new_n15012_ & ~new_n15050_;
  assign new_n15052_ = new_n2902_ & ~new_n13451_;
  assign new_n15053_ = ~new_n2902_ & new_n13451_;
  assign new_n15054_ = ~new_n15052_ & ~new_n15053_;
  assign new_n15055_ = ~new_n2882_ & ~new_n15054_;
  assign new_n15056_ = new_n3012_ & ~new_n13458_;
  assign new_n15057_ = ~new_n3012_ & new_n13458_;
  assign new_n15058_ = ~new_n15056_ & ~new_n15057_;
  assign new_n15059_ = ~new_n2992_ & ~new_n15058_;
  assign new_n15060_ = ~new_n15055_ & new_n15059_;
  assign new_n15061_ = new_n15055_ & ~new_n15059_;
  assign new_n15062_ = ~new_n15060_ & ~new_n15061_;
  assign new_n15063_ = new_n3125_ & ~new_n13468_;
  assign new_n15064_ = ~new_n3125_ & new_n13468_;
  assign new_n15065_ = ~new_n15063_ & ~new_n15064_;
  assign new_n15066_ = ~new_n3105_ & ~new_n15065_;
  assign new_n15067_ = new_n3235_ & ~new_n13475_;
  assign new_n15068_ = ~new_n3235_ & new_n13475_;
  assign new_n15069_ = ~new_n15067_ & ~new_n15068_;
  assign new_n15070_ = ~new_n3215_ & ~new_n15069_;
  assign new_n15071_ = new_n15062_ & ~new_n15070_;
  assign new_n15072_ = new_n3346_ & ~new_n13483_;
  assign new_n15073_ = ~new_n3346_ & new_n13483_;
  assign new_n15074_ = ~new_n15072_ & ~new_n15073_;
  assign new_n15075_ = ~new_n3326_ & ~new_n15074_;
  assign new_n15076_ = ~new_n15070_ & ~new_n15075_;
  assign new_n15077_ = ~new_n15071_ & ~new_n15076_;
  assign new_n15078_ = new_n15066_ & new_n15077_;
  assign new_n15079_ = ~new_n15066_ & ~new_n15077_;
  assign new_n15080_ = ~new_n15078_ & ~new_n15079_;
  assign A3574 = ~new_n15062_ & ~new_n15080_;
  assign new_n15082_ = ~new_n15059_ & ~new_n15078_;
  assign A3573 = ~new_n15062_ & ~new_n15082_;
  assign new_n15084_ = new_n15059_ & new_n15066_;
  assign new_n15085_ = ~new_n15062_ & ~new_n15084_;
  assign new_n15086_ = new_n15062_ & ~new_n15085_;
  assign new_n15087_ = new_n15062_ & new_n15084_;
  assign new_n15088_ = new_n15086_ & ~new_n15087_;
  assign new_n15089_ = new_n15066_ & ~new_n15088_;
  assign A3572 = new_n15077_ | new_n15089_;
  assign new_n15091_ = new_n15070_ & new_n15075_;
  assign new_n15092_ = ~new_n15076_ & ~new_n15091_;
  assign new_n15093_ = ~new_n15062_ & ~new_n15070_;
  assign new_n15094_ = new_n15062_ & new_n15070_;
  assign new_n15095_ = ~new_n15093_ & ~new_n15094_;
  assign new_n15096_ = new_n15092_ & ~new_n15095_;
  assign A3571 = new_n15089_ | new_n15096_;
  assign new_n15098_ = new_n15066_ & ~new_n15096_;
  assign new_n15099_ = ~new_n15066_ & new_n15096_;
  assign new_n15100_ = ~new_n15098_ & ~new_n15099_;
  assign A3570 = ~new_n15062_ & ~new_n15100_;
  assign new_n15102_ = new_n3553_ & ~new_n13516_;
  assign new_n15103_ = ~new_n3553_ & new_n13516_;
  assign new_n15104_ = ~new_n15102_ & ~new_n15103_;
  assign new_n15105_ = ~new_n3508_ & ~new_n15104_;
  assign new_n15106_ = new_n3788_ & ~new_n13523_;
  assign new_n15107_ = ~new_n3788_ & new_n13523_;
  assign new_n15108_ = ~new_n15106_ & ~new_n15107_;
  assign new_n15109_ = ~new_n3743_ & ~new_n15108_;
  assign new_n15110_ = ~new_n15105_ & new_n15109_;
  assign new_n15111_ = new_n15105_ & ~new_n15109_;
  assign new_n15112_ = ~new_n15110_ & ~new_n15111_;
  assign new_n15113_ = new_n4026_ & ~new_n13533_;
  assign new_n15114_ = ~new_n4026_ & new_n13533_;
  assign new_n15115_ = ~new_n15113_ & ~new_n15114_;
  assign new_n15116_ = ~new_n3981_ & ~new_n15115_;
  assign new_n15117_ = new_n4261_ & ~new_n13540_;
  assign new_n15118_ = ~new_n4261_ & new_n13540_;
  assign new_n15119_ = ~new_n15117_ & ~new_n15118_;
  assign new_n15120_ = ~new_n4216_ & ~new_n15119_;
  assign new_n15121_ = new_n15112_ & ~new_n15120_;
  assign new_n15122_ = new_n4497_ & ~new_n13548_;
  assign new_n15123_ = ~new_n4497_ & new_n13548_;
  assign new_n15124_ = ~new_n15122_ & ~new_n15123_;
  assign new_n15125_ = ~new_n4452_ & ~new_n15124_;
  assign new_n15126_ = ~new_n15120_ & ~new_n15125_;
  assign new_n15127_ = ~new_n15121_ & ~new_n15126_;
  assign new_n15128_ = new_n15116_ & new_n15127_;
  assign new_n15129_ = ~new_n15116_ & ~new_n15127_;
  assign new_n15130_ = ~new_n15128_ & ~new_n15129_;
  assign A3541 = ~new_n15112_ & ~new_n15130_;
  assign new_n15132_ = ~new_n15109_ & ~new_n15128_;
  assign A3540 = ~new_n15112_ & ~new_n15132_;
  assign new_n15134_ = new_n15109_ & new_n15116_;
  assign new_n15135_ = ~new_n15112_ & ~new_n15134_;
  assign new_n15136_ = new_n15112_ & ~new_n15135_;
  assign new_n15137_ = new_n15112_ & new_n15134_;
  assign new_n15138_ = new_n15136_ & ~new_n15137_;
  assign new_n15139_ = new_n15116_ & ~new_n15138_;
  assign A3539 = new_n15127_ | new_n15139_;
  assign new_n15141_ = new_n15120_ & new_n15125_;
  assign new_n15142_ = ~new_n15126_ & ~new_n15141_;
  assign new_n15143_ = ~new_n15112_ & ~new_n15120_;
  assign new_n15144_ = new_n15112_ & new_n15120_;
  assign new_n15145_ = ~new_n15143_ & ~new_n15144_;
  assign new_n15146_ = new_n15142_ & ~new_n15145_;
  assign A3538 = new_n15139_ | new_n15146_;
  assign new_n15148_ = new_n15116_ & ~new_n15146_;
  assign new_n15149_ = ~new_n15116_ & new_n15146_;
  assign new_n15150_ = ~new_n15148_ & ~new_n15149_;
  assign A3537 = ~new_n15112_ & ~new_n15150_;
  assign new_n15152_ = new_n4754_ & ~new_n13581_;
  assign new_n15153_ = ~new_n4754_ & new_n13581_;
  assign new_n15154_ = ~new_n15152_ & ~new_n15153_;
  assign new_n15155_ = ~new_n4709_ & ~new_n15154_;
  assign new_n15156_ = new_n4989_ & ~new_n13588_;
  assign new_n15157_ = ~new_n4989_ & new_n13588_;
  assign new_n15158_ = ~new_n15156_ & ~new_n15157_;
  assign new_n15159_ = ~new_n4944_ & ~new_n15158_;
  assign new_n15160_ = ~new_n15155_ & new_n15159_;
  assign new_n15161_ = new_n15155_ & ~new_n15159_;
  assign new_n15162_ = ~new_n15160_ & ~new_n15161_;
  assign new_n15163_ = new_n5227_ & ~new_n13598_;
  assign new_n15164_ = ~new_n5227_ & new_n13598_;
  assign new_n15165_ = ~new_n15163_ & ~new_n15164_;
  assign new_n15166_ = ~new_n5182_ & ~new_n15165_;
  assign new_n15167_ = new_n5462_ & ~new_n13605_;
  assign new_n15168_ = ~new_n5462_ & new_n13605_;
  assign new_n15169_ = ~new_n15167_ & ~new_n15168_;
  assign new_n15170_ = ~new_n5417_ & ~new_n15169_;
  assign new_n15171_ = new_n15162_ & ~new_n15170_;
  assign new_n15172_ = new_n5698_ & ~new_n13613_;
  assign new_n15173_ = ~new_n5698_ & new_n13613_;
  assign new_n15174_ = ~new_n15172_ & ~new_n15173_;
  assign new_n15175_ = ~new_n5653_ & ~new_n15174_;
  assign new_n15176_ = ~new_n15170_ & ~new_n15175_;
  assign new_n15177_ = ~new_n15171_ & ~new_n15176_;
  assign new_n15178_ = new_n15166_ & new_n15177_;
  assign new_n15179_ = ~new_n15166_ & ~new_n15177_;
  assign new_n15180_ = ~new_n15178_ & ~new_n15179_;
  assign A3508 = ~new_n15162_ & ~new_n15180_;
  assign new_n15182_ = ~new_n15159_ & ~new_n15178_;
  assign A3507 = ~new_n15162_ & ~new_n15182_;
  assign new_n15184_ = new_n15159_ & new_n15166_;
  assign new_n15185_ = ~new_n15162_ & ~new_n15184_;
  assign new_n15186_ = new_n15162_ & ~new_n15185_;
  assign new_n15187_ = new_n15162_ & new_n15184_;
  assign new_n15188_ = new_n15186_ & ~new_n15187_;
  assign new_n15189_ = new_n15166_ & ~new_n15188_;
  assign A3506 = new_n15177_ | new_n15189_;
  assign new_n15191_ = new_n15170_ & new_n15175_;
  assign new_n15192_ = ~new_n15176_ & ~new_n15191_;
  assign new_n15193_ = ~new_n15162_ & ~new_n15170_;
  assign new_n15194_ = new_n15162_ & new_n15170_;
  assign new_n15195_ = ~new_n15193_ & ~new_n15194_;
  assign new_n15196_ = new_n15192_ & ~new_n15195_;
  assign A3505 = new_n15189_ | new_n15196_;
  assign new_n15198_ = new_n15166_ & ~new_n15196_;
  assign new_n15199_ = ~new_n15166_ & new_n15196_;
  assign new_n15200_ = ~new_n15198_ & ~new_n15199_;
  assign A3504 = ~new_n15162_ & ~new_n15200_;
  assign new_n15202_ = new_n5917_ & ~new_n13646_;
  assign new_n15203_ = ~new_n5917_ & new_n13646_;
  assign new_n15204_ = ~new_n15202_ & ~new_n15203_;
  assign new_n15205_ = ~new_n5887_ & ~new_n15204_;
  assign new_n15206_ = new_n6077_ & ~new_n13653_;
  assign new_n15207_ = ~new_n6077_ & new_n13653_;
  assign new_n15208_ = ~new_n15206_ & ~new_n15207_;
  assign new_n15209_ = ~new_n6047_ & ~new_n15208_;
  assign new_n15210_ = ~new_n15205_ & new_n15209_;
  assign new_n15211_ = new_n15205_ & ~new_n15209_;
  assign new_n15212_ = ~new_n15210_ & ~new_n15211_;
  assign new_n15213_ = new_n6240_ & ~new_n13663_;
  assign new_n15214_ = ~new_n6240_ & new_n13663_;
  assign new_n15215_ = ~new_n15213_ & ~new_n15214_;
  assign new_n15216_ = ~new_n6210_ & ~new_n15215_;
  assign new_n15217_ = new_n6400_ & ~new_n13670_;
  assign new_n15218_ = ~new_n6400_ & new_n13670_;
  assign new_n15219_ = ~new_n15217_ & ~new_n15218_;
  assign new_n15220_ = ~new_n6370_ & ~new_n15219_;
  assign new_n15221_ = new_n15212_ & ~new_n15220_;
  assign new_n15222_ = new_n6561_ & ~new_n13678_;
  assign new_n15223_ = ~new_n6561_ & new_n13678_;
  assign new_n15224_ = ~new_n15222_ & ~new_n15223_;
  assign new_n15225_ = ~new_n6531_ & ~new_n15224_;
  assign new_n15226_ = ~new_n15220_ & ~new_n15225_;
  assign new_n15227_ = ~new_n15221_ & ~new_n15226_;
  assign new_n15228_ = new_n15216_ & new_n15227_;
  assign new_n15229_ = ~new_n15216_ & ~new_n15227_;
  assign new_n15230_ = ~new_n15228_ & ~new_n15229_;
  assign A3475 = ~new_n15212_ & ~new_n15230_;
  assign new_n15232_ = ~new_n15209_ & ~new_n15228_;
  assign A3474 = ~new_n15212_ & ~new_n15232_;
  assign new_n15234_ = new_n15209_ & new_n15216_;
  assign new_n15235_ = ~new_n15212_ & ~new_n15234_;
  assign new_n15236_ = new_n15212_ & ~new_n15235_;
  assign new_n15237_ = new_n15212_ & new_n15234_;
  assign new_n15238_ = new_n15236_ & ~new_n15237_;
  assign new_n15239_ = new_n15216_ & ~new_n15238_;
  assign A3473 = new_n15227_ | new_n15239_;
  assign new_n15241_ = new_n15220_ & new_n15225_;
  assign new_n15242_ = ~new_n15226_ & ~new_n15241_;
  assign new_n15243_ = ~new_n15212_ & ~new_n15220_;
  assign new_n15244_ = new_n15212_ & new_n15220_;
  assign new_n15245_ = ~new_n15243_ & ~new_n15244_;
  assign new_n15246_ = new_n15242_ & ~new_n15245_;
  assign A3472 = new_n15239_ | new_n15246_;
  assign new_n15248_ = new_n15216_ & ~new_n15246_;
  assign new_n15249_ = ~new_n15216_ & new_n15246_;
  assign new_n15250_ = ~new_n15248_ & ~new_n15249_;
  assign A3471 = ~new_n15212_ & ~new_n15250_;
  assign new_n15252_ = new_n6663_ & ~new_n13711_;
  assign new_n15253_ = ~new_n6663_ & new_n13711_;
  assign new_n15254_ = ~new_n15252_ & ~new_n15253_;
  assign new_n15255_ = ~new_n6661_ & ~new_n15254_;
  assign new_n15256_ = new_n6683_ & ~new_n13718_;
  assign new_n15257_ = ~new_n6683_ & new_n13718_;
  assign new_n15258_ = ~new_n15256_ & ~new_n15257_;
  assign new_n15259_ = ~new_n6681_ & ~new_n15258_;
  assign new_n15260_ = ~new_n15255_ & new_n15259_;
  assign new_n15261_ = new_n15255_ & ~new_n15259_;
  assign new_n15262_ = ~new_n15260_ & ~new_n15261_;
  assign new_n15263_ = new_n6706_ & ~new_n13728_;
  assign new_n15264_ = ~new_n6706_ & new_n13728_;
  assign new_n15265_ = ~new_n15263_ & ~new_n15264_;
  assign new_n15266_ = ~new_n6704_ & ~new_n15265_;
  assign new_n15267_ = new_n6726_ & ~new_n13735_;
  assign new_n15268_ = ~new_n6726_ & new_n13735_;
  assign new_n15269_ = ~new_n15267_ & ~new_n15268_;
  assign new_n15270_ = ~new_n6724_ & ~new_n15269_;
  assign new_n15271_ = new_n15262_ & ~new_n15270_;
  assign new_n15272_ = new_n6747_ & ~new_n13743_;
  assign new_n15273_ = ~new_n6747_ & new_n13743_;
  assign new_n15274_ = ~new_n15272_ & ~new_n15273_;
  assign new_n15275_ = ~new_n6745_ & ~new_n15274_;
  assign new_n15276_ = ~new_n15270_ & ~new_n15275_;
  assign new_n15277_ = ~new_n15271_ & ~new_n15276_;
  assign new_n15278_ = new_n15266_ & new_n15277_;
  assign new_n15279_ = ~new_n15266_ & ~new_n15277_;
  assign new_n15280_ = ~new_n15278_ & ~new_n15279_;
  assign A3442 = ~new_n15262_ & ~new_n15280_;
  assign new_n15282_ = ~new_n15259_ & ~new_n15278_;
  assign A3441 = ~new_n15262_ & ~new_n15282_;
  assign new_n15284_ = new_n15259_ & new_n15266_;
  assign new_n15285_ = ~new_n15262_ & ~new_n15284_;
  assign new_n15286_ = new_n15262_ & ~new_n15285_;
  assign new_n15287_ = new_n15262_ & new_n15284_;
  assign new_n15288_ = new_n15286_ & ~new_n15287_;
  assign new_n15289_ = new_n15266_ & ~new_n15288_;
  assign A3440 = new_n15277_ | new_n15289_;
  assign new_n15291_ = new_n15270_ & new_n15275_;
  assign new_n15292_ = ~new_n15276_ & ~new_n15291_;
  assign new_n15293_ = ~new_n15262_ & ~new_n15270_;
  assign new_n15294_ = new_n15262_ & new_n15270_;
  assign new_n15295_ = ~new_n15293_ & ~new_n15294_;
  assign new_n15296_ = new_n15292_ & ~new_n15295_;
  assign A3439 = new_n15289_ | new_n15296_;
  assign new_n15298_ = new_n15266_ & ~new_n15296_;
  assign new_n15299_ = ~new_n15266_ & new_n15296_;
  assign new_n15300_ = ~new_n15298_ & ~new_n15299_;
  assign A3438 = ~new_n15262_ & ~new_n15300_;
  assign new_n15302_ = new_n6793_ & ~new_n13776_;
  assign new_n15303_ = ~new_n6793_ & new_n13776_;
  assign new_n15304_ = ~new_n15302_ & ~new_n15303_;
  assign new_n15305_ = ~new_n6791_ & ~new_n15304_;
  assign new_n15306_ = new_n6813_ & ~new_n13783_;
  assign new_n15307_ = ~new_n6813_ & new_n13783_;
  assign new_n15308_ = ~new_n15306_ & ~new_n15307_;
  assign new_n15309_ = ~new_n6811_ & ~new_n15308_;
  assign new_n15310_ = ~new_n15305_ & new_n15309_;
  assign new_n15311_ = new_n15305_ & ~new_n15309_;
  assign new_n15312_ = ~new_n15310_ & ~new_n15311_;
  assign new_n15313_ = new_n6836_ & ~new_n13793_;
  assign new_n15314_ = ~new_n6836_ & new_n13793_;
  assign new_n15315_ = ~new_n15313_ & ~new_n15314_;
  assign new_n15316_ = ~new_n6834_ & ~new_n15315_;
  assign new_n15317_ = new_n6856_ & ~new_n13800_;
  assign new_n15318_ = ~new_n6856_ & new_n13800_;
  assign new_n15319_ = ~new_n15317_ & ~new_n15318_;
  assign new_n15320_ = ~new_n6854_ & ~new_n15319_;
  assign new_n15321_ = new_n15312_ & ~new_n15320_;
  assign new_n15322_ = new_n6877_ & ~new_n13808_;
  assign new_n15323_ = ~new_n6877_ & new_n13808_;
  assign new_n15324_ = ~new_n15322_ & ~new_n15323_;
  assign new_n15325_ = ~new_n6875_ & ~new_n15324_;
  assign new_n15326_ = ~new_n15320_ & ~new_n15325_;
  assign new_n15327_ = ~new_n15321_ & ~new_n15326_;
  assign new_n15328_ = new_n15316_ & new_n15327_;
  assign new_n15329_ = ~new_n15316_ & ~new_n15327_;
  assign new_n15330_ = ~new_n15328_ & ~new_n15329_;
  assign A3409 = ~new_n15312_ & ~new_n15330_;
  assign new_n15332_ = ~new_n15309_ & ~new_n15328_;
  assign A3408 = ~new_n15312_ & ~new_n15332_;
  assign new_n15334_ = new_n15309_ & new_n15316_;
  assign new_n15335_ = ~new_n15312_ & ~new_n15334_;
  assign new_n15336_ = new_n15312_ & ~new_n15335_;
  assign new_n15337_ = new_n15312_ & new_n15334_;
  assign new_n15338_ = new_n15336_ & ~new_n15337_;
  assign new_n15339_ = new_n15316_ & ~new_n15338_;
  assign A3407 = new_n15327_ | new_n15339_;
  assign new_n15341_ = new_n15320_ & new_n15325_;
  assign new_n15342_ = ~new_n15326_ & ~new_n15341_;
  assign new_n15343_ = ~new_n15312_ & ~new_n15320_;
  assign new_n15344_ = new_n15312_ & new_n15320_;
  assign new_n15345_ = ~new_n15343_ & ~new_n15344_;
  assign new_n15346_ = new_n15342_ & ~new_n15345_;
  assign A3406 = new_n15339_ | new_n15346_;
  assign new_n15348_ = new_n15316_ & ~new_n15346_;
  assign new_n15349_ = ~new_n15316_ & new_n15346_;
  assign new_n15350_ = ~new_n15348_ & ~new_n15349_;
  assign A3405 = ~new_n15312_ & ~new_n15350_;
  assign new_n15352_ = new_n6923_ & ~new_n13841_;
  assign new_n15353_ = ~new_n6923_ & new_n13841_;
  assign new_n15354_ = ~new_n15352_ & ~new_n15353_;
  assign new_n15355_ = ~new_n6921_ & ~new_n15354_;
  assign new_n15356_ = new_n6943_ & ~new_n13848_;
  assign new_n15357_ = ~new_n6943_ & new_n13848_;
  assign new_n15358_ = ~new_n15356_ & ~new_n15357_;
  assign new_n15359_ = ~new_n6941_ & ~new_n15358_;
  assign new_n15360_ = ~new_n15355_ & new_n15359_;
  assign new_n15361_ = new_n15355_ & ~new_n15359_;
  assign new_n15362_ = ~new_n15360_ & ~new_n15361_;
  assign new_n15363_ = new_n6966_ & ~new_n13858_;
  assign new_n15364_ = ~new_n6966_ & new_n13858_;
  assign new_n15365_ = ~new_n15363_ & ~new_n15364_;
  assign new_n15366_ = ~new_n6964_ & ~new_n15365_;
  assign new_n15367_ = new_n6986_ & ~new_n13865_;
  assign new_n15368_ = ~new_n6986_ & new_n13865_;
  assign new_n15369_ = ~new_n15367_ & ~new_n15368_;
  assign new_n15370_ = ~new_n6984_ & ~new_n15369_;
  assign new_n15371_ = new_n15362_ & ~new_n15370_;
  assign new_n15372_ = new_n7007_ & ~new_n13873_;
  assign new_n15373_ = ~new_n7007_ & new_n13873_;
  assign new_n15374_ = ~new_n15372_ & ~new_n15373_;
  assign new_n15375_ = ~new_n7005_ & ~new_n15374_;
  assign new_n15376_ = ~new_n15370_ & ~new_n15375_;
  assign new_n15377_ = ~new_n15371_ & ~new_n15376_;
  assign new_n15378_ = new_n15366_ & new_n15377_;
  assign new_n15379_ = ~new_n15366_ & ~new_n15377_;
  assign new_n15380_ = ~new_n15378_ & ~new_n15379_;
  assign A3376 = ~new_n15362_ & ~new_n15380_;
  assign new_n15382_ = ~new_n15359_ & ~new_n15378_;
  assign A3375 = ~new_n15362_ & ~new_n15382_;
  assign new_n15384_ = new_n15359_ & new_n15366_;
  assign new_n15385_ = ~new_n15362_ & ~new_n15384_;
  assign new_n15386_ = new_n15362_ & ~new_n15385_;
  assign new_n15387_ = new_n15362_ & new_n15384_;
  assign new_n15388_ = new_n15386_ & ~new_n15387_;
  assign new_n15389_ = new_n15366_ & ~new_n15388_;
  assign A3374 = new_n15377_ | new_n15389_;
  assign new_n15391_ = new_n15370_ & new_n15375_;
  assign new_n15392_ = ~new_n15376_ & ~new_n15391_;
  assign new_n15393_ = ~new_n15362_ & ~new_n15370_;
  assign new_n15394_ = new_n15362_ & new_n15370_;
  assign new_n15395_ = ~new_n15393_ & ~new_n15394_;
  assign new_n15396_ = new_n15392_ & ~new_n15395_;
  assign A3373 = new_n15389_ | new_n15396_;
  assign new_n15398_ = new_n15366_ & ~new_n15396_;
  assign new_n15399_ = ~new_n15366_ & new_n15396_;
  assign new_n15400_ = ~new_n15398_ & ~new_n15399_;
  assign A3372 = ~new_n15362_ & ~new_n15400_;
  assign new_n15402_ = new_n7053_ & ~new_n13906_;
  assign new_n15403_ = ~new_n7053_ & new_n13906_;
  assign new_n15404_ = ~new_n15402_ & ~new_n15403_;
  assign new_n15405_ = ~new_n7051_ & ~new_n15404_;
  assign new_n15406_ = new_n7073_ & ~new_n13913_;
  assign new_n15407_ = ~new_n7073_ & new_n13913_;
  assign new_n15408_ = ~new_n15406_ & ~new_n15407_;
  assign new_n15409_ = ~new_n7071_ & ~new_n15408_;
  assign new_n15410_ = ~new_n15405_ & new_n15409_;
  assign new_n15411_ = new_n15405_ & ~new_n15409_;
  assign new_n15412_ = ~new_n15410_ & ~new_n15411_;
  assign new_n15413_ = new_n7096_ & ~new_n13923_;
  assign new_n15414_ = ~new_n7096_ & new_n13923_;
  assign new_n15415_ = ~new_n15413_ & ~new_n15414_;
  assign new_n15416_ = ~new_n7094_ & ~new_n15415_;
  assign new_n15417_ = new_n7116_ & ~new_n13930_;
  assign new_n15418_ = ~new_n7116_ & new_n13930_;
  assign new_n15419_ = ~new_n15417_ & ~new_n15418_;
  assign new_n15420_ = ~new_n7114_ & ~new_n15419_;
  assign new_n15421_ = new_n15412_ & ~new_n15420_;
  assign new_n15422_ = new_n7137_ & ~new_n13938_;
  assign new_n15423_ = ~new_n7137_ & new_n13938_;
  assign new_n15424_ = ~new_n15422_ & ~new_n15423_;
  assign new_n15425_ = ~new_n7135_ & ~new_n15424_;
  assign new_n15426_ = ~new_n15420_ & ~new_n15425_;
  assign new_n15427_ = ~new_n15421_ & ~new_n15426_;
  assign new_n15428_ = new_n15416_ & new_n15427_;
  assign new_n15429_ = ~new_n15416_ & ~new_n15427_;
  assign new_n15430_ = ~new_n15428_ & ~new_n15429_;
  assign A3343 = ~new_n15412_ & ~new_n15430_;
  assign new_n15432_ = ~new_n15409_ & ~new_n15428_;
  assign A3342 = ~new_n15412_ & ~new_n15432_;
  assign new_n15434_ = new_n15409_ & new_n15416_;
  assign new_n15435_ = ~new_n15412_ & ~new_n15434_;
  assign new_n15436_ = new_n15412_ & ~new_n15435_;
  assign new_n15437_ = new_n15412_ & new_n15434_;
  assign new_n15438_ = new_n15436_ & ~new_n15437_;
  assign new_n15439_ = new_n15416_ & ~new_n15438_;
  assign A3341 = new_n15427_ | new_n15439_;
  assign new_n15441_ = new_n15420_ & new_n15425_;
  assign new_n15442_ = ~new_n15426_ & ~new_n15441_;
  assign new_n15443_ = ~new_n15412_ & ~new_n15420_;
  assign new_n15444_ = new_n15412_ & new_n15420_;
  assign new_n15445_ = ~new_n15443_ & ~new_n15444_;
  assign new_n15446_ = new_n15442_ & ~new_n15445_;
  assign A3340 = new_n15439_ | new_n15446_;
  assign new_n15448_ = new_n15416_ & ~new_n15446_;
  assign new_n15449_ = ~new_n15416_ & new_n15446_;
  assign new_n15450_ = ~new_n15448_ & ~new_n15449_;
  assign A3339 = ~new_n15412_ & ~new_n15450_;
  assign new_n15452_ = new_n7188_ & ~new_n13971_;
  assign new_n15453_ = ~new_n7188_ & new_n13971_;
  assign new_n15454_ = ~new_n15452_ & ~new_n15453_;
  assign new_n15455_ = ~new_n7186_ & ~new_n15454_;
  assign new_n15456_ = new_n7208_ & ~new_n13978_;
  assign new_n15457_ = ~new_n7208_ & new_n13978_;
  assign new_n15458_ = ~new_n15456_ & ~new_n15457_;
  assign new_n15459_ = ~new_n7206_ & ~new_n15458_;
  assign new_n15460_ = ~new_n15455_ & new_n15459_;
  assign new_n15461_ = new_n15455_ & ~new_n15459_;
  assign new_n15462_ = ~new_n15460_ & ~new_n15461_;
  assign new_n15463_ = new_n7231_ & ~new_n13988_;
  assign new_n15464_ = ~new_n7231_ & new_n13988_;
  assign new_n15465_ = ~new_n15463_ & ~new_n15464_;
  assign new_n15466_ = ~new_n7229_ & ~new_n15465_;
  assign new_n15467_ = new_n7251_ & ~new_n13995_;
  assign new_n15468_ = ~new_n7251_ & new_n13995_;
  assign new_n15469_ = ~new_n15467_ & ~new_n15468_;
  assign new_n15470_ = ~new_n7249_ & ~new_n15469_;
  assign new_n15471_ = new_n15462_ & ~new_n15470_;
  assign new_n15472_ = new_n7272_ & ~new_n14003_;
  assign new_n15473_ = ~new_n7272_ & new_n14003_;
  assign new_n15474_ = ~new_n15472_ & ~new_n15473_;
  assign new_n15475_ = ~new_n7270_ & ~new_n15474_;
  assign new_n15476_ = ~new_n15470_ & ~new_n15475_;
  assign new_n15477_ = ~new_n15471_ & ~new_n15476_;
  assign new_n15478_ = new_n15466_ & new_n15477_;
  assign new_n15479_ = ~new_n15466_ & ~new_n15477_;
  assign new_n15480_ = ~new_n15478_ & ~new_n15479_;
  assign A3310 = ~new_n15462_ & ~new_n15480_;
  assign new_n15482_ = ~new_n15459_ & ~new_n15478_;
  assign A3309 = ~new_n15462_ & ~new_n15482_;
  assign new_n15484_ = new_n15459_ & new_n15466_;
  assign new_n15485_ = ~new_n15462_ & ~new_n15484_;
  assign new_n15486_ = new_n15462_ & ~new_n15485_;
  assign new_n15487_ = new_n15462_ & new_n15484_;
  assign new_n15488_ = new_n15486_ & ~new_n15487_;
  assign new_n15489_ = new_n15466_ & ~new_n15488_;
  assign A3308 = new_n15477_ | new_n15489_;
  assign new_n15491_ = new_n15470_ & new_n15475_;
  assign new_n15492_ = ~new_n15476_ & ~new_n15491_;
  assign new_n15493_ = ~new_n15462_ & ~new_n15470_;
  assign new_n15494_ = new_n15462_ & new_n15470_;
  assign new_n15495_ = ~new_n15493_ & ~new_n15494_;
  assign new_n15496_ = new_n15492_ & ~new_n15495_;
  assign A3307 = new_n15489_ | new_n15496_;
  assign new_n15498_ = new_n15466_ & ~new_n15496_;
  assign new_n15499_ = ~new_n15466_ & new_n15496_;
  assign new_n15500_ = ~new_n15498_ & ~new_n15499_;
  assign A3306 = ~new_n15462_ & ~new_n15500_;
  assign new_n15502_ = ~new_n7333_ & ~new_n14036_;
  assign new_n15503_ = new_n7333_ & new_n14036_;
  assign new_n15504_ = ~new_n15502_ & ~new_n15503_;
  assign new_n15505_ = ~new_n7326_ & ~new_n15504_;
  assign new_n15506_ = ~new_n7378_ & ~new_n14043_;
  assign new_n15507_ = new_n7378_ & new_n14043_;
  assign new_n15508_ = ~new_n15506_ & ~new_n15507_;
  assign new_n15509_ = ~new_n7371_ & ~new_n15508_;
  assign new_n15510_ = ~new_n15505_ & new_n15509_;
  assign new_n15511_ = new_n15505_ & ~new_n15509_;
  assign new_n15512_ = ~new_n15510_ & ~new_n15511_;
  assign new_n15513_ = ~new_n7426_ & ~new_n14053_;
  assign new_n15514_ = new_n7426_ & new_n14053_;
  assign new_n15515_ = ~new_n15513_ & ~new_n15514_;
  assign new_n15516_ = ~new_n7419_ & ~new_n15515_;
  assign new_n15517_ = ~new_n7471_ & ~new_n14060_;
  assign new_n15518_ = new_n7471_ & new_n14060_;
  assign new_n15519_ = ~new_n15517_ & ~new_n15518_;
  assign new_n15520_ = ~new_n7464_ & ~new_n15519_;
  assign new_n15521_ = new_n15512_ & ~new_n15520_;
  assign new_n15522_ = ~new_n7517_ & ~new_n14068_;
  assign new_n15523_ = new_n7517_ & new_n14068_;
  assign new_n15524_ = ~new_n15522_ & ~new_n15523_;
  assign new_n15525_ = ~new_n7510_ & ~new_n15524_;
  assign new_n15526_ = ~new_n15520_ & ~new_n15525_;
  assign new_n15527_ = ~new_n15521_ & ~new_n15526_;
  assign new_n15528_ = new_n15516_ & new_n15527_;
  assign new_n15529_ = ~new_n15516_ & ~new_n15527_;
  assign new_n15530_ = ~new_n15528_ & ~new_n15529_;
  assign A3277 = ~new_n15512_ & ~new_n15530_;
  assign new_n15532_ = ~new_n15509_ & ~new_n15528_;
  assign A3276 = ~new_n15512_ & ~new_n15532_;
  assign new_n15534_ = new_n15509_ & new_n15516_;
  assign new_n15535_ = ~new_n15512_ & ~new_n15534_;
  assign new_n15536_ = new_n15512_ & ~new_n15535_;
  assign new_n15537_ = new_n15512_ & new_n15534_;
  assign new_n15538_ = new_n15536_ & ~new_n15537_;
  assign new_n15539_ = new_n15516_ & ~new_n15538_;
  assign A3275 = new_n15527_ | new_n15539_;
  assign new_n15541_ = new_n15520_ & new_n15525_;
  assign new_n15542_ = ~new_n15526_ & ~new_n15541_;
  assign new_n15543_ = ~new_n15512_ & ~new_n15520_;
  assign new_n15544_ = new_n15512_ & new_n15520_;
  assign new_n15545_ = ~new_n15543_ & ~new_n15544_;
  assign new_n15546_ = new_n15542_ & ~new_n15545_;
  assign A3274 = new_n15539_ | new_n15546_;
  assign new_n15548_ = new_n15516_ & ~new_n15546_;
  assign new_n15549_ = ~new_n15516_ & new_n15546_;
  assign new_n15550_ = ~new_n15548_ & ~new_n15549_;
  assign A3273 = ~new_n15512_ & ~new_n15550_;
  assign new_n15552_ = ~new_n7588_ & ~new_n14101_;
  assign new_n15553_ = new_n7588_ & new_n14101_;
  assign new_n15554_ = ~new_n15552_ & ~new_n15553_;
  assign new_n15555_ = ~new_n7581_ & ~new_n15554_;
  assign new_n15556_ = ~new_n7633_ & ~new_n14108_;
  assign new_n15557_ = new_n7633_ & new_n14108_;
  assign new_n15558_ = ~new_n15556_ & ~new_n15557_;
  assign new_n15559_ = ~new_n7626_ & ~new_n15558_;
  assign new_n15560_ = ~new_n15555_ & new_n15559_;
  assign new_n15561_ = new_n15555_ & ~new_n15559_;
  assign new_n15562_ = ~new_n15560_ & ~new_n15561_;
  assign new_n15563_ = ~new_n7681_ & ~new_n14118_;
  assign new_n15564_ = new_n7681_ & new_n14118_;
  assign new_n15565_ = ~new_n15563_ & ~new_n15564_;
  assign new_n15566_ = ~new_n7674_ & ~new_n15565_;
  assign new_n15567_ = ~new_n7726_ & ~new_n14125_;
  assign new_n15568_ = new_n7726_ & new_n14125_;
  assign new_n15569_ = ~new_n15567_ & ~new_n15568_;
  assign new_n15570_ = ~new_n7719_ & ~new_n15569_;
  assign new_n15571_ = new_n15562_ & ~new_n15570_;
  assign new_n15572_ = ~new_n7772_ & ~new_n14133_;
  assign new_n15573_ = new_n7772_ & new_n14133_;
  assign new_n15574_ = ~new_n15572_ & ~new_n15573_;
  assign new_n15575_ = ~new_n7765_ & ~new_n15574_;
  assign new_n15576_ = ~new_n15570_ & ~new_n15575_;
  assign new_n15577_ = ~new_n15571_ & ~new_n15576_;
  assign new_n15578_ = new_n15566_ & new_n15577_;
  assign new_n15579_ = ~new_n15566_ & ~new_n15577_;
  assign new_n15580_ = ~new_n15578_ & ~new_n15579_;
  assign A3244 = ~new_n15562_ & ~new_n15580_;
  assign new_n15582_ = ~new_n15559_ & ~new_n15578_;
  assign A3243 = ~new_n15562_ & ~new_n15582_;
  assign new_n15584_ = new_n15559_ & new_n15566_;
  assign new_n15585_ = ~new_n15562_ & ~new_n15584_;
  assign new_n15586_ = new_n15562_ & ~new_n15585_;
  assign new_n15587_ = new_n15562_ & new_n15584_;
  assign new_n15588_ = new_n15586_ & ~new_n15587_;
  assign new_n15589_ = new_n15566_ & ~new_n15588_;
  assign A3242 = new_n15577_ | new_n15589_;
  assign new_n15591_ = new_n15570_ & new_n15575_;
  assign new_n15592_ = ~new_n15576_ & ~new_n15591_;
  assign new_n15593_ = ~new_n15562_ & ~new_n15570_;
  assign new_n15594_ = new_n15562_ & new_n15570_;
  assign new_n15595_ = ~new_n15593_ & ~new_n15594_;
  assign new_n15596_ = new_n15592_ & ~new_n15595_;
  assign A3241 = new_n15589_ | new_n15596_;
  assign new_n15598_ = new_n15566_ & ~new_n15596_;
  assign new_n15599_ = ~new_n15566_ & new_n15596_;
  assign new_n15600_ = ~new_n15598_ & ~new_n15599_;
  assign A3240 = ~new_n15562_ & ~new_n15600_;
  assign new_n15602_ = ~new_n7843_ & ~new_n14166_;
  assign new_n15603_ = new_n7843_ & new_n14166_;
  assign new_n15604_ = ~new_n15602_ & ~new_n15603_;
  assign new_n15605_ = ~new_n7836_ & ~new_n15604_;
  assign new_n15606_ = ~new_n7888_ & ~new_n14173_;
  assign new_n15607_ = new_n7888_ & new_n14173_;
  assign new_n15608_ = ~new_n15606_ & ~new_n15607_;
  assign new_n15609_ = ~new_n7881_ & ~new_n15608_;
  assign new_n15610_ = ~new_n15605_ & new_n15609_;
  assign new_n15611_ = new_n15605_ & ~new_n15609_;
  assign new_n15612_ = ~new_n15610_ & ~new_n15611_;
  assign new_n15613_ = ~new_n7936_ & ~new_n14183_;
  assign new_n15614_ = new_n7936_ & new_n14183_;
  assign new_n15615_ = ~new_n15613_ & ~new_n15614_;
  assign new_n15616_ = ~new_n7929_ & ~new_n15615_;
  assign new_n15617_ = ~new_n7981_ & ~new_n14190_;
  assign new_n15618_ = new_n7981_ & new_n14190_;
  assign new_n15619_ = ~new_n15617_ & ~new_n15618_;
  assign new_n15620_ = ~new_n7974_ & ~new_n15619_;
  assign new_n15621_ = new_n15612_ & ~new_n15620_;
  assign new_n15622_ = ~new_n8027_ & ~new_n14198_;
  assign new_n15623_ = new_n8027_ & new_n14198_;
  assign new_n15624_ = ~new_n15622_ & ~new_n15623_;
  assign new_n15625_ = ~new_n8020_ & ~new_n15624_;
  assign new_n15626_ = ~new_n15620_ & ~new_n15625_;
  assign new_n15627_ = ~new_n15621_ & ~new_n15626_;
  assign new_n15628_ = new_n15616_ & new_n15627_;
  assign new_n15629_ = ~new_n15616_ & ~new_n15627_;
  assign new_n15630_ = ~new_n15628_ & ~new_n15629_;
  assign A3211 = ~new_n15612_ & ~new_n15630_;
  assign new_n15632_ = ~new_n15609_ & ~new_n15628_;
  assign A3210 = ~new_n15612_ & ~new_n15632_;
  assign new_n15634_ = new_n15609_ & new_n15616_;
  assign new_n15635_ = ~new_n15612_ & ~new_n15634_;
  assign new_n15636_ = new_n15612_ & ~new_n15635_;
  assign new_n15637_ = new_n15612_ & new_n15634_;
  assign new_n15638_ = new_n15636_ & ~new_n15637_;
  assign new_n15639_ = new_n15616_ & ~new_n15638_;
  assign A3209 = new_n15627_ | new_n15639_;
  assign new_n15641_ = new_n15620_ & new_n15625_;
  assign new_n15642_ = ~new_n15626_ & ~new_n15641_;
  assign new_n15643_ = ~new_n15612_ & ~new_n15620_;
  assign new_n15644_ = new_n15612_ & new_n15620_;
  assign new_n15645_ = ~new_n15643_ & ~new_n15644_;
  assign new_n15646_ = new_n15642_ & ~new_n15645_;
  assign A3208 = new_n15639_ | new_n15646_;
  assign new_n15648_ = new_n15616_ & ~new_n15646_;
  assign new_n15649_ = ~new_n15616_ & new_n15646_;
  assign new_n15650_ = ~new_n15648_ & ~new_n15649_;
  assign A3207 = ~new_n15612_ & ~new_n15650_;
  assign new_n15652_ = ~new_n8098_ & ~new_n14231_;
  assign new_n15653_ = new_n8098_ & new_n14231_;
  assign new_n15654_ = ~new_n15652_ & ~new_n15653_;
  assign new_n15655_ = ~new_n8091_ & ~new_n15654_;
  assign new_n15656_ = ~new_n8143_ & ~new_n14238_;
  assign new_n15657_ = new_n8143_ & new_n14238_;
  assign new_n15658_ = ~new_n15656_ & ~new_n15657_;
  assign new_n15659_ = ~new_n8136_ & ~new_n15658_;
  assign new_n15660_ = ~new_n15655_ & new_n15659_;
  assign new_n15661_ = new_n15655_ & ~new_n15659_;
  assign new_n15662_ = ~new_n15660_ & ~new_n15661_;
  assign new_n15663_ = ~new_n8191_ & ~new_n14248_;
  assign new_n15664_ = new_n8191_ & new_n14248_;
  assign new_n15665_ = ~new_n15663_ & ~new_n15664_;
  assign new_n15666_ = ~new_n8184_ & ~new_n15665_;
  assign new_n15667_ = ~new_n8236_ & ~new_n14255_;
  assign new_n15668_ = new_n8236_ & new_n14255_;
  assign new_n15669_ = ~new_n15667_ & ~new_n15668_;
  assign new_n15670_ = ~new_n8229_ & ~new_n15669_;
  assign new_n15671_ = new_n15662_ & ~new_n15670_;
  assign new_n15672_ = ~new_n8282_ & ~new_n14263_;
  assign new_n15673_ = new_n8282_ & new_n14263_;
  assign new_n15674_ = ~new_n15672_ & ~new_n15673_;
  assign new_n15675_ = ~new_n8275_ & ~new_n15674_;
  assign new_n15676_ = ~new_n15670_ & ~new_n15675_;
  assign new_n15677_ = ~new_n15671_ & ~new_n15676_;
  assign new_n15678_ = new_n15666_ & new_n15677_;
  assign new_n15679_ = ~new_n15666_ & ~new_n15677_;
  assign new_n15680_ = ~new_n15678_ & ~new_n15679_;
  assign A3178 = ~new_n15662_ & ~new_n15680_;
  assign new_n15682_ = ~new_n15659_ & ~new_n15678_;
  assign A3177 = ~new_n15662_ & ~new_n15682_;
  assign new_n15684_ = new_n15659_ & new_n15666_;
  assign new_n15685_ = ~new_n15662_ & ~new_n15684_;
  assign new_n15686_ = new_n15662_ & ~new_n15685_;
  assign new_n15687_ = new_n15662_ & new_n15684_;
  assign new_n15688_ = new_n15686_ & ~new_n15687_;
  assign new_n15689_ = new_n15666_ & ~new_n15688_;
  assign A3176 = new_n15677_ | new_n15689_;
  assign new_n15691_ = new_n15670_ & new_n15675_;
  assign new_n15692_ = ~new_n15676_ & ~new_n15691_;
  assign new_n15693_ = ~new_n15662_ & ~new_n15670_;
  assign new_n15694_ = new_n15662_ & new_n15670_;
  assign new_n15695_ = ~new_n15693_ & ~new_n15694_;
  assign new_n15696_ = new_n15692_ & ~new_n15695_;
  assign A3175 = new_n15689_ | new_n15696_;
  assign new_n15698_ = new_n15666_ & ~new_n15696_;
  assign new_n15699_ = ~new_n15666_ & new_n15696_;
  assign new_n15700_ = ~new_n15698_ & ~new_n15699_;
  assign A3174 = ~new_n15662_ & ~new_n15700_;
  assign new_n15702_ = ~new_n8349_ & ~new_n14296_;
  assign new_n15703_ = new_n8349_ & new_n14296_;
  assign new_n15704_ = ~new_n15702_ & ~new_n15703_;
  assign new_n15705_ = ~new_n8342_ & ~new_n15704_;
  assign new_n15706_ = ~new_n8394_ & ~new_n14303_;
  assign new_n15707_ = new_n8394_ & new_n14303_;
  assign new_n15708_ = ~new_n15706_ & ~new_n15707_;
  assign new_n15709_ = ~new_n8387_ & ~new_n15708_;
  assign new_n15710_ = ~new_n15705_ & new_n15709_;
  assign new_n15711_ = new_n15705_ & ~new_n15709_;
  assign new_n15712_ = ~new_n15710_ & ~new_n15711_;
  assign new_n15713_ = ~new_n8442_ & ~new_n14313_;
  assign new_n15714_ = new_n8442_ & new_n14313_;
  assign new_n15715_ = ~new_n15713_ & ~new_n15714_;
  assign new_n15716_ = ~new_n8435_ & ~new_n15715_;
  assign new_n15717_ = ~new_n8487_ & ~new_n14320_;
  assign new_n15718_ = new_n8487_ & new_n14320_;
  assign new_n15719_ = ~new_n15717_ & ~new_n15718_;
  assign new_n15720_ = ~new_n8480_ & ~new_n15719_;
  assign new_n15721_ = new_n15712_ & ~new_n15720_;
  assign new_n15722_ = ~new_n8533_ & ~new_n14328_;
  assign new_n15723_ = new_n8533_ & new_n14328_;
  assign new_n15724_ = ~new_n15722_ & ~new_n15723_;
  assign new_n15725_ = ~new_n8526_ & ~new_n15724_;
  assign new_n15726_ = ~new_n15720_ & ~new_n15725_;
  assign new_n15727_ = ~new_n15721_ & ~new_n15726_;
  assign new_n15728_ = new_n15716_ & new_n15727_;
  assign new_n15729_ = ~new_n15716_ & ~new_n15727_;
  assign new_n15730_ = ~new_n15728_ & ~new_n15729_;
  assign A3145 = ~new_n15712_ & ~new_n15730_;
  assign new_n15732_ = ~new_n15709_ & ~new_n15728_;
  assign A3144 = ~new_n15712_ & ~new_n15732_;
  assign new_n15734_ = new_n15709_ & new_n15716_;
  assign new_n15735_ = ~new_n15712_ & ~new_n15734_;
  assign new_n15736_ = new_n15712_ & ~new_n15735_;
  assign new_n15737_ = new_n15712_ & new_n15734_;
  assign new_n15738_ = new_n15736_ & ~new_n15737_;
  assign new_n15739_ = new_n15716_ & ~new_n15738_;
  assign A3143 = new_n15727_ | new_n15739_;
  assign new_n15741_ = new_n15720_ & new_n15725_;
  assign new_n15742_ = ~new_n15726_ & ~new_n15741_;
  assign new_n15743_ = ~new_n15712_ & ~new_n15720_;
  assign new_n15744_ = new_n15712_ & new_n15720_;
  assign new_n15745_ = ~new_n15743_ & ~new_n15744_;
  assign new_n15746_ = new_n15742_ & ~new_n15745_;
  assign A3142 = new_n15739_ | new_n15746_;
  assign new_n15748_ = new_n15716_ & ~new_n15746_;
  assign new_n15749_ = ~new_n15716_ & new_n15746_;
  assign new_n15750_ = ~new_n15748_ & ~new_n15749_;
  assign A3141 = ~new_n15712_ & ~new_n15750_;
  assign new_n15752_ = ~new_n8604_ & ~new_n14361_;
  assign new_n15753_ = new_n8604_ & new_n14361_;
  assign new_n15754_ = ~new_n15752_ & ~new_n15753_;
  assign new_n15755_ = ~new_n8597_ & ~new_n15754_;
  assign new_n15756_ = ~new_n8649_ & ~new_n14368_;
  assign new_n15757_ = new_n8649_ & new_n14368_;
  assign new_n15758_ = ~new_n15756_ & ~new_n15757_;
  assign new_n15759_ = ~new_n8642_ & ~new_n15758_;
  assign new_n15760_ = ~new_n15755_ & new_n15759_;
  assign new_n15761_ = new_n15755_ & ~new_n15759_;
  assign new_n15762_ = ~new_n15760_ & ~new_n15761_;
  assign new_n15763_ = ~new_n8697_ & ~new_n14378_;
  assign new_n15764_ = new_n8697_ & new_n14378_;
  assign new_n15765_ = ~new_n15763_ & ~new_n15764_;
  assign new_n15766_ = ~new_n8690_ & ~new_n15765_;
  assign new_n15767_ = ~new_n8742_ & ~new_n14385_;
  assign new_n15768_ = new_n8742_ & new_n14385_;
  assign new_n15769_ = ~new_n15767_ & ~new_n15768_;
  assign new_n15770_ = ~new_n8735_ & ~new_n15769_;
  assign new_n15771_ = new_n15762_ & ~new_n15770_;
  assign new_n15772_ = ~new_n8788_ & ~new_n14393_;
  assign new_n15773_ = new_n8788_ & new_n14393_;
  assign new_n15774_ = ~new_n15772_ & ~new_n15773_;
  assign new_n15775_ = ~new_n8781_ & ~new_n15774_;
  assign new_n15776_ = ~new_n15770_ & ~new_n15775_;
  assign new_n15777_ = ~new_n15771_ & ~new_n15776_;
  assign new_n15778_ = new_n15766_ & new_n15777_;
  assign new_n15779_ = ~new_n15766_ & ~new_n15777_;
  assign new_n15780_ = ~new_n15778_ & ~new_n15779_;
  assign A3112 = ~new_n15762_ & ~new_n15780_;
  assign new_n15782_ = ~new_n15759_ & ~new_n15778_;
  assign A3111 = ~new_n15762_ & ~new_n15782_;
  assign new_n15784_ = new_n15759_ & new_n15766_;
  assign new_n15785_ = ~new_n15762_ & ~new_n15784_;
  assign new_n15786_ = new_n15762_ & ~new_n15785_;
  assign new_n15787_ = new_n15762_ & new_n15784_;
  assign new_n15788_ = new_n15786_ & ~new_n15787_;
  assign new_n15789_ = new_n15766_ & ~new_n15788_;
  assign A3110 = new_n15777_ | new_n15789_;
  assign new_n15791_ = new_n15770_ & new_n15775_;
  assign new_n15792_ = ~new_n15776_ & ~new_n15791_;
  assign new_n15793_ = ~new_n15762_ & ~new_n15770_;
  assign new_n15794_ = new_n15762_ & new_n15770_;
  assign new_n15795_ = ~new_n15793_ & ~new_n15794_;
  assign new_n15796_ = new_n15792_ & ~new_n15795_;
  assign A3109 = new_n15789_ | new_n15796_;
  assign new_n15798_ = new_n15766_ & ~new_n15796_;
  assign new_n15799_ = ~new_n15766_ & new_n15796_;
  assign new_n15800_ = ~new_n15798_ & ~new_n15799_;
  assign A3108 = ~new_n15762_ & ~new_n15800_;
  assign new_n15802_ = ~new_n8859_ & ~new_n14426_;
  assign new_n15803_ = new_n8859_ & new_n14426_;
  assign new_n15804_ = ~new_n15802_ & ~new_n15803_;
  assign new_n15805_ = ~new_n8852_ & ~new_n15804_;
  assign new_n15806_ = ~new_n8904_ & ~new_n14433_;
  assign new_n15807_ = new_n8904_ & new_n14433_;
  assign new_n15808_ = ~new_n15806_ & ~new_n15807_;
  assign new_n15809_ = ~new_n8897_ & ~new_n15808_;
  assign new_n15810_ = ~new_n15805_ & new_n15809_;
  assign new_n15811_ = new_n15805_ & ~new_n15809_;
  assign new_n15812_ = ~new_n15810_ & ~new_n15811_;
  assign new_n15813_ = ~new_n8952_ & ~new_n14443_;
  assign new_n15814_ = new_n8952_ & new_n14443_;
  assign new_n15815_ = ~new_n15813_ & ~new_n15814_;
  assign new_n15816_ = ~new_n8945_ & ~new_n15815_;
  assign new_n15817_ = ~new_n8997_ & ~new_n14450_;
  assign new_n15818_ = new_n8997_ & new_n14450_;
  assign new_n15819_ = ~new_n15817_ & ~new_n15818_;
  assign new_n15820_ = ~new_n8990_ & ~new_n15819_;
  assign new_n15821_ = new_n15812_ & ~new_n15820_;
  assign new_n15822_ = ~new_n9043_ & ~new_n14458_;
  assign new_n15823_ = new_n9043_ & new_n14458_;
  assign new_n15824_ = ~new_n15822_ & ~new_n15823_;
  assign new_n15825_ = ~new_n9036_ & ~new_n15824_;
  assign new_n15826_ = ~new_n15820_ & ~new_n15825_;
  assign new_n15827_ = ~new_n15821_ & ~new_n15826_;
  assign new_n15828_ = new_n15816_ & new_n15827_;
  assign new_n15829_ = ~new_n15816_ & ~new_n15827_;
  assign new_n15830_ = ~new_n15828_ & ~new_n15829_;
  assign A3079 = ~new_n15812_ & ~new_n15830_;
  assign new_n15832_ = ~new_n15809_ & ~new_n15828_;
  assign A3078 = ~new_n15812_ & ~new_n15832_;
  assign new_n15834_ = new_n15809_ & new_n15816_;
  assign new_n15835_ = ~new_n15812_ & ~new_n15834_;
  assign new_n15836_ = new_n15812_ & ~new_n15835_;
  assign new_n15837_ = new_n15812_ & new_n15834_;
  assign new_n15838_ = new_n15836_ & ~new_n15837_;
  assign new_n15839_ = new_n15816_ & ~new_n15838_;
  assign A3077 = new_n15827_ | new_n15839_;
  assign new_n15841_ = new_n15820_ & new_n15825_;
  assign new_n15842_ = ~new_n15826_ & ~new_n15841_;
  assign new_n15843_ = ~new_n15812_ & ~new_n15820_;
  assign new_n15844_ = new_n15812_ & new_n15820_;
  assign new_n15845_ = ~new_n15843_ & ~new_n15844_;
  assign new_n15846_ = new_n15842_ & ~new_n15845_;
  assign A3076 = new_n15839_ | new_n15846_;
  assign new_n15848_ = new_n15816_ & ~new_n15846_;
  assign new_n15849_ = ~new_n15816_ & new_n15846_;
  assign new_n15850_ = ~new_n15848_ & ~new_n15849_;
  assign A3075 = ~new_n15812_ & ~new_n15850_;
  assign new_n15852_ = ~new_n9114_ & ~new_n14491_;
  assign new_n15853_ = new_n9114_ & new_n14491_;
  assign new_n15854_ = ~new_n15852_ & ~new_n15853_;
  assign new_n15855_ = ~new_n9107_ & ~new_n15854_;
  assign new_n15856_ = ~new_n9159_ & ~new_n14498_;
  assign new_n15857_ = new_n9159_ & new_n14498_;
  assign new_n15858_ = ~new_n15856_ & ~new_n15857_;
  assign new_n15859_ = ~new_n9152_ & ~new_n15858_;
  assign new_n15860_ = ~new_n15855_ & new_n15859_;
  assign new_n15861_ = new_n15855_ & ~new_n15859_;
  assign new_n15862_ = ~new_n15860_ & ~new_n15861_;
  assign new_n15863_ = ~new_n9207_ & ~new_n14508_;
  assign new_n15864_ = new_n9207_ & new_n14508_;
  assign new_n15865_ = ~new_n15863_ & ~new_n15864_;
  assign new_n15866_ = ~new_n9200_ & ~new_n15865_;
  assign new_n15867_ = ~new_n9252_ & ~new_n14515_;
  assign new_n15868_ = new_n9252_ & new_n14515_;
  assign new_n15869_ = ~new_n15867_ & ~new_n15868_;
  assign new_n15870_ = ~new_n9245_ & ~new_n15869_;
  assign new_n15871_ = new_n15862_ & ~new_n15870_;
  assign new_n15872_ = ~new_n9298_ & ~new_n14523_;
  assign new_n15873_ = new_n9298_ & new_n14523_;
  assign new_n15874_ = ~new_n15872_ & ~new_n15873_;
  assign new_n15875_ = ~new_n9291_ & ~new_n15874_;
  assign new_n15876_ = ~new_n15870_ & ~new_n15875_;
  assign new_n15877_ = ~new_n15871_ & ~new_n15876_;
  assign new_n15878_ = new_n15866_ & new_n15877_;
  assign new_n15879_ = ~new_n15866_ & ~new_n15877_;
  assign new_n15880_ = ~new_n15878_ & ~new_n15879_;
  assign A3046 = ~new_n15862_ & ~new_n15880_;
  assign new_n15882_ = ~new_n15859_ & ~new_n15878_;
  assign A3045 = ~new_n15862_ & ~new_n15882_;
  assign new_n15884_ = new_n15859_ & new_n15866_;
  assign new_n15885_ = ~new_n15862_ & ~new_n15884_;
  assign new_n15886_ = new_n15862_ & ~new_n15885_;
  assign new_n15887_ = new_n15862_ & new_n15884_;
  assign new_n15888_ = new_n15886_ & ~new_n15887_;
  assign new_n15889_ = new_n15866_ & ~new_n15888_;
  assign A3044 = new_n15877_ | new_n15889_;
  assign new_n15891_ = new_n15870_ & new_n15875_;
  assign new_n15892_ = ~new_n15876_ & ~new_n15891_;
  assign new_n15893_ = ~new_n15862_ & ~new_n15870_;
  assign new_n15894_ = new_n15862_ & new_n15870_;
  assign new_n15895_ = ~new_n15893_ & ~new_n15894_;
  assign new_n15896_ = new_n15892_ & ~new_n15895_;
  assign A3043 = new_n15889_ | new_n15896_;
  assign new_n15898_ = new_n15866_ & ~new_n15896_;
  assign new_n15899_ = ~new_n15866_ & new_n15896_;
  assign new_n15900_ = ~new_n15898_ & ~new_n15899_;
  assign A3042 = ~new_n15862_ & ~new_n15900_;
  assign new_n15902_ = ~new_n9369_ & ~new_n14556_;
  assign new_n15903_ = new_n9369_ & new_n14556_;
  assign new_n15904_ = ~new_n15902_ & ~new_n15903_;
  assign new_n15905_ = ~new_n9362_ & ~new_n15904_;
  assign new_n15906_ = ~new_n9414_ & ~new_n14563_;
  assign new_n15907_ = new_n9414_ & new_n14563_;
  assign new_n15908_ = ~new_n15906_ & ~new_n15907_;
  assign new_n15909_ = ~new_n9407_ & ~new_n15908_;
  assign new_n15910_ = ~new_n15905_ & new_n15909_;
  assign new_n15911_ = new_n15905_ & ~new_n15909_;
  assign new_n15912_ = ~new_n15910_ & ~new_n15911_;
  assign new_n15913_ = ~new_n9462_ & ~new_n14573_;
  assign new_n15914_ = new_n9462_ & new_n14573_;
  assign new_n15915_ = ~new_n15913_ & ~new_n15914_;
  assign new_n15916_ = ~new_n9455_ & ~new_n15915_;
  assign new_n15917_ = ~new_n9507_ & ~new_n14580_;
  assign new_n15918_ = new_n9507_ & new_n14580_;
  assign new_n15919_ = ~new_n15917_ & ~new_n15918_;
  assign new_n15920_ = ~new_n9500_ & ~new_n15919_;
  assign new_n15921_ = new_n15912_ & ~new_n15920_;
  assign new_n15922_ = ~new_n9553_ & ~new_n14588_;
  assign new_n15923_ = new_n9553_ & new_n14588_;
  assign new_n15924_ = ~new_n15922_ & ~new_n15923_;
  assign new_n15925_ = ~new_n9546_ & ~new_n15924_;
  assign new_n15926_ = ~new_n15920_ & ~new_n15925_;
  assign new_n15927_ = ~new_n15921_ & ~new_n15926_;
  assign new_n15928_ = new_n15916_ & new_n15927_;
  assign new_n15929_ = ~new_n15916_ & ~new_n15927_;
  assign new_n15930_ = ~new_n15928_ & ~new_n15929_;
  assign A3013 = ~new_n15912_ & ~new_n15930_;
  assign new_n15932_ = ~new_n15909_ & ~new_n15928_;
  assign A3012 = ~new_n15912_ & ~new_n15932_;
  assign new_n15934_ = new_n15909_ & new_n15916_;
  assign new_n15935_ = ~new_n15912_ & ~new_n15934_;
  assign new_n15936_ = new_n15912_ & ~new_n15935_;
  assign new_n15937_ = new_n15912_ & new_n15934_;
  assign new_n15938_ = new_n15936_ & ~new_n15937_;
  assign new_n15939_ = new_n15916_ & ~new_n15938_;
  assign A3011 = new_n15927_ | new_n15939_;
  assign new_n15941_ = new_n15920_ & new_n15925_;
  assign new_n15942_ = ~new_n15926_ & ~new_n15941_;
  assign new_n15943_ = ~new_n15912_ & ~new_n15920_;
  assign new_n15944_ = new_n15912_ & new_n15920_;
  assign new_n15945_ = ~new_n15943_ & ~new_n15944_;
  assign new_n15946_ = new_n15942_ & ~new_n15945_;
  assign A3010 = new_n15939_ | new_n15946_;
  assign new_n15948_ = new_n15916_ & ~new_n15946_;
  assign new_n15949_ = ~new_n15916_ & new_n15946_;
  assign new_n15950_ = ~new_n15948_ & ~new_n15949_;
  assign A3009 = ~new_n15912_ & ~new_n15950_;
  assign new_n15952_ = ~new_n9620_ & ~new_n14621_;
  assign new_n15953_ = new_n9620_ & new_n14621_;
  assign new_n15954_ = ~new_n15952_ & ~new_n15953_;
  assign new_n15955_ = ~new_n9613_ & ~new_n15954_;
  assign new_n15956_ = ~new_n9665_ & ~new_n14628_;
  assign new_n15957_ = new_n9665_ & new_n14628_;
  assign new_n15958_ = ~new_n15956_ & ~new_n15957_;
  assign new_n15959_ = ~new_n9658_ & ~new_n15958_;
  assign new_n15960_ = ~new_n15955_ & new_n15959_;
  assign new_n15961_ = new_n15955_ & ~new_n15959_;
  assign new_n15962_ = ~new_n15960_ & ~new_n15961_;
  assign new_n15963_ = ~new_n9713_ & ~new_n14638_;
  assign new_n15964_ = new_n9713_ & new_n14638_;
  assign new_n15965_ = ~new_n15963_ & ~new_n15964_;
  assign new_n15966_ = ~new_n9706_ & ~new_n15965_;
  assign new_n15967_ = ~new_n9758_ & ~new_n14645_;
  assign new_n15968_ = new_n9758_ & new_n14645_;
  assign new_n15969_ = ~new_n15967_ & ~new_n15968_;
  assign new_n15970_ = ~new_n9751_ & ~new_n15969_;
  assign new_n15971_ = new_n15962_ & ~new_n15970_;
  assign new_n15972_ = ~new_n9804_ & ~new_n14653_;
  assign new_n15973_ = new_n9804_ & new_n14653_;
  assign new_n15974_ = ~new_n15972_ & ~new_n15973_;
  assign new_n15975_ = ~new_n9797_ & ~new_n15974_;
  assign new_n15976_ = ~new_n15970_ & ~new_n15975_;
  assign new_n15977_ = ~new_n15971_ & ~new_n15976_;
  assign new_n15978_ = new_n15966_ & new_n15977_;
  assign new_n15979_ = ~new_n15966_ & ~new_n15977_;
  assign new_n15980_ = ~new_n15978_ & ~new_n15979_;
  assign A2980 = ~new_n15962_ & ~new_n15980_;
  assign new_n15982_ = ~new_n15959_ & ~new_n15978_;
  assign A2979 = ~new_n15962_ & ~new_n15982_;
  assign new_n15984_ = new_n15959_ & new_n15966_;
  assign new_n15985_ = ~new_n15962_ & ~new_n15984_;
  assign new_n15986_ = new_n15962_ & ~new_n15985_;
  assign new_n15987_ = new_n15962_ & new_n15984_;
  assign new_n15988_ = new_n15986_ & ~new_n15987_;
  assign new_n15989_ = new_n15966_ & ~new_n15988_;
  assign A2978 = new_n15977_ | new_n15989_;
  assign new_n15991_ = new_n15970_ & new_n15975_;
  assign new_n15992_ = ~new_n15976_ & ~new_n15991_;
  assign new_n15993_ = ~new_n15962_ & ~new_n15970_;
  assign new_n15994_ = new_n15962_ & new_n15970_;
  assign new_n15995_ = ~new_n15993_ & ~new_n15994_;
  assign new_n15996_ = new_n15992_ & ~new_n15995_;
  assign A2977 = new_n15989_ | new_n15996_;
  assign new_n15998_ = new_n15966_ & ~new_n15996_;
  assign new_n15999_ = ~new_n15966_ & new_n15996_;
  assign new_n16000_ = ~new_n15998_ & ~new_n15999_;
  assign A2976 = ~new_n15962_ & ~new_n16000_;
  assign new_n16002_ = new_n9866_ & ~new_n14686_;
  assign new_n16003_ = ~new_n9866_ & new_n14686_;
  assign new_n16004_ = ~new_n16002_ & ~new_n16003_;
  assign new_n16005_ = ~new_n9862_ & ~new_n16004_;
  assign new_n16006_ = new_n9896_ & ~new_n14693_;
  assign new_n16007_ = ~new_n9896_ & new_n14693_;
  assign new_n16008_ = ~new_n16006_ & ~new_n16007_;
  assign new_n16009_ = ~new_n9892_ & ~new_n16008_;
  assign new_n16010_ = ~new_n16005_ & new_n16009_;
  assign new_n16011_ = new_n16005_ & ~new_n16009_;
  assign new_n16012_ = ~new_n16010_ & ~new_n16011_;
  assign new_n16013_ = new_n9929_ & ~new_n14703_;
  assign new_n16014_ = ~new_n9929_ & new_n14703_;
  assign new_n16015_ = ~new_n16013_ & ~new_n16014_;
  assign new_n16016_ = ~new_n9925_ & ~new_n16015_;
  assign new_n16017_ = new_n9959_ & ~new_n14710_;
  assign new_n16018_ = ~new_n9959_ & new_n14710_;
  assign new_n16019_ = ~new_n16017_ & ~new_n16018_;
  assign new_n16020_ = ~new_n9955_ & ~new_n16019_;
  assign new_n16021_ = new_n16012_ & ~new_n16020_;
  assign new_n16022_ = new_n9990_ & ~new_n14718_;
  assign new_n16023_ = ~new_n9990_ & new_n14718_;
  assign new_n16024_ = ~new_n16022_ & ~new_n16023_;
  assign new_n16025_ = ~new_n9986_ & ~new_n16024_;
  assign new_n16026_ = ~new_n16020_ & ~new_n16025_;
  assign new_n16027_ = ~new_n16021_ & ~new_n16026_;
  assign new_n16028_ = new_n16016_ & new_n16027_;
  assign new_n16029_ = ~new_n16016_ & ~new_n16027_;
  assign new_n16030_ = ~new_n16028_ & ~new_n16029_;
  assign A2947 = ~new_n16012_ & ~new_n16030_;
  assign new_n16032_ = ~new_n16009_ & ~new_n16028_;
  assign A2946 = ~new_n16012_ & ~new_n16032_;
  assign new_n16034_ = new_n16009_ & new_n16016_;
  assign new_n16035_ = ~new_n16012_ & ~new_n16034_;
  assign new_n16036_ = new_n16012_ & ~new_n16035_;
  assign new_n16037_ = new_n16012_ & new_n16034_;
  assign new_n16038_ = new_n16036_ & ~new_n16037_;
  assign new_n16039_ = new_n16016_ & ~new_n16038_;
  assign A2945 = new_n16027_ | new_n16039_;
  assign new_n16041_ = new_n16020_ & new_n16025_;
  assign new_n16042_ = ~new_n16026_ & ~new_n16041_;
  assign new_n16043_ = ~new_n16012_ & ~new_n16020_;
  assign new_n16044_ = new_n16012_ & new_n16020_;
  assign new_n16045_ = ~new_n16043_ & ~new_n16044_;
  assign new_n16046_ = new_n16042_ & ~new_n16045_;
  assign A2944 = new_n16039_ | new_n16046_;
  assign new_n16048_ = new_n16016_ & ~new_n16046_;
  assign new_n16049_ = ~new_n16016_ & new_n16046_;
  assign new_n16050_ = ~new_n16048_ & ~new_n16049_;
  assign A2943 = ~new_n16012_ & ~new_n16050_;
  assign new_n16052_ = new_n10046_ & ~new_n14751_;
  assign new_n16053_ = ~new_n10046_ & new_n14751_;
  assign new_n16054_ = ~new_n16052_ & ~new_n16053_;
  assign new_n16055_ = ~new_n10042_ & ~new_n16054_;
  assign new_n16056_ = new_n10076_ & ~new_n14758_;
  assign new_n16057_ = ~new_n10076_ & new_n14758_;
  assign new_n16058_ = ~new_n16056_ & ~new_n16057_;
  assign new_n16059_ = ~new_n10072_ & ~new_n16058_;
  assign new_n16060_ = ~new_n16055_ & new_n16059_;
  assign new_n16061_ = new_n16055_ & ~new_n16059_;
  assign new_n16062_ = ~new_n16060_ & ~new_n16061_;
  assign new_n16063_ = new_n10109_ & ~new_n14768_;
  assign new_n16064_ = ~new_n10109_ & new_n14768_;
  assign new_n16065_ = ~new_n16063_ & ~new_n16064_;
  assign new_n16066_ = ~new_n10105_ & ~new_n16065_;
  assign new_n16067_ = new_n10139_ & ~new_n14775_;
  assign new_n16068_ = ~new_n10139_ & new_n14775_;
  assign new_n16069_ = ~new_n16067_ & ~new_n16068_;
  assign new_n16070_ = ~new_n10135_ & ~new_n16069_;
  assign new_n16071_ = new_n16062_ & ~new_n16070_;
  assign new_n16072_ = new_n10170_ & ~new_n14783_;
  assign new_n16073_ = ~new_n10170_ & new_n14783_;
  assign new_n16074_ = ~new_n16072_ & ~new_n16073_;
  assign new_n16075_ = ~new_n10166_ & ~new_n16074_;
  assign new_n16076_ = ~new_n16070_ & ~new_n16075_;
  assign new_n16077_ = ~new_n16071_ & ~new_n16076_;
  assign new_n16078_ = new_n16066_ & new_n16077_;
  assign new_n16079_ = ~new_n16066_ & ~new_n16077_;
  assign new_n16080_ = ~new_n16078_ & ~new_n16079_;
  assign A2914 = ~new_n16062_ & ~new_n16080_;
  assign new_n16082_ = ~new_n16059_ & ~new_n16078_;
  assign A2913 = ~new_n16062_ & ~new_n16082_;
  assign new_n16084_ = new_n16059_ & new_n16066_;
  assign new_n16085_ = ~new_n16062_ & ~new_n16084_;
  assign new_n16086_ = new_n16062_ & ~new_n16085_;
  assign new_n16087_ = new_n16062_ & new_n16084_;
  assign new_n16088_ = new_n16086_ & ~new_n16087_;
  assign new_n16089_ = new_n16066_ & ~new_n16088_;
  assign A2912 = new_n16077_ | new_n16089_;
  assign new_n16091_ = new_n16070_ & new_n16075_;
  assign new_n16092_ = ~new_n16076_ & ~new_n16091_;
  assign new_n16093_ = ~new_n16062_ & ~new_n16070_;
  assign new_n16094_ = new_n16062_ & new_n16070_;
  assign new_n16095_ = ~new_n16093_ & ~new_n16094_;
  assign new_n16096_ = new_n16092_ & ~new_n16095_;
  assign A2911 = new_n16089_ | new_n16096_;
  assign new_n16098_ = new_n16066_ & ~new_n16096_;
  assign new_n16099_ = ~new_n16066_ & new_n16096_;
  assign new_n16100_ = ~new_n16098_ & ~new_n16099_;
  assign A2910 = ~new_n16062_ & ~new_n16100_;
  assign new_n16102_ = new_n10226_ & ~new_n14816_;
  assign new_n16103_ = ~new_n10226_ & new_n14816_;
  assign new_n16104_ = ~new_n16102_ & ~new_n16103_;
  assign new_n16105_ = ~new_n10222_ & ~new_n16104_;
  assign new_n16106_ = new_n10256_ & ~new_n14823_;
  assign new_n16107_ = ~new_n10256_ & new_n14823_;
  assign new_n16108_ = ~new_n16106_ & ~new_n16107_;
  assign new_n16109_ = ~new_n10252_ & ~new_n16108_;
  assign new_n16110_ = ~new_n16105_ & new_n16109_;
  assign new_n16111_ = new_n16105_ & ~new_n16109_;
  assign new_n16112_ = ~new_n16110_ & ~new_n16111_;
  assign new_n16113_ = new_n10289_ & ~new_n14833_;
  assign new_n16114_ = ~new_n10289_ & new_n14833_;
  assign new_n16115_ = ~new_n16113_ & ~new_n16114_;
  assign new_n16116_ = ~new_n10285_ & ~new_n16115_;
  assign new_n16117_ = new_n10319_ & ~new_n14840_;
  assign new_n16118_ = ~new_n10319_ & new_n14840_;
  assign new_n16119_ = ~new_n16117_ & ~new_n16118_;
  assign new_n16120_ = ~new_n10315_ & ~new_n16119_;
  assign new_n16121_ = new_n16112_ & ~new_n16120_;
  assign new_n16122_ = new_n10350_ & ~new_n14848_;
  assign new_n16123_ = ~new_n10350_ & new_n14848_;
  assign new_n16124_ = ~new_n16122_ & ~new_n16123_;
  assign new_n16125_ = ~new_n10346_ & ~new_n16124_;
  assign new_n16126_ = ~new_n16120_ & ~new_n16125_;
  assign new_n16127_ = ~new_n16121_ & ~new_n16126_;
  assign new_n16128_ = new_n16116_ & new_n16127_;
  assign new_n16129_ = ~new_n16116_ & ~new_n16127_;
  assign new_n16130_ = ~new_n16128_ & ~new_n16129_;
  assign A2881 = ~new_n16112_ & ~new_n16130_;
  assign new_n16132_ = ~new_n16109_ & ~new_n16128_;
  assign A2880 = ~new_n16112_ & ~new_n16132_;
  assign new_n16134_ = new_n16109_ & new_n16116_;
  assign new_n16135_ = ~new_n16112_ & ~new_n16134_;
  assign new_n16136_ = new_n16112_ & ~new_n16135_;
  assign new_n16137_ = new_n16112_ & new_n16134_;
  assign new_n16138_ = new_n16136_ & ~new_n16137_;
  assign new_n16139_ = new_n16116_ & ~new_n16138_;
  assign A2879 = new_n16127_ | new_n16139_;
  assign new_n16141_ = new_n16120_ & new_n16125_;
  assign new_n16142_ = ~new_n16126_ & ~new_n16141_;
  assign new_n16143_ = ~new_n16112_ & ~new_n16120_;
  assign new_n16144_ = new_n16112_ & new_n16120_;
  assign new_n16145_ = ~new_n16143_ & ~new_n16144_;
  assign new_n16146_ = new_n16142_ & ~new_n16145_;
  assign A2878 = new_n16139_ | new_n16146_;
  assign new_n16148_ = new_n16116_ & ~new_n16146_;
  assign new_n16149_ = ~new_n16116_ & new_n16146_;
  assign new_n16150_ = ~new_n16148_ & ~new_n16149_;
  assign A2877 = ~new_n16112_ & ~new_n16150_;
  assign new_n16152_ = new_n10406_ & ~new_n14881_;
  assign new_n16153_ = ~new_n10406_ & new_n14881_;
  assign new_n16154_ = ~new_n16152_ & ~new_n16153_;
  assign new_n16155_ = ~new_n10402_ & ~new_n16154_;
  assign new_n16156_ = new_n10436_ & ~new_n14888_;
  assign new_n16157_ = ~new_n10436_ & new_n14888_;
  assign new_n16158_ = ~new_n16156_ & ~new_n16157_;
  assign new_n16159_ = ~new_n10432_ & ~new_n16158_;
  assign new_n16160_ = ~new_n16155_ & new_n16159_;
  assign new_n16161_ = new_n16155_ & ~new_n16159_;
  assign new_n16162_ = ~new_n16160_ & ~new_n16161_;
  assign new_n16163_ = new_n10469_ & ~new_n14898_;
  assign new_n16164_ = ~new_n10469_ & new_n14898_;
  assign new_n16165_ = ~new_n16163_ & ~new_n16164_;
  assign new_n16166_ = ~new_n10465_ & ~new_n16165_;
  assign new_n16167_ = new_n10499_ & ~new_n14905_;
  assign new_n16168_ = ~new_n10499_ & new_n14905_;
  assign new_n16169_ = ~new_n16167_ & ~new_n16168_;
  assign new_n16170_ = ~new_n10495_ & ~new_n16169_;
  assign new_n16171_ = new_n16162_ & ~new_n16170_;
  assign new_n16172_ = new_n10530_ & ~new_n14913_;
  assign new_n16173_ = ~new_n10530_ & new_n14913_;
  assign new_n16174_ = ~new_n16172_ & ~new_n16173_;
  assign new_n16175_ = ~new_n10526_ & ~new_n16174_;
  assign new_n16176_ = ~new_n16170_ & ~new_n16175_;
  assign new_n16177_ = ~new_n16171_ & ~new_n16176_;
  assign new_n16178_ = new_n16166_ & new_n16177_;
  assign new_n16179_ = ~new_n16166_ & ~new_n16177_;
  assign new_n16180_ = ~new_n16178_ & ~new_n16179_;
  assign A2848 = ~new_n16162_ & ~new_n16180_;
  assign new_n16182_ = ~new_n16159_ & ~new_n16178_;
  assign A2847 = ~new_n16162_ & ~new_n16182_;
  assign new_n16184_ = new_n16159_ & new_n16166_;
  assign new_n16185_ = ~new_n16162_ & ~new_n16184_;
  assign new_n16186_ = new_n16162_ & ~new_n16185_;
  assign new_n16187_ = new_n16162_ & new_n16184_;
  assign new_n16188_ = new_n16186_ & ~new_n16187_;
  assign new_n16189_ = new_n16166_ & ~new_n16188_;
  assign A2846 = new_n16177_ | new_n16189_;
  assign new_n16191_ = new_n16170_ & new_n16175_;
  assign new_n16192_ = ~new_n16176_ & ~new_n16191_;
  assign new_n16193_ = ~new_n16162_ & ~new_n16170_;
  assign new_n16194_ = new_n16162_ & new_n16170_;
  assign new_n16195_ = ~new_n16193_ & ~new_n16194_;
  assign new_n16196_ = new_n16192_ & ~new_n16195_;
  assign A2845 = new_n16189_ | new_n16196_;
  assign new_n16198_ = new_n16166_ & ~new_n16196_;
  assign new_n16199_ = ~new_n16166_ & new_n16196_;
  assign new_n16200_ = ~new_n16198_ & ~new_n16199_;
  assign A2844 = ~new_n16162_ & ~new_n16200_;
  assign new_n16202_ = new_n10619_ & ~new_n14949_;
  assign new_n16203_ = ~new_n10619_ & new_n14949_;
  assign new_n16204_ = ~new_n16202_ & ~new_n16203_;
  assign new_n16205_ = ~new_n10615_ & ~new_n16204_;
  assign new_n16206_ = ~new_n10600_ & ~new_n13321_;
  assign new_n16207_ = ~new_n14941_ & ~new_n16206_;
  assign new_n16208_ = ~new_n10592_ & ~new_n16207_;
  assign new_n16209_ = new_n16205_ & new_n16208_;
  assign new_n16210_ = ~new_n16205_ & ~new_n16208_;
  assign new_n16211_ = ~new_n16209_ & ~new_n16210_;
  assign new_n16212_ = new_n10713_ & ~new_n14974_;
  assign new_n16213_ = ~new_n10713_ & new_n14974_;
  assign new_n16214_ = ~new_n16212_ & ~new_n16213_;
  assign new_n16215_ = ~new_n10709_ & ~new_n16214_;
  assign new_n16216_ = new_n10682_ & ~new_n14966_;
  assign new_n16217_ = ~new_n10682_ & new_n14966_;
  assign new_n16218_ = ~new_n16216_ & ~new_n16217_;
  assign new_n16219_ = ~new_n10678_ & ~new_n16218_;
  assign new_n16220_ = ~new_n16215_ & new_n16219_;
  assign new_n16221_ = new_n16215_ & ~new_n16219_;
  assign new_n16222_ = ~new_n16220_ & ~new_n16221_;
  assign new_n16223_ = ~new_n16205_ & ~new_n16222_;
  assign new_n16224_ = new_n16205_ & new_n16222_;
  assign new_n16225_ = ~new_n16223_ & ~new_n16224_;
  assign new_n16226_ = new_n16211_ & ~new_n16225_;
  assign new_n16227_ = new_n10652_ & ~new_n14959_;
  assign new_n16228_ = ~new_n10652_ & new_n14959_;
  assign new_n16229_ = ~new_n16227_ & ~new_n16228_;
  assign new_n16230_ = ~new_n10648_ & ~new_n16229_;
  assign new_n16231_ = ~new_n16226_ & new_n16230_;
  assign new_n16232_ = new_n16226_ & ~new_n16230_;
  assign new_n16233_ = ~new_n16231_ & ~new_n16232_;
  assign A2811 = ~new_n16222_ & ~new_n16233_;
  assign new_n16235_ = new_n16219_ & new_n16230_;
  assign new_n16236_ = ~new_n16222_ & ~new_n16235_;
  assign new_n16237_ = new_n16222_ & ~new_n16236_;
  assign new_n16238_ = new_n16222_ & new_n16235_;
  assign new_n16239_ = new_n16237_ & ~new_n16238_;
  assign new_n16240_ = new_n16230_ & ~new_n16239_;
  assign A2812 = new_n16226_ | new_n16240_;
  assign new_n16242_ = ~new_n16205_ & new_n16222_;
  assign new_n16243_ = ~new_n16210_ & ~new_n16242_;
  assign A2813 = new_n16240_ | new_n16243_;
  assign new_n16245_ = new_n16230_ & new_n16243_;
  assign new_n16246_ = ~new_n16219_ & ~new_n16245_;
  assign A2814 = ~new_n16222_ & ~new_n16246_;
  assign new_n16248_ = ~new_n16230_ & ~new_n16243_;
  assign new_n16249_ = ~new_n16245_ & ~new_n16248_;
  assign A2815 = ~new_n16222_ & ~new_n16249_;
endmodule


