// Benchmark "b9" written by ABC on Fri Feb 25 15:12:38 2022

module b9 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1,
    h1, i1, j1  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0,
    o0;
  output p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1,
    g1, h1, i1, j1;
  wire new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n75_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n94_,
    new_n95_, new_n96_, new_n99_, new_n101_, new_n102_, new_n103_,
    new_n104_, new_n105_, new_n106_, new_n107_, new_n108_, new_n109_,
    new_n112_, new_n113_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n153_, new_n155_, new_n157_, new_n158_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_;
  assign new_n63_ = c0 & j0;
  assign new_n64_ = ~l0 & ~new_n63_;
  assign new_n65_ = b0 & ~new_n64_;
  assign new_n66_ = ~e & k;
  assign new_n67_ = ~c0 & j0;
  assign new_n68_ = ~k0 & ~new_n67_;
  assign new_n69_ = ~e & ~new_n68_;
  assign new_n70_ = b0 & new_n69_;
  assign new_n71_ = ~new_n66_ & ~new_n70_;
  assign new_n72_ = o0 & ~new_n71_;
  assign new_n73_ = n0 & new_n72_;
  assign b1 = ~new_n65_ & ~new_n73_;
  assign new_n75_ = ~p & ~b1;
  assign p0 = ~q | new_n75_;
  assign new_n77_ = e & b0;
  assign new_n78_ = k0 & new_n77_;
  assign new_n79_ = b0 & j0;
  assign new_n80_ = e & ~c0;
  assign new_n81_ = new_n79_ & new_n80_;
  assign new_n82_ = ~e0 & ~g0;
  assign new_n83_ = e & ~new_n82_;
  assign new_n84_ = ~new_n78_ & ~new_n81_;
  assign q0 = ~new_n83_ & new_n84_;
  assign new_n86_ = ~i & ~b0;
  assign new_n87_ = new_n67_ & ~new_n86_;
  assign new_n88_ = i & d0;
  assign new_n89_ = ~c & ~new_n88_;
  assign new_n90_ = e & ~new_n87_;
  assign new_n91_ = ~new_n89_ & ~new_n90_;
  assign new_n92_ = n0 & new_n91_;
  assign r0 = ~o0 | ~new_n92_;
  assign new_n94_ = ~b0 & l0;
  assign new_n95_ = b0 & new_n63_;
  assign new_n96_ = ~new_n94_ & ~new_n95_;
  assign s0 = ~v | new_n96_;
  assign t0 = v | new_n96_;
  assign new_n99_ = b0 & c0;
  assign v0 = ~l0 & ~new_n99_;
  assign new_n101_ = ~p & r;
  assign new_n102_ = ~f0 & ~new_n101_;
  assign new_n103_ = ~h0 & new_n102_;
  assign new_n104_ = o & ~new_n103_;
  assign new_n105_ = d & ~new_n104_;
  assign new_n106_ = ~o & z;
  assign new_n107_ = a & ~z;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = m0 & new_n108_;
  assign w0 = new_n105_ & ~new_n109_;
  assign x0 = n0 & o0;
  assign new_n112_ = a0 & i0;
  assign new_n113_ = l & b0;
  assign y0 = new_n112_ & new_n113_;
  assign new_n115_ = g & b0;
  assign new_n116_ = l0 & new_n115_;
  assign new_n117_ = o0 & ~new_n68_;
  assign new_n118_ = b0 & new_n117_;
  assign new_n119_ = o0 & ~new_n82_;
  assign new_n120_ = ~new_n118_ & ~new_n119_;
  assign new_n121_ = ~e & n0;
  assign new_n122_ = f & ~new_n120_;
  assign new_n123_ = new_n121_ & new_n122_;
  assign new_n124_ = ~e & h;
  assign new_n125_ = b0 & ~new_n68_;
  assign new_n126_ = new_n124_ & new_n125_;
  assign new_n127_ = ~x0 & new_n126_;
  assign new_n128_ = ~new_n116_ & ~new_n123_;
  assign z0 = new_n127_ | ~new_n128_;
  assign new_n130_ = ~j & ~e0;
  assign new_n131_ = ~e & b0;
  assign new_n132_ = new_n67_ & new_n131_;
  assign new_n133_ = i & j0;
  assign new_n134_ = ~c0 & new_n133_;
  assign new_n135_ = ~b0 & new_n134_;
  assign new_n136_ = new_n130_ & ~new_n132_;
  assign new_n137_ = ~new_n135_ & new_n136_;
  assign new_n138_ = o0 & new_n88_;
  assign new_n139_ = n0 & new_n138_;
  assign a1 = new_n137_ & ~new_n139_;
  assign new_n141_ = ~t & u;
  assign new_n142_ = ~s & new_n141_;
  assign new_n143_ = new_n65_ & new_n142_;
  assign new_n144_ = ~e & o0;
  assign new_n145_ = j0 & k0;
  assign new_n146_ = c0 & ~new_n145_;
  assign new_n147_ = b0 & ~new_n146_;
  assign new_n148_ = new_n82_ & ~new_n147_;
  assign new_n149_ = ~n & new_n144_;
  assign new_n150_ = ~new_n148_ & new_n149_;
  assign new_n151_ = n0 & new_n150_;
  assign d1 = ~new_n143_ & ~new_n151_;
  assign new_n153_ = m & b0;
  assign e1 = new_n112_ & new_n153_;
  assign new_n155_ = w & ~x;
  assign f1 = b & new_n155_;
  assign new_n157_ = x & ~y;
  assign new_n158_ = b & w;
  assign g1 = new_n157_ & new_n158_;
  assign new_n160_ = i & ~c0;
  assign new_n161_ = j0 & new_n160_;
  assign new_n162_ = ~new_n79_ & ~new_n161_;
  assign new_n163_ = new_n130_ & new_n162_;
  assign new_n164_ = i & o0;
  assign new_n165_ = d0 & new_n164_;
  assign new_n166_ = n0 & new_n165_;
  assign j1 = new_n163_ & ~new_n166_;
  assign u0 = ~v0;
  assign c1 = ~d1;
  assign h1 = ~a1;
  assign i1 = a1;
endmodule


