// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:33 2022

module in2  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18,
    \v19.0 , \v19.1 , \v19.2 , \v19.3 , \v19.4 , \v19.5 , \v19.6 , \v19.7 ,
    \v19.8 , \v19.9   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18;
  output \v19.0 , \v19.1 , \v19.2 , \v19.3 , \v19.4 , \v19.5 , \v19.6 ,
    \v19.7 , \v19.8 , \v19.9 ;
  wire new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_;
  assign new_n30_ = v12 & ~v13;
  assign new_n31_ = v12 & ~new_n30_;
  assign new_n32_ = ~v18 & ~new_n31_;
  assign new_n33_ = ~v15 & new_n32_;
  assign new_n34_ = ~v11 & new_n33_;
  assign new_n35_ = v1 & new_n34_;
  assign new_n36_ = v15 & v18;
  assign new_n37_ = ~new_n35_ & ~new_n36_;
  assign new_n38_ = v10 & ~new_n37_;
  assign new_n39_ = v8 & v9;
  assign new_n40_ = v18 & ~new_n39_;
  assign new_n41_ = v15 & new_n40_;
  assign new_n42_ = ~v10 & new_n41_;
  assign new_n43_ = ~v7 & new_n42_;
  assign new_n44_ = ~v6 & new_n43_;
  assign new_n45_ = ~v2 & new_n44_;
  assign new_n46_ = ~new_n38_ & ~new_n45_;
  assign new_n47_ = ~v17 & ~new_n46_;
  assign new_n48_ = v9 & ~v18;
  assign new_n49_ = ~v8 & ~new_n48_;
  assign new_n50_ = ~v9 & v18;
  assign new_n51_ = ~new_n49_ & ~new_n50_;
  assign new_n52_ = v7 & ~new_n51_;
  assign new_n53_ = v8 & ~v18;
  assign new_n54_ = ~v7 & new_n53_;
  assign new_n55_ = ~new_n52_ & ~new_n54_;
  assign new_n56_ = ~v10 & ~new_n55_;
  assign new_n57_ = ~v6 & new_n56_;
  assign new_n58_ = ~v2 & new_n57_;
  assign new_n59_ = v10 & ~v18;
  assign new_n60_ = ~new_n58_ & ~new_n59_;
  assign new_n61_ = v17 & ~new_n60_;
  assign new_n62_ = v15 & new_n61_;
  assign new_n63_ = ~new_n47_ & ~new_n62_;
  assign new_n64_ = ~v16 & ~new_n63_;
  assign new_n65_ = ~v7 & v17;
  assign new_n66_ = v6 & new_n65_;
  assign new_n67_ = v7 & ~v17;
  assign new_n68_ = ~v6 & new_n67_;
  assign new_n69_ = ~new_n66_ & ~new_n68_;
  assign new_n70_ = ~v18 & ~new_n69_;
  assign new_n71_ = v8 & new_n70_;
  assign new_n72_ = v7 & v17;
  assign new_n73_ = ~v7 & ~v17;
  assign new_n74_ = ~new_n72_ & ~new_n73_;
  assign new_n75_ = ~new_n51_ & ~new_n74_;
  assign new_n76_ = v6 & new_n75_;
  assign new_n77_ = ~new_n71_ & ~new_n76_;
  assign new_n78_ = v16 & ~new_n77_;
  assign new_n79_ = v15 & new_n78_;
  assign new_n80_ = ~v10 & new_n79_;
  assign new_n81_ = ~v2 & new_n80_;
  assign new_n82_ = ~new_n64_ & ~new_n81_;
  assign new_n83_ = ~v14 & ~new_n82_;
  assign new_n84_ = ~v17 & v18;
  assign new_n85_ = ~v8 & new_n84_;
  assign new_n86_ = v17 & ~v18;
  assign new_n87_ = v8 & new_n86_;
  assign new_n88_ = ~new_n85_ & ~new_n87_;
  assign new_n89_ = ~v7 & ~new_n88_;
  assign new_n90_ = v7 & ~v8;
  assign new_n91_ = v17 & v18;
  assign new_n92_ = new_n90_ & new_n91_;
  assign new_n93_ = ~new_n89_ & ~new_n92_;
  assign new_n94_ = v6 & v16;
  assign new_n95_ = ~v6 & ~v16;
  assign new_n96_ = ~new_n94_ & ~new_n95_;
  assign new_n97_ = ~new_n93_ & ~new_n96_;
  assign new_n98_ = v7 & v8;
  assign new_n99_ = ~v6 & new_n98_;
  assign new_n100_ = ~v17 & ~v18;
  assign new_n101_ = v16 & new_n100_;
  assign new_n102_ = new_n99_ & new_n101_;
  assign new_n103_ = ~new_n97_ & ~new_n102_;
  assign new_n104_ = ~v15 & ~new_n103_;
  assign new_n105_ = v14 & new_n104_;
  assign new_n106_ = ~new_n83_ & ~new_n105_;
  assign \v19.0  = ~v0 & ~new_n106_;
  assign new_n108_ = ~v16 & v17;
  assign new_n109_ = ~v7 & new_n108_;
  assign new_n110_ = v16 & ~v17;
  assign new_n111_ = v7 & new_n110_;
  assign new_n112_ = ~new_n109_ & ~new_n111_;
  assign new_n113_ = ~v18 & ~new_n112_;
  assign new_n114_ = v8 & new_n113_;
  assign new_n115_ = ~new_n39_ & ~new_n74_;
  assign new_n116_ = v18 & new_n115_;
  assign new_n117_ = ~v9 & v17;
  assign new_n118_ = new_n90_ & new_n117_;
  assign new_n119_ = ~new_n116_ & ~new_n118_;
  assign new_n120_ = ~v16 & ~new_n119_;
  assign new_n121_ = ~new_n114_ & ~new_n120_;
  assign new_n122_ = ~v6 & ~new_n121_;
  assign new_n123_ = ~v7 & v8;
  assign new_n124_ = new_n86_ & new_n123_;
  assign new_n125_ = ~new_n75_ & ~new_n124_;
  assign new_n126_ = v16 & ~new_n125_;
  assign new_n127_ = v6 & new_n126_;
  assign new_n128_ = ~new_n122_ & ~new_n127_;
  assign new_n129_ = ~v10 & ~new_n128_;
  assign new_n130_ = ~v2 & new_n129_;
  assign new_n131_ = ~v0 & new_n130_;
  assign new_n132_ = ~v16 & new_n100_;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign new_n134_ = v15 & ~new_n133_;
  assign new_n135_ = ~v14 & new_n134_;
  assign \v19.1  = v0 | new_n135_;
  assign new_n137_ = v3 & v9;
  assign new_n138_ = v4 & ~v9;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = ~new_n96_ & ~new_n139_;
  assign new_n141_ = ~new_n93_ & new_n140_;
  assign new_n142_ = v8 & v18;
  assign new_n143_ = ~v8 & ~v18;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = v16 & ~new_n74_;
  assign new_n146_ = v6 & new_n145_;
  assign new_n147_ = ~v6 & v7;
  assign new_n148_ = new_n108_ & new_n147_;
  assign new_n149_ = ~new_n146_ & ~new_n148_;
  assign new_n150_ = ~new_n144_ & ~new_n149_;
  assign new_n151_ = ~v6 & new_n123_;
  assign new_n152_ = ~v16 & new_n84_;
  assign new_n153_ = new_n151_ & new_n152_;
  assign new_n154_ = ~new_n150_ & ~new_n153_;
  assign new_n155_ = ~v9 & ~new_n154_;
  assign new_n156_ = v9 & v16;
  assign new_n157_ = new_n100_ & new_n156_;
  assign new_n158_ = new_n99_ & new_n157_;
  assign new_n159_ = ~new_n155_ & ~new_n158_;
  assign new_n160_ = v3 & ~new_n159_;
  assign new_n161_ = v4 & new_n147_;
  assign new_n162_ = ~v9 & v16;
  assign new_n163_ = v8 & new_n162_;
  assign new_n164_ = new_n161_ & new_n163_;
  assign new_n165_ = v1 & ~v3;
  assign new_n166_ = ~v10 & ~v16;
  assign new_n167_ = new_n165_ & new_n166_;
  assign new_n168_ = ~new_n164_ & ~new_n167_;
  assign new_n169_ = ~v18 & ~new_n168_;
  assign new_n170_ = ~v17 & new_n169_;
  assign new_n171_ = ~new_n160_ & ~new_n170_;
  assign new_n172_ = ~new_n141_ & new_n171_;
  assign new_n173_ = ~v15 & ~new_n172_;
  assign new_n174_ = ~v14 & new_n173_;
  assign \v19.2  = ~v0 & new_n174_;
  assign new_n176_ = ~v18 & ~new_n100_;
  assign new_n177_ = v16 & ~new_n176_;
  assign new_n178_ = v5 & ~v10;
  assign new_n179_ = v1 & new_n178_;
  assign new_n180_ = ~new_n152_ & ~new_n179_;
  assign new_n181_ = ~v17 & new_n180_;
  assign new_n182_ = ~new_n177_ & new_n181_;
  assign new_n183_ = v3 & ~new_n182_;
  assign new_n184_ = v4 & ~v5;
  assign new_n185_ = ~v2 & ~new_n184_;
  assign new_n186_ = ~v18 & ~new_n185_;
  assign new_n187_ = ~v17 & new_n186_;
  assign new_n188_ = ~v16 & new_n187_;
  assign new_n189_ = ~v10 & new_n188_;
  assign new_n190_ = v1 & new_n189_;
  assign new_n191_ = ~new_n183_ & ~new_n190_;
  assign new_n192_ = ~v15 & ~new_n191_;
  assign new_n193_ = ~v14 & new_n192_;
  assign \v19.3  = ~v0 & new_n193_;
  assign new_n195_ = ~v14 & v15;
  assign new_n196_ = v14 & ~v15;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = ~v6 & ~v7;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = ~v7 & ~v8;
  assign new_n201_ = ~v6 & new_n200_;
  assign new_n202_ = v4 & new_n201_;
  assign new_n203_ = ~v3 & ~new_n202_;
  assign new_n204_ = ~v15 & ~new_n203_;
  assign new_n205_ = ~v10 & ~new_n39_;
  assign new_n206_ = ~v2 & new_n205_;
  assign new_n207_ = v15 & ~new_n206_;
  assign new_n208_ = ~new_n204_ & ~new_n207_;
  assign new_n209_ = ~v14 & ~new_n208_;
  assign new_n210_ = v4 & ~v6;
  assign new_n211_ = ~v7 & ~v9;
  assign new_n212_ = new_n210_ & new_n211_;
  assign new_n213_ = ~v14 & ~new_n212_;
  assign new_n214_ = ~v15 & ~new_n213_;
  assign new_n215_ = v8 & new_n214_;
  assign new_n216_ = ~new_n209_ & ~new_n215_;
  assign new_n217_ = ~new_n199_ & new_n216_;
  assign new_n218_ = v18 & ~new_n217_;
  assign new_n219_ = ~v5 & ~v10;
  assign new_n220_ = v3 & new_n219_;
  assign new_n221_ = ~v18 & ~new_n220_;
  assign new_n222_ = ~v15 & new_n221_;
  assign new_n223_ = ~v14 & new_n222_;
  assign new_n224_ = ~v12 & new_n223_;
  assign new_n225_ = ~v11 & new_n224_;
  assign new_n226_ = v1 & new_n225_;
  assign new_n227_ = ~new_n218_ & ~new_n226_;
  assign new_n228_ = ~v17 & ~new_n227_;
  assign new_n229_ = ~v16 & new_n228_;
  assign \v19.4  = ~v0 & new_n229_;
  assign new_n231_ = v8 & ~v9;
  assign new_n232_ = v9 & ~v14;
  assign new_n233_ = ~v8 & new_n232_;
  assign new_n234_ = ~new_n231_ & ~new_n233_;
  assign new_n235_ = ~v7 & ~new_n234_;
  assign new_n236_ = ~v6 & new_n235_;
  assign new_n237_ = v4 & new_n236_;
  assign new_n238_ = v14 & ~new_n201_;
  assign new_n239_ = ~new_n237_ & ~new_n238_;
  assign new_n240_ = v18 & ~new_n239_;
  assign new_n241_ = ~v12 & v13;
  assign new_n242_ = v13 & ~new_n241_;
  assign new_n243_ = v11 & ~new_n242_;
  assign new_n244_ = ~v11 & v13;
  assign new_n245_ = v13 & ~new_n244_;
  assign new_n246_ = v12 & ~new_n245_;
  assign new_n247_ = ~new_n243_ & ~new_n246_;
  assign new_n248_ = ~v18 & ~new_n247_;
  assign new_n249_ = ~v14 & new_n248_;
  assign new_n250_ = ~v10 & new_n249_;
  assign new_n251_ = ~v5 & new_n250_;
  assign new_n252_ = v3 & new_n251_;
  assign new_n253_ = v1 & new_n252_;
  assign new_n254_ = ~new_n240_ & ~new_n253_;
  assign new_n255_ = ~v16 & ~new_n254_;
  assign new_n256_ = v14 & v18;
  assign new_n257_ = ~v6 & v8;
  assign new_n258_ = v4 & new_n257_;
  assign new_n259_ = ~v14 & ~v18;
  assign new_n260_ = v9 & new_n259_;
  assign new_n261_ = new_n258_ & new_n260_;
  assign new_n262_ = ~new_n256_ & ~new_n261_;
  assign new_n263_ = v7 & ~new_n262_;
  assign new_n264_ = ~v14 & v18;
  assign new_n265_ = v9 & new_n264_;
  assign new_n266_ = ~v9 & ~v18;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign new_n268_ = ~v8 & ~new_n267_;
  assign new_n269_ = v8 & new_n50_;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = ~v7 & ~new_n270_;
  assign new_n272_ = v4 & new_n271_;
  assign new_n273_ = v14 & ~v18;
  assign new_n274_ = ~new_n272_ & ~new_n273_;
  assign new_n275_ = v6 & ~new_n274_;
  assign new_n276_ = ~v18 & ~new_n98_;
  assign new_n277_ = v14 & new_n276_;
  assign new_n278_ = ~new_n275_ & ~new_n277_;
  assign new_n279_ = ~new_n263_ & new_n278_;
  assign new_n280_ = v16 & ~new_n279_;
  assign new_n281_ = ~new_n255_ & ~new_n280_;
  assign new_n282_ = ~v17 & ~new_n281_;
  assign new_n283_ = v7 & new_n50_;
  assign new_n284_ = ~v7 & v9;
  assign new_n285_ = new_n259_ & new_n284_;
  assign new_n286_ = ~new_n283_ & ~new_n285_;
  assign new_n287_ = v8 & ~new_n286_;
  assign new_n288_ = v7 & new_n268_;
  assign new_n289_ = ~new_n287_ & ~new_n288_;
  assign new_n290_ = ~new_n96_ & ~new_n289_;
  assign new_n291_ = v4 & new_n290_;
  assign new_n292_ = v6 & ~v16;
  assign new_n293_ = v18 & ~new_n90_;
  assign new_n294_ = ~v6 & v16;
  assign new_n295_ = v8 & ~new_n294_;
  assign new_n296_ = ~v7 & new_n295_;
  assign new_n297_ = ~v18 & ~new_n296_;
  assign new_n298_ = ~new_n293_ & ~new_n297_;
  assign new_n299_ = ~new_n292_ & new_n298_;
  assign new_n300_ = v14 & ~new_n299_;
  assign new_n301_ = ~new_n291_ & ~new_n300_;
  assign new_n302_ = v17 & ~new_n301_;
  assign new_n303_ = v6 & ~v8;
  assign new_n304_ = v18 & ~new_n303_;
  assign new_n305_ = v16 & new_n304_;
  assign new_n306_ = v14 & new_n305_;
  assign new_n307_ = ~new_n302_ & ~new_n306_;
  assign new_n308_ = ~new_n282_ & new_n307_;
  assign new_n309_ = ~v15 & ~new_n308_;
  assign \v19.5  = ~v0 & new_n309_;
  assign new_n311_ = ~v17 & ~new_n152_;
  assign new_n312_ = ~new_n177_ & new_n311_;
  assign new_n313_ = ~v2 & ~v10;
  assign new_n314_ = v15 & ~new_n313_;
  assign new_n315_ = v3 & ~v15;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = ~new_n312_ & ~new_n316_;
  assign new_n318_ = ~new_n108_ & ~new_n111_;
  assign new_n319_ = v6 & ~new_n318_;
  assign new_n320_ = ~v8 & ~v17;
  assign new_n321_ = ~v17 & ~new_n320_;
  assign new_n322_ = ~v6 & ~new_n321_;
  assign new_n323_ = ~v8 & v9;
  assign new_n324_ = ~new_n123_ & ~new_n323_;
  assign new_n325_ = ~v17 & ~new_n324_;
  assign new_n326_ = ~new_n322_ & ~new_n325_;
  assign new_n327_ = v16 & ~new_n326_;
  assign new_n328_ = v7 & ~v9;
  assign new_n329_ = ~v8 & ~new_n328_;
  assign new_n330_ = ~new_n98_ & ~new_n329_;
  assign new_n331_ = v17 & ~new_n330_;
  assign new_n332_ = ~new_n327_ & ~new_n331_;
  assign new_n333_ = ~new_n319_ & new_n332_;
  assign new_n334_ = v15 & ~new_n333_;
  assign new_n335_ = ~v6 & ~new_n112_;
  assign new_n336_ = v6 & ~v7;
  assign new_n337_ = v16 & v17;
  assign new_n338_ = new_n336_ & new_n337_;
  assign new_n339_ = ~new_n335_ & ~new_n338_;
  assign new_n340_ = ~v9 & ~new_n339_;
  assign new_n341_ = v8 & new_n340_;
  assign new_n342_ = v4 & new_n341_;
  assign new_n343_ = v12 & v13;
  assign new_n344_ = v12 & ~new_n343_;
  assign new_n345_ = ~v11 & ~new_n344_;
  assign new_n346_ = ~new_n243_ & ~new_n345_;
  assign new_n347_ = ~new_n220_ & ~new_n346_;
  assign new_n348_ = ~v11 & ~new_n219_;
  assign new_n349_ = v3 & ~new_n348_;
  assign new_n350_ = ~v13 & ~new_n349_;
  assign new_n351_ = v12 & new_n350_;
  assign new_n352_ = ~new_n347_ & ~new_n351_;
  assign new_n353_ = ~v17 & ~new_n352_;
  assign new_n354_ = ~v16 & new_n353_;
  assign new_n355_ = v1 & new_n354_;
  assign new_n356_ = ~new_n342_ & ~new_n355_;
  assign new_n357_ = ~v15 & ~new_n356_;
  assign new_n358_ = ~new_n334_ & ~new_n357_;
  assign new_n359_ = ~v18 & ~new_n358_;
  assign new_n360_ = ~new_n74_ & ~new_n96_;
  assign new_n361_ = ~v15 & new_n360_;
  assign new_n362_ = ~v9 & new_n361_;
  assign new_n363_ = ~v8 & new_n362_;
  assign new_n364_ = v4 & new_n363_;
  assign new_n365_ = ~v7 & ~new_n39_;
  assign new_n366_ = ~v17 & ~new_n365_;
  assign new_n367_ = ~v6 & ~new_n366_;
  assign new_n368_ = ~v16 & ~new_n367_;
  assign new_n369_ = ~v16 & ~v17;
  assign new_n370_ = v9 & ~new_n369_;
  assign new_n371_ = v8 & new_n370_;
  assign new_n372_ = v6 & ~new_n67_;
  assign new_n373_ = v16 & ~new_n372_;
  assign new_n374_ = ~new_n65_ & ~new_n373_;
  assign new_n375_ = ~new_n371_ & new_n374_;
  assign new_n376_ = ~new_n368_ & new_n375_;
  assign new_n377_ = v15 & ~new_n376_;
  assign new_n378_ = ~new_n364_ & ~new_n377_;
  assign new_n379_ = v18 & ~new_n378_;
  assign new_n380_ = ~new_n359_ & ~new_n379_;
  assign new_n381_ = ~new_n317_ & new_n380_;
  assign new_n382_ = ~v14 & ~new_n381_;
  assign \v19.6  = ~v0 & new_n382_;
  assign new_n384_ = v16 & v18;
  assign new_n385_ = ~v10 & v11;
  assign new_n386_ = v1 & ~v5;
  assign new_n387_ = new_n385_ & new_n386_;
  assign new_n388_ = new_n132_ & new_n241_;
  assign new_n389_ = new_n387_ & new_n388_;
  assign new_n390_ = ~new_n384_ & ~new_n389_;
  assign new_n391_ = v3 & ~new_n390_;
  assign new_n392_ = v16 & ~new_n93_;
  assign new_n393_ = v6 & new_n392_;
  assign new_n394_ = v4 & new_n393_;
  assign new_n395_ = v13 & ~new_n220_;
  assign new_n396_ = ~v12 & new_n395_;
  assign new_n397_ = ~new_n30_ & ~new_n396_;
  assign new_n398_ = ~v18 & ~new_n397_;
  assign new_n399_ = ~v17 & new_n398_;
  assign new_n400_ = ~v16 & new_n399_;
  assign new_n401_ = v11 & new_n400_;
  assign new_n402_ = v1 & new_n401_;
  assign new_n403_ = ~new_n394_ & ~new_n402_;
  assign new_n404_ = ~new_n391_ & new_n403_;
  assign new_n405_ = ~v15 & ~new_n404_;
  assign new_n406_ = ~v2 & new_n98_;
  assign new_n407_ = ~v10 & new_n100_;
  assign new_n408_ = new_n406_ & new_n407_;
  assign new_n409_ = ~v18 & ~new_n408_;
  assign new_n410_ = ~v6 & ~new_n409_;
  assign new_n411_ = ~v10 & ~new_n51_;
  assign new_n412_ = ~v7 & new_n411_;
  assign new_n413_ = v6 & new_n412_;
  assign new_n414_ = ~v2 & new_n413_;
  assign new_n415_ = v7 & v18;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = ~v17 & ~new_n416_;
  assign new_n418_ = v18 & ~new_n206_;
  assign new_n419_ = ~v17 & ~new_n418_;
  assign new_n420_ = ~new_n417_ & new_n419_;
  assign new_n421_ = ~new_n410_ & new_n420_;
  assign new_n422_ = v16 & ~new_n421_;
  assign new_n423_ = v15 & new_n422_;
  assign new_n424_ = ~new_n405_ & ~new_n423_;
  assign new_n425_ = ~v14 & ~new_n424_;
  assign new_n426_ = new_n98_ & new_n100_;
  assign new_n427_ = ~v18 & ~new_n426_;
  assign new_n428_ = ~v6 & ~new_n427_;
  assign new_n429_ = v6 & new_n200_;
  assign new_n430_ = ~v7 & ~new_n429_;
  assign new_n431_ = ~v17 & ~new_n430_;
  assign new_n432_ = ~v8 & ~new_n431_;
  assign new_n433_ = v18 & ~new_n432_;
  assign new_n434_ = ~v17 & ~new_n433_;
  assign new_n435_ = ~new_n428_ & new_n434_;
  assign new_n436_ = v14 & ~new_n435_;
  assign new_n437_ = v17 & ~new_n144_;
  assign new_n438_ = v7 & new_n437_;
  assign new_n439_ = new_n84_ & new_n123_;
  assign new_n440_ = ~new_n438_ & ~new_n439_;
  assign new_n441_ = ~v9 & ~new_n440_;
  assign new_n442_ = v6 & new_n441_;
  assign new_n443_ = v4 & new_n442_;
  assign new_n444_ = v3 & v17;
  assign new_n445_ = ~new_n443_ & ~new_n444_;
  assign new_n446_ = ~new_n436_ & new_n445_;
  assign new_n447_ = v16 & ~new_n446_;
  assign new_n448_ = ~v15 & new_n447_;
  assign new_n449_ = ~new_n425_ & ~new_n448_;
  assign \v19.7  = ~v0 & ~new_n449_;
  assign new_n451_ = v17 & ~new_n96_;
  assign new_n452_ = ~v10 & new_n451_;
  assign new_n453_ = ~v2 & new_n452_;
  assign new_n454_ = ~new_n110_ & ~new_n453_;
  assign new_n455_ = v8 & ~new_n454_;
  assign new_n456_ = ~v7 & new_n455_;
  assign new_n457_ = v6 & ~v9;
  assign new_n458_ = ~v8 & ~new_n457_;
  assign new_n459_ = v6 & v7;
  assign new_n460_ = ~v10 & ~new_n459_;
  assign new_n461_ = ~v2 & new_n460_;
  assign new_n462_ = ~new_n458_ & new_n461_;
  assign new_n463_ = ~v17 & ~new_n462_;
  assign new_n464_ = v16 & new_n463_;
  assign new_n465_ = ~new_n456_ & ~new_n464_;
  assign new_n466_ = v15 & ~new_n465_;
  assign new_n467_ = ~v11 & new_n343_;
  assign new_n468_ = v11 & ~v13;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_ = v3 & ~v5;
  assign new_n471_ = ~v10 & ~new_n220_;
  assign new_n472_ = new_n470_ & new_n471_;
  assign new_n473_ = ~new_n469_ & ~new_n472_;
  assign new_n474_ = ~v16 & new_n473_;
  assign new_n475_ = v1 & new_n474_;
  assign new_n476_ = v4 & new_n99_;
  assign new_n477_ = ~v3 & ~new_n476_;
  assign new_n478_ = v16 & ~new_n477_;
  assign new_n479_ = ~new_n475_ & ~new_n478_;
  assign new_n480_ = ~v17 & ~new_n479_;
  assign new_n481_ = ~v15 & new_n480_;
  assign new_n482_ = ~new_n466_ & ~new_n481_;
  assign new_n483_ = ~v18 & ~new_n482_;
  assign new_n484_ = ~v15 & v18;
  assign new_n485_ = v4 & new_n484_;
  assign new_n486_ = ~v2 & ~v9;
  assign new_n487_ = ~v10 & v15;
  assign new_n488_ = new_n486_ & new_n487_;
  assign new_n489_ = ~new_n485_ & ~new_n488_;
  assign new_n490_ = ~new_n96_ & ~new_n489_;
  assign new_n491_ = ~v8 & new_n490_;
  assign new_n492_ = v7 & new_n491_;
  assign new_n493_ = ~v15 & ~new_n315_;
  assign new_n494_ = v18 & ~new_n493_;
  assign new_n495_ = ~new_n492_ & ~new_n494_;
  assign new_n496_ = v17 & ~new_n495_;
  assign new_n497_ = ~new_n483_ & ~new_n496_;
  assign new_n498_ = ~v14 & ~new_n497_;
  assign new_n499_ = v4 & v7;
  assign new_n500_ = new_n50_ & new_n499_;
  assign new_n501_ = ~v7 & new_n273_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~new_n96_ & ~new_n502_;
  assign new_n504_ = v8 & new_n503_;
  assign new_n505_ = ~new_n256_ & ~new_n504_;
  assign new_n506_ = v17 & ~new_n505_;
  assign new_n507_ = v4 & ~v7;
  assign new_n508_ = ~v8 & ~v9;
  assign new_n509_ = new_n507_ & new_n508_;
  assign new_n510_ = ~v14 & ~new_n509_;
  assign new_n511_ = v6 & ~new_n510_;
  assign new_n512_ = v14 & ~new_n98_;
  assign new_n513_ = ~new_n511_ & ~new_n512_;
  assign new_n514_ = ~v18 & ~new_n513_;
  assign new_n515_ = ~v17 & new_n514_;
  assign new_n516_ = v16 & new_n515_;
  assign new_n517_ = ~new_n506_ & ~new_n516_;
  assign new_n518_ = ~v15 & ~new_n517_;
  assign new_n519_ = ~new_n498_ & ~new_n518_;
  assign \v19.8  = ~v0 & ~new_n519_;
  assign new_n521_ = ~v17 & ~new_n110_;
  assign new_n522_ = v9 & new_n195_;
  assign new_n523_ = ~new_n196_ & ~new_n522_;
  assign new_n524_ = ~v8 & ~new_n523_;
  assign new_n525_ = ~v14 & ~new_n316_;
  assign new_n526_ = ~new_n524_ & ~new_n525_;
  assign new_n527_ = ~new_n521_ & ~new_n526_;
  assign new_n528_ = ~v11 & ~v12;
  assign new_n529_ = v3 & ~new_n220_;
  assign new_n530_ = ~new_n528_ & ~new_n529_;
  assign new_n531_ = ~v11 & v12;
  assign new_n532_ = ~v11 & ~new_n531_;
  assign new_n533_ = ~new_n219_ & ~new_n532_;
  assign new_n534_ = ~new_n530_ & ~new_n533_;
  assign new_n535_ = ~v17 & ~new_n534_;
  assign new_n536_ = ~v13 & new_n535_;
  assign new_n537_ = v1 & new_n536_;
  assign new_n538_ = v8 & v17;
  assign new_n539_ = ~v7 & new_n538_;
  assign new_n540_ = ~v6 & new_n539_;
  assign new_n541_ = v4 & new_n540_;
  assign new_n542_ = ~new_n537_ & ~new_n541_;
  assign new_n543_ = ~v16 & ~new_n542_;
  assign new_n544_ = v16 & ~new_n69_;
  assign new_n545_ = v8 & new_n544_;
  assign new_n546_ = v4 & new_n545_;
  assign new_n547_ = ~new_n543_ & ~new_n546_;
  assign new_n548_ = ~v14 & ~new_n547_;
  assign new_n549_ = ~v9 & ~new_n96_;
  assign new_n550_ = ~v8 & new_n549_;
  assign new_n551_ = v4 & new_n550_;
  assign new_n552_ = ~v14 & ~new_n551_;
  assign new_n553_ = v7 & ~new_n552_;
  assign new_n554_ = ~new_n292_ & ~new_n294_;
  assign new_n555_ = v14 & ~new_n554_;
  assign new_n556_ = ~new_n553_ & ~new_n555_;
  assign new_n557_ = v17 & ~new_n556_;
  assign new_n558_ = ~v7 & v14;
  assign new_n559_ = ~new_n511_ & ~new_n558_;
  assign new_n560_ = ~v17 & ~new_n559_;
  assign new_n561_ = v16 & new_n560_;
  assign new_n562_ = ~new_n557_ & ~new_n561_;
  assign new_n563_ = ~new_n548_ & new_n562_;
  assign new_n564_ = ~v15 & ~new_n563_;
  assign new_n565_ = v8 & ~v17;
  assign new_n566_ = ~v7 & new_n565_;
  assign new_n567_ = ~new_n322_ & ~new_n566_;
  assign new_n568_ = v16 & ~new_n567_;
  assign new_n569_ = ~new_n98_ & ~new_n200_;
  assign new_n570_ = v17 & ~new_n569_;
  assign new_n571_ = ~new_n568_ & ~new_n570_;
  assign new_n572_ = ~new_n319_ & new_n571_;
  assign new_n573_ = v15 & ~new_n572_;
  assign new_n574_ = ~v14 & new_n573_;
  assign new_n575_ = ~new_n564_ & ~new_n574_;
  assign new_n576_ = ~new_n527_ & new_n575_;
  assign new_n577_ = ~v18 & ~new_n576_;
  assign new_n578_ = v15 & ~new_n39_;
  assign new_n579_ = ~v14 & new_n578_;
  assign new_n580_ = ~v10 & new_n579_;
  assign new_n581_ = ~v2 & new_n580_;
  assign new_n582_ = ~v8 & new_n196_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = ~new_n96_ & ~new_n583_;
  assign new_n585_ = ~new_n74_ & new_n584_;
  assign new_n586_ = v18 & new_n585_;
  assign new_n587_ = ~new_n577_ & ~new_n586_;
  assign \v19.9  = ~v0 & ~new_n587_;
endmodule


