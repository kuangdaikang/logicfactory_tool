// Benchmark "sqrt" written by ABC on Fri Sep 15 11:24:10 2023

module sqrt ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] ,
    \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] , \asqrt[5] ,
    \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] , \asqrt[10] ,
    \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] , \asqrt[15] ,
    \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] , \asqrt[20] ,
    \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] , \asqrt[25] ,
    \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] , \asqrt[30] ,
    \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] , \asqrt[35] ,
    \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] , \asqrt[40] ,
    \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] , \asqrt[45] ,
    \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] , \asqrt[50] ,
    \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] , \asqrt[55] ,
    \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] , \asqrt[60] ,
    \asqrt[61] , \asqrt[62] , \asqrt[63]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] ;
  output \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] ,
    \asqrt[5] , \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] ,
    \asqrt[10] , \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] ,
    \asqrt[15] , \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] ,
    \asqrt[20] , \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] ,
    \asqrt[25] , \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] ,
    \asqrt[30] , \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] ,
    \asqrt[35] , \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] ,
    \asqrt[40] , \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] ,
    \asqrt[45] , \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] ,
    \asqrt[50] , \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] ,
    \asqrt[55] , \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] ,
    \asqrt[60] , \asqrt[61] , \asqrt[62] , \asqrt[63] ;
  wire new_n193_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_,
    new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_,
    new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_,
    new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_,
    new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_,
    new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_,
    new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_,
    new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_,
    new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_,
    new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_,
    new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_,
    new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_,
    new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_,
    new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_,
    new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_,
    new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_,
    new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_,
    new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_,
    new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_,
    new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_,
    new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_,
    new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_,
    new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_,
    new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_,
    new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_,
    new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_,
    new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_,
    new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_,
    new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_,
    new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_,
    new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_,
    new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_,
    new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_,
    new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_,
    new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_,
    new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_,
    new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_,
    new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_,
    new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_,
    new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_,
    new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_,
    new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_,
    new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_,
    new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_,
    new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_,
    new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_,
    new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_,
    new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_,
    new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_,
    new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_,
    new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_,
    new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_,
    new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_,
    new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_,
    new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_,
    new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_,
    new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_,
    new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_,
    new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_,
    new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_,
    new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_,
    new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_,
    new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_,
    new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_,
    new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_,
    new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_,
    new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_,
    new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_,
    new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_,
    new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_,
    new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_,
    new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_,
    new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_,
    new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_,
    new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_,
    new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_,
    new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_,
    new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5419_, new_n5420_,
    new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_,
    new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_,
    new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_,
    new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_,
    new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_,
    new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_,
    new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_,
    new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_,
    new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_,
    new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_,
    new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_,
    new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_,
    new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_,
    new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_,
    new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_,
    new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_,
    new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_,
    new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_,
    new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_,
    new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_,
    new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_,
    new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_,
    new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_,
    new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_,
    new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_,
    new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_,
    new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_,
    new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_,
    new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_,
    new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_,
    new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_,
    new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_,
    new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_,
    new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_,
    new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_,
    new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_,
    new_n5763_, new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_,
    new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_,
    new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_,
    new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_,
    new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_,
    new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_,
    new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_,
    new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_,
    new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_,
    new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_,
    new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_,
    new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_,
    new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_,
    new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_,
    new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_,
    new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_,
    new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_,
    new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_,
    new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_,
    new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_,
    new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_,
    new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_,
    new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_,
    new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6087_, new_n6088_,
    new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_,
    new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_,
    new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_,
    new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_,
    new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_,
    new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_,
    new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_,
    new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_,
    new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_,
    new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_,
    new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_,
    new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_,
    new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_,
    new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_,
    new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_,
    new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_,
    new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_,
    new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_,
    new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_,
    new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_,
    new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_,
    new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_,
    new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_,
    new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_,
    new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_,
    new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_,
    new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_,
    new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6434_, new_n6435_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_,
    new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_,
    new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_,
    new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_,
    new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_,
    new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_,
    new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_,
    new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_,
    new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_,
    new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_,
    new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_,
    new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_,
    new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_,
    new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_,
    new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_,
    new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_,
    new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_,
    new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_,
    new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_,
    new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_,
    new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_,
    new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_,
    new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_,
    new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_,
    new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_,
    new_n7947_, new_n7948_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_,
    new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_,
    new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_,
    new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_,
    new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_,
    new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_,
    new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_,
    new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_,
    new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_,
    new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_,
    new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_,
    new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_,
    new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_,
    new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_,
    new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_,
    new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_,
    new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_,
    new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_,
    new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_,
    new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_,
    new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_,
    new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_,
    new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_,
    new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_,
    new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_,
    new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_,
    new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_,
    new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_,
    new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_,
    new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_,
    new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_,
    new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_,
    new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_,
    new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_,
    new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_,
    new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_,
    new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_,
    new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_,
    new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_,
    new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_,
    new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_,
    new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_,
    new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_,
    new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_,
    new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_,
    new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_,
    new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_,
    new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_,
    new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_,
    new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_,
    new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_,
    new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_,
    new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_,
    new_n9156_, new_n9157_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_,
    new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_,
    new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_,
    new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_,
    new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_,
    new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_,
    new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_,
    new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_,
    new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_,
    new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_,
    new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_,
    new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_,
    new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_,
    new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_,
    new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_,
    new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_,
    new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_,
    new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_,
    new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_,
    new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_,
    new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_,
    new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_,
    new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_,
    new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_,
    new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_,
    new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_,
    new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10027_, new_n10028_,
    new_n10029_, new_n10030_, new_n10031_, new_n10032_, new_n10033_,
    new_n10034_, new_n10035_, new_n10036_, new_n10037_, new_n10038_,
    new_n10039_, new_n10040_, new_n10041_, new_n10042_, new_n10043_,
    new_n10044_, new_n10045_, new_n10046_, new_n10047_, new_n10048_,
    new_n10049_, new_n10050_, new_n10051_, new_n10052_, new_n10053_,
    new_n10054_, new_n10055_, new_n10056_, new_n10057_, new_n10058_,
    new_n10059_, new_n10060_, new_n10061_, new_n10062_, new_n10063_,
    new_n10064_, new_n10065_, new_n10066_, new_n10067_, new_n10068_,
    new_n10069_, new_n10070_, new_n10071_, new_n10072_, new_n10073_,
    new_n10074_, new_n10075_, new_n10076_, new_n10077_, new_n10078_,
    new_n10079_, new_n10080_, new_n10081_, new_n10082_, new_n10083_,
    new_n10084_, new_n10085_, new_n10086_, new_n10087_, new_n10088_,
    new_n10089_, new_n10090_, new_n10091_, new_n10092_, new_n10093_,
    new_n10094_, new_n10095_, new_n10096_, new_n10097_, new_n10098_,
    new_n10099_, new_n10100_, new_n10101_, new_n10102_, new_n10103_,
    new_n10104_, new_n10105_, new_n10106_, new_n10107_, new_n10108_,
    new_n10109_, new_n10110_, new_n10111_, new_n10112_, new_n10113_,
    new_n10114_, new_n10115_, new_n10116_, new_n10117_, new_n10118_,
    new_n10119_, new_n10120_, new_n10121_, new_n10122_, new_n10123_,
    new_n10124_, new_n10125_, new_n10126_, new_n10127_, new_n10128_,
    new_n10129_, new_n10130_, new_n10131_, new_n10132_, new_n10133_,
    new_n10134_, new_n10135_, new_n10136_, new_n10137_, new_n10138_,
    new_n10139_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10146_, new_n10147_, new_n10148_,
    new_n10149_, new_n10150_, new_n10151_, new_n10152_, new_n10153_,
    new_n10154_, new_n10155_, new_n10156_, new_n10157_, new_n10158_,
    new_n10159_, new_n10160_, new_n10161_, new_n10162_, new_n10163_,
    new_n10164_, new_n10165_, new_n10166_, new_n10167_, new_n10168_,
    new_n10169_, new_n10170_, new_n10171_, new_n10172_, new_n10173_,
    new_n10174_, new_n10175_, new_n10176_, new_n10177_, new_n10178_,
    new_n10179_, new_n10180_, new_n10181_, new_n10182_, new_n10183_,
    new_n10184_, new_n10185_, new_n10186_, new_n10187_, new_n10188_,
    new_n10189_, new_n10190_, new_n10191_, new_n10192_, new_n10193_,
    new_n10194_, new_n10195_, new_n10196_, new_n10197_, new_n10198_,
    new_n10199_, new_n10200_, new_n10201_, new_n10202_, new_n10203_,
    new_n10204_, new_n10205_, new_n10206_, new_n10207_, new_n10208_,
    new_n10209_, new_n10210_, new_n10211_, new_n10212_, new_n10213_,
    new_n10214_, new_n10215_, new_n10216_, new_n10217_, new_n10218_,
    new_n10219_, new_n10220_, new_n10221_, new_n10222_, new_n10223_,
    new_n10224_, new_n10225_, new_n10226_, new_n10227_, new_n10228_,
    new_n10229_, new_n10230_, new_n10231_, new_n10232_, new_n10233_,
    new_n10234_, new_n10235_, new_n10236_, new_n10237_, new_n10238_,
    new_n10239_, new_n10240_, new_n10241_, new_n10242_, new_n10243_,
    new_n10244_, new_n10245_, new_n10246_, new_n10247_, new_n10248_,
    new_n10249_, new_n10250_, new_n10251_, new_n10252_, new_n10253_,
    new_n10254_, new_n10255_, new_n10256_, new_n10257_, new_n10258_,
    new_n10259_, new_n10260_, new_n10261_, new_n10262_, new_n10263_,
    new_n10264_, new_n10265_, new_n10266_, new_n10267_, new_n10268_,
    new_n10269_, new_n10270_, new_n10271_, new_n10272_, new_n10273_,
    new_n10274_, new_n10275_, new_n10276_, new_n10277_, new_n10278_,
    new_n10279_, new_n10280_, new_n10281_, new_n10282_, new_n10283_,
    new_n10284_, new_n10285_, new_n10286_, new_n10287_, new_n10288_,
    new_n10289_, new_n10290_, new_n10291_, new_n10292_, new_n10293_,
    new_n10294_, new_n10295_, new_n10296_, new_n10297_, new_n10298_,
    new_n10299_, new_n10300_, new_n10301_, new_n10302_, new_n10303_,
    new_n10304_, new_n10305_, new_n10306_, new_n10307_, new_n10308_,
    new_n10309_, new_n10310_, new_n10311_, new_n10312_, new_n10313_,
    new_n10314_, new_n10315_, new_n10316_, new_n10317_, new_n10318_,
    new_n10319_, new_n10320_, new_n10321_, new_n10322_, new_n10323_,
    new_n10324_, new_n10325_, new_n10326_, new_n10327_, new_n10328_,
    new_n10329_, new_n10330_, new_n10331_, new_n10332_, new_n10333_,
    new_n10334_, new_n10335_, new_n10336_, new_n10337_, new_n10338_,
    new_n10339_, new_n10340_, new_n10341_, new_n10342_, new_n10343_,
    new_n10344_, new_n10345_, new_n10346_, new_n10347_, new_n10348_,
    new_n10349_, new_n10350_, new_n10351_, new_n10352_, new_n10353_,
    new_n10354_, new_n10355_, new_n10356_, new_n10357_, new_n10358_,
    new_n10359_, new_n10360_, new_n10361_, new_n10362_, new_n10363_,
    new_n10364_, new_n10365_, new_n10366_, new_n10367_, new_n10368_,
    new_n10369_, new_n10370_, new_n10371_, new_n10372_, new_n10373_,
    new_n10374_, new_n10375_, new_n10376_, new_n10377_, new_n10378_,
    new_n10379_, new_n10380_, new_n10381_, new_n10382_, new_n10383_,
    new_n10384_, new_n10385_, new_n10386_, new_n10387_, new_n10388_,
    new_n10389_, new_n10390_, new_n10391_, new_n10392_, new_n10393_,
    new_n10394_, new_n10395_, new_n10396_, new_n10397_, new_n10398_,
    new_n10399_, new_n10400_, new_n10401_, new_n10402_, new_n10403_,
    new_n10404_, new_n10405_, new_n10406_, new_n10407_, new_n10408_,
    new_n10409_, new_n10410_, new_n10411_, new_n10412_, new_n10413_,
    new_n10414_, new_n10415_, new_n10416_, new_n10417_, new_n10418_,
    new_n10419_, new_n10420_, new_n10421_, new_n10422_, new_n10423_,
    new_n10424_, new_n10425_, new_n10426_, new_n10427_, new_n10428_,
    new_n10429_, new_n10430_, new_n10431_, new_n10432_, new_n10433_,
    new_n10434_, new_n10435_, new_n10436_, new_n10437_, new_n10438_,
    new_n10439_, new_n10440_, new_n10441_, new_n10442_, new_n10443_,
    new_n10444_, new_n10445_, new_n10446_, new_n10447_, new_n10448_,
    new_n10449_, new_n10450_, new_n10451_, new_n10452_, new_n10453_,
    new_n10454_, new_n10455_, new_n10456_, new_n10457_, new_n10458_,
    new_n10459_, new_n10460_, new_n10461_, new_n10462_, new_n10463_,
    new_n10464_, new_n10465_, new_n10466_, new_n10467_, new_n10468_,
    new_n10469_, new_n10470_, new_n10471_, new_n10472_, new_n10473_,
    new_n10474_, new_n10475_, new_n10476_, new_n10477_, new_n10478_,
    new_n10479_, new_n10480_, new_n10481_, new_n10482_, new_n10483_,
    new_n10484_, new_n10485_, new_n10486_, new_n10487_, new_n10488_,
    new_n10489_, new_n10490_, new_n10491_, new_n10492_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10914_,
    new_n10915_, new_n10916_, new_n10917_, new_n10918_, new_n10919_,
    new_n10920_, new_n10921_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11422_, new_n11423_, new_n11424_, new_n11425_, new_n11426_,
    new_n11427_, new_n11428_, new_n11429_, new_n11430_, new_n11431_,
    new_n11432_, new_n11433_, new_n11434_, new_n11435_, new_n11436_,
    new_n11437_, new_n11438_, new_n11439_, new_n11440_, new_n11441_,
    new_n11442_, new_n11443_, new_n11444_, new_n11445_, new_n11446_,
    new_n11447_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11454_, new_n11455_, new_n11456_,
    new_n11457_, new_n11458_, new_n11459_, new_n11460_, new_n11461_,
    new_n11462_, new_n11463_, new_n11464_, new_n11465_, new_n11466_,
    new_n11467_, new_n11468_, new_n11469_, new_n11470_, new_n11471_,
    new_n11472_, new_n11473_, new_n11474_, new_n11475_, new_n11476_,
    new_n11477_, new_n11478_, new_n11479_, new_n11480_, new_n11481_,
    new_n11482_, new_n11483_, new_n11484_, new_n11485_, new_n11486_,
    new_n11487_, new_n11488_, new_n11489_, new_n11490_, new_n11491_,
    new_n11492_, new_n11493_, new_n11494_, new_n11495_, new_n11496_,
    new_n11497_, new_n11498_, new_n11499_, new_n11500_, new_n11501_,
    new_n11502_, new_n11503_, new_n11504_, new_n11505_, new_n11506_,
    new_n11507_, new_n11508_, new_n11509_, new_n11510_, new_n11511_,
    new_n11512_, new_n11513_, new_n11514_, new_n11515_, new_n11516_,
    new_n11517_, new_n11518_, new_n11519_, new_n11520_, new_n11521_,
    new_n11522_, new_n11523_, new_n11524_, new_n11525_, new_n11526_,
    new_n11527_, new_n11528_, new_n11529_, new_n11530_, new_n11531_,
    new_n11532_, new_n11533_, new_n11534_, new_n11535_, new_n11536_,
    new_n11537_, new_n11538_, new_n11539_, new_n11540_, new_n11541_,
    new_n11542_, new_n11543_, new_n11544_, new_n11545_, new_n11546_,
    new_n11547_, new_n11548_, new_n11549_, new_n11550_, new_n11551_,
    new_n11552_, new_n11553_, new_n11554_, new_n11555_, new_n11556_,
    new_n11557_, new_n11558_, new_n11559_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11796_,
    new_n11797_, new_n11798_, new_n11799_, new_n11800_, new_n11801_,
    new_n11802_, new_n11803_, new_n11804_, new_n11805_, new_n11806_,
    new_n11807_, new_n11808_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11830_, new_n11831_,
    new_n11832_, new_n11833_, new_n11834_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11966_, new_n11967_,
    new_n11968_, new_n11969_, new_n11970_, new_n11971_, new_n11972_,
    new_n11973_, new_n11974_, new_n11975_, new_n11976_, new_n11977_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11988_, new_n11989_, new_n11990_, new_n11991_, new_n11992_,
    new_n11993_, new_n11994_, new_n11995_, new_n11996_, new_n11997_,
    new_n11998_, new_n11999_, new_n12000_, new_n12001_, new_n12002_,
    new_n12003_, new_n12004_, new_n12005_, new_n12006_, new_n12007_,
    new_n12008_, new_n12009_, new_n12010_, new_n12011_, new_n12012_,
    new_n12013_, new_n12014_, new_n12015_, new_n12016_, new_n12017_,
    new_n12018_, new_n12019_, new_n12020_, new_n12021_, new_n12022_,
    new_n12023_, new_n12024_, new_n12025_, new_n12026_, new_n12027_,
    new_n12028_, new_n12029_, new_n12030_, new_n12031_, new_n12032_,
    new_n12033_, new_n12034_, new_n12035_, new_n12036_, new_n12037_,
    new_n12038_, new_n12039_, new_n12040_, new_n12041_, new_n12042_,
    new_n12043_, new_n12044_, new_n12045_, new_n12046_, new_n12047_,
    new_n12048_, new_n12049_, new_n12050_, new_n12051_, new_n12052_,
    new_n12053_, new_n12054_, new_n12055_, new_n12056_, new_n12057_,
    new_n12058_, new_n12059_, new_n12060_, new_n12061_, new_n12062_,
    new_n12063_, new_n12064_, new_n12065_, new_n12066_, new_n12067_,
    new_n12068_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12073_, new_n12074_, new_n12075_, new_n12076_, new_n12077_,
    new_n12078_, new_n12079_, new_n12080_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12164_, new_n12165_, new_n12166_, new_n12167_,
    new_n12168_, new_n12169_, new_n12170_, new_n12171_, new_n12172_,
    new_n12173_, new_n12174_, new_n12175_, new_n12176_, new_n12177_,
    new_n12178_, new_n12179_, new_n12180_, new_n12181_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12226_, new_n12227_,
    new_n12228_, new_n12229_, new_n12230_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12238_, new_n12239_, new_n12240_, new_n12241_, new_n12242_,
    new_n12243_, new_n12244_, new_n12245_, new_n12246_, new_n12247_,
    new_n12248_, new_n12249_, new_n12250_, new_n12251_, new_n12252_,
    new_n12253_, new_n12254_, new_n12255_, new_n12256_, new_n12257_,
    new_n12258_, new_n12259_, new_n12260_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12290_, new_n12291_, new_n12292_,
    new_n12293_, new_n12294_, new_n12295_, new_n12296_, new_n12297_,
    new_n12298_, new_n12299_, new_n12300_, new_n12301_, new_n12302_,
    new_n12303_, new_n12304_, new_n12305_, new_n12306_, new_n12307_,
    new_n12308_, new_n12309_, new_n12310_, new_n12311_, new_n12312_,
    new_n12313_, new_n12314_, new_n12315_, new_n12316_, new_n12317_,
    new_n12318_, new_n12319_, new_n12320_, new_n12321_, new_n12322_,
    new_n12323_, new_n12324_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12390_, new_n12391_, new_n12392_, new_n12393_,
    new_n12394_, new_n12395_, new_n12396_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12417_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12483_,
    new_n12484_, new_n12485_, new_n12486_, new_n12487_, new_n12488_,
    new_n12489_, new_n12490_, new_n12491_, new_n12492_, new_n12493_,
    new_n12494_, new_n12495_, new_n12496_, new_n12497_, new_n12498_,
    new_n12499_, new_n12500_, new_n12501_, new_n12502_, new_n12503_,
    new_n12504_, new_n12505_, new_n12506_, new_n12507_, new_n12508_,
    new_n12509_, new_n12510_, new_n12511_, new_n12512_, new_n12513_,
    new_n12514_, new_n12515_, new_n12516_, new_n12517_, new_n12518_,
    new_n12519_, new_n12520_, new_n12521_, new_n12522_, new_n12523_,
    new_n12524_, new_n12525_, new_n12526_, new_n12527_, new_n12528_,
    new_n12529_, new_n12530_, new_n12531_, new_n12532_, new_n12533_,
    new_n12534_, new_n12535_, new_n12536_, new_n12537_, new_n12538_,
    new_n12539_, new_n12540_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12567_, new_n12568_,
    new_n12569_, new_n12570_, new_n12571_, new_n12572_, new_n12573_,
    new_n12574_, new_n12575_, new_n12576_, new_n12577_, new_n12578_,
    new_n12579_, new_n12580_, new_n12581_, new_n12582_, new_n12583_,
    new_n12584_, new_n12585_, new_n12586_, new_n12587_, new_n12588_,
    new_n12589_, new_n12590_, new_n12591_, new_n12592_, new_n12593_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12610_, new_n12611_, new_n12612_, new_n12613_,
    new_n12614_, new_n12615_, new_n12616_, new_n12617_, new_n12618_,
    new_n12619_, new_n12620_, new_n12621_, new_n12622_, new_n12623_,
    new_n12624_, new_n12625_, new_n12626_, new_n12627_, new_n12628_,
    new_n12629_, new_n12630_, new_n12631_, new_n12632_, new_n12633_,
    new_n12634_, new_n12635_, new_n12636_, new_n12637_, new_n12638_,
    new_n12639_, new_n12640_, new_n12641_, new_n12642_, new_n12643_,
    new_n12644_, new_n12645_, new_n12646_, new_n12647_, new_n12648_,
    new_n12649_, new_n12650_, new_n12651_, new_n12652_, new_n12653_,
    new_n12654_, new_n12655_, new_n12656_, new_n12657_, new_n12658_,
    new_n12659_, new_n12660_, new_n12661_, new_n12662_, new_n12663_,
    new_n12664_, new_n12665_, new_n12666_, new_n12667_, new_n12668_,
    new_n12669_, new_n12670_, new_n12671_, new_n12672_, new_n12673_,
    new_n12674_, new_n12675_, new_n12676_, new_n12677_, new_n12678_,
    new_n12679_, new_n12680_, new_n12681_, new_n12682_, new_n12683_,
    new_n12684_, new_n12685_, new_n12686_, new_n12687_, new_n12688_,
    new_n12689_, new_n12690_, new_n12691_, new_n12692_, new_n12693_,
    new_n12694_, new_n12695_, new_n12696_, new_n12697_, new_n12698_,
    new_n12699_, new_n12700_, new_n12701_, new_n12702_, new_n12703_,
    new_n12704_, new_n12705_, new_n12706_, new_n12707_, new_n12708_,
    new_n12709_, new_n12710_, new_n12711_, new_n12712_, new_n12713_,
    new_n12714_, new_n12715_, new_n12716_, new_n12717_, new_n12718_,
    new_n12719_, new_n12720_, new_n12721_, new_n12722_, new_n12723_,
    new_n12724_, new_n12725_, new_n12726_, new_n12727_, new_n12728_,
    new_n12729_, new_n12730_, new_n12731_, new_n12732_, new_n12733_,
    new_n12734_, new_n12735_, new_n12736_, new_n12737_, new_n12738_,
    new_n12739_, new_n12740_, new_n12741_, new_n12742_, new_n12743_,
    new_n12744_, new_n12745_, new_n12746_, new_n12747_, new_n12748_,
    new_n12749_, new_n12750_, new_n12751_, new_n12752_, new_n12753_,
    new_n12754_, new_n12755_, new_n12756_, new_n12757_, new_n12758_,
    new_n12759_, new_n12760_, new_n12761_, new_n12762_, new_n12763_,
    new_n12764_, new_n12765_, new_n12766_, new_n12767_, new_n12768_,
    new_n12769_, new_n12770_, new_n12771_, new_n12772_, new_n12773_,
    new_n12774_, new_n12775_, new_n12776_, new_n12777_, new_n12778_,
    new_n12779_, new_n12780_, new_n12781_, new_n12782_, new_n12783_,
    new_n12784_, new_n12785_, new_n12786_, new_n12787_, new_n12788_,
    new_n12789_, new_n12790_, new_n12791_, new_n12792_, new_n12793_,
    new_n12794_, new_n12795_, new_n12796_, new_n12797_, new_n12798_,
    new_n12799_, new_n12800_, new_n12801_, new_n12802_, new_n12803_,
    new_n12804_, new_n12805_, new_n12806_, new_n12807_, new_n12808_,
    new_n12809_, new_n12810_, new_n12811_, new_n12812_, new_n12813_,
    new_n12814_, new_n12815_, new_n12816_, new_n12817_, new_n12818_,
    new_n12819_, new_n12820_, new_n12821_, new_n12822_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12833_,
    new_n12834_, new_n12835_, new_n12836_, new_n12837_, new_n12838_,
    new_n12839_, new_n12840_, new_n12841_, new_n12842_, new_n12843_,
    new_n12844_, new_n12845_, new_n12846_, new_n12847_, new_n12848_,
    new_n12849_, new_n12850_, new_n12851_, new_n12852_, new_n12853_,
    new_n12854_, new_n12855_, new_n12856_, new_n12857_, new_n12858_,
    new_n12859_, new_n12860_, new_n12861_, new_n12862_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12868_,
    new_n12869_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13102_, new_n13103_, new_n13104_,
    new_n13105_, new_n13106_, new_n13107_, new_n13108_, new_n13109_,
    new_n13110_, new_n13111_, new_n13112_, new_n13113_, new_n13114_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13121_, new_n13122_, new_n13123_, new_n13124_,
    new_n13125_, new_n13126_, new_n13127_, new_n13128_, new_n13129_,
    new_n13130_, new_n13131_, new_n13132_, new_n13133_, new_n13134_,
    new_n13135_, new_n13136_, new_n13137_, new_n13138_, new_n13139_,
    new_n13140_, new_n13141_, new_n13142_, new_n13143_, new_n13144_,
    new_n13145_, new_n13146_, new_n13147_, new_n13148_, new_n13149_,
    new_n13150_, new_n13151_, new_n13152_, new_n13153_, new_n13154_,
    new_n13155_, new_n13156_, new_n13157_, new_n13158_, new_n13159_,
    new_n13160_, new_n13161_, new_n13162_, new_n13163_, new_n13164_,
    new_n13165_, new_n13166_, new_n13167_, new_n13168_, new_n13169_,
    new_n13170_, new_n13171_, new_n13172_, new_n13173_, new_n13174_,
    new_n13175_, new_n13176_, new_n13177_, new_n13178_, new_n13179_,
    new_n13180_, new_n13181_, new_n13182_, new_n13183_, new_n13184_,
    new_n13185_, new_n13186_, new_n13187_, new_n13188_, new_n13189_,
    new_n13190_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13200_, new_n13201_, new_n13202_, new_n13203_, new_n13204_,
    new_n13205_, new_n13206_, new_n13207_, new_n13208_, new_n13209_,
    new_n13210_, new_n13211_, new_n13212_, new_n13213_, new_n13214_,
    new_n13215_, new_n13216_, new_n13217_, new_n13218_, new_n13219_,
    new_n13220_, new_n13221_, new_n13222_, new_n13223_, new_n13224_,
    new_n13225_, new_n13226_, new_n13227_, new_n13228_, new_n13229_,
    new_n13230_, new_n13231_, new_n13232_, new_n13233_, new_n13234_,
    new_n13235_, new_n13236_, new_n13237_, new_n13238_, new_n13239_,
    new_n13240_, new_n13241_, new_n13242_, new_n13243_, new_n13244_,
    new_n13245_, new_n13246_, new_n13247_, new_n13248_, new_n13249_,
    new_n13250_, new_n13251_, new_n13252_, new_n13253_, new_n13254_,
    new_n13255_, new_n13256_, new_n13257_, new_n13258_, new_n13259_,
    new_n13260_, new_n13261_, new_n13262_, new_n13263_, new_n13264_,
    new_n13265_, new_n13266_, new_n13267_, new_n13268_, new_n13269_,
    new_n13270_, new_n13271_, new_n13272_, new_n13273_, new_n13274_,
    new_n13275_, new_n13276_, new_n13277_, new_n13278_, new_n13279_,
    new_n13280_, new_n13281_, new_n13282_, new_n13283_, new_n13284_,
    new_n13285_, new_n13286_, new_n13287_, new_n13288_, new_n13289_,
    new_n13290_, new_n13291_, new_n13292_, new_n13293_, new_n13294_,
    new_n13295_, new_n13296_, new_n13297_, new_n13298_, new_n13299_,
    new_n13300_, new_n13301_, new_n13302_, new_n13303_, new_n13304_,
    new_n13305_, new_n13306_, new_n13307_, new_n13308_, new_n13309_,
    new_n13310_, new_n13311_, new_n13312_, new_n13313_, new_n13314_,
    new_n13315_, new_n13316_, new_n13317_, new_n13318_, new_n13319_,
    new_n13320_, new_n13321_, new_n13322_, new_n13323_, new_n13324_,
    new_n13325_, new_n13326_, new_n13327_, new_n13328_, new_n13329_,
    new_n13330_, new_n13331_, new_n13332_, new_n13333_, new_n13334_,
    new_n13335_, new_n13336_, new_n13337_, new_n13338_, new_n13339_,
    new_n13340_, new_n13341_, new_n13342_, new_n13343_, new_n13344_,
    new_n13345_, new_n13346_, new_n13347_, new_n13348_, new_n13349_,
    new_n13350_, new_n13351_, new_n13352_, new_n13353_, new_n13354_,
    new_n13355_, new_n13356_, new_n13357_, new_n13358_, new_n13359_,
    new_n13360_, new_n13361_, new_n13362_, new_n13363_, new_n13364_,
    new_n13365_, new_n13366_, new_n13367_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13375_, new_n13376_, new_n13377_, new_n13378_, new_n13379_,
    new_n13380_, new_n13381_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14280_, new_n14281_,
    new_n14282_, new_n14283_, new_n14284_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14290_, new_n14291_,
    new_n14292_, new_n14293_, new_n14294_, new_n14295_, new_n14296_,
    new_n14297_, new_n14298_, new_n14299_, new_n14300_, new_n14301_,
    new_n14302_, new_n14303_, new_n14304_, new_n14305_, new_n14306_,
    new_n14307_, new_n14308_, new_n14309_, new_n14310_, new_n14311_,
    new_n14312_, new_n14313_, new_n14314_, new_n14315_, new_n14316_,
    new_n14317_, new_n14318_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14325_, new_n14326_,
    new_n14327_, new_n14328_, new_n14329_, new_n14330_, new_n14331_,
    new_n14332_, new_n14333_, new_n14334_, new_n14335_, new_n14336_,
    new_n14337_, new_n14338_, new_n14339_, new_n14340_, new_n14341_,
    new_n14342_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14350_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14356_,
    new_n14357_, new_n14358_, new_n14359_, new_n14360_, new_n14361_,
    new_n14362_, new_n14363_, new_n14364_, new_n14365_, new_n14366_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14379_, new_n14380_, new_n14381_,
    new_n14382_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14387_, new_n14388_, new_n14389_, new_n14390_, new_n14391_,
    new_n14392_, new_n14393_, new_n14394_, new_n14395_, new_n14396_,
    new_n14397_, new_n14398_, new_n14399_, new_n14400_, new_n14401_,
    new_n14402_, new_n14403_, new_n14404_, new_n14405_, new_n14406_,
    new_n14407_, new_n14408_, new_n14409_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14416_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14424_, new_n14425_, new_n14426_,
    new_n14427_, new_n14428_, new_n14429_, new_n14430_, new_n14431_,
    new_n14432_, new_n14433_, new_n14434_, new_n14435_, new_n14436_,
    new_n14437_, new_n14438_, new_n14439_, new_n14440_, new_n14441_,
    new_n14442_, new_n14443_, new_n14444_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14551_, new_n14552_,
    new_n14553_, new_n14554_, new_n14555_, new_n14556_, new_n14557_,
    new_n14558_, new_n14559_, new_n14560_, new_n14561_, new_n14562_,
    new_n14563_, new_n14564_, new_n14565_, new_n14566_, new_n14567_,
    new_n14568_, new_n14569_, new_n14570_, new_n14571_, new_n14572_,
    new_n14573_, new_n14574_, new_n14575_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14712_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14719_, new_n14720_, new_n14721_, new_n14722_,
    new_n14723_, new_n14724_, new_n14725_, new_n14726_, new_n14727_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14734_, new_n14735_, new_n14736_, new_n14737_,
    new_n14738_, new_n14739_, new_n14740_, new_n14741_, new_n14742_,
    new_n14743_, new_n14744_, new_n14745_, new_n14746_, new_n14747_,
    new_n14748_, new_n14749_, new_n14750_, new_n14751_, new_n14752_,
    new_n14753_, new_n14754_, new_n14755_, new_n14756_, new_n14757_,
    new_n14758_, new_n14759_, new_n14760_, new_n14761_, new_n14762_,
    new_n14763_, new_n14764_, new_n14765_, new_n14766_, new_n14767_,
    new_n14768_, new_n14769_, new_n14770_, new_n14771_, new_n14772_,
    new_n14773_, new_n14774_, new_n14775_, new_n14776_, new_n14777_,
    new_n14778_, new_n14779_, new_n14780_, new_n14781_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14818_, new_n14819_, new_n14820_, new_n14821_, new_n14822_,
    new_n14823_, new_n14824_, new_n14825_, new_n14826_, new_n14827_,
    new_n14828_, new_n14829_, new_n14830_, new_n14831_, new_n14832_,
    new_n14833_, new_n14834_, new_n14835_, new_n14836_, new_n14837_,
    new_n14838_, new_n14839_, new_n14840_, new_n14841_, new_n14842_,
    new_n14843_, new_n14844_, new_n14845_, new_n14846_, new_n14847_,
    new_n14848_, new_n14849_, new_n14850_, new_n14851_, new_n14852_,
    new_n14853_, new_n14854_, new_n14855_, new_n14856_, new_n14857_,
    new_n14858_, new_n14859_, new_n14860_, new_n14861_, new_n14862_,
    new_n14863_, new_n14864_, new_n14865_, new_n14866_, new_n14867_,
    new_n14868_, new_n14869_, new_n14870_, new_n14871_, new_n14872_,
    new_n14873_, new_n14874_, new_n14875_, new_n14876_, new_n14877_,
    new_n14878_, new_n14879_, new_n14880_, new_n14881_, new_n14882_,
    new_n14883_, new_n14884_, new_n14885_, new_n14886_, new_n14887_,
    new_n14888_, new_n14889_, new_n14890_, new_n14891_, new_n14892_,
    new_n14893_, new_n14894_, new_n14895_, new_n14896_, new_n14897_,
    new_n14898_, new_n14899_, new_n14900_, new_n14901_, new_n14902_,
    new_n14903_, new_n14904_, new_n14905_, new_n14906_, new_n14907_,
    new_n14908_, new_n14909_, new_n14910_, new_n14911_, new_n14912_,
    new_n14913_, new_n14914_, new_n14915_, new_n14916_, new_n14917_,
    new_n14918_, new_n14919_, new_n14920_, new_n14921_, new_n14922_,
    new_n14923_, new_n14924_, new_n14925_, new_n14926_, new_n14927_,
    new_n14928_, new_n14929_, new_n14930_, new_n14931_, new_n14932_,
    new_n14933_, new_n14934_, new_n14935_, new_n14936_, new_n14937_,
    new_n14938_, new_n14939_, new_n14940_, new_n14941_, new_n14942_,
    new_n14943_, new_n14944_, new_n14945_, new_n14946_, new_n14947_,
    new_n14948_, new_n14949_, new_n14950_, new_n14951_, new_n14952_,
    new_n14953_, new_n14954_, new_n14955_, new_n14956_, new_n14957_,
    new_n14958_, new_n14959_, new_n14960_, new_n14961_, new_n14962_,
    new_n14963_, new_n14964_, new_n14965_, new_n14967_, new_n14968_,
    new_n14969_, new_n14970_, new_n14971_, new_n14972_, new_n14973_,
    new_n14974_, new_n14975_, new_n14976_, new_n14977_, new_n14978_,
    new_n14979_, new_n14980_, new_n14981_, new_n14982_, new_n14983_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15007_, new_n15008_,
    new_n15009_, new_n15010_, new_n15011_, new_n15012_, new_n15013_,
    new_n15014_, new_n15015_, new_n15016_, new_n15017_, new_n15018_,
    new_n15019_, new_n15020_, new_n15021_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15026_, new_n15027_, new_n15028_,
    new_n15029_, new_n15030_, new_n15031_, new_n15032_, new_n15033_,
    new_n15034_, new_n15035_, new_n15036_, new_n15037_, new_n15038_,
    new_n15039_, new_n15040_, new_n15041_, new_n15042_, new_n15043_,
    new_n15044_, new_n15045_, new_n15046_, new_n15047_, new_n15048_,
    new_n15049_, new_n15050_, new_n15051_, new_n15052_, new_n15053_,
    new_n15054_, new_n15055_, new_n15056_, new_n15057_, new_n15058_,
    new_n15059_, new_n15060_, new_n15061_, new_n15062_, new_n15063_,
    new_n15064_, new_n15065_, new_n15066_, new_n15067_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15074_, new_n15075_, new_n15076_, new_n15077_, new_n15078_,
    new_n15079_, new_n15080_, new_n15081_, new_n15082_, new_n15083_,
    new_n15084_, new_n15085_, new_n15086_, new_n15087_, new_n15088_,
    new_n15089_, new_n15090_, new_n15091_, new_n15092_, new_n15093_,
    new_n15094_, new_n15095_, new_n15096_, new_n15097_, new_n15098_,
    new_n15099_, new_n15100_, new_n15101_, new_n15102_, new_n15103_,
    new_n15104_, new_n15105_, new_n15106_, new_n15107_, new_n15108_,
    new_n15109_, new_n15110_, new_n15111_, new_n15112_, new_n15113_,
    new_n15114_, new_n15115_, new_n15116_, new_n15117_, new_n15118_,
    new_n15119_, new_n15120_, new_n15121_, new_n15122_, new_n15123_,
    new_n15124_, new_n15125_, new_n15126_, new_n15127_, new_n15128_,
    new_n15129_, new_n15130_, new_n15131_, new_n15132_, new_n15133_,
    new_n15134_, new_n15135_, new_n15136_, new_n15137_, new_n15138_,
    new_n15139_, new_n15140_, new_n15141_, new_n15142_, new_n15143_,
    new_n15144_, new_n15145_, new_n15146_, new_n15147_, new_n15148_,
    new_n15149_, new_n15150_, new_n15151_, new_n15152_, new_n15153_,
    new_n15154_, new_n15155_, new_n15156_, new_n15157_, new_n15158_,
    new_n15159_, new_n15160_, new_n15161_, new_n15162_, new_n15163_,
    new_n15164_, new_n15165_, new_n15166_, new_n15167_, new_n15168_,
    new_n15169_, new_n15170_, new_n15171_, new_n15172_, new_n15173_,
    new_n15174_, new_n15175_, new_n15176_, new_n15177_, new_n15178_,
    new_n15179_, new_n15180_, new_n15181_, new_n15182_, new_n15183_,
    new_n15184_, new_n15185_, new_n15186_, new_n15187_, new_n15188_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15197_, new_n15198_,
    new_n15199_, new_n15200_, new_n15201_, new_n15202_, new_n15203_,
    new_n15204_, new_n15205_, new_n15206_, new_n15207_, new_n15208_,
    new_n15209_, new_n15210_, new_n15211_, new_n15212_, new_n15213_,
    new_n15214_, new_n15215_, new_n15216_, new_n15217_, new_n15218_,
    new_n15219_, new_n15220_, new_n15221_, new_n15222_, new_n15223_,
    new_n15224_, new_n15225_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15232_, new_n15233_,
    new_n15234_, new_n15235_, new_n15236_, new_n15237_, new_n15238_,
    new_n15239_, new_n15240_, new_n15241_, new_n15242_, new_n15243_,
    new_n15244_, new_n15245_, new_n15246_, new_n15247_, new_n15248_,
    new_n15249_, new_n15250_, new_n15251_, new_n15252_, new_n15253_,
    new_n15254_, new_n15255_, new_n15256_, new_n15257_, new_n15258_,
    new_n15259_, new_n15260_, new_n15261_, new_n15262_, new_n15263_,
    new_n15264_, new_n15265_, new_n15266_, new_n15267_, new_n15268_,
    new_n15269_, new_n15270_, new_n15271_, new_n15272_, new_n15273_,
    new_n15274_, new_n15275_, new_n15276_, new_n15277_, new_n15278_,
    new_n15279_, new_n15280_, new_n15281_, new_n15282_, new_n15283_,
    new_n15284_, new_n15285_, new_n15286_, new_n15287_, new_n15288_,
    new_n15289_, new_n15290_, new_n15291_, new_n15292_, new_n15293_,
    new_n15294_, new_n15295_, new_n15296_, new_n15297_, new_n15298_,
    new_n15299_, new_n15300_, new_n15301_, new_n15302_, new_n15303_,
    new_n15304_, new_n15305_, new_n15306_, new_n15307_, new_n15308_,
    new_n15309_, new_n15310_, new_n15311_, new_n15312_, new_n15313_,
    new_n15314_, new_n15315_, new_n15316_, new_n15317_, new_n15318_,
    new_n15319_, new_n15320_, new_n15321_, new_n15322_, new_n15323_,
    new_n15324_, new_n15325_, new_n15326_, new_n15327_, new_n15328_,
    new_n15329_, new_n15330_, new_n15331_, new_n15332_, new_n15333_,
    new_n15334_, new_n15335_, new_n15336_, new_n15337_, new_n15338_,
    new_n15339_, new_n15340_, new_n15341_, new_n15342_, new_n15343_,
    new_n15344_, new_n15345_, new_n15346_, new_n15347_, new_n15348_,
    new_n15349_, new_n15350_, new_n15351_, new_n15352_, new_n15353_,
    new_n15354_, new_n15355_, new_n15356_, new_n15357_, new_n15358_,
    new_n15359_, new_n15360_, new_n15361_, new_n15362_, new_n15363_,
    new_n15364_, new_n15365_, new_n15366_, new_n15367_, new_n15368_,
    new_n15369_, new_n15370_, new_n15371_, new_n15372_, new_n15373_,
    new_n15374_, new_n15375_, new_n15376_, new_n15377_, new_n15378_,
    new_n15379_, new_n15380_, new_n15381_, new_n15382_, new_n15383_,
    new_n15384_, new_n15385_, new_n15386_, new_n15387_, new_n15388_,
    new_n15389_, new_n15390_, new_n15391_, new_n15392_, new_n15393_,
    new_n15394_, new_n15395_, new_n15396_, new_n15397_, new_n15398_,
    new_n15399_, new_n15400_, new_n15401_, new_n15402_, new_n15403_,
    new_n15404_, new_n15405_, new_n15406_, new_n15407_, new_n15408_,
    new_n15409_, new_n15410_, new_n15411_, new_n15412_, new_n15413_,
    new_n15414_, new_n15415_, new_n15416_, new_n15417_, new_n15418_,
    new_n15419_, new_n15420_, new_n15421_, new_n15422_, new_n15423_,
    new_n15424_, new_n15425_, new_n15426_, new_n15427_, new_n15428_,
    new_n15429_, new_n15430_, new_n15431_, new_n15432_, new_n15433_,
    new_n15434_, new_n15435_, new_n15436_, new_n15437_, new_n15438_,
    new_n15439_, new_n15440_, new_n15441_, new_n15442_, new_n15443_,
    new_n15444_, new_n15445_, new_n15446_, new_n15447_, new_n15448_,
    new_n15449_, new_n15450_, new_n15451_, new_n15452_, new_n15453_,
    new_n15454_, new_n15455_, new_n15456_, new_n15457_, new_n15458_,
    new_n15459_, new_n15460_, new_n15461_, new_n15462_, new_n15463_,
    new_n15464_, new_n15465_, new_n15466_, new_n15467_, new_n15468_,
    new_n15469_, new_n15470_, new_n15471_, new_n15472_, new_n15473_,
    new_n15474_, new_n15475_, new_n15476_, new_n15477_, new_n15478_,
    new_n15479_, new_n15480_, new_n15481_, new_n15482_, new_n15483_,
    new_n15484_, new_n15485_, new_n15486_, new_n15487_, new_n15488_,
    new_n15489_, new_n15490_, new_n15491_, new_n15492_, new_n15493_,
    new_n15494_, new_n15495_, new_n15496_, new_n15497_, new_n15498_,
    new_n15499_, new_n15500_, new_n15501_, new_n15502_, new_n15503_,
    new_n15504_, new_n15505_, new_n15506_, new_n15507_, new_n15508_,
    new_n15509_, new_n15510_, new_n15511_, new_n15512_, new_n15513_,
    new_n15514_, new_n15515_, new_n15516_, new_n15517_, new_n15518_,
    new_n15519_, new_n15520_, new_n15521_, new_n15522_, new_n15523_,
    new_n15524_, new_n15525_, new_n15526_, new_n15527_, new_n15528_,
    new_n15529_, new_n15530_, new_n15531_, new_n15532_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15633_, new_n15634_,
    new_n15635_, new_n15636_, new_n15637_, new_n15638_, new_n15639_,
    new_n15640_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15690_, new_n15691_, new_n15692_, new_n15693_, new_n15694_,
    new_n15695_, new_n15696_, new_n15697_, new_n15698_, new_n15699_,
    new_n15700_, new_n15701_, new_n15702_, new_n15703_, new_n15704_,
    new_n15705_, new_n15706_, new_n15707_, new_n15708_, new_n15709_,
    new_n15710_, new_n15711_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15808_, new_n15809_,
    new_n15810_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15897_, new_n15898_, new_n15899_,
    new_n15900_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15910_, new_n15911_, new_n15912_, new_n15913_, new_n15914_,
    new_n15915_, new_n15916_, new_n15917_, new_n15918_, new_n15919_,
    new_n15920_, new_n15921_, new_n15922_, new_n15923_, new_n15924_,
    new_n15925_, new_n15926_, new_n15927_, new_n15928_, new_n15929_,
    new_n15930_, new_n15931_, new_n15932_, new_n15933_, new_n15934_,
    new_n15935_, new_n15936_, new_n15937_, new_n15938_, new_n15939_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15945_, new_n15946_, new_n15947_, new_n15948_, new_n15949_,
    new_n15950_, new_n15951_, new_n15952_, new_n15953_, new_n15954_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16001_, new_n16002_, new_n16003_, new_n16004_,
    new_n16005_, new_n16006_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16067_, new_n16068_, new_n16069_,
    new_n16070_, new_n16071_, new_n16072_, new_n16073_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16349_, new_n16350_,
    new_n16351_, new_n16352_, new_n16353_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16361_, new_n16362_, new_n16363_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16489_, new_n16490_,
    new_n16491_, new_n16492_, new_n16493_, new_n16494_, new_n16495_,
    new_n16496_, new_n16497_, new_n16498_, new_n16499_, new_n16500_,
    new_n16501_, new_n16502_, new_n16503_, new_n16504_, new_n16505_,
    new_n16506_, new_n16507_, new_n16508_, new_n16509_, new_n16510_,
    new_n16511_, new_n16512_, new_n16513_, new_n16514_, new_n16515_,
    new_n16516_, new_n16517_, new_n16518_, new_n16519_, new_n16520_,
    new_n16521_, new_n16522_, new_n16523_, new_n16524_, new_n16525_,
    new_n16526_, new_n16527_, new_n16528_, new_n16529_, new_n16530_,
    new_n16531_, new_n16532_, new_n16533_, new_n16534_, new_n16535_,
    new_n16536_, new_n16537_, new_n16538_, new_n16539_, new_n16540_,
    new_n16541_, new_n16542_, new_n16543_, new_n16544_, new_n16545_,
    new_n16546_, new_n16547_, new_n16548_, new_n16549_, new_n16550_,
    new_n16551_, new_n16552_, new_n16553_, new_n16554_, new_n16555_,
    new_n16556_, new_n16557_, new_n16558_, new_n16559_, new_n16560_,
    new_n16561_, new_n16562_, new_n16563_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16618_, new_n16619_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16933_, new_n16934_, new_n16935_, new_n16936_,
    new_n16937_, new_n16938_, new_n16939_, new_n16940_, new_n16941_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16955_, new_n16956_,
    new_n16957_, new_n16958_, new_n16959_, new_n16960_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16980_, new_n16981_,
    new_n16982_, new_n16983_, new_n16984_, new_n16985_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16992_, new_n16993_, new_n16994_, new_n16995_, new_n16996_,
    new_n16997_, new_n16998_, new_n16999_, new_n17000_, new_n17001_,
    new_n17002_, new_n17003_, new_n17004_, new_n17005_, new_n17006_,
    new_n17007_, new_n17008_, new_n17009_, new_n17010_, new_n17011_,
    new_n17012_, new_n17013_, new_n17014_, new_n17015_, new_n17016_,
    new_n17017_, new_n17018_, new_n17019_, new_n17020_, new_n17021_,
    new_n17022_, new_n17023_, new_n17024_, new_n17025_, new_n17026_,
    new_n17027_, new_n17028_, new_n17029_, new_n17030_, new_n17031_,
    new_n17032_, new_n17033_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17106_,
    new_n17107_, new_n17108_, new_n17109_, new_n17110_, new_n17111_,
    new_n17112_, new_n17113_, new_n17114_, new_n17115_, new_n17116_,
    new_n17117_, new_n17118_, new_n17119_, new_n17120_, new_n17121_,
    new_n17122_, new_n17123_, new_n17124_, new_n17125_, new_n17126_,
    new_n17127_, new_n17128_, new_n17129_, new_n17130_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17226_, new_n17227_,
    new_n17228_, new_n17229_, new_n17230_, new_n17231_, new_n17232_,
    new_n17233_, new_n17234_, new_n17235_, new_n17236_, new_n17237_,
    new_n17238_, new_n17239_, new_n17240_, new_n17241_, new_n17242_,
    new_n17243_, new_n17244_, new_n17245_, new_n17246_, new_n17247_,
    new_n17248_, new_n17249_, new_n17250_, new_n17251_, new_n17252_,
    new_n17253_, new_n17254_, new_n17255_, new_n17256_, new_n17257_,
    new_n17258_, new_n17259_, new_n17260_, new_n17261_, new_n17262_,
    new_n17263_, new_n17264_, new_n17265_, new_n17266_, new_n17267_,
    new_n17268_, new_n17269_, new_n17270_, new_n17271_, new_n17272_,
    new_n17273_, new_n17274_, new_n17275_, new_n17276_, new_n17277_,
    new_n17278_, new_n17279_, new_n17280_, new_n17281_, new_n17282_,
    new_n17283_, new_n17284_, new_n17285_, new_n17286_, new_n17287_,
    new_n17288_, new_n17289_, new_n17290_, new_n17291_, new_n17292_,
    new_n17293_, new_n17294_, new_n17295_, new_n17296_, new_n17297_,
    new_n17298_, new_n17299_, new_n17300_, new_n17301_, new_n17302_,
    new_n17303_, new_n17304_, new_n17305_, new_n17306_, new_n17307_,
    new_n17308_, new_n17309_, new_n17310_, new_n17311_, new_n17312_,
    new_n17313_, new_n17314_, new_n17315_, new_n17316_, new_n17317_,
    new_n17318_, new_n17319_, new_n17320_, new_n17321_, new_n17322_,
    new_n17323_, new_n17324_, new_n17325_, new_n17326_, new_n17327_,
    new_n17328_, new_n17329_, new_n17330_, new_n17331_, new_n17332_,
    new_n17333_, new_n17334_, new_n17335_, new_n17336_, new_n17337_,
    new_n17338_, new_n17339_, new_n17340_, new_n17341_, new_n17342_,
    new_n17343_, new_n17344_, new_n17345_, new_n17346_, new_n17347_,
    new_n17348_, new_n17349_, new_n17350_, new_n17351_, new_n17352_,
    new_n17353_, new_n17354_, new_n17355_, new_n17356_, new_n17357_,
    new_n17358_, new_n17359_, new_n17360_, new_n17361_, new_n17362_,
    new_n17363_, new_n17364_, new_n17365_, new_n17366_, new_n17367_,
    new_n17368_, new_n17369_, new_n17370_, new_n17371_, new_n17372_,
    new_n17373_, new_n17374_, new_n17375_, new_n17376_, new_n17377_,
    new_n17378_, new_n17379_, new_n17380_, new_n17381_, new_n17382_,
    new_n17383_, new_n17384_, new_n17385_, new_n17386_, new_n17387_,
    new_n17388_, new_n17389_, new_n17390_, new_n17391_, new_n17392_,
    new_n17393_, new_n17394_, new_n17395_, new_n17396_, new_n17397_,
    new_n17398_, new_n17399_, new_n17400_, new_n17401_, new_n17402_,
    new_n17403_, new_n17404_, new_n17405_, new_n17406_, new_n17407_,
    new_n17408_, new_n17409_, new_n17410_, new_n17411_, new_n17412_,
    new_n17413_, new_n17414_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17450_, new_n17451_, new_n17452_,
    new_n17453_, new_n17454_, new_n17455_, new_n17456_, new_n17457_,
    new_n17458_, new_n17459_, new_n17460_, new_n17461_, new_n17462_,
    new_n17463_, new_n17464_, new_n17465_, new_n17466_, new_n17467_,
    new_n17468_, new_n17469_, new_n17470_, new_n17471_, new_n17472_,
    new_n17473_, new_n17474_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17480_, new_n17481_, new_n17482_,
    new_n17483_, new_n17484_, new_n17485_, new_n17486_, new_n17487_,
    new_n17488_, new_n17489_, new_n17490_, new_n17491_, new_n17492_,
    new_n17493_, new_n17494_, new_n17495_, new_n17496_, new_n17497_,
    new_n17498_, new_n17499_, new_n17500_, new_n17501_, new_n17502_,
    new_n17503_, new_n17504_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17510_, new_n17511_, new_n17512_,
    new_n17513_, new_n17514_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17563_, new_n17564_, new_n17565_, new_n17566_, new_n17567_,
    new_n17568_, new_n17569_, new_n17570_, new_n17571_, new_n17572_,
    new_n17573_, new_n17574_, new_n17575_, new_n17576_, new_n17577_,
    new_n17578_, new_n17579_, new_n17580_, new_n17581_, new_n17582_,
    new_n17583_, new_n17584_, new_n17585_, new_n17586_, new_n17587_,
    new_n17588_, new_n17589_, new_n17590_, new_n17591_, new_n17592_,
    new_n17593_, new_n17594_, new_n17595_, new_n17596_, new_n17597_,
    new_n17598_, new_n17599_, new_n17600_, new_n17601_, new_n17602_,
    new_n17603_, new_n17604_, new_n17605_, new_n17606_, new_n17607_,
    new_n17608_, new_n17609_, new_n17610_, new_n17611_, new_n17612_,
    new_n17613_, new_n17614_, new_n17615_, new_n17616_, new_n17617_,
    new_n17618_, new_n17619_, new_n17620_, new_n17621_, new_n17622_,
    new_n17623_, new_n17624_, new_n17625_, new_n17626_, new_n17627_,
    new_n17628_, new_n17629_, new_n17630_, new_n17631_, new_n17632_,
    new_n17633_, new_n17634_, new_n17635_, new_n17636_, new_n17637_,
    new_n17638_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17653_, new_n17654_, new_n17655_, new_n17656_, new_n17657_,
    new_n17658_, new_n17659_, new_n17660_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17680_, new_n17681_, new_n17682_,
    new_n17683_, new_n17684_, new_n17685_, new_n17686_, new_n17687_,
    new_n17688_, new_n17689_, new_n17690_, new_n17691_, new_n17692_,
    new_n17693_, new_n17694_, new_n17695_, new_n17696_, new_n17697_,
    new_n17698_, new_n17699_, new_n17700_, new_n17701_, new_n17702_,
    new_n17703_, new_n17704_, new_n17705_, new_n17706_, new_n17707_,
    new_n17708_, new_n17709_, new_n17710_, new_n17711_, new_n17712_,
    new_n17713_, new_n17714_, new_n17715_, new_n17716_, new_n17717_,
    new_n17718_, new_n17719_, new_n17720_, new_n17721_, new_n17722_,
    new_n17723_, new_n17724_, new_n17725_, new_n17726_, new_n17727_,
    new_n17728_, new_n17729_, new_n17730_, new_n17731_, new_n17732_,
    new_n17733_, new_n17734_, new_n17735_, new_n17736_, new_n17737_,
    new_n17738_, new_n17739_, new_n17740_, new_n17741_, new_n17742_,
    new_n17743_, new_n17744_, new_n17745_, new_n17746_, new_n17747_,
    new_n17748_, new_n17749_, new_n17750_, new_n17751_, new_n17752_,
    new_n17753_, new_n17754_, new_n17755_, new_n17756_, new_n17757_,
    new_n17758_, new_n17759_, new_n17760_, new_n17761_, new_n17762_,
    new_n17763_, new_n17764_, new_n17765_, new_n17766_, new_n17767_,
    new_n17768_, new_n17769_, new_n17770_, new_n17771_, new_n17772_,
    new_n17773_, new_n17774_, new_n17775_, new_n17776_, new_n17777_,
    new_n17778_, new_n17779_, new_n17780_, new_n17781_, new_n17782_,
    new_n17783_, new_n17784_, new_n17785_, new_n17786_, new_n17787_,
    new_n17788_, new_n17789_, new_n17790_, new_n17791_, new_n17792_,
    new_n17793_, new_n17794_, new_n17795_, new_n17796_, new_n17797_,
    new_n17798_, new_n17799_, new_n17800_, new_n17801_, new_n17802_,
    new_n17803_, new_n17804_, new_n17805_, new_n17806_, new_n17807_,
    new_n17808_, new_n17809_, new_n17810_, new_n17811_, new_n17812_,
    new_n17813_, new_n17814_, new_n17815_, new_n17816_, new_n17817_,
    new_n17818_, new_n17819_, new_n17820_, new_n17821_, new_n17822_,
    new_n17823_, new_n17824_, new_n17825_, new_n17826_, new_n17827_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17834_, new_n17835_, new_n17836_, new_n17837_, new_n17838_,
    new_n17839_, new_n17840_, new_n17841_, new_n17842_, new_n17843_,
    new_n17844_, new_n17845_, new_n17846_, new_n17847_, new_n17848_,
    new_n17849_, new_n17850_, new_n17851_, new_n17852_, new_n17853_,
    new_n17854_, new_n17855_, new_n17856_, new_n17857_, new_n17858_,
    new_n17859_, new_n17860_, new_n17861_, new_n17862_, new_n17863_,
    new_n17864_, new_n17865_, new_n17866_, new_n17867_, new_n17868_,
    new_n17869_, new_n17870_, new_n17871_, new_n17872_, new_n17873_,
    new_n17874_, new_n17875_, new_n17876_, new_n17877_, new_n17878_,
    new_n17879_, new_n17880_, new_n17881_, new_n17882_, new_n17883_,
    new_n17884_, new_n17885_, new_n17886_, new_n17887_, new_n17888_,
    new_n17889_, new_n17890_, new_n17891_, new_n17892_, new_n17893_,
    new_n17894_, new_n17895_, new_n17896_, new_n17897_, new_n17898_,
    new_n17899_, new_n17900_, new_n17901_, new_n17902_, new_n17903_,
    new_n17904_, new_n17905_, new_n17906_, new_n17907_, new_n17908_,
    new_n17909_, new_n17910_, new_n17911_, new_n17912_, new_n17913_,
    new_n17914_, new_n17915_, new_n17916_, new_n17917_, new_n17918_,
    new_n17919_, new_n17920_, new_n17921_, new_n17922_, new_n17923_,
    new_n17924_, new_n17925_, new_n17926_, new_n17927_, new_n17928_,
    new_n17929_, new_n17930_, new_n17931_, new_n17932_, new_n17933_,
    new_n17934_, new_n17935_, new_n17936_, new_n17937_, new_n17938_,
    new_n17939_, new_n17940_, new_n17941_, new_n17942_, new_n17943_,
    new_n17944_, new_n17945_, new_n17946_, new_n17947_, new_n17948_,
    new_n17949_, new_n17950_, new_n17951_, new_n17952_, new_n17953_,
    new_n17954_, new_n17955_, new_n17956_, new_n17957_, new_n17958_,
    new_n17959_, new_n17960_, new_n17961_, new_n17962_, new_n17963_,
    new_n17964_, new_n17965_, new_n17966_, new_n17967_, new_n17968_,
    new_n17969_, new_n17970_, new_n17971_, new_n17972_, new_n17973_,
    new_n17974_, new_n17975_, new_n17976_, new_n17977_, new_n17978_,
    new_n17979_, new_n17980_, new_n17981_, new_n17982_, new_n17983_,
    new_n17984_, new_n17985_, new_n17986_, new_n17987_, new_n17988_,
    new_n17989_, new_n17990_, new_n17991_, new_n17992_, new_n17993_,
    new_n17994_, new_n17995_, new_n17996_, new_n17997_, new_n17998_,
    new_n17999_, new_n18000_, new_n18001_, new_n18002_, new_n18003_,
    new_n18004_, new_n18005_, new_n18006_, new_n18007_, new_n18008_,
    new_n18009_, new_n18010_, new_n18011_, new_n18012_, new_n18013_,
    new_n18014_, new_n18015_, new_n18016_, new_n18017_, new_n18018_,
    new_n18019_, new_n18020_, new_n18021_, new_n18022_, new_n18023_,
    new_n18024_, new_n18025_, new_n18026_, new_n18027_, new_n18028_,
    new_n18029_, new_n18030_, new_n18031_, new_n18032_, new_n18033_,
    new_n18034_, new_n18035_, new_n18036_, new_n18037_, new_n18038_,
    new_n18039_, new_n18040_, new_n18041_, new_n18042_, new_n18043_,
    new_n18044_, new_n18045_, new_n18046_, new_n18047_, new_n18048_,
    new_n18049_, new_n18050_, new_n18051_, new_n18052_, new_n18053_,
    new_n18054_, new_n18055_, new_n18056_, new_n18057_, new_n18058_,
    new_n18059_, new_n18060_, new_n18061_, new_n18062_, new_n18063_,
    new_n18064_, new_n18065_, new_n18066_, new_n18067_, new_n18068_,
    new_n18069_, new_n18070_, new_n18071_, new_n18072_, new_n18073_,
    new_n18074_, new_n18075_, new_n18076_, new_n18077_, new_n18078_,
    new_n18079_, new_n18080_, new_n18081_, new_n18082_, new_n18083_,
    new_n18084_, new_n18085_, new_n18086_, new_n18087_, new_n18088_,
    new_n18089_, new_n18090_, new_n18091_, new_n18092_, new_n18093_,
    new_n18094_, new_n18095_, new_n18096_, new_n18097_, new_n18098_,
    new_n18099_, new_n18100_, new_n18101_, new_n18102_, new_n18103_,
    new_n18104_, new_n18105_, new_n18106_, new_n18107_, new_n18108_,
    new_n18109_, new_n18110_, new_n18111_, new_n18112_, new_n18113_,
    new_n18114_, new_n18115_, new_n18116_, new_n18117_, new_n18118_,
    new_n18119_, new_n18120_, new_n18121_, new_n18122_, new_n18123_,
    new_n18124_, new_n18125_, new_n18126_, new_n18127_, new_n18128_,
    new_n18129_, new_n18130_, new_n18131_, new_n18132_, new_n18133_,
    new_n18134_, new_n18135_, new_n18136_, new_n18137_, new_n18138_,
    new_n18139_, new_n18140_, new_n18141_, new_n18142_, new_n18143_,
    new_n18144_, new_n18145_, new_n18146_, new_n18147_, new_n18148_,
    new_n18149_, new_n18150_, new_n18151_, new_n18152_, new_n18153_,
    new_n18154_, new_n18155_, new_n18156_, new_n18157_, new_n18158_,
    new_n18159_, new_n18160_, new_n18161_, new_n18162_, new_n18163_,
    new_n18164_, new_n18165_, new_n18166_, new_n18167_, new_n18168_,
    new_n18169_, new_n18170_, new_n18171_, new_n18172_, new_n18173_,
    new_n18174_, new_n18175_, new_n18176_, new_n18177_, new_n18178_,
    new_n18179_, new_n18180_, new_n18181_, new_n18182_, new_n18183_,
    new_n18184_, new_n18185_, new_n18186_, new_n18187_, new_n18188_,
    new_n18189_, new_n18190_, new_n18191_, new_n18192_, new_n18193_,
    new_n18194_, new_n18195_, new_n18196_, new_n18197_, new_n18198_,
    new_n18199_, new_n18200_, new_n18201_, new_n18202_, new_n18203_,
    new_n18204_, new_n18205_, new_n18206_, new_n18207_, new_n18208_,
    new_n18209_, new_n18210_, new_n18211_, new_n18212_, new_n18213_,
    new_n18214_, new_n18215_, new_n18216_, new_n18217_, new_n18218_,
    new_n18219_, new_n18220_, new_n18221_, new_n18222_, new_n18223_,
    new_n18224_, new_n18225_, new_n18226_, new_n18227_, new_n18228_,
    new_n18229_, new_n18230_, new_n18231_, new_n18232_, new_n18233_,
    new_n18234_, new_n18235_, new_n18236_, new_n18237_, new_n18238_,
    new_n18239_, new_n18240_, new_n18241_, new_n18242_, new_n18243_,
    new_n18244_, new_n18245_, new_n18246_, new_n18247_, new_n18248_,
    new_n18249_, new_n18250_, new_n18251_, new_n18252_, new_n18253_,
    new_n18254_, new_n18255_, new_n18256_, new_n18257_, new_n18258_,
    new_n18259_, new_n18260_, new_n18261_, new_n18262_, new_n18263_,
    new_n18264_, new_n18265_, new_n18266_, new_n18267_, new_n18268_,
    new_n18269_, new_n18270_, new_n18271_, new_n18272_, new_n18273_,
    new_n18274_, new_n18275_, new_n18276_, new_n18277_, new_n18278_,
    new_n18279_, new_n18280_, new_n18281_, new_n18282_, new_n18283_,
    new_n18284_, new_n18285_, new_n18286_, new_n18287_, new_n18288_,
    new_n18289_, new_n18290_, new_n18291_, new_n18292_, new_n18293_,
    new_n18294_, new_n18295_, new_n18296_, new_n18297_, new_n18298_,
    new_n18299_, new_n18300_, new_n18301_, new_n18302_, new_n18303_,
    new_n18304_, new_n18305_, new_n18306_, new_n18307_, new_n18308_,
    new_n18309_, new_n18310_, new_n18311_, new_n18312_, new_n18313_,
    new_n18314_, new_n18315_, new_n18316_, new_n18317_, new_n18318_,
    new_n18319_, new_n18320_, new_n18321_, new_n18322_, new_n18323_,
    new_n18324_, new_n18325_, new_n18326_, new_n18327_, new_n18328_,
    new_n18329_, new_n18330_, new_n18331_, new_n18332_, new_n18333_,
    new_n18334_, new_n18335_, new_n18336_, new_n18337_, new_n18338_,
    new_n18339_, new_n18340_, new_n18341_, new_n18342_, new_n18343_,
    new_n18344_, new_n18345_, new_n18346_, new_n18347_, new_n18348_,
    new_n18349_, new_n18350_, new_n18351_, new_n18352_, new_n18353_,
    new_n18354_, new_n18355_, new_n18356_, new_n18357_, new_n18358_,
    new_n18359_, new_n18360_, new_n18361_, new_n18362_, new_n18363_,
    new_n18364_, new_n18365_, new_n18366_, new_n18367_, new_n18368_,
    new_n18369_, new_n18370_, new_n18371_, new_n18372_, new_n18373_,
    new_n18374_, new_n18375_, new_n18376_, new_n18377_, new_n18378_,
    new_n18379_, new_n18380_, new_n18381_, new_n18382_, new_n18383_,
    new_n18384_, new_n18385_, new_n18386_, new_n18387_, new_n18388_,
    new_n18389_, new_n18390_, new_n18391_, new_n18392_, new_n18393_,
    new_n18394_, new_n18395_, new_n18396_, new_n18397_, new_n18398_,
    new_n18399_, new_n18400_, new_n18401_, new_n18402_, new_n18403_,
    new_n18404_, new_n18405_, new_n18406_, new_n18407_, new_n18409_,
    new_n18410_, new_n18411_, new_n18412_, new_n18413_, new_n18414_,
    new_n18415_, new_n18416_, new_n18417_, new_n18418_, new_n18419_,
    new_n18420_, new_n18421_, new_n18422_, new_n18423_, new_n18424_,
    new_n18425_, new_n18426_, new_n18427_, new_n18428_, new_n18429_,
    new_n18430_, new_n18431_, new_n18432_, new_n18433_, new_n18434_,
    new_n18435_, new_n18436_, new_n18437_, new_n18438_, new_n18439_,
    new_n18440_, new_n18441_, new_n18442_, new_n18443_, new_n18444_,
    new_n18445_, new_n18446_, new_n18447_, new_n18448_, new_n18449_,
    new_n18450_, new_n18451_, new_n18452_, new_n18453_, new_n18454_,
    new_n18455_, new_n18456_, new_n18457_, new_n18458_, new_n18459_,
    new_n18460_, new_n18461_, new_n18462_, new_n18463_, new_n18464_,
    new_n18465_, new_n18466_, new_n18467_, new_n18468_, new_n18469_,
    new_n18470_, new_n18471_, new_n18472_, new_n18473_, new_n18474_,
    new_n18475_, new_n18476_, new_n18477_, new_n18478_, new_n18479_,
    new_n18480_, new_n18481_, new_n18482_, new_n18483_, new_n18484_,
    new_n18485_, new_n18486_, new_n18487_, new_n18488_, new_n18489_,
    new_n18490_, new_n18491_, new_n18492_, new_n18493_, new_n18494_,
    new_n18495_, new_n18496_, new_n18497_, new_n18498_, new_n18499_,
    new_n18500_, new_n18501_, new_n18502_, new_n18503_, new_n18504_,
    new_n18505_, new_n18506_, new_n18507_, new_n18508_, new_n18509_,
    new_n18510_, new_n18511_, new_n18512_, new_n18513_, new_n18514_,
    new_n18515_, new_n18516_, new_n18517_, new_n18518_, new_n18519_,
    new_n18520_, new_n18521_, new_n18522_, new_n18523_, new_n18524_,
    new_n18525_, new_n18526_, new_n18527_, new_n18528_, new_n18529_,
    new_n18530_, new_n18531_, new_n18532_, new_n18533_, new_n18534_,
    new_n18535_, new_n18536_, new_n18537_, new_n18538_, new_n18539_,
    new_n18540_, new_n18541_, new_n18542_, new_n18543_, new_n18544_,
    new_n18545_, new_n18546_, new_n18547_, new_n18548_, new_n18549_,
    new_n18550_, new_n18551_, new_n18552_, new_n18553_, new_n18554_,
    new_n18555_, new_n18556_, new_n18557_, new_n18558_, new_n18559_,
    new_n18560_, new_n18561_, new_n18562_, new_n18563_, new_n18564_,
    new_n18565_, new_n18566_, new_n18567_, new_n18568_, new_n18569_,
    new_n18570_, new_n18571_, new_n18572_, new_n18573_, new_n18574_,
    new_n18575_, new_n18576_, new_n18577_, new_n18578_, new_n18579_,
    new_n18580_, new_n18581_, new_n18582_, new_n18583_, new_n18584_,
    new_n18585_, new_n18586_, new_n18587_, new_n18588_, new_n18589_,
    new_n18590_, new_n18591_, new_n18592_, new_n18593_, new_n18594_,
    new_n18595_, new_n18596_, new_n18597_, new_n18598_, new_n18599_,
    new_n18600_, new_n18601_, new_n18602_, new_n18603_, new_n18604_,
    new_n18605_, new_n18606_, new_n18607_, new_n18608_, new_n18609_,
    new_n18610_, new_n18611_, new_n18612_, new_n18613_, new_n18614_,
    new_n18615_, new_n18616_, new_n18617_, new_n18618_, new_n18619_,
    new_n18620_, new_n18621_, new_n18622_, new_n18623_, new_n18624_,
    new_n18625_, new_n18626_, new_n18627_, new_n18628_, new_n18629_,
    new_n18630_, new_n18631_, new_n18632_, new_n18633_, new_n18634_,
    new_n18635_, new_n18636_, new_n18637_, new_n18638_, new_n18639_,
    new_n18640_, new_n18641_, new_n18642_, new_n18643_, new_n18644_,
    new_n18645_, new_n18646_, new_n18647_, new_n18648_, new_n18649_,
    new_n18650_, new_n18651_, new_n18652_, new_n18653_, new_n18654_,
    new_n18655_, new_n18656_, new_n18657_, new_n18658_, new_n18659_,
    new_n18660_, new_n18661_, new_n18662_, new_n18663_, new_n18664_,
    new_n18665_, new_n18666_, new_n18667_, new_n18668_, new_n18669_,
    new_n18670_, new_n18671_, new_n18672_, new_n18673_, new_n18674_,
    new_n18675_, new_n18676_, new_n18677_, new_n18678_, new_n18679_,
    new_n18680_, new_n18681_, new_n18682_, new_n18683_, new_n18684_,
    new_n18685_, new_n18686_, new_n18687_, new_n18688_, new_n18689_,
    new_n18690_, new_n18691_, new_n18692_, new_n18693_, new_n18694_,
    new_n18695_, new_n18696_, new_n18697_, new_n18698_, new_n18699_,
    new_n18700_, new_n18701_, new_n18702_, new_n18703_, new_n18704_,
    new_n18705_, new_n18706_, new_n18707_, new_n18708_, new_n18709_,
    new_n18710_, new_n18711_, new_n18712_, new_n18713_, new_n18714_,
    new_n18715_, new_n18716_, new_n18717_, new_n18718_, new_n18719_,
    new_n18720_, new_n18721_, new_n18722_, new_n18723_, new_n18724_,
    new_n18725_, new_n18726_, new_n18727_, new_n18728_, new_n18729_,
    new_n18730_, new_n18731_, new_n18732_, new_n18733_, new_n18734_,
    new_n18735_, new_n18736_, new_n18737_, new_n18738_, new_n18739_,
    new_n18740_, new_n18741_, new_n18742_, new_n18743_, new_n18744_,
    new_n18745_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18752_, new_n18753_, new_n18754_,
    new_n18755_, new_n18756_, new_n18757_, new_n18758_, new_n18759_,
    new_n18760_, new_n18761_, new_n18762_, new_n18763_, new_n18764_,
    new_n18765_, new_n18766_, new_n18767_, new_n18768_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18773_, new_n18774_,
    new_n18775_, new_n18776_, new_n18777_, new_n18778_, new_n18779_,
    new_n18780_, new_n18781_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18794_,
    new_n18795_, new_n18796_, new_n18797_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18951_, new_n18952_, new_n18953_, new_n18954_,
    new_n18955_, new_n18956_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18962_, new_n18963_, new_n18964_,
    new_n18965_, new_n18966_, new_n18967_, new_n18968_, new_n18969_,
    new_n18970_, new_n18971_, new_n18972_, new_n18973_, new_n18974_,
    new_n18975_, new_n18976_, new_n18977_, new_n18978_, new_n18979_,
    new_n18980_, new_n18981_, new_n18982_, new_n18983_, new_n18984_,
    new_n18985_, new_n18986_, new_n18987_, new_n18988_, new_n18989_,
    new_n18990_, new_n18991_, new_n18992_, new_n18993_, new_n18994_,
    new_n18995_, new_n18996_, new_n18997_, new_n18998_, new_n18999_,
    new_n19000_, new_n19001_, new_n19002_, new_n19003_, new_n19004_,
    new_n19005_, new_n19006_, new_n19007_, new_n19008_, new_n19009_,
    new_n19010_, new_n19011_, new_n19012_, new_n19013_, new_n19014_,
    new_n19015_, new_n19016_, new_n19017_, new_n19018_, new_n19019_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19107_, new_n19108_, new_n19109_, new_n19110_,
    new_n19111_, new_n19112_, new_n19113_, new_n19114_, new_n19115_,
    new_n19116_, new_n19117_, new_n19118_, new_n19119_, new_n19120_,
    new_n19121_, new_n19122_, new_n19123_, new_n19124_, new_n19125_,
    new_n19126_, new_n19127_, new_n19128_, new_n19129_, new_n19130_,
    new_n19131_, new_n19132_, new_n19133_, new_n19134_, new_n19135_,
    new_n19136_, new_n19137_, new_n19138_, new_n19139_, new_n19140_,
    new_n19141_, new_n19142_, new_n19143_, new_n19144_, new_n19145_,
    new_n19146_, new_n19147_, new_n19148_, new_n19149_, new_n19150_,
    new_n19151_, new_n19152_, new_n19153_, new_n19154_, new_n19155_,
    new_n19156_, new_n19157_, new_n19158_, new_n19159_, new_n19160_,
    new_n19161_, new_n19162_, new_n19163_, new_n19164_, new_n19165_,
    new_n19166_, new_n19167_, new_n19168_, new_n19169_, new_n19170_,
    new_n19171_, new_n19172_, new_n19173_, new_n19174_, new_n19175_,
    new_n19176_, new_n19177_, new_n19178_, new_n19179_, new_n19180_,
    new_n19181_, new_n19182_, new_n19183_, new_n19184_, new_n19185_,
    new_n19186_, new_n19187_, new_n19188_, new_n19189_, new_n19190_,
    new_n19191_, new_n19192_, new_n19193_, new_n19194_, new_n19195_,
    new_n19196_, new_n19197_, new_n19198_, new_n19199_, new_n19200_,
    new_n19201_, new_n19202_, new_n19203_, new_n19204_, new_n19205_,
    new_n19206_, new_n19207_, new_n19208_, new_n19209_, new_n19210_,
    new_n19211_, new_n19212_, new_n19213_, new_n19214_, new_n19215_,
    new_n19216_, new_n19217_, new_n19218_, new_n19219_, new_n19220_,
    new_n19221_, new_n19222_, new_n19223_, new_n19224_, new_n19225_,
    new_n19226_, new_n19227_, new_n19228_, new_n19229_, new_n19230_,
    new_n19231_, new_n19232_, new_n19233_, new_n19234_, new_n19235_,
    new_n19236_, new_n19237_, new_n19238_, new_n19239_, new_n19240_,
    new_n19241_, new_n19242_, new_n19243_, new_n19244_, new_n19245_,
    new_n19246_, new_n19247_, new_n19248_, new_n19249_, new_n19250_,
    new_n19251_, new_n19252_, new_n19253_, new_n19254_, new_n19255_,
    new_n19256_, new_n19257_, new_n19258_, new_n19259_, new_n19260_,
    new_n19261_, new_n19262_, new_n19263_, new_n19264_, new_n19265_,
    new_n19266_, new_n19267_, new_n19268_, new_n19269_, new_n19270_,
    new_n19271_, new_n19272_, new_n19273_, new_n19274_, new_n19275_,
    new_n19276_, new_n19277_, new_n19278_, new_n19279_, new_n19280_,
    new_n19281_, new_n19282_, new_n19283_, new_n19284_, new_n19285_,
    new_n19286_, new_n19287_, new_n19288_, new_n19289_, new_n19290_,
    new_n19291_, new_n19292_, new_n19293_, new_n19294_, new_n19295_,
    new_n19296_, new_n19297_, new_n19298_, new_n19299_, new_n19300_,
    new_n19301_, new_n19302_, new_n19303_, new_n19304_, new_n19305_,
    new_n19306_, new_n19307_, new_n19308_, new_n19309_, new_n19310_,
    new_n19311_, new_n19312_, new_n19313_, new_n19314_, new_n19315_,
    new_n19316_, new_n19317_, new_n19318_, new_n19319_, new_n19320_,
    new_n19321_, new_n19322_, new_n19323_, new_n19324_, new_n19325_,
    new_n19326_, new_n19327_, new_n19328_, new_n19329_, new_n19330_,
    new_n19331_, new_n19332_, new_n19333_, new_n19334_, new_n19335_,
    new_n19336_, new_n19337_, new_n19338_, new_n19339_, new_n19340_,
    new_n19341_, new_n19342_, new_n19343_, new_n19344_, new_n19345_,
    new_n19346_, new_n19347_, new_n19348_, new_n19349_, new_n19350_,
    new_n19351_, new_n19352_, new_n19353_, new_n19354_, new_n19355_,
    new_n19356_, new_n19357_, new_n19358_, new_n19359_, new_n19360_,
    new_n19361_, new_n19362_, new_n19363_, new_n19364_, new_n19365_,
    new_n19366_, new_n19367_, new_n19368_, new_n19369_, new_n19370_,
    new_n19371_, new_n19372_, new_n19373_, new_n19374_, new_n19375_,
    new_n19376_, new_n19377_, new_n19378_, new_n19379_, new_n19380_,
    new_n19381_, new_n19382_, new_n19383_, new_n19384_, new_n19385_,
    new_n19386_, new_n19387_, new_n19388_, new_n19389_, new_n19390_,
    new_n19391_, new_n19392_, new_n19393_, new_n19394_, new_n19395_,
    new_n19396_, new_n19397_, new_n19398_, new_n19399_, new_n19400_,
    new_n19401_, new_n19402_, new_n19403_, new_n19404_, new_n19405_,
    new_n19406_, new_n19407_, new_n19408_, new_n19409_, new_n19410_,
    new_n19411_, new_n19412_, new_n19413_, new_n19414_, new_n19415_,
    new_n19416_, new_n19417_, new_n19418_, new_n19419_, new_n19420_,
    new_n19421_, new_n19422_, new_n19423_, new_n19424_, new_n19425_,
    new_n19426_, new_n19427_, new_n19428_, new_n19429_, new_n19430_,
    new_n19431_, new_n19432_, new_n19433_, new_n19434_, new_n19435_,
    new_n19436_, new_n19437_, new_n19438_, new_n19439_, new_n19440_,
    new_n19441_, new_n19442_, new_n19443_, new_n19444_, new_n19445_,
    new_n19446_, new_n19447_, new_n19448_, new_n19449_, new_n19450_,
    new_n19451_, new_n19452_, new_n19453_, new_n19454_, new_n19455_,
    new_n19456_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19513_, new_n19514_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19640_, new_n19641_,
    new_n19642_, new_n19643_, new_n19644_, new_n19645_, new_n19646_,
    new_n19647_, new_n19648_, new_n19649_, new_n19650_, new_n19651_,
    new_n19652_, new_n19653_, new_n19654_, new_n19655_, new_n19656_,
    new_n19657_, new_n19658_, new_n19659_, new_n19660_, new_n19661_,
    new_n19662_, new_n19663_, new_n19664_, new_n19665_, new_n19666_,
    new_n19667_, new_n19668_, new_n19669_, new_n19670_, new_n19671_,
    new_n19672_, new_n19673_, new_n19674_, new_n19675_, new_n19676_,
    new_n19677_, new_n19678_, new_n19679_, new_n19680_, new_n19681_,
    new_n19682_, new_n19683_, new_n19684_, new_n19685_, new_n19686_,
    new_n19687_, new_n19688_, new_n19689_, new_n19690_, new_n19691_,
    new_n19692_, new_n19693_, new_n19694_, new_n19695_, new_n19696_,
    new_n19697_, new_n19698_, new_n19699_, new_n19700_, new_n19701_,
    new_n19702_, new_n19703_, new_n19704_, new_n19705_, new_n19706_,
    new_n19707_, new_n19708_, new_n19709_, new_n19710_, new_n19711_,
    new_n19712_, new_n19713_, new_n19714_, new_n19715_, new_n19716_,
    new_n19717_, new_n19718_, new_n19719_, new_n19720_, new_n19721_,
    new_n19722_, new_n19723_, new_n19724_, new_n19725_, new_n19726_,
    new_n19727_, new_n19728_, new_n19729_, new_n19730_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19842_, new_n19843_, new_n19844_, new_n19845_, new_n19846_,
    new_n19847_, new_n19848_, new_n19849_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20153_, new_n20154_, new_n20155_, new_n20156_,
    new_n20157_, new_n20158_, new_n20159_, new_n20160_, new_n20161_,
    new_n20162_, new_n20163_, new_n20164_, new_n20165_, new_n20166_,
    new_n20167_, new_n20168_, new_n20169_, new_n20170_, new_n20171_,
    new_n20172_, new_n20173_, new_n20174_, new_n20175_, new_n20176_,
    new_n20177_, new_n20178_, new_n20179_, new_n20180_, new_n20181_,
    new_n20182_, new_n20183_, new_n20184_, new_n20185_, new_n20186_,
    new_n20187_, new_n20188_, new_n20189_, new_n20190_, new_n20191_,
    new_n20192_, new_n20193_, new_n20194_, new_n20195_, new_n20196_,
    new_n20197_, new_n20198_, new_n20199_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20247_,
    new_n20248_, new_n20249_, new_n20250_, new_n20251_, new_n20252_,
    new_n20253_, new_n20254_, new_n20255_, new_n20256_, new_n20257_,
    new_n20258_, new_n20259_, new_n20260_, new_n20261_, new_n20262_,
    new_n20263_, new_n20264_, new_n20265_, new_n20266_, new_n20267_,
    new_n20268_, new_n20269_, new_n20270_, new_n20271_, new_n20272_,
    new_n20273_, new_n20274_, new_n20275_, new_n20276_, new_n20277_,
    new_n20278_, new_n20279_, new_n20280_, new_n20281_, new_n20282_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20290_, new_n20291_, new_n20292_,
    new_n20293_, new_n20294_, new_n20295_, new_n20296_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20376_, new_n20377_,
    new_n20378_, new_n20379_, new_n20380_, new_n20381_, new_n20382_,
    new_n20383_, new_n20384_, new_n20385_, new_n20386_, new_n20387_,
    new_n20388_, new_n20389_, new_n20390_, new_n20391_, new_n20392_,
    new_n20393_, new_n20394_, new_n20395_, new_n20396_, new_n20397_,
    new_n20398_, new_n20399_, new_n20400_, new_n20401_, new_n20402_,
    new_n20403_, new_n20404_, new_n20405_, new_n20406_, new_n20407_,
    new_n20408_, new_n20409_, new_n20410_, new_n20411_, new_n20412_,
    new_n20413_, new_n20414_, new_n20415_, new_n20416_, new_n20417_,
    new_n20418_, new_n20419_, new_n20420_, new_n20421_, new_n20422_,
    new_n20423_, new_n20424_, new_n20425_, new_n20426_, new_n20427_,
    new_n20428_, new_n20429_, new_n20430_, new_n20431_, new_n20432_,
    new_n20433_, new_n20434_, new_n20435_, new_n20436_, new_n20437_,
    new_n20438_, new_n20439_, new_n20440_, new_n20441_, new_n20442_,
    new_n20443_, new_n20444_, new_n20445_, new_n20446_, new_n20447_,
    new_n20448_, new_n20449_, new_n20450_, new_n20451_, new_n20452_,
    new_n20453_, new_n20454_, new_n20455_, new_n20456_, new_n20457_,
    new_n20458_, new_n20459_, new_n20460_, new_n20461_, new_n20462_,
    new_n20463_, new_n20464_, new_n20465_, new_n20466_, new_n20467_,
    new_n20468_, new_n20469_, new_n20470_, new_n20471_, new_n20472_,
    new_n20473_, new_n20474_, new_n20475_, new_n20476_, new_n20477_,
    new_n20478_, new_n20479_, new_n20480_, new_n20481_, new_n20482_,
    new_n20483_, new_n20484_, new_n20485_, new_n20486_, new_n20487_,
    new_n20488_, new_n20489_, new_n20490_, new_n20491_, new_n20492_,
    new_n20493_, new_n20494_, new_n20495_, new_n20496_, new_n20497_,
    new_n20498_, new_n20499_, new_n20500_, new_n20501_, new_n20502_,
    new_n20503_, new_n20504_, new_n20505_, new_n20506_, new_n20507_,
    new_n20508_, new_n20509_, new_n20510_, new_n20511_, new_n20512_,
    new_n20513_, new_n20514_, new_n20515_, new_n20516_, new_n20517_,
    new_n20518_, new_n20519_, new_n20520_, new_n20521_, new_n20522_,
    new_n20523_, new_n20524_, new_n20525_, new_n20526_, new_n20527_,
    new_n20528_, new_n20529_, new_n20530_, new_n20531_, new_n20532_,
    new_n20533_, new_n20534_, new_n20535_, new_n20536_, new_n20537_,
    new_n20538_, new_n20539_, new_n20540_, new_n20541_, new_n20542_,
    new_n20543_, new_n20544_, new_n20545_, new_n20546_, new_n20547_,
    new_n20548_, new_n20549_, new_n20550_, new_n20551_, new_n20552_,
    new_n20553_, new_n20554_, new_n20555_, new_n20556_, new_n20557_,
    new_n20558_, new_n20559_, new_n20560_, new_n20561_, new_n20562_,
    new_n20563_, new_n20564_, new_n20565_, new_n20566_, new_n20567_,
    new_n20568_, new_n20569_, new_n20570_, new_n20571_, new_n20572_,
    new_n20573_, new_n20574_, new_n20575_, new_n20576_, new_n20577_,
    new_n20578_, new_n20579_, new_n20580_, new_n20581_, new_n20582_,
    new_n20583_, new_n20584_, new_n20585_, new_n20586_, new_n20587_,
    new_n20588_, new_n20589_, new_n20590_, new_n20591_, new_n20592_,
    new_n20593_, new_n20594_, new_n20595_, new_n20596_, new_n20597_,
    new_n20598_, new_n20599_, new_n20600_, new_n20601_, new_n20602_,
    new_n20603_, new_n20604_, new_n20605_, new_n20606_, new_n20607_,
    new_n20608_, new_n20609_, new_n20610_, new_n20611_, new_n20612_,
    new_n20613_, new_n20614_, new_n20615_, new_n20616_, new_n20617_,
    new_n20618_, new_n20619_, new_n20620_, new_n20621_, new_n20622_,
    new_n20623_, new_n20624_, new_n20625_, new_n20626_, new_n20627_,
    new_n20628_, new_n20629_, new_n20630_, new_n20631_, new_n20632_,
    new_n20633_, new_n20634_, new_n20635_, new_n20636_, new_n20637_,
    new_n20638_, new_n20639_, new_n20640_, new_n20641_, new_n20642_,
    new_n20643_, new_n20644_, new_n20645_, new_n20646_, new_n20647_,
    new_n20648_, new_n20649_, new_n20650_, new_n20651_, new_n20652_;
  NOR2_X1    g00000(.A1(\a[126] ), .A2(\a[127] ), .ZN(new_n193_));
  INV_X1     g00001(.I(new_n193_), .ZN(\asqrt[63] ));
  INV_X1     g00002(.I(\a[64] ), .ZN(new_n195_));
  INV_X1     g00003(.I(\a[65] ), .ZN(new_n196_));
  INV_X1     g00004(.I(\a[96] ), .ZN(new_n197_));
  INV_X1     g00005(.I(\a[97] ), .ZN(new_n198_));
  INV_X1     g00006(.I(\a[112] ), .ZN(new_n199_));
  INV_X1     g00007(.I(\a[113] ), .ZN(new_n200_));
  INV_X1     g00008(.I(\a[120] ), .ZN(new_n201_));
  INV_X1     g00009(.I(\a[121] ), .ZN(new_n202_));
  INV_X1     g00010(.I(\a[127] ), .ZN(new_n203_));
  INV_X1     g00011(.I(\a[124] ), .ZN(new_n204_));
  INV_X1     g00012(.I(\a[125] ), .ZN(new_n205_));
  AOI21_X1   g00013(.A1(new_n204_), .A2(new_n205_), .B(\a[126] ), .ZN(new_n206_));
  INV_X1     g00014(.I(\a[126] ), .ZN(new_n207_));
  NOR3_X1    g00015(.A1(new_n207_), .A2(\a[124] ), .A3(\a[125] ), .ZN(new_n208_));
  NOR3_X1    g00016(.A1(new_n206_), .A2(new_n208_), .A3(new_n203_), .ZN(new_n209_));
  NAND2_X1   g00017(.A1(\a[124] ), .A2(\a[125] ), .ZN(new_n210_));
  INV_X1     g00018(.I(new_n210_), .ZN(new_n211_));
  OAI21_X1   g00019(.A1(\a[124] ), .A2(\a[125] ), .B(\a[127] ), .ZN(new_n212_));
  OAI21_X1   g00020(.A1(\a[125] ), .A2(\a[127] ), .B(\a[126] ), .ZN(new_n213_));
  INV_X1     g00021(.I(new_n213_), .ZN(new_n214_));
  AOI21_X1   g00022(.A1(new_n214_), .A2(new_n212_), .B(new_n211_), .ZN(new_n215_));
  NAND2_X1   g00023(.A1(new_n203_), .A2(\a[126] ), .ZN(new_n216_));
  NOR3_X1    g00024(.A1(\a[122] ), .A2(\a[123] ), .A3(\a[124] ), .ZN(new_n217_));
  AOI21_X1   g00025(.A1(new_n216_), .A2(\a[124] ), .B(new_n217_), .ZN(new_n218_));
  NOR2_X1    g00026(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1     g00027(.I(new_n219_), .ZN(new_n220_));
  NOR3_X1    g00028(.A1(new_n220_), .A2(new_n193_), .A3(new_n209_), .ZN(new_n221_));
  INV_X1     g00029(.I(new_n221_), .ZN(new_n222_));
  OAI21_X1   g00030(.A1(\a[124] ), .A2(\a[125] ), .B(new_n207_), .ZN(new_n223_));
  NOR2_X1    g00031(.A1(\a[124] ), .A2(\a[125] ), .ZN(new_n224_));
  NAND2_X1   g00032(.A1(new_n224_), .A2(\a[126] ), .ZN(new_n225_));
  NAND3_X1   g00033(.A1(new_n223_), .A2(new_n225_), .A3(\a[127] ), .ZN(new_n226_));
  INV_X1     g00034(.I(new_n212_), .ZN(new_n227_));
  OAI21_X1   g00035(.A1(new_n227_), .A2(new_n213_), .B(new_n210_), .ZN(new_n228_));
  OAI21_X1   g00036(.A1(new_n207_), .A2(\a[127] ), .B(\a[124] ), .ZN(new_n229_));
  OR3_X2     g00037(.A1(\a[122] ), .A2(\a[123] ), .A3(\a[124] ), .Z(new_n230_));
  NAND2_X1   g00038(.A1(new_n230_), .A2(new_n229_), .ZN(new_n231_));
  NOR3_X1    g00039(.A1(new_n226_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n232_));
  OAI21_X1   g00040(.A1(new_n232_), .A2(new_n219_), .B(\asqrt[63] ), .ZN(new_n233_));
  AOI21_X1   g00041(.A1(\a[126] ), .A2(\a[127] ), .B(new_n206_), .ZN(new_n234_));
  OAI21_X1   g00042(.A1(new_n228_), .A2(new_n218_), .B(new_n193_), .ZN(new_n235_));
  NAND2_X1   g00043(.A1(new_n228_), .A2(new_n218_), .ZN(new_n236_));
  NAND3_X1   g00044(.A1(new_n235_), .A2(new_n236_), .A3(new_n226_), .ZN(new_n237_));
  NOR2_X1    g00045(.A1(new_n237_), .A2(new_n234_), .ZN(new_n238_));
  AOI21_X1   g00046(.A1(new_n215_), .A2(new_n231_), .B(\asqrt[63] ), .ZN(new_n239_));
  NAND3_X1   g00047(.A1(new_n214_), .A2(new_n230_), .A3(new_n212_), .ZN(new_n240_));
  NAND2_X1   g00048(.A1(new_n226_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1    g00049(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NOR3_X1    g00050(.A1(new_n242_), .A2(\a[122] ), .A3(\a[123] ), .ZN(new_n243_));
  OAI21_X1   g00051(.A1(new_n243_), .A2(new_n238_), .B(new_n204_), .ZN(new_n244_));
  INV_X1     g00052(.I(new_n234_), .ZN(\asqrt[62] ));
  NOR2_X1    g00053(.A1(new_n215_), .A2(new_n231_), .ZN(new_n246_));
  NOR3_X1    g00054(.A1(new_n239_), .A2(new_n246_), .A3(new_n209_), .ZN(new_n247_));
  NAND2_X1   g00055(.A1(new_n247_), .A2(\asqrt[62] ), .ZN(new_n248_));
  NOR2_X1    g00056(.A1(\a[122] ), .A2(\a[123] ), .ZN(new_n249_));
  NOR3_X1    g00057(.A1(new_n227_), .A2(new_n213_), .A3(new_n217_), .ZN(new_n250_));
  NOR2_X1    g00058(.A1(new_n250_), .A2(new_n209_), .ZN(new_n251_));
  NAND2_X1   g00059(.A1(new_n235_), .A2(new_n251_), .ZN(\asqrt[61] ));
  NAND2_X1   g00060(.A1(\asqrt[61] ), .A2(new_n249_), .ZN(new_n253_));
  NAND3_X1   g00061(.A1(new_n248_), .A2(new_n253_), .A3(\a[124] ), .ZN(new_n254_));
  NAND2_X1   g00062(.A1(new_n244_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1    g00063(.A1(\a[120] ), .A2(\a[121] ), .ZN(new_n256_));
  NOR2_X1    g00064(.A1(new_n256_), .A2(\a[122] ), .ZN(new_n257_));
  INV_X1     g00065(.I(new_n257_), .ZN(new_n258_));
  NAND3_X1   g00066(.A1(new_n235_), .A2(new_n251_), .A3(\a[122] ), .ZN(new_n259_));
  NAND3_X1   g00067(.A1(new_n259_), .A2(\asqrt[62] ), .A3(new_n258_), .ZN(new_n260_));
  INV_X1     g00068(.I(new_n260_), .ZN(new_n261_));
  NAND2_X1   g00069(.A1(new_n259_), .A2(new_n258_), .ZN(new_n262_));
  INV_X1     g00070(.I(\a[123] ), .ZN(new_n263_));
  OAI21_X1   g00071(.A1(new_n242_), .A2(\a[122] ), .B(new_n263_), .ZN(new_n264_));
  INV_X1     g00072(.I(\a[122] ), .ZN(new_n265_));
  NAND3_X1   g00073(.A1(\asqrt[61] ), .A2(new_n265_), .A3(\a[123] ), .ZN(new_n266_));
  AOI22_X1   g00074(.A1(new_n264_), .A2(new_n266_), .B1(new_n262_), .B2(new_n234_), .ZN(new_n267_));
  NOR2_X1    g00075(.A1(new_n228_), .A2(new_n218_), .ZN(new_n268_));
  AOI21_X1   g00076(.A1(\asqrt[61] ), .A2(new_n268_), .B(new_n246_), .ZN(new_n269_));
  OAI21_X1   g00077(.A1(new_n267_), .A2(new_n261_), .B(new_n269_), .ZN(new_n270_));
  OAI21_X1   g00078(.A1(new_n270_), .A2(new_n255_), .B(new_n193_), .ZN(new_n271_));
  AOI21_X1   g00079(.A1(\asqrt[61] ), .A2(new_n265_), .B(\a[123] ), .ZN(new_n272_));
  NOR3_X1    g00080(.A1(new_n242_), .A2(\a[122] ), .A3(new_n263_), .ZN(new_n273_));
  NOR3_X1    g00081(.A1(new_n239_), .A2(new_n241_), .A3(new_n265_), .ZN(new_n274_));
  OAI21_X1   g00082(.A1(new_n274_), .A2(new_n257_), .B(new_n234_), .ZN(new_n275_));
  OAI21_X1   g00083(.A1(new_n272_), .A2(new_n273_), .B(new_n275_), .ZN(new_n276_));
  NAND3_X1   g00084(.A1(new_n255_), .A2(new_n260_), .A3(new_n276_), .ZN(new_n277_));
  NAND4_X1   g00085(.A1(new_n271_), .A2(new_n222_), .A3(new_n233_), .A4(new_n277_), .ZN(\asqrt[60] ));
  AOI21_X1   g00086(.A1(\asqrt[60] ), .A2(new_n201_), .B(new_n202_), .ZN(new_n279_));
  INV_X1     g00087(.I(new_n233_), .ZN(new_n280_));
  AOI21_X1   g00088(.A1(new_n248_), .A2(new_n253_), .B(\a[124] ), .ZN(new_n281_));
  NOR3_X1    g00089(.A1(new_n243_), .A2(new_n238_), .A3(new_n204_), .ZN(new_n282_));
  NOR2_X1    g00090(.A1(new_n282_), .A2(new_n281_), .ZN(new_n283_));
  INV_X1     g00091(.I(new_n269_), .ZN(new_n284_));
  AOI21_X1   g00092(.A1(new_n276_), .A2(new_n260_), .B(new_n284_), .ZN(new_n285_));
  AOI21_X1   g00093(.A1(new_n285_), .A2(new_n283_), .B(\asqrt[63] ), .ZN(new_n286_));
  NOR3_X1    g00094(.A1(new_n283_), .A2(new_n261_), .A3(new_n267_), .ZN(new_n287_));
  NOR4_X1    g00095(.A1(new_n286_), .A2(new_n221_), .A3(new_n280_), .A4(new_n287_), .ZN(new_n288_));
  NOR3_X1    g00096(.A1(new_n288_), .A2(\a[120] ), .A3(\a[121] ), .ZN(new_n289_));
  NOR2_X1    g00097(.A1(new_n289_), .A2(new_n279_), .ZN(new_n290_));
  NAND2_X1   g00098(.A1(\asqrt[60] ), .A2(\a[120] ), .ZN(new_n291_));
  INV_X1     g00099(.I(\a[118] ), .ZN(new_n292_));
  INV_X1     g00100(.I(\a[119] ), .ZN(new_n293_));
  NAND3_X1   g00101(.A1(new_n292_), .A2(new_n293_), .A3(new_n201_), .ZN(new_n294_));
  AOI21_X1   g00102(.A1(new_n291_), .A2(new_n294_), .B(new_n242_), .ZN(new_n295_));
  OAI21_X1   g00103(.A1(new_n288_), .A2(new_n201_), .B(new_n294_), .ZN(new_n296_));
  NOR2_X1    g00104(.A1(new_n296_), .A2(new_n237_), .ZN(new_n297_));
  NOR2_X1    g00105(.A1(new_n267_), .A2(new_n261_), .ZN(new_n298_));
  NOR2_X1    g00106(.A1(new_n298_), .A2(new_n283_), .ZN(new_n299_));
  INV_X1     g00107(.I(new_n299_), .ZN(new_n300_));
  NAND3_X1   g00108(.A1(\asqrt[60] ), .A2(new_n283_), .A3(new_n298_), .ZN(new_n301_));
  AOI21_X1   g00109(.A1(new_n301_), .A2(new_n300_), .B(new_n193_), .ZN(new_n302_));
  NOR2_X1    g00110(.A1(new_n273_), .A2(new_n272_), .ZN(new_n303_));
  INV_X1     g00111(.I(new_n303_), .ZN(new_n304_));
  NAND2_X1   g00112(.A1(new_n275_), .A2(new_n260_), .ZN(new_n305_));
  INV_X1     g00113(.I(new_n305_), .ZN(new_n306_));
  NAND2_X1   g00114(.A1(\asqrt[60] ), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1    g00115(.A1(new_n307_), .A2(new_n304_), .Z(new_n308_));
  OAI21_X1   g00116(.A1(new_n261_), .A2(new_n267_), .B(\asqrt[60] ), .ZN(new_n309_));
  AOI21_X1   g00117(.A1(new_n309_), .A2(new_n283_), .B(new_n299_), .ZN(new_n310_));
  NOR2_X1    g00118(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1   g00119(.A1(new_n288_), .A2(\a[120] ), .B(\a[121] ), .ZN(new_n312_));
  NAND3_X1   g00120(.A1(\asqrt[60] ), .A2(new_n201_), .A3(new_n202_), .ZN(new_n313_));
  NAND2_X1   g00121(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1   g00122(.A1(new_n296_), .A2(\asqrt[61] ), .ZN(new_n315_));
  OAI21_X1   g00123(.A1(new_n314_), .A2(new_n297_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1   g00124(.A1(new_n316_), .A2(\asqrt[62] ), .ZN(new_n317_));
  NAND2_X1   g00125(.A1(\asqrt[60] ), .A2(new_n256_), .ZN(new_n318_));
  NAND4_X1   g00126(.A1(new_n271_), .A2(new_n233_), .A3(\asqrt[61] ), .A4(new_n277_), .ZN(new_n319_));
  AOI21_X1   g00127(.A1(new_n318_), .A2(new_n319_), .B(\a[122] ), .ZN(new_n320_));
  INV_X1     g00128(.I(new_n256_), .ZN(new_n321_));
  NOR2_X1    g00129(.A1(new_n288_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1     g00130(.I(new_n319_), .ZN(new_n323_));
  NOR3_X1    g00131(.A1(new_n322_), .A2(new_n265_), .A3(new_n323_), .ZN(new_n324_));
  NOR2_X1    g00132(.A1(new_n324_), .A2(new_n320_), .ZN(new_n325_));
  OAI21_X1   g00133(.A1(new_n316_), .A2(\asqrt[62] ), .B(new_n325_), .ZN(new_n326_));
  NAND2_X1   g00134(.A1(new_n326_), .A2(new_n317_), .ZN(new_n327_));
  AOI21_X1   g00135(.A1(new_n327_), .A2(new_n311_), .B(\asqrt[63] ), .ZN(new_n328_));
  INV_X1     g00136(.I(new_n308_), .ZN(new_n329_));
  NAND3_X1   g00137(.A1(new_n291_), .A2(new_n247_), .A3(new_n294_), .ZN(new_n330_));
  AOI21_X1   g00138(.A1(new_n290_), .A2(new_n330_), .B(new_n295_), .ZN(new_n331_));
  NOR2_X1    g00139(.A1(new_n331_), .A2(new_n234_), .ZN(new_n332_));
  OAI21_X1   g00140(.A1(new_n322_), .A2(new_n323_), .B(new_n265_), .ZN(new_n333_));
  NAND3_X1   g00141(.A1(new_n318_), .A2(\a[122] ), .A3(new_n319_), .ZN(new_n334_));
  NAND2_X1   g00142(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1   g00143(.A1(new_n331_), .A2(new_n234_), .B(new_n335_), .ZN(new_n336_));
  NOR3_X1    g00144(.A1(new_n336_), .A2(new_n332_), .A3(new_n329_), .ZN(new_n337_));
  NOR2_X1    g00145(.A1(\asqrt[60] ), .A2(new_n283_), .ZN(new_n338_));
  NOR4_X1    g00146(.A1(new_n328_), .A2(new_n302_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  NOR3_X1    g00147(.A1(new_n339_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n340_));
  XOR2_X1    g00148(.A1(new_n340_), .A2(new_n290_), .Z(new_n341_));
  INV_X1     g00149(.I(\a[116] ), .ZN(new_n342_));
  INV_X1     g00150(.I(\a[117] ), .ZN(new_n343_));
  NAND3_X1   g00151(.A1(new_n342_), .A2(new_n343_), .A3(new_n292_), .ZN(new_n344_));
  OAI21_X1   g00152(.A1(new_n339_), .A2(new_n292_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1   g00153(.A1(new_n345_), .A2(\asqrt[60] ), .ZN(new_n346_));
  INV_X1     g00154(.I(new_n302_), .ZN(new_n347_));
  OAI21_X1   g00155(.A1(new_n336_), .A2(new_n332_), .B(new_n311_), .ZN(new_n348_));
  NAND2_X1   g00156(.A1(new_n348_), .A2(new_n193_), .ZN(new_n349_));
  NAND3_X1   g00157(.A1(new_n326_), .A2(new_n317_), .A3(new_n308_), .ZN(new_n350_));
  INV_X1     g00158(.I(new_n338_), .ZN(new_n351_));
  NAND4_X1   g00159(.A1(new_n349_), .A2(new_n347_), .A3(new_n350_), .A4(new_n351_), .ZN(\asqrt[59] ));
  NAND3_X1   g00160(.A1(\asqrt[59] ), .A2(new_n292_), .A3(new_n293_), .ZN(new_n353_));
  OAI21_X1   g00161(.A1(new_n339_), .A2(\a[118] ), .B(\a[119] ), .ZN(new_n354_));
  NAND2_X1   g00162(.A1(\asqrt[59] ), .A2(\a[118] ), .ZN(new_n355_));
  NAND3_X1   g00163(.A1(new_n355_), .A2(new_n288_), .A3(new_n344_), .ZN(new_n356_));
  NAND3_X1   g00164(.A1(new_n356_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n357_));
  AOI21_X1   g00165(.A1(new_n357_), .A2(new_n346_), .B(new_n242_), .ZN(new_n358_));
  NOR4_X1    g00166(.A1(new_n328_), .A2(new_n288_), .A3(new_n337_), .A4(new_n302_), .ZN(new_n359_));
  INV_X1     g00167(.I(new_n359_), .ZN(new_n360_));
  AOI21_X1   g00168(.A1(new_n353_), .A2(new_n360_), .B(\a[120] ), .ZN(new_n361_));
  NOR3_X1    g00169(.A1(new_n339_), .A2(\a[118] ), .A3(\a[119] ), .ZN(new_n362_));
  NOR3_X1    g00170(.A1(new_n362_), .A2(new_n201_), .A3(new_n359_), .ZN(new_n363_));
  NOR2_X1    g00171(.A1(new_n363_), .A2(new_n361_), .ZN(new_n364_));
  INV_X1     g00172(.I(new_n364_), .ZN(new_n365_));
  NAND2_X1   g00173(.A1(new_n354_), .A2(new_n353_), .ZN(new_n366_));
  NOR2_X1    g00174(.A1(new_n345_), .A2(\asqrt[60] ), .ZN(new_n367_));
  OAI21_X1   g00175(.A1(new_n366_), .A2(new_n367_), .B(new_n346_), .ZN(new_n368_));
  NOR2_X1    g00176(.A1(new_n368_), .A2(\asqrt[61] ), .ZN(new_n369_));
  NOR2_X1    g00177(.A1(new_n369_), .A2(new_n365_), .ZN(new_n370_));
  OAI21_X1   g00178(.A1(new_n370_), .A2(new_n358_), .B(\asqrt[62] ), .ZN(new_n371_));
  NAND2_X1   g00179(.A1(new_n368_), .A2(\asqrt[61] ), .ZN(new_n372_));
  OAI21_X1   g00180(.A1(new_n368_), .A2(\asqrt[61] ), .B(new_n364_), .ZN(new_n373_));
  NAND3_X1   g00181(.A1(new_n373_), .A2(new_n372_), .A3(new_n234_), .ZN(new_n374_));
  OAI21_X1   g00182(.A1(new_n339_), .A2(new_n327_), .B(new_n329_), .ZN(new_n375_));
  NAND3_X1   g00183(.A1(new_n375_), .A2(\asqrt[63] ), .A3(new_n350_), .ZN(new_n376_));
  NAND2_X1   g00184(.A1(new_n331_), .A2(new_n234_), .ZN(new_n377_));
  NAND3_X1   g00185(.A1(\asqrt[59] ), .A2(new_n317_), .A3(new_n377_), .ZN(new_n378_));
  XOR2_X1    g00186(.A1(new_n378_), .A2(new_n325_), .Z(new_n379_));
  NAND3_X1   g00187(.A1(new_n357_), .A2(new_n242_), .A3(new_n346_), .ZN(new_n380_));
  AOI21_X1   g00188(.A1(new_n364_), .A2(new_n380_), .B(new_n358_), .ZN(new_n381_));
  NOR2_X1    g00189(.A1(new_n381_), .A2(new_n234_), .ZN(new_n382_));
  NOR2_X1    g00190(.A1(new_n339_), .A2(new_n308_), .ZN(new_n383_));
  AOI21_X1   g00191(.A1(new_n383_), .A2(new_n327_), .B(new_n337_), .ZN(new_n384_));
  INV_X1     g00192(.I(new_n341_), .ZN(new_n385_));
  AOI21_X1   g00193(.A1(new_n381_), .A2(new_n234_), .B(new_n385_), .ZN(new_n386_));
  OAI21_X1   g00194(.A1(new_n386_), .A2(new_n382_), .B(new_n384_), .ZN(new_n387_));
  OAI21_X1   g00195(.A1(new_n387_), .A2(new_n379_), .B(new_n193_), .ZN(new_n388_));
  NAND2_X1   g00196(.A1(new_n374_), .A2(new_n341_), .ZN(new_n389_));
  NAND3_X1   g00197(.A1(new_n389_), .A2(new_n371_), .A3(new_n379_), .ZN(new_n390_));
  NOR2_X1    g00198(.A1(\asqrt[59] ), .A2(new_n329_), .ZN(new_n391_));
  INV_X1     g00199(.I(new_n391_), .ZN(new_n392_));
  NAND4_X1   g00200(.A1(new_n388_), .A2(new_n376_), .A3(new_n390_), .A4(new_n392_), .ZN(\asqrt[58] ));
  NAND3_X1   g00201(.A1(\asqrt[58] ), .A2(new_n371_), .A3(new_n374_), .ZN(new_n394_));
  XOR2_X1    g00202(.A1(new_n394_), .A2(new_n341_), .Z(new_n395_));
  INV_X1     g00203(.I(new_n395_), .ZN(new_n396_));
  INV_X1     g00204(.I(new_n376_), .ZN(new_n397_));
  INV_X1     g00205(.I(new_n379_), .ZN(new_n398_));
  INV_X1     g00206(.I(new_n384_), .ZN(new_n399_));
  AOI21_X1   g00207(.A1(new_n389_), .A2(new_n371_), .B(new_n399_), .ZN(new_n400_));
  AOI21_X1   g00208(.A1(new_n400_), .A2(new_n398_), .B(\asqrt[63] ), .ZN(new_n401_));
  INV_X1     g00209(.I(new_n390_), .ZN(new_n402_));
  NOR4_X1    g00210(.A1(new_n401_), .A2(new_n397_), .A3(new_n402_), .A4(new_n391_), .ZN(new_n403_));
  NOR3_X1    g00211(.A1(new_n403_), .A2(\a[116] ), .A3(\a[117] ), .ZN(new_n404_));
  NOR4_X1    g00212(.A1(new_n401_), .A2(new_n339_), .A3(new_n397_), .A4(new_n402_), .ZN(new_n405_));
  OAI21_X1   g00213(.A1(new_n404_), .A2(new_n405_), .B(new_n292_), .ZN(new_n406_));
  NAND3_X1   g00214(.A1(\asqrt[58] ), .A2(new_n342_), .A3(new_n343_), .ZN(new_n407_));
  INV_X1     g00215(.I(new_n405_), .ZN(new_n408_));
  NAND3_X1   g00216(.A1(new_n407_), .A2(new_n408_), .A3(\a[118] ), .ZN(new_n409_));
  NAND2_X1   g00217(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1     g00218(.I(\a[114] ), .ZN(new_n411_));
  INV_X1     g00219(.I(\a[115] ), .ZN(new_n412_));
  NAND3_X1   g00220(.A1(new_n411_), .A2(new_n412_), .A3(new_n342_), .ZN(new_n413_));
  NAND2_X1   g00221(.A1(\asqrt[58] ), .A2(\a[116] ), .ZN(new_n414_));
  AOI21_X1   g00222(.A1(new_n414_), .A2(new_n413_), .B(new_n339_), .ZN(new_n415_));
  AOI21_X1   g00223(.A1(\asqrt[58] ), .A2(new_n342_), .B(new_n343_), .ZN(new_n416_));
  NOR2_X1    g00224(.A1(new_n404_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1   g00225(.A1(new_n414_), .A2(new_n339_), .A3(new_n413_), .ZN(new_n418_));
  AOI21_X1   g00226(.A1(new_n417_), .A2(new_n418_), .B(new_n415_), .ZN(new_n419_));
  AOI21_X1   g00227(.A1(new_n419_), .A2(new_n288_), .B(new_n410_), .ZN(new_n420_));
  NOR2_X1    g00228(.A1(new_n419_), .A2(new_n288_), .ZN(new_n421_));
  OAI21_X1   g00229(.A1(new_n420_), .A2(new_n421_), .B(\asqrt[61] ), .ZN(new_n422_));
  NOR3_X1    g00230(.A1(new_n420_), .A2(\asqrt[61] ), .A3(new_n421_), .ZN(new_n423_));
  NAND3_X1   g00231(.A1(\asqrt[58] ), .A2(new_n346_), .A3(new_n356_), .ZN(new_n424_));
  XOR2_X1    g00232(.A1(new_n424_), .A2(new_n366_), .Z(new_n425_));
  INV_X1     g00233(.I(new_n425_), .ZN(new_n426_));
  OAI21_X1   g00234(.A1(new_n423_), .A2(new_n426_), .B(new_n422_), .ZN(new_n427_));
  NAND2_X1   g00235(.A1(new_n427_), .A2(\asqrt[62] ), .ZN(new_n428_));
  NOR3_X1    g00236(.A1(new_n403_), .A2(new_n358_), .A3(new_n369_), .ZN(new_n429_));
  XOR2_X1    g00237(.A1(new_n429_), .A2(new_n364_), .Z(new_n430_));
  OAI21_X1   g00238(.A1(new_n427_), .A2(\asqrt[62] ), .B(new_n430_), .ZN(new_n431_));
  NAND2_X1   g00239(.A1(new_n431_), .A2(new_n428_), .ZN(new_n432_));
  INV_X1     g00240(.I(new_n432_), .ZN(new_n433_));
  NOR2_X1    g00241(.A1(new_n433_), .A2(new_n396_), .ZN(new_n434_));
  INV_X1     g00242(.I(new_n434_), .ZN(new_n435_));
  NAND2_X1   g00243(.A1(new_n389_), .A2(new_n371_), .ZN(new_n436_));
  INV_X1     g00244(.I(new_n436_), .ZN(new_n437_));
  NOR2_X1    g00245(.A1(new_n437_), .A2(new_n398_), .ZN(new_n438_));
  INV_X1     g00246(.I(new_n438_), .ZN(new_n439_));
  NOR2_X1    g00247(.A1(new_n403_), .A2(new_n379_), .ZN(new_n440_));
  NAND2_X1   g00248(.A1(new_n440_), .A2(new_n437_), .ZN(new_n441_));
  AOI21_X1   g00249(.A1(new_n441_), .A2(new_n439_), .B(new_n193_), .ZN(new_n442_));
  AOI21_X1   g00250(.A1(new_n440_), .A2(new_n436_), .B(new_n402_), .ZN(new_n443_));
  INV_X1     g00251(.I(new_n443_), .ZN(new_n444_));
  AOI21_X1   g00252(.A1(new_n431_), .A2(new_n428_), .B(new_n444_), .ZN(new_n445_));
  AOI21_X1   g00253(.A1(new_n445_), .A2(new_n396_), .B(\asqrt[63] ), .ZN(new_n446_));
  NAND3_X1   g00254(.A1(new_n431_), .A2(new_n428_), .A3(new_n395_), .ZN(new_n447_));
  INV_X1     g00255(.I(new_n447_), .ZN(new_n448_));
  NOR2_X1    g00256(.A1(\asqrt[58] ), .A2(new_n398_), .ZN(new_n449_));
  NOR4_X1    g00257(.A1(new_n446_), .A2(new_n442_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NOR2_X1    g00258(.A1(new_n450_), .A2(new_n395_), .ZN(new_n451_));
  NAND2_X1   g00259(.A1(new_n451_), .A2(new_n433_), .ZN(new_n452_));
  AOI21_X1   g00260(.A1(new_n452_), .A2(new_n435_), .B(new_n193_), .ZN(new_n453_));
  INV_X1     g00261(.I(new_n453_), .ZN(new_n454_));
  AOI21_X1   g00262(.A1(new_n407_), .A2(new_n408_), .B(\a[118] ), .ZN(new_n455_));
  NOR3_X1    g00263(.A1(new_n404_), .A2(new_n292_), .A3(new_n405_), .ZN(new_n456_));
  NOR2_X1    g00264(.A1(new_n456_), .A2(new_n455_), .ZN(new_n457_));
  OAI21_X1   g00265(.A1(new_n403_), .A2(new_n342_), .B(new_n413_), .ZN(new_n458_));
  NAND2_X1   g00266(.A1(new_n458_), .A2(\asqrt[59] ), .ZN(new_n459_));
  OAI21_X1   g00267(.A1(new_n403_), .A2(\a[116] ), .B(\a[117] ), .ZN(new_n460_));
  NAND2_X1   g00268(.A1(new_n460_), .A2(new_n407_), .ZN(new_n461_));
  NOR2_X1    g00269(.A1(new_n458_), .A2(\asqrt[59] ), .ZN(new_n462_));
  OAI21_X1   g00270(.A1(new_n461_), .A2(new_n462_), .B(new_n459_), .ZN(new_n463_));
  OAI21_X1   g00271(.A1(new_n463_), .A2(\asqrt[60] ), .B(new_n457_), .ZN(new_n464_));
  NAND2_X1   g00272(.A1(new_n463_), .A2(\asqrt[60] ), .ZN(new_n465_));
  AOI21_X1   g00273(.A1(new_n464_), .A2(new_n465_), .B(new_n242_), .ZN(new_n466_));
  NAND3_X1   g00274(.A1(new_n464_), .A2(new_n465_), .A3(new_n242_), .ZN(new_n467_));
  AOI21_X1   g00275(.A1(new_n467_), .A2(new_n425_), .B(new_n466_), .ZN(new_n468_));
  NAND2_X1   g00276(.A1(new_n468_), .A2(new_n234_), .ZN(new_n469_));
  INV_X1     g00277(.I(new_n442_), .ZN(new_n470_));
  NOR2_X1    g00278(.A1(new_n468_), .A2(new_n234_), .ZN(new_n471_));
  INV_X1     g00279(.I(new_n430_), .ZN(new_n472_));
  AOI21_X1   g00280(.A1(new_n468_), .A2(new_n234_), .B(new_n472_), .ZN(new_n473_));
  OAI21_X1   g00281(.A1(new_n473_), .A2(new_n471_), .B(new_n443_), .ZN(new_n474_));
  OAI21_X1   g00282(.A1(new_n474_), .A2(new_n395_), .B(new_n193_), .ZN(new_n475_));
  INV_X1     g00283(.I(new_n449_), .ZN(new_n476_));
  NAND4_X1   g00284(.A1(new_n475_), .A2(new_n470_), .A3(new_n447_), .A4(new_n476_), .ZN(\asqrt[57] ));
  NAND3_X1   g00285(.A1(\asqrt[57] ), .A2(new_n428_), .A3(new_n469_), .ZN(new_n478_));
  XOR2_X1    g00286(.A1(new_n478_), .A2(new_n430_), .Z(new_n479_));
  NAND3_X1   g00287(.A1(\asqrt[57] ), .A2(new_n411_), .A3(new_n412_), .ZN(new_n480_));
  NOR4_X1    g00288(.A1(new_n446_), .A2(new_n403_), .A3(new_n442_), .A4(new_n448_), .ZN(new_n481_));
  INV_X1     g00289(.I(new_n481_), .ZN(new_n482_));
  AOI21_X1   g00290(.A1(new_n480_), .A2(new_n482_), .B(\a[116] ), .ZN(new_n483_));
  NOR3_X1    g00291(.A1(new_n450_), .A2(\a[114] ), .A3(\a[115] ), .ZN(new_n484_));
  NOR3_X1    g00292(.A1(new_n484_), .A2(new_n342_), .A3(new_n481_), .ZN(new_n485_));
  NOR2_X1    g00293(.A1(new_n485_), .A2(new_n483_), .ZN(new_n486_));
  NAND3_X1   g00294(.A1(new_n199_), .A2(new_n200_), .A3(new_n411_), .ZN(new_n487_));
  OAI21_X1   g00295(.A1(new_n450_), .A2(new_n411_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1   g00296(.A1(new_n488_), .A2(\asqrt[58] ), .ZN(new_n489_));
  OAI21_X1   g00297(.A1(new_n450_), .A2(\a[114] ), .B(\a[115] ), .ZN(new_n490_));
  NAND2_X1   g00298(.A1(new_n490_), .A2(new_n480_), .ZN(new_n491_));
  NOR2_X1    g00299(.A1(new_n488_), .A2(\asqrt[58] ), .ZN(new_n492_));
  OAI21_X1   g00300(.A1(new_n491_), .A2(new_n492_), .B(new_n489_), .ZN(new_n493_));
  OAI21_X1   g00301(.A1(new_n493_), .A2(\asqrt[59] ), .B(new_n486_), .ZN(new_n494_));
  NAND2_X1   g00302(.A1(new_n493_), .A2(\asqrt[59] ), .ZN(new_n495_));
  NAND3_X1   g00303(.A1(new_n494_), .A2(new_n288_), .A3(new_n495_), .ZN(new_n496_));
  NAND3_X1   g00304(.A1(\asqrt[57] ), .A2(new_n459_), .A3(new_n418_), .ZN(new_n497_));
  XOR2_X1    g00305(.A1(new_n497_), .A2(new_n461_), .Z(new_n498_));
  NAND2_X1   g00306(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1   g00307(.A1(new_n484_), .A2(new_n481_), .B(new_n342_), .ZN(new_n500_));
  NAND3_X1   g00308(.A1(new_n480_), .A2(\a[116] ), .A3(new_n482_), .ZN(new_n501_));
  NAND2_X1   g00309(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1   g00310(.A1(\asqrt[57] ), .A2(\a[114] ), .ZN(new_n503_));
  AOI21_X1   g00311(.A1(new_n503_), .A2(new_n487_), .B(new_n403_), .ZN(new_n504_));
  AOI21_X1   g00312(.A1(\asqrt[57] ), .A2(new_n411_), .B(new_n412_), .ZN(new_n505_));
  NOR2_X1    g00313(.A1(new_n484_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1   g00314(.A1(new_n503_), .A2(new_n403_), .A3(new_n487_), .ZN(new_n507_));
  AOI21_X1   g00315(.A1(new_n506_), .A2(new_n507_), .B(new_n504_), .ZN(new_n508_));
  AOI21_X1   g00316(.A1(new_n508_), .A2(new_n339_), .B(new_n502_), .ZN(new_n509_));
  NOR2_X1    g00317(.A1(new_n508_), .A2(new_n339_), .ZN(new_n510_));
  OAI21_X1   g00318(.A1(new_n509_), .A2(new_n510_), .B(\asqrt[60] ), .ZN(new_n511_));
  AOI21_X1   g00319(.A1(new_n499_), .A2(new_n511_), .B(new_n242_), .ZN(new_n512_));
  NAND2_X1   g00320(.A1(new_n419_), .A2(new_n288_), .ZN(new_n513_));
  NAND3_X1   g00321(.A1(\asqrt[57] ), .A2(new_n513_), .A3(new_n465_), .ZN(new_n514_));
  XOR2_X1    g00322(.A1(new_n514_), .A2(new_n410_), .Z(new_n515_));
  NAND3_X1   g00323(.A1(new_n499_), .A2(new_n242_), .A3(new_n511_), .ZN(new_n516_));
  AOI21_X1   g00324(.A1(new_n515_), .A2(new_n516_), .B(new_n512_), .ZN(new_n517_));
  NOR2_X1    g00325(.A1(new_n517_), .A2(new_n234_), .ZN(new_n518_));
  NOR3_X1    g00326(.A1(new_n450_), .A2(new_n466_), .A3(new_n423_), .ZN(new_n519_));
  XOR2_X1    g00327(.A1(new_n519_), .A2(new_n425_), .Z(new_n520_));
  INV_X1     g00328(.I(new_n520_), .ZN(new_n521_));
  AOI21_X1   g00329(.A1(new_n517_), .A2(new_n234_), .B(new_n521_), .ZN(new_n522_));
  AOI21_X1   g00330(.A1(new_n451_), .A2(new_n432_), .B(new_n448_), .ZN(new_n523_));
  OAI21_X1   g00331(.A1(new_n522_), .A2(new_n518_), .B(new_n523_), .ZN(new_n524_));
  OAI21_X1   g00332(.A1(new_n524_), .A2(new_n479_), .B(new_n193_), .ZN(new_n525_));
  NOR3_X1    g00333(.A1(new_n509_), .A2(\asqrt[60] ), .A3(new_n510_), .ZN(new_n526_));
  INV_X1     g00334(.I(new_n498_), .ZN(new_n527_));
  OAI21_X1   g00335(.A1(new_n526_), .A2(new_n527_), .B(new_n511_), .ZN(new_n528_));
  OAI21_X1   g00336(.A1(new_n528_), .A2(\asqrt[61] ), .B(new_n515_), .ZN(new_n529_));
  INV_X1     g00337(.I(new_n529_), .ZN(new_n530_));
  OAI21_X1   g00338(.A1(new_n530_), .A2(new_n512_), .B(\asqrt[62] ), .ZN(new_n531_));
  NAND2_X1   g00339(.A1(new_n528_), .A2(\asqrt[61] ), .ZN(new_n532_));
  NAND3_X1   g00340(.A1(new_n529_), .A2(new_n532_), .A3(new_n234_), .ZN(new_n533_));
  NAND2_X1   g00341(.A1(new_n533_), .A2(new_n520_), .ZN(new_n534_));
  NAND3_X1   g00342(.A1(new_n534_), .A2(new_n531_), .A3(new_n479_), .ZN(new_n535_));
  NOR2_X1    g00343(.A1(\asqrt[57] ), .A2(new_n396_), .ZN(new_n536_));
  INV_X1     g00344(.I(new_n536_), .ZN(new_n537_));
  NAND4_X1   g00345(.A1(new_n525_), .A2(new_n454_), .A3(new_n535_), .A4(new_n537_), .ZN(\asqrt[56] ));
  NAND3_X1   g00346(.A1(\asqrt[56] ), .A2(new_n199_), .A3(new_n200_), .ZN(new_n539_));
  INV_X1     g00347(.I(new_n479_), .ZN(new_n540_));
  INV_X1     g00348(.I(new_n523_), .ZN(new_n541_));
  AOI21_X1   g00349(.A1(new_n534_), .A2(new_n531_), .B(new_n541_), .ZN(new_n542_));
  AOI21_X1   g00350(.A1(new_n542_), .A2(new_n540_), .B(\asqrt[63] ), .ZN(new_n543_));
  INV_X1     g00351(.I(new_n535_), .ZN(new_n544_));
  NOR4_X1    g00352(.A1(new_n543_), .A2(new_n453_), .A3(new_n544_), .A4(new_n536_), .ZN(new_n545_));
  OAI21_X1   g00353(.A1(new_n545_), .A2(\a[112] ), .B(\a[113] ), .ZN(new_n546_));
  NAND2_X1   g00354(.A1(new_n546_), .A2(new_n539_), .ZN(new_n547_));
  INV_X1     g00355(.I(\a[110] ), .ZN(new_n548_));
  INV_X1     g00356(.I(\a[111] ), .ZN(new_n549_));
  NAND3_X1   g00357(.A1(new_n548_), .A2(new_n549_), .A3(new_n199_), .ZN(new_n550_));
  OAI21_X1   g00358(.A1(new_n545_), .A2(new_n199_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1   g00359(.A1(new_n551_), .A2(\asqrt[57] ), .ZN(new_n552_));
  NAND2_X1   g00360(.A1(\asqrt[56] ), .A2(\a[112] ), .ZN(new_n553_));
  NAND3_X1   g00361(.A1(new_n553_), .A2(new_n450_), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1   g00362(.A1(new_n534_), .A2(new_n531_), .ZN(new_n555_));
  NAND2_X1   g00363(.A1(new_n555_), .A2(new_n479_), .ZN(new_n556_));
  NOR2_X1    g00364(.A1(new_n545_), .A2(new_n479_), .ZN(new_n557_));
  NAND3_X1   g00365(.A1(new_n557_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n558_));
  AOI21_X1   g00366(.A1(new_n558_), .A2(new_n556_), .B(new_n193_), .ZN(new_n559_));
  INV_X1     g00367(.I(new_n559_), .ZN(new_n560_));
  NAND3_X1   g00368(.A1(\asqrt[56] ), .A2(new_n531_), .A3(new_n533_), .ZN(new_n561_));
  XOR2_X1    g00369(.A1(new_n561_), .A2(new_n520_), .Z(new_n562_));
  AOI21_X1   g00370(.A1(new_n557_), .A2(new_n555_), .B(new_n544_), .ZN(new_n563_));
  NOR2_X1    g00371(.A1(new_n493_), .A2(\asqrt[59] ), .ZN(new_n564_));
  NOR3_X1    g00372(.A1(new_n545_), .A2(new_n564_), .A3(new_n510_), .ZN(new_n565_));
  XOR2_X1    g00373(.A1(new_n565_), .A2(new_n486_), .Z(new_n566_));
  NOR3_X1    g00374(.A1(new_n545_), .A2(\a[112] ), .A3(\a[113] ), .ZN(new_n567_));
  NOR4_X1    g00375(.A1(new_n543_), .A2(new_n450_), .A3(new_n453_), .A4(new_n544_), .ZN(new_n568_));
  OAI21_X1   g00376(.A1(new_n567_), .A2(new_n568_), .B(new_n411_), .ZN(new_n569_));
  INV_X1     g00377(.I(new_n568_), .ZN(new_n570_));
  NAND3_X1   g00378(.A1(new_n539_), .A2(\a[114] ), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1   g00379(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1   g00380(.A1(\asqrt[56] ), .A2(new_n199_), .B(new_n200_), .ZN(new_n573_));
  NOR2_X1    g00381(.A1(new_n567_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1   g00382(.A1(new_n553_), .A2(new_n550_), .B(new_n450_), .ZN(new_n575_));
  AOI21_X1   g00383(.A1(new_n574_), .A2(new_n554_), .B(new_n575_), .ZN(new_n576_));
  AOI21_X1   g00384(.A1(new_n576_), .A2(new_n403_), .B(new_n572_), .ZN(new_n577_));
  NOR2_X1    g00385(.A1(new_n576_), .A2(new_n403_), .ZN(new_n578_));
  NOR3_X1    g00386(.A1(new_n577_), .A2(\asqrt[59] ), .A3(new_n578_), .ZN(new_n579_));
  NOR3_X1    g00387(.A1(new_n545_), .A2(new_n504_), .A3(new_n492_), .ZN(new_n580_));
  XOR2_X1    g00388(.A1(new_n580_), .A2(new_n506_), .Z(new_n581_));
  INV_X1     g00389(.I(new_n581_), .ZN(new_n582_));
  OAI21_X1   g00390(.A1(new_n577_), .A2(new_n578_), .B(\asqrt[59] ), .ZN(new_n583_));
  OAI21_X1   g00391(.A1(new_n579_), .A2(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OAI21_X1   g00392(.A1(new_n584_), .A2(\asqrt[60] ), .B(new_n566_), .ZN(new_n585_));
  NAND2_X1   g00393(.A1(new_n584_), .A2(\asqrt[60] ), .ZN(new_n586_));
  AOI21_X1   g00394(.A1(new_n585_), .A2(new_n586_), .B(new_n242_), .ZN(new_n587_));
  AND3_X2    g00395(.A1(\asqrt[56] ), .A2(new_n496_), .A3(new_n511_), .Z(new_n588_));
  XOR2_X1    g00396(.A1(new_n588_), .A2(new_n498_), .Z(new_n589_));
  NAND3_X1   g00397(.A1(new_n585_), .A2(new_n586_), .A3(new_n242_), .ZN(new_n590_));
  AOI21_X1   g00398(.A1(new_n589_), .A2(new_n590_), .B(new_n587_), .ZN(new_n591_));
  NOR2_X1    g00399(.A1(new_n591_), .A2(new_n234_), .ZN(new_n592_));
  AND3_X2    g00400(.A1(\asqrt[56] ), .A2(new_n532_), .A3(new_n516_), .Z(new_n593_));
  XOR2_X1    g00401(.A1(new_n593_), .A2(new_n515_), .Z(new_n594_));
  INV_X1     g00402(.I(new_n594_), .ZN(new_n595_));
  AOI21_X1   g00403(.A1(new_n591_), .A2(new_n234_), .B(new_n595_), .ZN(new_n596_));
  OAI21_X1   g00404(.A1(new_n596_), .A2(new_n592_), .B(new_n563_), .ZN(new_n597_));
  OAI21_X1   g00405(.A1(new_n597_), .A2(new_n562_), .B(new_n193_), .ZN(new_n598_));
  INV_X1     g00406(.I(new_n562_), .ZN(new_n599_));
  NOR3_X1    g00407(.A1(new_n596_), .A2(new_n592_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1     g00408(.I(new_n600_), .ZN(new_n601_));
  NOR2_X1    g00409(.A1(\asqrt[56] ), .A2(new_n540_), .ZN(new_n602_));
  INV_X1     g00410(.I(new_n602_), .ZN(new_n603_));
  NAND4_X1   g00411(.A1(new_n598_), .A2(new_n560_), .A3(new_n601_), .A4(new_n603_), .ZN(\asqrt[55] ));
  NAND3_X1   g00412(.A1(\asqrt[55] ), .A2(new_n552_), .A3(new_n554_), .ZN(new_n605_));
  XOR2_X1    g00413(.A1(new_n605_), .A2(new_n547_), .Z(new_n606_));
  INV_X1     g00414(.I(new_n563_), .ZN(new_n607_));
  INV_X1     g00415(.I(new_n566_), .ZN(new_n608_));
  AOI21_X1   g00416(.A1(new_n539_), .A2(new_n570_), .B(\a[114] ), .ZN(new_n609_));
  NOR3_X1    g00417(.A1(new_n567_), .A2(new_n411_), .A3(new_n568_), .ZN(new_n610_));
  NOR2_X1    g00418(.A1(new_n610_), .A2(new_n609_), .ZN(new_n611_));
  NOR2_X1    g00419(.A1(new_n551_), .A2(\asqrt[57] ), .ZN(new_n612_));
  OAI21_X1   g00420(.A1(new_n547_), .A2(new_n612_), .B(new_n552_), .ZN(new_n613_));
  OAI21_X1   g00421(.A1(new_n613_), .A2(\asqrt[58] ), .B(new_n611_), .ZN(new_n614_));
  NAND2_X1   g00422(.A1(new_n613_), .A2(\asqrt[58] ), .ZN(new_n615_));
  NAND3_X1   g00423(.A1(new_n614_), .A2(new_n339_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1   g00424(.A1(new_n614_), .A2(new_n615_), .B(new_n339_), .ZN(new_n617_));
  AOI21_X1   g00425(.A1(new_n616_), .A2(new_n581_), .B(new_n617_), .ZN(new_n618_));
  AOI21_X1   g00426(.A1(new_n618_), .A2(new_n288_), .B(new_n608_), .ZN(new_n619_));
  NAND2_X1   g00427(.A1(new_n616_), .A2(new_n581_), .ZN(new_n620_));
  AOI21_X1   g00428(.A1(new_n620_), .A2(new_n583_), .B(new_n288_), .ZN(new_n621_));
  OAI21_X1   g00429(.A1(new_n619_), .A2(new_n621_), .B(\asqrt[61] ), .ZN(new_n622_));
  INV_X1     g00430(.I(new_n589_), .ZN(new_n623_));
  NOR3_X1    g00431(.A1(new_n619_), .A2(\asqrt[61] ), .A3(new_n621_), .ZN(new_n624_));
  OAI21_X1   g00432(.A1(new_n623_), .A2(new_n624_), .B(new_n622_), .ZN(new_n625_));
  NAND2_X1   g00433(.A1(new_n625_), .A2(\asqrt[62] ), .ZN(new_n626_));
  OAI21_X1   g00434(.A1(new_n625_), .A2(\asqrt[62] ), .B(new_n594_), .ZN(new_n627_));
  AOI21_X1   g00435(.A1(new_n627_), .A2(new_n626_), .B(new_n607_), .ZN(new_n628_));
  AOI21_X1   g00436(.A1(new_n628_), .A2(new_n599_), .B(\asqrt[63] ), .ZN(new_n629_));
  NOR4_X1    g00437(.A1(new_n629_), .A2(new_n559_), .A3(new_n600_), .A4(new_n602_), .ZN(new_n630_));
  NOR3_X1    g00438(.A1(new_n630_), .A2(\a[110] ), .A3(\a[111] ), .ZN(new_n631_));
  NAND4_X1   g00439(.A1(new_n598_), .A2(\asqrt[56] ), .A3(new_n601_), .A4(new_n560_), .ZN(new_n632_));
  INV_X1     g00440(.I(new_n632_), .ZN(new_n633_));
  OAI21_X1   g00441(.A1(new_n631_), .A2(new_n633_), .B(new_n199_), .ZN(new_n634_));
  NAND3_X1   g00442(.A1(\asqrt[55] ), .A2(new_n548_), .A3(new_n549_), .ZN(new_n635_));
  NAND3_X1   g00443(.A1(new_n635_), .A2(\a[112] ), .A3(new_n632_), .ZN(new_n636_));
  NAND2_X1   g00444(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1     g00445(.I(\a[108] ), .ZN(new_n638_));
  INV_X1     g00446(.I(\a[109] ), .ZN(new_n639_));
  NAND3_X1   g00447(.A1(new_n638_), .A2(new_n639_), .A3(new_n548_), .ZN(new_n640_));
  NAND2_X1   g00448(.A1(\asqrt[55] ), .A2(\a[110] ), .ZN(new_n641_));
  AOI21_X1   g00449(.A1(new_n641_), .A2(new_n640_), .B(new_n545_), .ZN(new_n642_));
  AOI21_X1   g00450(.A1(\asqrt[55] ), .A2(new_n548_), .B(new_n549_), .ZN(new_n643_));
  NOR2_X1    g00451(.A1(new_n631_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1   g00452(.A1(new_n641_), .A2(new_n545_), .A3(new_n640_), .ZN(new_n645_));
  AOI21_X1   g00453(.A1(new_n644_), .A2(new_n645_), .B(new_n642_), .ZN(new_n646_));
  AOI21_X1   g00454(.A1(new_n646_), .A2(new_n450_), .B(new_n637_), .ZN(new_n647_));
  NOR2_X1    g00455(.A1(new_n646_), .A2(new_n450_), .ZN(new_n648_));
  NOR3_X1    g00456(.A1(new_n647_), .A2(\asqrt[58] ), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1   g00457(.A1(new_n647_), .A2(new_n648_), .B(\asqrt[58] ), .ZN(new_n650_));
  INV_X1     g00458(.I(new_n650_), .ZN(new_n651_));
  NOR2_X1    g00459(.A1(new_n596_), .A2(new_n592_), .ZN(new_n652_));
  INV_X1     g00460(.I(new_n652_), .ZN(new_n653_));
  NAND2_X1   g00461(.A1(new_n653_), .A2(new_n562_), .ZN(new_n654_));
  NOR2_X1    g00462(.A1(new_n630_), .A2(new_n562_), .ZN(new_n655_));
  NAND2_X1   g00463(.A1(new_n655_), .A2(new_n652_), .ZN(new_n656_));
  AOI21_X1   g00464(.A1(new_n656_), .A2(new_n654_), .B(new_n193_), .ZN(new_n657_));
  NOR2_X1    g00465(.A1(new_n625_), .A2(\asqrt[62] ), .ZN(new_n658_));
  OR3_X2     g00466(.A1(new_n630_), .A2(new_n592_), .A3(new_n658_), .Z(new_n659_));
  XOR2_X1    g00467(.A1(new_n659_), .A2(new_n594_), .Z(new_n660_));
  INV_X1     g00468(.I(new_n660_), .ZN(new_n661_));
  AOI21_X1   g00469(.A1(new_n655_), .A2(new_n653_), .B(new_n600_), .ZN(new_n662_));
  INV_X1     g00470(.I(new_n662_), .ZN(new_n663_));
  NOR3_X1    g00471(.A1(new_n630_), .A2(new_n579_), .A3(new_n617_), .ZN(new_n664_));
  XOR2_X1    g00472(.A1(new_n664_), .A2(new_n581_), .Z(new_n665_));
  NAND2_X1   g00473(.A1(new_n576_), .A2(new_n403_), .ZN(new_n666_));
  NAND3_X1   g00474(.A1(\asqrt[55] ), .A2(new_n666_), .A3(new_n615_), .ZN(new_n667_));
  XOR2_X1    g00475(.A1(new_n667_), .A2(new_n572_), .Z(new_n668_));
  INV_X1     g00476(.I(new_n606_), .ZN(new_n669_));
  OAI21_X1   g00477(.A1(new_n669_), .A2(new_n649_), .B(new_n650_), .ZN(new_n670_));
  OAI21_X1   g00478(.A1(new_n670_), .A2(\asqrt[59] ), .B(new_n668_), .ZN(new_n671_));
  NOR2_X1    g00479(.A1(new_n649_), .A2(new_n669_), .ZN(new_n672_));
  OAI21_X1   g00480(.A1(new_n672_), .A2(new_n651_), .B(\asqrt[59] ), .ZN(new_n673_));
  NAND3_X1   g00481(.A1(new_n671_), .A2(new_n288_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1   g00482(.A1(new_n674_), .A2(new_n665_), .ZN(new_n675_));
  INV_X1     g00483(.I(new_n668_), .ZN(new_n676_));
  NOR2_X1    g00484(.A1(new_n672_), .A2(new_n651_), .ZN(new_n677_));
  AOI21_X1   g00485(.A1(new_n677_), .A2(new_n339_), .B(new_n676_), .ZN(new_n678_));
  AOI21_X1   g00486(.A1(new_n635_), .A2(new_n632_), .B(\a[112] ), .ZN(new_n679_));
  NOR3_X1    g00487(.A1(new_n631_), .A2(new_n199_), .A3(new_n633_), .ZN(new_n680_));
  NOR2_X1    g00488(.A1(new_n680_), .A2(new_n679_), .ZN(new_n681_));
  OAI21_X1   g00489(.A1(new_n630_), .A2(new_n548_), .B(new_n640_), .ZN(new_n682_));
  NAND2_X1   g00490(.A1(new_n682_), .A2(\asqrt[56] ), .ZN(new_n683_));
  OAI21_X1   g00491(.A1(new_n630_), .A2(\a[110] ), .B(\a[111] ), .ZN(new_n684_));
  NAND2_X1   g00492(.A1(new_n684_), .A2(new_n635_), .ZN(new_n685_));
  NOR2_X1    g00493(.A1(new_n682_), .A2(\asqrt[56] ), .ZN(new_n686_));
  OAI21_X1   g00494(.A1(new_n685_), .A2(new_n686_), .B(new_n683_), .ZN(new_n687_));
  OAI21_X1   g00495(.A1(new_n687_), .A2(\asqrt[57] ), .B(new_n681_), .ZN(new_n688_));
  NAND2_X1   g00496(.A1(new_n687_), .A2(\asqrt[57] ), .ZN(new_n689_));
  NAND3_X1   g00497(.A1(new_n688_), .A2(new_n689_), .A3(new_n403_), .ZN(new_n690_));
  NAND2_X1   g00498(.A1(new_n690_), .A2(new_n606_), .ZN(new_n691_));
  AOI21_X1   g00499(.A1(new_n691_), .A2(new_n650_), .B(new_n339_), .ZN(new_n692_));
  OAI21_X1   g00500(.A1(new_n678_), .A2(new_n692_), .B(\asqrt[60] ), .ZN(new_n693_));
  AOI21_X1   g00501(.A1(new_n675_), .A2(new_n693_), .B(new_n242_), .ZN(new_n694_));
  NOR2_X1    g00502(.A1(new_n584_), .A2(\asqrt[60] ), .ZN(new_n695_));
  NOR3_X1    g00503(.A1(new_n630_), .A2(new_n695_), .A3(new_n621_), .ZN(new_n696_));
  XOR2_X1    g00504(.A1(new_n696_), .A2(new_n566_), .Z(new_n697_));
  INV_X1     g00505(.I(new_n697_), .ZN(new_n698_));
  NAND2_X1   g00506(.A1(new_n671_), .A2(new_n673_), .ZN(new_n699_));
  AOI21_X1   g00507(.A1(new_n699_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n700_));
  AOI21_X1   g00508(.A1(new_n700_), .A2(new_n675_), .B(new_n698_), .ZN(new_n701_));
  OAI21_X1   g00509(.A1(new_n701_), .A2(new_n694_), .B(\asqrt[62] ), .ZN(new_n702_));
  NOR3_X1    g00510(.A1(new_n630_), .A2(new_n587_), .A3(new_n624_), .ZN(new_n703_));
  XOR2_X1    g00511(.A1(new_n703_), .A2(new_n589_), .Z(new_n704_));
  INV_X1     g00512(.I(new_n665_), .ZN(new_n705_));
  NAND3_X1   g00513(.A1(new_n691_), .A2(new_n339_), .A3(new_n650_), .ZN(new_n706_));
  AOI21_X1   g00514(.A1(new_n668_), .A2(new_n706_), .B(new_n692_), .ZN(new_n707_));
  AOI21_X1   g00515(.A1(new_n707_), .A2(new_n288_), .B(new_n705_), .ZN(new_n708_));
  NOR2_X1    g00516(.A1(new_n707_), .A2(new_n288_), .ZN(new_n709_));
  OAI21_X1   g00517(.A1(new_n708_), .A2(new_n709_), .B(\asqrt[61] ), .ZN(new_n710_));
  OAI21_X1   g00518(.A1(new_n707_), .A2(new_n288_), .B(new_n242_), .ZN(new_n711_));
  OAI21_X1   g00519(.A1(new_n708_), .A2(new_n711_), .B(new_n697_), .ZN(new_n712_));
  NAND3_X1   g00520(.A1(new_n712_), .A2(new_n710_), .A3(new_n234_), .ZN(new_n713_));
  NAND2_X1   g00521(.A1(new_n713_), .A2(new_n704_), .ZN(new_n714_));
  AOI21_X1   g00522(.A1(new_n714_), .A2(new_n702_), .B(new_n663_), .ZN(new_n715_));
  AOI21_X1   g00523(.A1(new_n715_), .A2(new_n661_), .B(\asqrt[63] ), .ZN(new_n716_));
  NAND2_X1   g00524(.A1(new_n714_), .A2(new_n702_), .ZN(new_n717_));
  NOR2_X1    g00525(.A1(new_n717_), .A2(new_n661_), .ZN(new_n718_));
  NOR2_X1    g00526(.A1(\asqrt[55] ), .A2(new_n599_), .ZN(new_n719_));
  NOR4_X1    g00527(.A1(new_n716_), .A2(new_n657_), .A3(new_n718_), .A4(new_n719_), .ZN(new_n720_));
  NOR3_X1    g00528(.A1(new_n720_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n721_));
  XOR2_X1    g00529(.A1(new_n721_), .A2(new_n606_), .Z(new_n722_));
  INV_X1     g00530(.I(new_n722_), .ZN(new_n723_));
  NAND2_X1   g00531(.A1(new_n717_), .A2(new_n660_), .ZN(new_n724_));
  INV_X1     g00532(.I(new_n702_), .ZN(new_n725_));
  NOR2_X1    g00533(.A1(new_n701_), .A2(new_n694_), .ZN(new_n726_));
  INV_X1     g00534(.I(new_n704_), .ZN(new_n727_));
  AOI21_X1   g00535(.A1(new_n726_), .A2(new_n234_), .B(new_n727_), .ZN(new_n728_));
  NOR2_X1    g00536(.A1(new_n728_), .A2(new_n725_), .ZN(new_n729_));
  NOR2_X1    g00537(.A1(new_n720_), .A2(new_n660_), .ZN(new_n730_));
  NAND2_X1   g00538(.A1(new_n730_), .A2(new_n729_), .ZN(new_n731_));
  AOI21_X1   g00539(.A1(new_n731_), .A2(new_n724_), .B(new_n193_), .ZN(new_n732_));
  INV_X1     g00540(.I(new_n732_), .ZN(new_n733_));
  INV_X1     g00541(.I(new_n657_), .ZN(new_n734_));
  OAI21_X1   g00542(.A1(new_n728_), .A2(new_n725_), .B(new_n662_), .ZN(new_n735_));
  OAI21_X1   g00543(.A1(new_n735_), .A2(new_n660_), .B(new_n193_), .ZN(new_n736_));
  NAND2_X1   g00544(.A1(new_n729_), .A2(new_n660_), .ZN(new_n737_));
  INV_X1     g00545(.I(new_n719_), .ZN(new_n738_));
  NAND4_X1   g00546(.A1(new_n736_), .A2(new_n734_), .A3(new_n737_), .A4(new_n738_), .ZN(\asqrt[54] ));
  NAND3_X1   g00547(.A1(\asqrt[54] ), .A2(new_n702_), .A3(new_n713_), .ZN(new_n740_));
  XOR2_X1    g00548(.A1(new_n740_), .A2(new_n704_), .Z(new_n741_));
  AOI21_X1   g00549(.A1(new_n730_), .A2(new_n717_), .B(new_n718_), .ZN(new_n742_));
  AND3_X2    g00550(.A1(\asqrt[54] ), .A2(new_n706_), .A3(new_n673_), .Z(new_n743_));
  XOR2_X1    g00551(.A1(new_n743_), .A2(new_n668_), .Z(new_n744_));
  NOR2_X1    g00552(.A1(new_n687_), .A2(\asqrt[57] ), .ZN(new_n745_));
  NOR3_X1    g00553(.A1(new_n720_), .A2(new_n745_), .A3(new_n648_), .ZN(new_n746_));
  XOR2_X1    g00554(.A1(new_n746_), .A2(new_n681_), .Z(new_n747_));
  INV_X1     g00555(.I(new_n747_), .ZN(new_n748_));
  NAND3_X1   g00556(.A1(\asqrt[54] ), .A2(new_n638_), .A3(new_n639_), .ZN(new_n749_));
  NOR4_X1    g00557(.A1(new_n716_), .A2(new_n630_), .A3(new_n657_), .A4(new_n718_), .ZN(new_n750_));
  INV_X1     g00558(.I(new_n750_), .ZN(new_n751_));
  AOI21_X1   g00559(.A1(new_n749_), .A2(new_n751_), .B(\a[110] ), .ZN(new_n752_));
  NOR3_X1    g00560(.A1(new_n720_), .A2(\a[108] ), .A3(\a[109] ), .ZN(new_n753_));
  NOR3_X1    g00561(.A1(new_n753_), .A2(new_n548_), .A3(new_n750_), .ZN(new_n754_));
  NOR2_X1    g00562(.A1(new_n754_), .A2(new_n752_), .ZN(new_n755_));
  INV_X1     g00563(.I(\a[106] ), .ZN(new_n756_));
  INV_X1     g00564(.I(\a[107] ), .ZN(new_n757_));
  NAND3_X1   g00565(.A1(new_n756_), .A2(new_n757_), .A3(new_n638_), .ZN(new_n758_));
  OAI21_X1   g00566(.A1(new_n720_), .A2(new_n638_), .B(new_n758_), .ZN(new_n759_));
  NAND2_X1   g00567(.A1(new_n759_), .A2(\asqrt[55] ), .ZN(new_n760_));
  OAI21_X1   g00568(.A1(new_n720_), .A2(\a[108] ), .B(\a[109] ), .ZN(new_n761_));
  NAND2_X1   g00569(.A1(new_n761_), .A2(new_n749_), .ZN(new_n762_));
  NOR2_X1    g00570(.A1(new_n759_), .A2(\asqrt[55] ), .ZN(new_n763_));
  OAI21_X1   g00571(.A1(new_n762_), .A2(new_n763_), .B(new_n760_), .ZN(new_n764_));
  OAI21_X1   g00572(.A1(new_n764_), .A2(\asqrt[56] ), .B(new_n755_), .ZN(new_n765_));
  NAND2_X1   g00573(.A1(new_n764_), .A2(\asqrt[56] ), .ZN(new_n766_));
  NAND3_X1   g00574(.A1(new_n765_), .A2(new_n450_), .A3(new_n766_), .ZN(new_n767_));
  NOR3_X1    g00575(.A1(new_n720_), .A2(new_n642_), .A3(new_n686_), .ZN(new_n768_));
  XOR2_X1    g00576(.A1(new_n768_), .A2(new_n644_), .Z(new_n769_));
  AOI21_X1   g00577(.A1(new_n765_), .A2(new_n766_), .B(new_n450_), .ZN(new_n770_));
  AOI21_X1   g00578(.A1(new_n767_), .A2(new_n769_), .B(new_n770_), .ZN(new_n771_));
  AOI21_X1   g00579(.A1(new_n771_), .A2(new_n403_), .B(new_n748_), .ZN(new_n772_));
  OAI21_X1   g00580(.A1(new_n771_), .A2(new_n403_), .B(new_n339_), .ZN(new_n773_));
  OAI21_X1   g00581(.A1(new_n772_), .A2(new_n773_), .B(new_n722_), .ZN(new_n774_));
  NOR2_X1    g00582(.A1(new_n771_), .A2(new_n403_), .ZN(new_n775_));
  OAI21_X1   g00583(.A1(new_n772_), .A2(new_n775_), .B(\asqrt[59] ), .ZN(new_n776_));
  NAND3_X1   g00584(.A1(new_n774_), .A2(new_n776_), .A3(new_n288_), .ZN(new_n777_));
  NAND2_X1   g00585(.A1(new_n777_), .A2(new_n744_), .ZN(new_n778_));
  OAI21_X1   g00586(.A1(new_n753_), .A2(new_n750_), .B(new_n548_), .ZN(new_n779_));
  NAND3_X1   g00587(.A1(new_n749_), .A2(new_n751_), .A3(\a[110] ), .ZN(new_n780_));
  NAND2_X1   g00588(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1   g00589(.A1(\asqrt[54] ), .A2(\a[108] ), .ZN(new_n782_));
  AOI21_X1   g00590(.A1(new_n782_), .A2(new_n758_), .B(new_n630_), .ZN(new_n783_));
  AOI21_X1   g00591(.A1(\asqrt[54] ), .A2(new_n638_), .B(new_n639_), .ZN(new_n784_));
  NOR2_X1    g00592(.A1(new_n753_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1   g00593(.A1(new_n782_), .A2(new_n630_), .A3(new_n758_), .ZN(new_n786_));
  AOI21_X1   g00594(.A1(new_n785_), .A2(new_n786_), .B(new_n783_), .ZN(new_n787_));
  AOI21_X1   g00595(.A1(new_n787_), .A2(new_n545_), .B(new_n781_), .ZN(new_n788_));
  NOR2_X1    g00596(.A1(new_n787_), .A2(new_n545_), .ZN(new_n789_));
  NOR3_X1    g00597(.A1(new_n788_), .A2(\asqrt[57] ), .A3(new_n789_), .ZN(new_n790_));
  INV_X1     g00598(.I(new_n769_), .ZN(new_n791_));
  OAI21_X1   g00599(.A1(new_n788_), .A2(new_n789_), .B(\asqrt[57] ), .ZN(new_n792_));
  OAI21_X1   g00600(.A1(new_n790_), .A2(new_n791_), .B(new_n792_), .ZN(new_n793_));
  OAI21_X1   g00601(.A1(new_n793_), .A2(\asqrt[58] ), .B(new_n747_), .ZN(new_n794_));
  AOI21_X1   g00602(.A1(new_n793_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n795_));
  AOI21_X1   g00603(.A1(new_n795_), .A2(new_n794_), .B(new_n723_), .ZN(new_n796_));
  NAND2_X1   g00604(.A1(new_n793_), .A2(\asqrt[58] ), .ZN(new_n797_));
  AOI21_X1   g00605(.A1(new_n794_), .A2(new_n797_), .B(new_n339_), .ZN(new_n798_));
  OAI21_X1   g00606(.A1(new_n796_), .A2(new_n798_), .B(\asqrt[60] ), .ZN(new_n799_));
  AOI21_X1   g00607(.A1(new_n778_), .A2(new_n799_), .B(new_n242_), .ZN(new_n800_));
  NAND3_X1   g00608(.A1(\asqrt[54] ), .A2(new_n674_), .A3(new_n693_), .ZN(new_n801_));
  XOR2_X1    g00609(.A1(new_n801_), .A2(new_n705_), .Z(new_n802_));
  INV_X1     g00610(.I(new_n802_), .ZN(new_n803_));
  NAND2_X1   g00611(.A1(new_n774_), .A2(new_n776_), .ZN(new_n804_));
  AOI21_X1   g00612(.A1(new_n804_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n805_));
  AOI21_X1   g00613(.A1(new_n805_), .A2(new_n778_), .B(new_n803_), .ZN(new_n806_));
  OAI21_X1   g00614(.A1(new_n806_), .A2(new_n800_), .B(\asqrt[62] ), .ZN(new_n807_));
  INV_X1     g00615(.I(new_n807_), .ZN(new_n808_));
  NOR2_X1    g00616(.A1(new_n806_), .A2(new_n800_), .ZN(new_n809_));
  OAI21_X1   g00617(.A1(new_n708_), .A2(new_n711_), .B(new_n710_), .ZN(new_n810_));
  NOR2_X1    g00618(.A1(new_n720_), .A2(new_n810_), .ZN(new_n811_));
  XOR2_X1    g00619(.A1(new_n811_), .A2(new_n697_), .Z(new_n812_));
  INV_X1     g00620(.I(new_n812_), .ZN(new_n813_));
  AOI21_X1   g00621(.A1(new_n809_), .A2(new_n234_), .B(new_n813_), .ZN(new_n814_));
  OAI21_X1   g00622(.A1(new_n814_), .A2(new_n808_), .B(new_n742_), .ZN(new_n815_));
  OAI21_X1   g00623(.A1(new_n815_), .A2(new_n741_), .B(new_n193_), .ZN(new_n816_));
  NOR2_X1    g00624(.A1(new_n814_), .A2(new_n808_), .ZN(new_n817_));
  NAND2_X1   g00625(.A1(new_n817_), .A2(new_n741_), .ZN(new_n818_));
  NOR2_X1    g00626(.A1(\asqrt[54] ), .A2(new_n661_), .ZN(new_n819_));
  INV_X1     g00627(.I(new_n819_), .ZN(new_n820_));
  NAND4_X1   g00628(.A1(new_n816_), .A2(new_n733_), .A3(new_n818_), .A4(new_n820_), .ZN(\asqrt[53] ));
  AOI21_X1   g00629(.A1(new_n794_), .A2(new_n795_), .B(new_n798_), .ZN(new_n822_));
  NAND2_X1   g00630(.A1(\asqrt[53] ), .A2(new_n822_), .ZN(new_n823_));
  XOR2_X1    g00631(.A1(new_n823_), .A2(new_n723_), .Z(new_n824_));
  INV_X1     g00632(.I(new_n824_), .ZN(new_n825_));
  NOR2_X1    g00633(.A1(new_n793_), .A2(\asqrt[58] ), .ZN(new_n826_));
  INV_X1     g00634(.I(new_n741_), .ZN(new_n827_));
  INV_X1     g00635(.I(new_n742_), .ZN(new_n828_));
  INV_X1     g00636(.I(new_n744_), .ZN(new_n829_));
  NOR2_X1    g00637(.A1(new_n796_), .A2(new_n798_), .ZN(new_n830_));
  AOI21_X1   g00638(.A1(new_n830_), .A2(new_n288_), .B(new_n829_), .ZN(new_n831_));
  INV_X1     g00639(.I(new_n799_), .ZN(new_n832_));
  OAI21_X1   g00640(.A1(new_n831_), .A2(new_n832_), .B(\asqrt[61] ), .ZN(new_n833_));
  NAND2_X1   g00641(.A1(new_n799_), .A2(new_n242_), .ZN(new_n834_));
  OAI21_X1   g00642(.A1(new_n831_), .A2(new_n834_), .B(new_n802_), .ZN(new_n835_));
  NAND3_X1   g00643(.A1(new_n835_), .A2(new_n833_), .A3(new_n234_), .ZN(new_n836_));
  NAND2_X1   g00644(.A1(new_n836_), .A2(new_n812_), .ZN(new_n837_));
  AOI21_X1   g00645(.A1(new_n837_), .A2(new_n807_), .B(new_n828_), .ZN(new_n838_));
  AOI21_X1   g00646(.A1(new_n838_), .A2(new_n827_), .B(\asqrt[63] ), .ZN(new_n839_));
  NAND2_X1   g00647(.A1(new_n837_), .A2(new_n807_), .ZN(new_n840_));
  NOR2_X1    g00648(.A1(new_n840_), .A2(new_n827_), .ZN(new_n841_));
  NOR4_X1    g00649(.A1(new_n839_), .A2(new_n732_), .A3(new_n841_), .A4(new_n819_), .ZN(new_n842_));
  NOR3_X1    g00650(.A1(new_n842_), .A2(new_n826_), .A3(new_n775_), .ZN(new_n843_));
  XOR2_X1    g00651(.A1(new_n843_), .A2(new_n747_), .Z(new_n844_));
  NOR3_X1    g00652(.A1(new_n842_), .A2(new_n790_), .A3(new_n770_), .ZN(new_n845_));
  XOR2_X1    g00653(.A1(new_n845_), .A2(new_n769_), .Z(new_n846_));
  INV_X1     g00654(.I(new_n846_), .ZN(new_n847_));
  NOR2_X1    g00655(.A1(new_n764_), .A2(\asqrt[56] ), .ZN(new_n848_));
  NOR3_X1    g00656(.A1(new_n842_), .A2(new_n848_), .A3(new_n789_), .ZN(new_n849_));
  XOR2_X1    g00657(.A1(new_n849_), .A2(new_n755_), .Z(new_n850_));
  INV_X1     g00658(.I(new_n850_), .ZN(new_n851_));
  NAND3_X1   g00659(.A1(\asqrt[53] ), .A2(new_n756_), .A3(new_n757_), .ZN(new_n852_));
  NOR4_X1    g00660(.A1(new_n839_), .A2(new_n720_), .A3(new_n732_), .A4(new_n841_), .ZN(new_n853_));
  INV_X1     g00661(.I(new_n853_), .ZN(new_n854_));
  AOI21_X1   g00662(.A1(new_n852_), .A2(new_n854_), .B(\a[108] ), .ZN(new_n855_));
  NOR3_X1    g00663(.A1(new_n842_), .A2(\a[106] ), .A3(\a[107] ), .ZN(new_n856_));
  NOR3_X1    g00664(.A1(new_n856_), .A2(new_n638_), .A3(new_n853_), .ZN(new_n857_));
  NOR2_X1    g00665(.A1(new_n857_), .A2(new_n855_), .ZN(new_n858_));
  INV_X1     g00666(.I(\a[104] ), .ZN(new_n859_));
  INV_X1     g00667(.I(\a[105] ), .ZN(new_n860_));
  NAND3_X1   g00668(.A1(new_n859_), .A2(new_n860_), .A3(new_n756_), .ZN(new_n861_));
  OAI21_X1   g00669(.A1(new_n842_), .A2(new_n756_), .B(new_n861_), .ZN(new_n862_));
  NAND2_X1   g00670(.A1(new_n862_), .A2(\asqrt[54] ), .ZN(new_n863_));
  OAI21_X1   g00671(.A1(new_n842_), .A2(\a[106] ), .B(\a[107] ), .ZN(new_n864_));
  NAND2_X1   g00672(.A1(new_n864_), .A2(new_n852_), .ZN(new_n865_));
  NOR2_X1    g00673(.A1(new_n862_), .A2(\asqrt[54] ), .ZN(new_n866_));
  OAI21_X1   g00674(.A1(new_n865_), .A2(new_n866_), .B(new_n863_), .ZN(new_n867_));
  OAI21_X1   g00675(.A1(\asqrt[55] ), .A2(new_n867_), .B(new_n858_), .ZN(new_n868_));
  NAND2_X1   g00676(.A1(new_n867_), .A2(\asqrt[55] ), .ZN(new_n869_));
  NAND3_X1   g00677(.A1(new_n868_), .A2(new_n545_), .A3(new_n869_), .ZN(new_n870_));
  NOR3_X1    g00678(.A1(new_n842_), .A2(new_n783_), .A3(new_n763_), .ZN(new_n871_));
  XOR2_X1    g00679(.A1(new_n871_), .A2(new_n785_), .Z(new_n872_));
  NAND2_X1   g00680(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1   g00681(.A1(new_n868_), .A2(new_n869_), .ZN(new_n874_));
  AOI21_X1   g00682(.A1(new_n874_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n875_));
  AOI21_X1   g00683(.A1(new_n875_), .A2(new_n873_), .B(new_n851_), .ZN(new_n876_));
  OAI21_X1   g00684(.A1(new_n856_), .A2(new_n853_), .B(new_n638_), .ZN(new_n877_));
  NAND3_X1   g00685(.A1(new_n852_), .A2(\a[108] ), .A3(new_n854_), .ZN(new_n878_));
  NAND2_X1   g00686(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1   g00687(.A1(\asqrt[53] ), .A2(\a[106] ), .ZN(new_n880_));
  AOI21_X1   g00688(.A1(new_n880_), .A2(new_n861_), .B(new_n720_), .ZN(new_n881_));
  AOI21_X1   g00689(.A1(\asqrt[53] ), .A2(new_n756_), .B(new_n757_), .ZN(new_n882_));
  NOR2_X1    g00690(.A1(new_n882_), .A2(new_n856_), .ZN(new_n883_));
  NAND3_X1   g00691(.A1(new_n880_), .A2(new_n720_), .A3(new_n861_), .ZN(new_n884_));
  AOI21_X1   g00692(.A1(new_n883_), .A2(new_n884_), .B(new_n881_), .ZN(new_n885_));
  AOI21_X1   g00693(.A1(new_n885_), .A2(new_n630_), .B(new_n879_), .ZN(new_n886_));
  NOR2_X1    g00694(.A1(new_n885_), .A2(new_n630_), .ZN(new_n887_));
  OAI21_X1   g00695(.A1(new_n886_), .A2(new_n887_), .B(\asqrt[56] ), .ZN(new_n888_));
  AOI21_X1   g00696(.A1(new_n873_), .A2(new_n888_), .B(new_n450_), .ZN(new_n889_));
  NOR2_X1    g00697(.A1(new_n876_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1   g00698(.A1(new_n890_), .A2(new_n403_), .B(new_n847_), .ZN(new_n891_));
  OAI21_X1   g00699(.A1(new_n876_), .A2(new_n889_), .B(\asqrt[58] ), .ZN(new_n892_));
  NAND2_X1   g00700(.A1(new_n892_), .A2(new_n339_), .ZN(new_n893_));
  OAI21_X1   g00701(.A1(new_n891_), .A2(new_n893_), .B(new_n844_), .ZN(new_n894_));
  INV_X1     g00702(.I(new_n892_), .ZN(new_n895_));
  OAI21_X1   g00703(.A1(new_n891_), .A2(new_n895_), .B(\asqrt[59] ), .ZN(new_n896_));
  NAND3_X1   g00704(.A1(new_n894_), .A2(new_n896_), .A3(new_n288_), .ZN(new_n897_));
  INV_X1     g00705(.I(new_n844_), .ZN(new_n898_));
  NOR2_X1    g00706(.A1(new_n886_), .A2(new_n887_), .ZN(new_n899_));
  INV_X1     g00707(.I(new_n872_), .ZN(new_n900_));
  AOI21_X1   g00708(.A1(new_n899_), .A2(new_n545_), .B(new_n900_), .ZN(new_n901_));
  NAND2_X1   g00709(.A1(new_n888_), .A2(new_n450_), .ZN(new_n902_));
  OAI21_X1   g00710(.A1(new_n901_), .A2(new_n902_), .B(new_n850_), .ZN(new_n903_));
  INV_X1     g00711(.I(new_n888_), .ZN(new_n904_));
  OAI21_X1   g00712(.A1(new_n901_), .A2(new_n904_), .B(\asqrt[57] ), .ZN(new_n905_));
  NAND3_X1   g00713(.A1(new_n903_), .A2(new_n905_), .A3(new_n403_), .ZN(new_n906_));
  NAND2_X1   g00714(.A1(new_n906_), .A2(new_n846_), .ZN(new_n907_));
  NAND2_X1   g00715(.A1(new_n903_), .A2(new_n905_), .ZN(new_n908_));
  AOI21_X1   g00716(.A1(new_n908_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n909_));
  AOI21_X1   g00717(.A1(new_n909_), .A2(new_n907_), .B(new_n898_), .ZN(new_n910_));
  AOI21_X1   g00718(.A1(new_n907_), .A2(new_n892_), .B(new_n339_), .ZN(new_n911_));
  OAI21_X1   g00719(.A1(new_n910_), .A2(new_n911_), .B(\asqrt[60] ), .ZN(new_n912_));
  NAND2_X1   g00720(.A1(new_n840_), .A2(new_n741_), .ZN(new_n913_));
  NOR2_X1    g00721(.A1(new_n842_), .A2(new_n741_), .ZN(new_n914_));
  NAND2_X1   g00722(.A1(new_n914_), .A2(new_n817_), .ZN(new_n915_));
  AOI21_X1   g00723(.A1(new_n915_), .A2(new_n913_), .B(new_n193_), .ZN(new_n916_));
  INV_X1     g00724(.I(new_n916_), .ZN(new_n917_));
  NAND3_X1   g00725(.A1(\asqrt[53] ), .A2(new_n807_), .A3(new_n836_), .ZN(new_n918_));
  XOR2_X1    g00726(.A1(new_n918_), .A2(new_n812_), .Z(new_n919_));
  AOI21_X1   g00727(.A1(new_n914_), .A2(new_n840_), .B(new_n841_), .ZN(new_n920_));
  NAND2_X1   g00728(.A1(new_n897_), .A2(new_n824_), .ZN(new_n921_));
  AOI21_X1   g00729(.A1(new_n921_), .A2(new_n912_), .B(new_n242_), .ZN(new_n922_));
  NAND3_X1   g00730(.A1(\asqrt[53] ), .A2(new_n777_), .A3(new_n799_), .ZN(new_n923_));
  XOR2_X1    g00731(.A1(new_n923_), .A2(new_n829_), .Z(new_n924_));
  INV_X1     g00732(.I(new_n924_), .ZN(new_n925_));
  NAND2_X1   g00733(.A1(new_n894_), .A2(new_n896_), .ZN(new_n926_));
  AOI21_X1   g00734(.A1(new_n926_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n927_));
  AOI21_X1   g00735(.A1(new_n927_), .A2(new_n921_), .B(new_n925_), .ZN(new_n928_));
  OAI21_X1   g00736(.A1(new_n928_), .A2(new_n922_), .B(\asqrt[62] ), .ZN(new_n929_));
  INV_X1     g00737(.I(new_n929_), .ZN(new_n930_));
  NOR2_X1    g00738(.A1(new_n928_), .A2(new_n922_), .ZN(new_n931_));
  AOI21_X1   g00739(.A1(new_n778_), .A2(new_n805_), .B(new_n800_), .ZN(new_n932_));
  NAND2_X1   g00740(.A1(\asqrt[53] ), .A2(new_n932_), .ZN(new_n933_));
  XOR2_X1    g00741(.A1(new_n933_), .A2(new_n803_), .Z(new_n934_));
  INV_X1     g00742(.I(new_n934_), .ZN(new_n935_));
  AOI21_X1   g00743(.A1(new_n931_), .A2(new_n234_), .B(new_n935_), .ZN(new_n936_));
  OAI21_X1   g00744(.A1(new_n936_), .A2(new_n930_), .B(new_n920_), .ZN(new_n937_));
  OAI21_X1   g00745(.A1(new_n937_), .A2(new_n919_), .B(new_n193_), .ZN(new_n938_));
  NOR2_X1    g00746(.A1(new_n936_), .A2(new_n930_), .ZN(new_n939_));
  NAND2_X1   g00747(.A1(new_n939_), .A2(new_n919_), .ZN(new_n940_));
  NOR2_X1    g00748(.A1(\asqrt[53] ), .A2(new_n827_), .ZN(new_n941_));
  INV_X1     g00749(.I(new_n941_), .ZN(new_n942_));
  NAND4_X1   g00750(.A1(new_n938_), .A2(new_n917_), .A3(new_n940_), .A4(new_n942_), .ZN(\asqrt[52] ));
  NAND3_X1   g00751(.A1(\asqrt[52] ), .A2(new_n897_), .A3(new_n912_), .ZN(new_n944_));
  XOR2_X1    g00752(.A1(new_n944_), .A2(new_n825_), .Z(new_n945_));
  INV_X1     g00753(.I(new_n945_), .ZN(new_n946_));
  NOR2_X1    g00754(.A1(new_n910_), .A2(new_n911_), .ZN(new_n947_));
  AOI21_X1   g00755(.A1(new_n947_), .A2(new_n288_), .B(new_n825_), .ZN(new_n948_));
  INV_X1     g00756(.I(new_n912_), .ZN(new_n949_));
  OAI21_X1   g00757(.A1(new_n948_), .A2(new_n949_), .B(\asqrt[61] ), .ZN(new_n950_));
  NAND2_X1   g00758(.A1(new_n912_), .A2(new_n242_), .ZN(new_n951_));
  OAI21_X1   g00759(.A1(new_n948_), .A2(new_n951_), .B(new_n924_), .ZN(new_n952_));
  NAND3_X1   g00760(.A1(new_n952_), .A2(new_n950_), .A3(new_n234_), .ZN(new_n953_));
  NAND2_X1   g00761(.A1(new_n953_), .A2(new_n934_), .ZN(new_n954_));
  NAND2_X1   g00762(.A1(new_n954_), .A2(new_n929_), .ZN(new_n955_));
  NAND2_X1   g00763(.A1(new_n955_), .A2(new_n919_), .ZN(new_n956_));
  INV_X1     g00764(.I(new_n919_), .ZN(new_n957_));
  INV_X1     g00765(.I(new_n920_), .ZN(new_n958_));
  AOI21_X1   g00766(.A1(new_n954_), .A2(new_n929_), .B(new_n958_), .ZN(new_n959_));
  AOI21_X1   g00767(.A1(new_n959_), .A2(new_n957_), .B(\asqrt[63] ), .ZN(new_n960_));
  NOR2_X1    g00768(.A1(new_n955_), .A2(new_n957_), .ZN(new_n961_));
  NOR4_X1    g00769(.A1(new_n960_), .A2(new_n916_), .A3(new_n961_), .A4(new_n941_), .ZN(new_n962_));
  NOR2_X1    g00770(.A1(new_n962_), .A2(new_n919_), .ZN(new_n963_));
  NAND2_X1   g00771(.A1(new_n963_), .A2(new_n939_), .ZN(new_n964_));
  AOI21_X1   g00772(.A1(new_n964_), .A2(new_n956_), .B(new_n193_), .ZN(new_n965_));
  INV_X1     g00773(.I(new_n965_), .ZN(new_n966_));
  NAND3_X1   g00774(.A1(\asqrt[52] ), .A2(new_n929_), .A3(new_n953_), .ZN(new_n967_));
  XOR2_X1    g00775(.A1(new_n967_), .A2(new_n934_), .Z(new_n968_));
  AOI21_X1   g00776(.A1(new_n963_), .A2(new_n955_), .B(new_n961_), .ZN(new_n969_));
  OAI21_X1   g00777(.A1(new_n891_), .A2(new_n893_), .B(new_n896_), .ZN(new_n970_));
  NOR2_X1    g00778(.A1(new_n962_), .A2(new_n970_), .ZN(new_n971_));
  XOR2_X1    g00779(.A1(new_n971_), .A2(new_n844_), .Z(new_n972_));
  NAND3_X1   g00780(.A1(\asqrt[52] ), .A2(new_n906_), .A3(new_n892_), .ZN(new_n973_));
  XOR2_X1    g00781(.A1(new_n973_), .A2(new_n847_), .Z(new_n974_));
  OAI21_X1   g00782(.A1(new_n901_), .A2(new_n902_), .B(new_n905_), .ZN(new_n975_));
  NOR2_X1    g00783(.A1(new_n962_), .A2(new_n975_), .ZN(new_n976_));
  XOR2_X1    g00784(.A1(new_n976_), .A2(new_n850_), .Z(new_n977_));
  INV_X1     g00785(.I(new_n977_), .ZN(new_n978_));
  NAND3_X1   g00786(.A1(\asqrt[52] ), .A2(new_n870_), .A3(new_n888_), .ZN(new_n979_));
  XOR2_X1    g00787(.A1(new_n979_), .A2(new_n900_), .Z(new_n980_));
  INV_X1     g00788(.I(new_n980_), .ZN(new_n981_));
  NAND2_X1   g00789(.A1(new_n885_), .A2(new_n630_), .ZN(new_n982_));
  NAND3_X1   g00790(.A1(\asqrt[52] ), .A2(new_n982_), .A3(new_n869_), .ZN(new_n983_));
  XOR2_X1    g00791(.A1(new_n983_), .A2(new_n879_), .Z(new_n984_));
  NOR3_X1    g00792(.A1(new_n962_), .A2(\a[104] ), .A3(\a[105] ), .ZN(new_n985_));
  NOR4_X1    g00793(.A1(new_n960_), .A2(new_n842_), .A3(new_n916_), .A4(new_n961_), .ZN(new_n986_));
  OAI21_X1   g00794(.A1(new_n985_), .A2(new_n986_), .B(new_n756_), .ZN(new_n987_));
  NAND3_X1   g00795(.A1(\asqrt[52] ), .A2(new_n859_), .A3(new_n860_), .ZN(new_n988_));
  INV_X1     g00796(.I(new_n986_), .ZN(new_n989_));
  NAND3_X1   g00797(.A1(new_n988_), .A2(\a[106] ), .A3(new_n989_), .ZN(new_n990_));
  NAND2_X1   g00798(.A1(new_n987_), .A2(new_n990_), .ZN(new_n991_));
  INV_X1     g00799(.I(\a[102] ), .ZN(new_n992_));
  INV_X1     g00800(.I(\a[103] ), .ZN(new_n993_));
  NAND3_X1   g00801(.A1(new_n992_), .A2(new_n993_), .A3(new_n859_), .ZN(new_n994_));
  NAND2_X1   g00802(.A1(\asqrt[52] ), .A2(\a[104] ), .ZN(new_n995_));
  AOI21_X1   g00803(.A1(new_n995_), .A2(new_n994_), .B(new_n842_), .ZN(new_n996_));
  AOI21_X1   g00804(.A1(\asqrt[52] ), .A2(new_n859_), .B(new_n860_), .ZN(new_n997_));
  NOR2_X1    g00805(.A1(new_n985_), .A2(new_n997_), .ZN(new_n998_));
  NAND3_X1   g00806(.A1(new_n995_), .A2(new_n842_), .A3(new_n994_), .ZN(new_n999_));
  AOI21_X1   g00807(.A1(new_n998_), .A2(new_n999_), .B(new_n996_), .ZN(new_n1000_));
  AOI21_X1   g00808(.A1(new_n1000_), .A2(new_n720_), .B(new_n991_), .ZN(new_n1001_));
  NOR2_X1    g00809(.A1(new_n1000_), .A2(new_n720_), .ZN(new_n1002_));
  NOR3_X1    g00810(.A1(new_n1001_), .A2(\asqrt[55] ), .A3(new_n1002_), .ZN(new_n1003_));
  NOR3_X1    g00811(.A1(new_n962_), .A2(new_n881_), .A3(new_n866_), .ZN(new_n1004_));
  XOR2_X1    g00812(.A1(new_n1004_), .A2(new_n883_), .Z(new_n1005_));
  INV_X1     g00813(.I(new_n1005_), .ZN(new_n1006_));
  OAI21_X1   g00814(.A1(new_n1001_), .A2(new_n1002_), .B(\asqrt[55] ), .ZN(new_n1007_));
  OAI21_X1   g00815(.A1(new_n1003_), .A2(new_n1006_), .B(new_n1007_), .ZN(new_n1008_));
  OAI21_X1   g00816(.A1(new_n1008_), .A2(\asqrt[56] ), .B(new_n984_), .ZN(new_n1009_));
  AOI21_X1   g00817(.A1(new_n1008_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1010_));
  AOI21_X1   g00818(.A1(new_n1010_), .A2(new_n1009_), .B(new_n981_), .ZN(new_n1011_));
  NAND2_X1   g00819(.A1(new_n1008_), .A2(\asqrt[56] ), .ZN(new_n1012_));
  AOI21_X1   g00820(.A1(new_n1009_), .A2(new_n1012_), .B(new_n450_), .ZN(new_n1013_));
  NOR2_X1    g00821(.A1(new_n1011_), .A2(new_n1013_), .ZN(new_n1014_));
  AOI21_X1   g00822(.A1(new_n1014_), .A2(new_n403_), .B(new_n978_), .ZN(new_n1015_));
  OAI21_X1   g00823(.A1(new_n1011_), .A2(new_n1013_), .B(\asqrt[58] ), .ZN(new_n1016_));
  NAND2_X1   g00824(.A1(new_n1016_), .A2(new_n339_), .ZN(new_n1017_));
  OAI21_X1   g00825(.A1(new_n1015_), .A2(new_n1017_), .B(new_n974_), .ZN(new_n1018_));
  INV_X1     g00826(.I(new_n1016_), .ZN(new_n1019_));
  OAI21_X1   g00827(.A1(new_n1015_), .A2(new_n1019_), .B(\asqrt[59] ), .ZN(new_n1020_));
  NAND3_X1   g00828(.A1(new_n1018_), .A2(new_n1020_), .A3(new_n288_), .ZN(new_n1021_));
  NAND2_X1   g00829(.A1(new_n1021_), .A2(new_n972_), .ZN(new_n1022_));
  INV_X1     g00830(.I(new_n974_), .ZN(new_n1023_));
  INV_X1     g00831(.I(new_n984_), .ZN(new_n1024_));
  AOI21_X1   g00832(.A1(new_n988_), .A2(new_n989_), .B(\a[106] ), .ZN(new_n1025_));
  NOR3_X1    g00833(.A1(new_n985_), .A2(new_n756_), .A3(new_n986_), .ZN(new_n1026_));
  NOR2_X1    g00834(.A1(new_n1026_), .A2(new_n1025_), .ZN(new_n1027_));
  OAI21_X1   g00835(.A1(new_n962_), .A2(new_n859_), .B(new_n994_), .ZN(new_n1028_));
  NAND2_X1   g00836(.A1(new_n1028_), .A2(\asqrt[53] ), .ZN(new_n1029_));
  OAI21_X1   g00837(.A1(new_n962_), .A2(\a[104] ), .B(\a[105] ), .ZN(new_n1030_));
  NAND2_X1   g00838(.A1(new_n1030_), .A2(new_n988_), .ZN(new_n1031_));
  NOR2_X1    g00839(.A1(new_n1028_), .A2(\asqrt[53] ), .ZN(new_n1032_));
  OAI21_X1   g00840(.A1(new_n1031_), .A2(new_n1032_), .B(new_n1029_), .ZN(new_n1033_));
  OAI21_X1   g00841(.A1(\asqrt[54] ), .A2(new_n1033_), .B(new_n1027_), .ZN(new_n1034_));
  NAND2_X1   g00842(.A1(new_n1033_), .A2(\asqrt[54] ), .ZN(new_n1035_));
  NAND3_X1   g00843(.A1(new_n1034_), .A2(new_n630_), .A3(new_n1035_), .ZN(new_n1036_));
  AOI21_X1   g00844(.A1(new_n1034_), .A2(new_n1035_), .B(new_n630_), .ZN(new_n1037_));
  AOI21_X1   g00845(.A1(new_n1036_), .A2(new_n1005_), .B(new_n1037_), .ZN(new_n1038_));
  AOI21_X1   g00846(.A1(new_n1038_), .A2(new_n545_), .B(new_n1024_), .ZN(new_n1039_));
  OAI21_X1   g00847(.A1(new_n1038_), .A2(new_n545_), .B(new_n450_), .ZN(new_n1040_));
  OAI21_X1   g00848(.A1(new_n1039_), .A2(new_n1040_), .B(new_n980_), .ZN(new_n1041_));
  NOR2_X1    g00849(.A1(new_n1038_), .A2(new_n545_), .ZN(new_n1042_));
  OAI21_X1   g00850(.A1(new_n1039_), .A2(new_n1042_), .B(\asqrt[57] ), .ZN(new_n1043_));
  NAND3_X1   g00851(.A1(new_n1041_), .A2(new_n1043_), .A3(new_n403_), .ZN(new_n1044_));
  NAND2_X1   g00852(.A1(new_n1044_), .A2(new_n977_), .ZN(new_n1045_));
  NAND2_X1   g00853(.A1(new_n1041_), .A2(new_n1043_), .ZN(new_n1046_));
  AOI21_X1   g00854(.A1(new_n1046_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1047_));
  AOI21_X1   g00855(.A1(new_n1047_), .A2(new_n1045_), .B(new_n1023_), .ZN(new_n1048_));
  AOI21_X1   g00856(.A1(new_n1045_), .A2(new_n1016_), .B(new_n339_), .ZN(new_n1049_));
  OAI21_X1   g00857(.A1(new_n1048_), .A2(new_n1049_), .B(\asqrt[60] ), .ZN(new_n1050_));
  AOI21_X1   g00858(.A1(new_n1022_), .A2(new_n1050_), .B(new_n242_), .ZN(new_n1051_));
  NAND2_X1   g00859(.A1(new_n1018_), .A2(new_n1020_), .ZN(new_n1052_));
  AOI21_X1   g00860(.A1(new_n1052_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1053_));
  AOI21_X1   g00861(.A1(new_n1053_), .A2(new_n1022_), .B(new_n946_), .ZN(new_n1054_));
  OAI21_X1   g00862(.A1(new_n1054_), .A2(new_n1051_), .B(\asqrt[62] ), .ZN(new_n1055_));
  INV_X1     g00863(.I(new_n1055_), .ZN(new_n1056_));
  NOR2_X1    g00864(.A1(new_n1054_), .A2(new_n1051_), .ZN(new_n1057_));
  AOI21_X1   g00865(.A1(new_n921_), .A2(new_n927_), .B(new_n922_), .ZN(new_n1058_));
  NAND2_X1   g00866(.A1(\asqrt[52] ), .A2(new_n1058_), .ZN(new_n1059_));
  XOR2_X1    g00867(.A1(new_n1059_), .A2(new_n925_), .Z(new_n1060_));
  INV_X1     g00868(.I(new_n1060_), .ZN(new_n1061_));
  AOI21_X1   g00869(.A1(new_n1057_), .A2(new_n234_), .B(new_n1061_), .ZN(new_n1062_));
  OAI21_X1   g00870(.A1(new_n1062_), .A2(new_n1056_), .B(new_n969_), .ZN(new_n1063_));
  OAI21_X1   g00871(.A1(new_n1063_), .A2(new_n968_), .B(new_n193_), .ZN(new_n1064_));
  NOR2_X1    g00872(.A1(new_n1062_), .A2(new_n1056_), .ZN(new_n1065_));
  NAND2_X1   g00873(.A1(new_n1065_), .A2(new_n968_), .ZN(new_n1066_));
  NOR2_X1    g00874(.A1(\asqrt[52] ), .A2(new_n957_), .ZN(new_n1067_));
  INV_X1     g00875(.I(new_n1067_), .ZN(new_n1068_));
  NAND4_X1   g00876(.A1(new_n1064_), .A2(new_n966_), .A3(new_n1066_), .A4(new_n1068_), .ZN(\asqrt[51] ));
  AOI21_X1   g00877(.A1(new_n1022_), .A2(new_n1053_), .B(new_n1051_), .ZN(new_n1070_));
  NAND2_X1   g00878(.A1(\asqrt[51] ), .A2(new_n1070_), .ZN(new_n1071_));
  XOR2_X1    g00879(.A1(new_n1071_), .A2(new_n946_), .Z(new_n1072_));
  INV_X1     g00880(.I(new_n968_), .ZN(new_n1073_));
  INV_X1     g00881(.I(new_n969_), .ZN(new_n1074_));
  INV_X1     g00882(.I(new_n972_), .ZN(new_n1075_));
  NOR2_X1    g00883(.A1(new_n1048_), .A2(new_n1049_), .ZN(new_n1076_));
  AOI21_X1   g00884(.A1(new_n1076_), .A2(new_n288_), .B(new_n1075_), .ZN(new_n1077_));
  INV_X1     g00885(.I(new_n1050_), .ZN(new_n1078_));
  OAI21_X1   g00886(.A1(new_n1077_), .A2(new_n1078_), .B(\asqrt[61] ), .ZN(new_n1079_));
  NAND2_X1   g00887(.A1(new_n1050_), .A2(new_n242_), .ZN(new_n1080_));
  OAI21_X1   g00888(.A1(new_n1077_), .A2(new_n1080_), .B(new_n945_), .ZN(new_n1081_));
  NAND3_X1   g00889(.A1(new_n1081_), .A2(new_n1079_), .A3(new_n234_), .ZN(new_n1082_));
  NAND2_X1   g00890(.A1(new_n1082_), .A2(new_n1060_), .ZN(new_n1083_));
  AOI21_X1   g00891(.A1(new_n1083_), .A2(new_n1055_), .B(new_n1074_), .ZN(new_n1084_));
  AOI21_X1   g00892(.A1(new_n1084_), .A2(new_n1073_), .B(\asqrt[63] ), .ZN(new_n1085_));
  NAND2_X1   g00893(.A1(new_n1083_), .A2(new_n1055_), .ZN(new_n1086_));
  NOR2_X1    g00894(.A1(new_n1086_), .A2(new_n1073_), .ZN(new_n1087_));
  NOR4_X1    g00895(.A1(new_n1085_), .A2(new_n965_), .A3(new_n1087_), .A4(new_n1067_), .ZN(new_n1088_));
  OAI21_X1   g00896(.A1(new_n1015_), .A2(new_n1017_), .B(new_n1020_), .ZN(new_n1089_));
  NOR2_X1    g00897(.A1(new_n1088_), .A2(new_n1089_), .ZN(new_n1090_));
  XOR2_X1    g00898(.A1(new_n1090_), .A2(new_n974_), .Z(new_n1091_));
  NAND3_X1   g00899(.A1(\asqrt[51] ), .A2(new_n1044_), .A3(new_n1016_), .ZN(new_n1092_));
  XOR2_X1    g00900(.A1(new_n1092_), .A2(new_n978_), .Z(new_n1093_));
  AOI21_X1   g00901(.A1(new_n1009_), .A2(new_n1010_), .B(new_n1013_), .ZN(new_n1094_));
  NAND2_X1   g00902(.A1(\asqrt[51] ), .A2(new_n1094_), .ZN(new_n1095_));
  XOR2_X1    g00903(.A1(new_n1095_), .A2(new_n981_), .Z(new_n1096_));
  INV_X1     g00904(.I(new_n1096_), .ZN(new_n1097_));
  NOR2_X1    g00905(.A1(new_n1008_), .A2(\asqrt[56] ), .ZN(new_n1098_));
  NOR3_X1    g00906(.A1(new_n1088_), .A2(new_n1098_), .A3(new_n1042_), .ZN(new_n1099_));
  XOR2_X1    g00907(.A1(new_n1099_), .A2(new_n984_), .Z(new_n1100_));
  INV_X1     g00908(.I(new_n1100_), .ZN(new_n1101_));
  NOR3_X1    g00909(.A1(new_n1088_), .A2(new_n1003_), .A3(new_n1037_), .ZN(new_n1102_));
  XOR2_X1    g00910(.A1(new_n1102_), .A2(new_n1005_), .Z(new_n1103_));
  NAND2_X1   g00911(.A1(new_n1000_), .A2(new_n720_), .ZN(new_n1104_));
  NAND3_X1   g00912(.A1(\asqrt[51] ), .A2(new_n1104_), .A3(new_n1035_), .ZN(new_n1105_));
  XOR2_X1    g00913(.A1(new_n1105_), .A2(new_n991_), .Z(new_n1106_));
  NOR3_X1    g00914(.A1(new_n1088_), .A2(\a[102] ), .A3(\a[103] ), .ZN(new_n1107_));
  NAND4_X1   g00915(.A1(new_n1064_), .A2(\asqrt[52] ), .A3(new_n1066_), .A4(new_n966_), .ZN(new_n1108_));
  INV_X1     g00916(.I(new_n1108_), .ZN(new_n1109_));
  OAI21_X1   g00917(.A1(new_n1107_), .A2(new_n1109_), .B(new_n859_), .ZN(new_n1110_));
  NAND3_X1   g00918(.A1(\asqrt[51] ), .A2(new_n992_), .A3(new_n993_), .ZN(new_n1111_));
  NAND3_X1   g00919(.A1(new_n1111_), .A2(\a[104] ), .A3(new_n1108_), .ZN(new_n1112_));
  NAND2_X1   g00920(.A1(new_n1110_), .A2(new_n1112_), .ZN(new_n1113_));
  INV_X1     g00921(.I(\a[100] ), .ZN(new_n1114_));
  INV_X1     g00922(.I(\a[101] ), .ZN(new_n1115_));
  NAND3_X1   g00923(.A1(new_n1114_), .A2(new_n1115_), .A3(new_n992_), .ZN(new_n1116_));
  NAND2_X1   g00924(.A1(\asqrt[51] ), .A2(\a[102] ), .ZN(new_n1117_));
  AOI21_X1   g00925(.A1(new_n1117_), .A2(new_n1116_), .B(new_n962_), .ZN(new_n1118_));
  AOI21_X1   g00926(.A1(\asqrt[51] ), .A2(new_n992_), .B(new_n993_), .ZN(new_n1119_));
  NOR2_X1    g00927(.A1(new_n1107_), .A2(new_n1119_), .ZN(new_n1120_));
  NAND3_X1   g00928(.A1(new_n1117_), .A2(new_n962_), .A3(new_n1116_), .ZN(new_n1121_));
  AOI21_X1   g00929(.A1(new_n1120_), .A2(new_n1121_), .B(new_n1118_), .ZN(new_n1122_));
  AOI21_X1   g00930(.A1(new_n1122_), .A2(new_n842_), .B(new_n1113_), .ZN(new_n1123_));
  NOR2_X1    g00931(.A1(new_n1122_), .A2(new_n842_), .ZN(new_n1124_));
  NOR2_X1    g00932(.A1(new_n1123_), .A2(new_n1124_), .ZN(new_n1125_));
  NOR3_X1    g00933(.A1(new_n1088_), .A2(new_n996_), .A3(new_n1032_), .ZN(new_n1126_));
  XOR2_X1    g00934(.A1(new_n1126_), .A2(new_n998_), .Z(new_n1127_));
  INV_X1     g00935(.I(new_n1127_), .ZN(new_n1128_));
  AOI21_X1   g00936(.A1(new_n1125_), .A2(new_n720_), .B(new_n1128_), .ZN(new_n1129_));
  OAI21_X1   g00937(.A1(new_n1123_), .A2(new_n1124_), .B(\asqrt[54] ), .ZN(new_n1130_));
  NAND2_X1   g00938(.A1(new_n1130_), .A2(new_n630_), .ZN(new_n1131_));
  OAI21_X1   g00939(.A1(new_n1129_), .A2(new_n1131_), .B(new_n1106_), .ZN(new_n1132_));
  INV_X1     g00940(.I(new_n1130_), .ZN(new_n1133_));
  OAI21_X1   g00941(.A1(new_n1129_), .A2(new_n1133_), .B(\asqrt[55] ), .ZN(new_n1134_));
  NAND3_X1   g00942(.A1(new_n1132_), .A2(new_n1134_), .A3(new_n545_), .ZN(new_n1135_));
  NAND2_X1   g00943(.A1(new_n1135_), .A2(new_n1103_), .ZN(new_n1136_));
  NAND2_X1   g00944(.A1(new_n1132_), .A2(new_n1134_), .ZN(new_n1137_));
  AOI21_X1   g00945(.A1(new_n1137_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1138_));
  AOI21_X1   g00946(.A1(new_n1138_), .A2(new_n1136_), .B(new_n1101_), .ZN(new_n1139_));
  INV_X1     g00947(.I(new_n1106_), .ZN(new_n1140_));
  AOI21_X1   g00948(.A1(new_n1111_), .A2(new_n1108_), .B(\a[104] ), .ZN(new_n1141_));
  NOR3_X1    g00949(.A1(new_n1107_), .A2(new_n859_), .A3(new_n1109_), .ZN(new_n1142_));
  NOR2_X1    g00950(.A1(new_n1142_), .A2(new_n1141_), .ZN(new_n1143_));
  OAI21_X1   g00951(.A1(new_n1088_), .A2(new_n992_), .B(new_n1116_), .ZN(new_n1144_));
  NAND2_X1   g00952(.A1(new_n1144_), .A2(\asqrt[52] ), .ZN(new_n1145_));
  OAI21_X1   g00953(.A1(new_n1088_), .A2(\a[102] ), .B(\a[103] ), .ZN(new_n1146_));
  NAND2_X1   g00954(.A1(new_n1146_), .A2(new_n1111_), .ZN(new_n1147_));
  NOR2_X1    g00955(.A1(new_n1144_), .A2(\asqrt[52] ), .ZN(new_n1148_));
  OAI21_X1   g00956(.A1(new_n1147_), .A2(new_n1148_), .B(new_n1145_), .ZN(new_n1149_));
  OAI21_X1   g00957(.A1(new_n1149_), .A2(\asqrt[53] ), .B(new_n1143_), .ZN(new_n1150_));
  NAND2_X1   g00958(.A1(new_n1149_), .A2(\asqrt[53] ), .ZN(new_n1151_));
  NAND3_X1   g00959(.A1(new_n1150_), .A2(new_n720_), .A3(new_n1151_), .ZN(new_n1152_));
  NAND2_X1   g00960(.A1(new_n1152_), .A2(new_n1127_), .ZN(new_n1153_));
  NAND2_X1   g00961(.A1(new_n1150_), .A2(new_n1151_), .ZN(new_n1154_));
  AOI21_X1   g00962(.A1(new_n1154_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1155_));
  AOI21_X1   g00963(.A1(new_n1155_), .A2(new_n1153_), .B(new_n1140_), .ZN(new_n1156_));
  AOI21_X1   g00964(.A1(new_n1153_), .A2(new_n1130_), .B(new_n630_), .ZN(new_n1157_));
  OAI21_X1   g00965(.A1(new_n1156_), .A2(new_n1157_), .B(\asqrt[56] ), .ZN(new_n1158_));
  AOI21_X1   g00966(.A1(new_n1136_), .A2(new_n1158_), .B(new_n450_), .ZN(new_n1159_));
  NOR2_X1    g00967(.A1(new_n1139_), .A2(new_n1159_), .ZN(new_n1160_));
  AOI21_X1   g00968(.A1(new_n1160_), .A2(new_n403_), .B(new_n1097_), .ZN(new_n1161_));
  OAI21_X1   g00969(.A1(new_n1139_), .A2(new_n1159_), .B(\asqrt[58] ), .ZN(new_n1162_));
  NAND2_X1   g00970(.A1(new_n1162_), .A2(new_n339_), .ZN(new_n1163_));
  OAI21_X1   g00971(.A1(new_n1161_), .A2(new_n1163_), .B(new_n1093_), .ZN(new_n1164_));
  INV_X1     g00972(.I(new_n1162_), .ZN(new_n1165_));
  OAI21_X1   g00973(.A1(new_n1161_), .A2(new_n1165_), .B(\asqrt[59] ), .ZN(new_n1166_));
  NAND3_X1   g00974(.A1(new_n1164_), .A2(new_n1166_), .A3(new_n288_), .ZN(new_n1167_));
  NAND2_X1   g00975(.A1(new_n1167_), .A2(new_n1091_), .ZN(new_n1168_));
  INV_X1     g00976(.I(new_n1093_), .ZN(new_n1169_));
  INV_X1     g00977(.I(new_n1103_), .ZN(new_n1170_));
  NOR2_X1    g00978(.A1(new_n1156_), .A2(new_n1157_), .ZN(new_n1171_));
  AOI21_X1   g00979(.A1(new_n1171_), .A2(new_n545_), .B(new_n1170_), .ZN(new_n1172_));
  NAND2_X1   g00980(.A1(new_n1158_), .A2(new_n450_), .ZN(new_n1173_));
  OAI21_X1   g00981(.A1(new_n1172_), .A2(new_n1173_), .B(new_n1100_), .ZN(new_n1174_));
  INV_X1     g00982(.I(new_n1158_), .ZN(new_n1175_));
  OAI21_X1   g00983(.A1(new_n1172_), .A2(new_n1175_), .B(\asqrt[57] ), .ZN(new_n1176_));
  NAND3_X1   g00984(.A1(new_n1174_), .A2(new_n1176_), .A3(new_n403_), .ZN(new_n1177_));
  NAND2_X1   g00985(.A1(new_n1177_), .A2(new_n1096_), .ZN(new_n1178_));
  NAND2_X1   g00986(.A1(new_n1174_), .A2(new_n1176_), .ZN(new_n1179_));
  AOI21_X1   g00987(.A1(new_n1179_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1180_));
  AOI21_X1   g00988(.A1(new_n1180_), .A2(new_n1178_), .B(new_n1169_), .ZN(new_n1181_));
  AOI21_X1   g00989(.A1(new_n1178_), .A2(new_n1162_), .B(new_n339_), .ZN(new_n1182_));
  OAI21_X1   g00990(.A1(new_n1181_), .A2(new_n1182_), .B(\asqrt[60] ), .ZN(new_n1183_));
  AOI21_X1   g00991(.A1(new_n1168_), .A2(new_n1183_), .B(new_n242_), .ZN(new_n1184_));
  NAND3_X1   g00992(.A1(\asqrt[51] ), .A2(new_n1021_), .A3(new_n1050_), .ZN(new_n1185_));
  XOR2_X1    g00993(.A1(new_n1185_), .A2(new_n1075_), .Z(new_n1186_));
  INV_X1     g00994(.I(new_n1186_), .ZN(new_n1187_));
  NAND2_X1   g00995(.A1(new_n1164_), .A2(new_n1166_), .ZN(new_n1188_));
  AOI21_X1   g00996(.A1(new_n1188_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1189_));
  AOI21_X1   g00997(.A1(new_n1189_), .A2(new_n1168_), .B(new_n1187_), .ZN(new_n1190_));
  OAI21_X1   g00998(.A1(new_n1190_), .A2(new_n1184_), .B(\asqrt[62] ), .ZN(new_n1191_));
  INV_X1     g00999(.I(new_n1091_), .ZN(new_n1192_));
  NOR2_X1    g01000(.A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1193_));
  AOI21_X1   g01001(.A1(new_n1193_), .A2(new_n288_), .B(new_n1192_), .ZN(new_n1194_));
  INV_X1     g01002(.I(new_n1183_), .ZN(new_n1195_));
  OAI21_X1   g01003(.A1(new_n1194_), .A2(new_n1195_), .B(\asqrt[61] ), .ZN(new_n1196_));
  NAND2_X1   g01004(.A1(new_n1183_), .A2(new_n242_), .ZN(new_n1197_));
  OAI21_X1   g01005(.A1(new_n1194_), .A2(new_n1197_), .B(new_n1186_), .ZN(new_n1198_));
  NAND3_X1   g01006(.A1(new_n1198_), .A2(new_n1196_), .A3(new_n234_), .ZN(new_n1199_));
  NAND2_X1   g01007(.A1(new_n1086_), .A2(new_n968_), .ZN(new_n1200_));
  NOR2_X1    g01008(.A1(new_n1088_), .A2(new_n968_), .ZN(new_n1201_));
  NAND2_X1   g01009(.A1(new_n1201_), .A2(new_n1065_), .ZN(new_n1202_));
  AOI21_X1   g01010(.A1(new_n1202_), .A2(new_n1200_), .B(new_n193_), .ZN(new_n1203_));
  INV_X1     g01011(.I(new_n1203_), .ZN(new_n1204_));
  NAND3_X1   g01012(.A1(\asqrt[51] ), .A2(new_n1055_), .A3(new_n1082_), .ZN(new_n1205_));
  XOR2_X1    g01013(.A1(new_n1205_), .A2(new_n1060_), .Z(new_n1206_));
  INV_X1     g01014(.I(new_n1191_), .ZN(new_n1207_));
  AOI21_X1   g01015(.A1(new_n1201_), .A2(new_n1086_), .B(new_n1087_), .ZN(new_n1208_));
  INV_X1     g01016(.I(new_n1072_), .ZN(new_n1209_));
  NOR2_X1    g01017(.A1(new_n1190_), .A2(new_n1184_), .ZN(new_n1210_));
  AOI21_X1   g01018(.A1(new_n1210_), .A2(new_n234_), .B(new_n1209_), .ZN(new_n1211_));
  OAI21_X1   g01019(.A1(new_n1211_), .A2(new_n1207_), .B(new_n1208_), .ZN(new_n1212_));
  OAI21_X1   g01020(.A1(new_n1212_), .A2(new_n1206_), .B(new_n193_), .ZN(new_n1213_));
  NOR2_X1    g01021(.A1(new_n1211_), .A2(new_n1207_), .ZN(new_n1214_));
  NAND2_X1   g01022(.A1(new_n1214_), .A2(new_n1206_), .ZN(new_n1215_));
  NOR2_X1    g01023(.A1(\asqrt[51] ), .A2(new_n1073_), .ZN(new_n1216_));
  INV_X1     g01024(.I(new_n1216_), .ZN(new_n1217_));
  NAND4_X1   g01025(.A1(new_n1213_), .A2(new_n1204_), .A3(new_n1215_), .A4(new_n1217_), .ZN(\asqrt[50] ));
  NAND3_X1   g01026(.A1(\asqrt[50] ), .A2(new_n1191_), .A3(new_n1199_), .ZN(new_n1219_));
  XOR2_X1    g01027(.A1(new_n1219_), .A2(new_n1072_), .Z(new_n1220_));
  INV_X1     g01028(.I(new_n1206_), .ZN(new_n1221_));
  INV_X1     g01029(.I(new_n1208_), .ZN(new_n1222_));
  NAND2_X1   g01030(.A1(new_n1199_), .A2(new_n1072_), .ZN(new_n1223_));
  AOI21_X1   g01031(.A1(new_n1223_), .A2(new_n1191_), .B(new_n1222_), .ZN(new_n1224_));
  AOI21_X1   g01032(.A1(new_n1224_), .A2(new_n1221_), .B(\asqrt[63] ), .ZN(new_n1225_));
  NAND2_X1   g01033(.A1(new_n1223_), .A2(new_n1191_), .ZN(new_n1226_));
  NOR2_X1    g01034(.A1(new_n1226_), .A2(new_n1221_), .ZN(new_n1227_));
  NOR4_X1    g01035(.A1(new_n1225_), .A2(new_n1203_), .A3(new_n1227_), .A4(new_n1216_), .ZN(new_n1228_));
  OAI21_X1   g01036(.A1(new_n1161_), .A2(new_n1163_), .B(new_n1166_), .ZN(new_n1229_));
  NOR2_X1    g01037(.A1(new_n1228_), .A2(new_n1229_), .ZN(new_n1230_));
  XOR2_X1    g01038(.A1(new_n1230_), .A2(new_n1093_), .Z(new_n1231_));
  NAND3_X1   g01039(.A1(\asqrt[50] ), .A2(new_n1177_), .A3(new_n1162_), .ZN(new_n1232_));
  XOR2_X1    g01040(.A1(new_n1232_), .A2(new_n1097_), .Z(new_n1233_));
  OAI21_X1   g01041(.A1(new_n1172_), .A2(new_n1173_), .B(new_n1176_), .ZN(new_n1234_));
  NOR2_X1    g01042(.A1(new_n1228_), .A2(new_n1234_), .ZN(new_n1235_));
  XOR2_X1    g01043(.A1(new_n1235_), .A2(new_n1100_), .Z(new_n1236_));
  INV_X1     g01044(.I(new_n1236_), .ZN(new_n1237_));
  NAND3_X1   g01045(.A1(\asqrt[50] ), .A2(new_n1135_), .A3(new_n1158_), .ZN(new_n1238_));
  XOR2_X1    g01046(.A1(new_n1238_), .A2(new_n1170_), .Z(new_n1239_));
  INV_X1     g01047(.I(new_n1239_), .ZN(new_n1240_));
  OAI21_X1   g01048(.A1(new_n1129_), .A2(new_n1131_), .B(new_n1134_), .ZN(new_n1241_));
  NOR2_X1    g01049(.A1(new_n1228_), .A2(new_n1241_), .ZN(new_n1242_));
  XOR2_X1    g01050(.A1(new_n1242_), .A2(new_n1106_), .Z(new_n1243_));
  NAND3_X1   g01051(.A1(\asqrt[50] ), .A2(new_n1152_), .A3(new_n1130_), .ZN(new_n1244_));
  XOR2_X1    g01052(.A1(new_n1244_), .A2(new_n1128_), .Z(new_n1245_));
  NAND2_X1   g01053(.A1(new_n1122_), .A2(new_n842_), .ZN(new_n1246_));
  NAND3_X1   g01054(.A1(\asqrt[50] ), .A2(new_n1246_), .A3(new_n1151_), .ZN(new_n1247_));
  XOR2_X1    g01055(.A1(new_n1247_), .A2(new_n1113_), .Z(new_n1248_));
  INV_X1     g01056(.I(new_n1248_), .ZN(new_n1249_));
  NAND3_X1   g01057(.A1(\asqrt[50] ), .A2(new_n1114_), .A3(new_n1115_), .ZN(new_n1250_));
  NOR4_X1    g01058(.A1(new_n1225_), .A2(new_n1088_), .A3(new_n1203_), .A4(new_n1227_), .ZN(new_n1251_));
  INV_X1     g01059(.I(new_n1251_), .ZN(new_n1252_));
  AOI21_X1   g01060(.A1(new_n1250_), .A2(new_n1252_), .B(\a[102] ), .ZN(new_n1253_));
  NOR3_X1    g01061(.A1(new_n1228_), .A2(\a[100] ), .A3(\a[101] ), .ZN(new_n1254_));
  NOR3_X1    g01062(.A1(new_n1254_), .A2(new_n992_), .A3(new_n1251_), .ZN(new_n1255_));
  NOR2_X1    g01063(.A1(new_n1255_), .A2(new_n1253_), .ZN(new_n1256_));
  INV_X1     g01064(.I(\a[98] ), .ZN(new_n1257_));
  INV_X1     g01065(.I(\a[99] ), .ZN(new_n1258_));
  NAND3_X1   g01066(.A1(new_n1257_), .A2(new_n1258_), .A3(new_n1114_), .ZN(new_n1259_));
  OAI21_X1   g01067(.A1(new_n1228_), .A2(new_n1114_), .B(new_n1259_), .ZN(new_n1260_));
  NAND2_X1   g01068(.A1(new_n1260_), .A2(\asqrt[51] ), .ZN(new_n1261_));
  OAI21_X1   g01069(.A1(new_n1228_), .A2(\a[100] ), .B(\a[101] ), .ZN(new_n1262_));
  NAND2_X1   g01070(.A1(new_n1262_), .A2(new_n1250_), .ZN(new_n1263_));
  NOR2_X1    g01071(.A1(new_n1260_), .A2(\asqrt[51] ), .ZN(new_n1264_));
  OAI21_X1   g01072(.A1(new_n1263_), .A2(new_n1264_), .B(new_n1261_), .ZN(new_n1265_));
  OAI21_X1   g01073(.A1(new_n1265_), .A2(\asqrt[52] ), .B(new_n1256_), .ZN(new_n1266_));
  NAND2_X1   g01074(.A1(new_n1265_), .A2(\asqrt[52] ), .ZN(new_n1267_));
  NAND3_X1   g01075(.A1(new_n1266_), .A2(new_n842_), .A3(new_n1267_), .ZN(new_n1268_));
  NOR3_X1    g01076(.A1(new_n1228_), .A2(new_n1118_), .A3(new_n1148_), .ZN(new_n1269_));
  XOR2_X1    g01077(.A1(new_n1269_), .A2(new_n1120_), .Z(new_n1270_));
  AOI21_X1   g01078(.A1(new_n1266_), .A2(new_n1267_), .B(new_n842_), .ZN(new_n1271_));
  AOI21_X1   g01079(.A1(new_n1268_), .A2(new_n1270_), .B(new_n1271_), .ZN(new_n1272_));
  AOI21_X1   g01080(.A1(new_n1272_), .A2(new_n720_), .B(new_n1249_), .ZN(new_n1273_));
  OAI21_X1   g01081(.A1(new_n1272_), .A2(new_n720_), .B(new_n630_), .ZN(new_n1274_));
  OAI21_X1   g01082(.A1(new_n1273_), .A2(new_n1274_), .B(new_n1245_), .ZN(new_n1275_));
  NOR2_X1    g01083(.A1(new_n1272_), .A2(new_n720_), .ZN(new_n1276_));
  OAI21_X1   g01084(.A1(new_n1273_), .A2(new_n1276_), .B(\asqrt[55] ), .ZN(new_n1277_));
  NAND3_X1   g01085(.A1(new_n1275_), .A2(new_n1277_), .A3(new_n545_), .ZN(new_n1278_));
  NAND2_X1   g01086(.A1(new_n1278_), .A2(new_n1243_), .ZN(new_n1279_));
  NAND2_X1   g01087(.A1(new_n1275_), .A2(new_n1277_), .ZN(new_n1280_));
  AOI21_X1   g01088(.A1(new_n1280_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1281_));
  AOI21_X1   g01089(.A1(new_n1281_), .A2(new_n1279_), .B(new_n1240_), .ZN(new_n1282_));
  INV_X1     g01090(.I(new_n1245_), .ZN(new_n1283_));
  OAI21_X1   g01091(.A1(new_n1254_), .A2(new_n1251_), .B(new_n992_), .ZN(new_n1284_));
  NAND3_X1   g01092(.A1(new_n1250_), .A2(new_n1252_), .A3(\a[102] ), .ZN(new_n1285_));
  NAND2_X1   g01093(.A1(new_n1284_), .A2(new_n1285_), .ZN(new_n1286_));
  NAND2_X1   g01094(.A1(\asqrt[50] ), .A2(\a[100] ), .ZN(new_n1287_));
  AOI21_X1   g01095(.A1(new_n1287_), .A2(new_n1259_), .B(new_n1088_), .ZN(new_n1288_));
  AOI21_X1   g01096(.A1(\asqrt[50] ), .A2(new_n1114_), .B(new_n1115_), .ZN(new_n1289_));
  NOR2_X1    g01097(.A1(new_n1254_), .A2(new_n1289_), .ZN(new_n1290_));
  NAND3_X1   g01098(.A1(new_n1287_), .A2(new_n1088_), .A3(new_n1259_), .ZN(new_n1291_));
  AOI21_X1   g01099(.A1(new_n1290_), .A2(new_n1291_), .B(new_n1288_), .ZN(new_n1292_));
  AOI21_X1   g01100(.A1(new_n1292_), .A2(new_n962_), .B(new_n1286_), .ZN(new_n1293_));
  NOR2_X1    g01101(.A1(new_n1292_), .A2(new_n962_), .ZN(new_n1294_));
  NOR3_X1    g01102(.A1(new_n1293_), .A2(\asqrt[53] ), .A3(new_n1294_), .ZN(new_n1295_));
  INV_X1     g01103(.I(new_n1270_), .ZN(new_n1296_));
  OAI21_X1   g01104(.A1(new_n1293_), .A2(new_n1294_), .B(\asqrt[53] ), .ZN(new_n1297_));
  OAI21_X1   g01105(.A1(new_n1295_), .A2(new_n1296_), .B(new_n1297_), .ZN(new_n1298_));
  OAI21_X1   g01106(.A1(new_n1298_), .A2(\asqrt[54] ), .B(new_n1248_), .ZN(new_n1299_));
  AOI21_X1   g01107(.A1(new_n1298_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1300_));
  AOI21_X1   g01108(.A1(new_n1300_), .A2(new_n1299_), .B(new_n1283_), .ZN(new_n1301_));
  NAND2_X1   g01109(.A1(new_n1298_), .A2(\asqrt[54] ), .ZN(new_n1302_));
  AOI21_X1   g01110(.A1(new_n1299_), .A2(new_n1302_), .B(new_n630_), .ZN(new_n1303_));
  OAI21_X1   g01111(.A1(new_n1301_), .A2(new_n1303_), .B(\asqrt[56] ), .ZN(new_n1304_));
  AOI21_X1   g01112(.A1(new_n1279_), .A2(new_n1304_), .B(new_n450_), .ZN(new_n1305_));
  NOR2_X1    g01113(.A1(new_n1282_), .A2(new_n1305_), .ZN(new_n1306_));
  AOI21_X1   g01114(.A1(new_n1306_), .A2(new_n403_), .B(new_n1237_), .ZN(new_n1307_));
  OAI21_X1   g01115(.A1(new_n1282_), .A2(new_n1305_), .B(\asqrt[58] ), .ZN(new_n1308_));
  NAND2_X1   g01116(.A1(new_n1308_), .A2(new_n339_), .ZN(new_n1309_));
  OAI21_X1   g01117(.A1(new_n1307_), .A2(new_n1309_), .B(new_n1233_), .ZN(new_n1310_));
  INV_X1     g01118(.I(new_n1308_), .ZN(new_n1311_));
  OAI21_X1   g01119(.A1(new_n1307_), .A2(new_n1311_), .B(\asqrt[59] ), .ZN(new_n1312_));
  NAND3_X1   g01120(.A1(new_n1310_), .A2(new_n1312_), .A3(new_n288_), .ZN(new_n1313_));
  NAND2_X1   g01121(.A1(new_n1313_), .A2(new_n1231_), .ZN(new_n1314_));
  INV_X1     g01122(.I(new_n1233_), .ZN(new_n1315_));
  INV_X1     g01123(.I(new_n1243_), .ZN(new_n1316_));
  NOR2_X1    g01124(.A1(new_n1301_), .A2(new_n1303_), .ZN(new_n1317_));
  AOI21_X1   g01125(.A1(new_n1317_), .A2(new_n545_), .B(new_n1316_), .ZN(new_n1318_));
  NAND2_X1   g01126(.A1(new_n1304_), .A2(new_n450_), .ZN(new_n1319_));
  OAI21_X1   g01127(.A1(new_n1318_), .A2(new_n1319_), .B(new_n1239_), .ZN(new_n1320_));
  INV_X1     g01128(.I(new_n1304_), .ZN(new_n1321_));
  OAI21_X1   g01129(.A1(new_n1318_), .A2(new_n1321_), .B(\asqrt[57] ), .ZN(new_n1322_));
  NAND3_X1   g01130(.A1(new_n1320_), .A2(new_n1322_), .A3(new_n403_), .ZN(new_n1323_));
  NAND2_X1   g01131(.A1(new_n1323_), .A2(new_n1236_), .ZN(new_n1324_));
  NAND2_X1   g01132(.A1(new_n1320_), .A2(new_n1322_), .ZN(new_n1325_));
  AOI21_X1   g01133(.A1(new_n1325_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1326_));
  AOI21_X1   g01134(.A1(new_n1326_), .A2(new_n1324_), .B(new_n1315_), .ZN(new_n1327_));
  AOI21_X1   g01135(.A1(new_n1324_), .A2(new_n1308_), .B(new_n339_), .ZN(new_n1328_));
  OAI21_X1   g01136(.A1(new_n1327_), .A2(new_n1328_), .B(\asqrt[60] ), .ZN(new_n1329_));
  AOI21_X1   g01137(.A1(new_n1314_), .A2(new_n1329_), .B(new_n242_), .ZN(new_n1330_));
  NAND3_X1   g01138(.A1(\asqrt[50] ), .A2(new_n1167_), .A3(new_n1183_), .ZN(new_n1331_));
  XOR2_X1    g01139(.A1(new_n1331_), .A2(new_n1192_), .Z(new_n1332_));
  INV_X1     g01140(.I(new_n1332_), .ZN(new_n1333_));
  NAND2_X1   g01141(.A1(new_n1310_), .A2(new_n1312_), .ZN(new_n1334_));
  AOI21_X1   g01142(.A1(new_n1334_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1335_));
  AOI21_X1   g01143(.A1(new_n1335_), .A2(new_n1314_), .B(new_n1333_), .ZN(new_n1336_));
  OAI21_X1   g01144(.A1(new_n1336_), .A2(new_n1330_), .B(\asqrt[62] ), .ZN(new_n1337_));
  AOI21_X1   g01145(.A1(new_n1168_), .A2(new_n1189_), .B(new_n1184_), .ZN(new_n1338_));
  NAND2_X1   g01146(.A1(\asqrt[50] ), .A2(new_n1338_), .ZN(new_n1339_));
  XOR2_X1    g01147(.A1(new_n1339_), .A2(new_n1187_), .Z(new_n1340_));
  INV_X1     g01148(.I(new_n1231_), .ZN(new_n1341_));
  NOR2_X1    g01149(.A1(new_n1327_), .A2(new_n1328_), .ZN(new_n1342_));
  AOI21_X1   g01150(.A1(new_n1342_), .A2(new_n288_), .B(new_n1341_), .ZN(new_n1343_));
  INV_X1     g01151(.I(new_n1329_), .ZN(new_n1344_));
  OAI21_X1   g01152(.A1(new_n1343_), .A2(new_n1344_), .B(\asqrt[61] ), .ZN(new_n1345_));
  NAND2_X1   g01153(.A1(new_n1329_), .A2(new_n242_), .ZN(new_n1346_));
  OAI21_X1   g01154(.A1(new_n1343_), .A2(new_n1346_), .B(new_n1332_), .ZN(new_n1347_));
  NAND3_X1   g01155(.A1(new_n1347_), .A2(new_n1345_), .A3(new_n234_), .ZN(new_n1348_));
  NAND2_X1   g01156(.A1(new_n1348_), .A2(new_n1340_), .ZN(new_n1349_));
  NAND2_X1   g01157(.A1(new_n1349_), .A2(new_n1337_), .ZN(new_n1350_));
  NAND2_X1   g01158(.A1(new_n1350_), .A2(new_n1220_), .ZN(new_n1351_));
  INV_X1     g01159(.I(new_n1337_), .ZN(new_n1352_));
  NOR2_X1    g01160(.A1(new_n1336_), .A2(new_n1330_), .ZN(new_n1353_));
  INV_X1     g01161(.I(new_n1340_), .ZN(new_n1354_));
  AOI21_X1   g01162(.A1(new_n1353_), .A2(new_n234_), .B(new_n1354_), .ZN(new_n1355_));
  NOR2_X1    g01163(.A1(new_n1355_), .A2(new_n1352_), .ZN(new_n1356_));
  NAND2_X1   g01164(.A1(new_n1226_), .A2(new_n1206_), .ZN(new_n1357_));
  NOR2_X1    g01165(.A1(new_n1228_), .A2(new_n1206_), .ZN(new_n1358_));
  NAND2_X1   g01166(.A1(new_n1358_), .A2(new_n1214_), .ZN(new_n1359_));
  AOI21_X1   g01167(.A1(new_n1359_), .A2(new_n1357_), .B(new_n193_), .ZN(new_n1360_));
  INV_X1     g01168(.I(new_n1220_), .ZN(new_n1361_));
  AOI21_X1   g01169(.A1(new_n1358_), .A2(new_n1226_), .B(new_n1227_), .ZN(new_n1362_));
  INV_X1     g01170(.I(new_n1362_), .ZN(new_n1363_));
  AOI21_X1   g01171(.A1(new_n1349_), .A2(new_n1337_), .B(new_n1363_), .ZN(new_n1364_));
  AOI21_X1   g01172(.A1(new_n1364_), .A2(new_n1361_), .B(\asqrt[63] ), .ZN(new_n1365_));
  NOR2_X1    g01173(.A1(new_n1350_), .A2(new_n1361_), .ZN(new_n1366_));
  NOR2_X1    g01174(.A1(\asqrt[50] ), .A2(new_n1221_), .ZN(new_n1367_));
  NOR4_X1    g01175(.A1(new_n1365_), .A2(new_n1360_), .A3(new_n1366_), .A4(new_n1367_), .ZN(new_n1368_));
  NOR2_X1    g01176(.A1(new_n1368_), .A2(new_n1220_), .ZN(new_n1369_));
  NAND2_X1   g01177(.A1(new_n1369_), .A2(new_n1356_), .ZN(new_n1370_));
  AOI21_X1   g01178(.A1(new_n1370_), .A2(new_n1351_), .B(new_n193_), .ZN(new_n1371_));
  INV_X1     g01179(.I(new_n1371_), .ZN(new_n1372_));
  INV_X1     g01180(.I(new_n1360_), .ZN(new_n1373_));
  OAI21_X1   g01181(.A1(new_n1355_), .A2(new_n1352_), .B(new_n1362_), .ZN(new_n1374_));
  OAI21_X1   g01182(.A1(new_n1374_), .A2(new_n1220_), .B(new_n193_), .ZN(new_n1375_));
  NAND2_X1   g01183(.A1(new_n1356_), .A2(new_n1220_), .ZN(new_n1376_));
  INV_X1     g01184(.I(new_n1367_), .ZN(new_n1377_));
  NAND4_X1   g01185(.A1(new_n1375_), .A2(new_n1373_), .A3(new_n1376_), .A4(new_n1377_), .ZN(\asqrt[49] ));
  NAND3_X1   g01186(.A1(\asqrt[49] ), .A2(new_n1337_), .A3(new_n1348_), .ZN(new_n1379_));
  XOR2_X1    g01187(.A1(new_n1379_), .A2(new_n1340_), .Z(new_n1380_));
  AOI21_X1   g01188(.A1(new_n1369_), .A2(new_n1350_), .B(new_n1366_), .ZN(new_n1381_));
  OAI21_X1   g01189(.A1(new_n1307_), .A2(new_n1309_), .B(new_n1312_), .ZN(new_n1382_));
  NOR2_X1    g01190(.A1(new_n1368_), .A2(new_n1382_), .ZN(new_n1383_));
  XOR2_X1    g01191(.A1(new_n1383_), .A2(new_n1233_), .Z(new_n1384_));
  NAND3_X1   g01192(.A1(\asqrt[49] ), .A2(new_n1323_), .A3(new_n1308_), .ZN(new_n1385_));
  XOR2_X1    g01193(.A1(new_n1385_), .A2(new_n1237_), .Z(new_n1386_));
  OAI21_X1   g01194(.A1(new_n1318_), .A2(new_n1319_), .B(new_n1322_), .ZN(new_n1387_));
  NOR2_X1    g01195(.A1(new_n1368_), .A2(new_n1387_), .ZN(new_n1388_));
  XOR2_X1    g01196(.A1(new_n1388_), .A2(new_n1239_), .Z(new_n1389_));
  INV_X1     g01197(.I(new_n1389_), .ZN(new_n1390_));
  NAND3_X1   g01198(.A1(\asqrt[49] ), .A2(new_n1278_), .A3(new_n1304_), .ZN(new_n1391_));
  XOR2_X1    g01199(.A1(new_n1391_), .A2(new_n1316_), .Z(new_n1392_));
  INV_X1     g01200(.I(new_n1392_), .ZN(new_n1393_));
  AOI21_X1   g01201(.A1(new_n1299_), .A2(new_n1300_), .B(new_n1303_), .ZN(new_n1394_));
  NAND2_X1   g01202(.A1(\asqrt[49] ), .A2(new_n1394_), .ZN(new_n1395_));
  XOR2_X1    g01203(.A1(new_n1395_), .A2(new_n1283_), .Z(new_n1396_));
  NOR2_X1    g01204(.A1(new_n1298_), .A2(\asqrt[54] ), .ZN(new_n1397_));
  NOR3_X1    g01205(.A1(new_n1368_), .A2(new_n1397_), .A3(new_n1276_), .ZN(new_n1398_));
  XOR2_X1    g01206(.A1(new_n1398_), .A2(new_n1248_), .Z(new_n1399_));
  NOR3_X1    g01207(.A1(new_n1368_), .A2(new_n1295_), .A3(new_n1271_), .ZN(new_n1400_));
  XOR2_X1    g01208(.A1(new_n1400_), .A2(new_n1270_), .Z(new_n1401_));
  INV_X1     g01209(.I(new_n1401_), .ZN(new_n1402_));
  NAND2_X1   g01210(.A1(new_n1292_), .A2(new_n962_), .ZN(new_n1403_));
  NAND3_X1   g01211(.A1(\asqrt[49] ), .A2(new_n1403_), .A3(new_n1267_), .ZN(new_n1404_));
  XOR2_X1    g01212(.A1(new_n1404_), .A2(new_n1286_), .Z(new_n1405_));
  INV_X1     g01213(.I(new_n1405_), .ZN(new_n1406_));
  NAND3_X1   g01214(.A1(\asqrt[49] ), .A2(new_n1257_), .A3(new_n1258_), .ZN(new_n1407_));
  NOR4_X1    g01215(.A1(new_n1365_), .A2(new_n1228_), .A3(new_n1360_), .A4(new_n1366_), .ZN(new_n1408_));
  INV_X1     g01216(.I(new_n1408_), .ZN(new_n1409_));
  AOI21_X1   g01217(.A1(new_n1407_), .A2(new_n1409_), .B(\a[100] ), .ZN(new_n1410_));
  NOR3_X1    g01218(.A1(new_n1368_), .A2(\a[98] ), .A3(\a[99] ), .ZN(new_n1411_));
  NOR3_X1    g01219(.A1(new_n1411_), .A2(new_n1114_), .A3(new_n1408_), .ZN(new_n1412_));
  NOR2_X1    g01220(.A1(new_n1412_), .A2(new_n1410_), .ZN(new_n1413_));
  NAND3_X1   g01221(.A1(new_n197_), .A2(new_n198_), .A3(new_n1257_), .ZN(new_n1414_));
  OAI21_X1   g01222(.A1(new_n1368_), .A2(new_n1257_), .B(new_n1414_), .ZN(new_n1415_));
  NAND2_X1   g01223(.A1(new_n1415_), .A2(\asqrt[50] ), .ZN(new_n1416_));
  OAI21_X1   g01224(.A1(new_n1368_), .A2(\a[98] ), .B(\a[99] ), .ZN(new_n1417_));
  NAND2_X1   g01225(.A1(new_n1417_), .A2(new_n1407_), .ZN(new_n1418_));
  NOR2_X1    g01226(.A1(new_n1415_), .A2(\asqrt[50] ), .ZN(new_n1419_));
  OAI21_X1   g01227(.A1(new_n1418_), .A2(new_n1419_), .B(new_n1416_), .ZN(new_n1420_));
  OAI21_X1   g01228(.A1(\asqrt[51] ), .A2(new_n1420_), .B(new_n1413_), .ZN(new_n1421_));
  NAND2_X1   g01229(.A1(new_n1420_), .A2(\asqrt[51] ), .ZN(new_n1422_));
  NAND3_X1   g01230(.A1(new_n1421_), .A2(new_n962_), .A3(new_n1422_), .ZN(new_n1423_));
  NOR3_X1    g01231(.A1(new_n1368_), .A2(new_n1288_), .A3(new_n1264_), .ZN(new_n1424_));
  XOR2_X1    g01232(.A1(new_n1424_), .A2(new_n1290_), .Z(new_n1425_));
  NAND2_X1   g01233(.A1(new_n1423_), .A2(new_n1425_), .ZN(new_n1426_));
  NAND2_X1   g01234(.A1(new_n1421_), .A2(new_n1422_), .ZN(new_n1427_));
  AOI21_X1   g01235(.A1(new_n1427_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n1428_));
  AOI21_X1   g01236(.A1(new_n1428_), .A2(new_n1426_), .B(new_n1406_), .ZN(new_n1429_));
  OAI21_X1   g01237(.A1(new_n1411_), .A2(new_n1408_), .B(new_n1114_), .ZN(new_n1430_));
  NAND3_X1   g01238(.A1(new_n1407_), .A2(\a[100] ), .A3(new_n1409_), .ZN(new_n1431_));
  NAND2_X1   g01239(.A1(new_n1430_), .A2(new_n1431_), .ZN(new_n1432_));
  NAND2_X1   g01240(.A1(\asqrt[49] ), .A2(\a[98] ), .ZN(new_n1433_));
  AOI21_X1   g01241(.A1(new_n1433_), .A2(new_n1414_), .B(new_n1228_), .ZN(new_n1434_));
  AOI21_X1   g01242(.A1(\asqrt[49] ), .A2(new_n1257_), .B(new_n1258_), .ZN(new_n1435_));
  NOR2_X1    g01243(.A1(new_n1435_), .A2(new_n1411_), .ZN(new_n1436_));
  NAND3_X1   g01244(.A1(new_n1433_), .A2(new_n1228_), .A3(new_n1414_), .ZN(new_n1437_));
  AOI21_X1   g01245(.A1(new_n1436_), .A2(new_n1437_), .B(new_n1434_), .ZN(new_n1438_));
  AOI21_X1   g01246(.A1(new_n1438_), .A2(new_n1088_), .B(new_n1432_), .ZN(new_n1439_));
  NOR2_X1    g01247(.A1(new_n1438_), .A2(new_n1088_), .ZN(new_n1440_));
  OAI21_X1   g01248(.A1(new_n1439_), .A2(new_n1440_), .B(\asqrt[52] ), .ZN(new_n1441_));
  AOI21_X1   g01249(.A1(new_n1426_), .A2(new_n1441_), .B(new_n842_), .ZN(new_n1442_));
  NOR2_X1    g01250(.A1(new_n1429_), .A2(new_n1442_), .ZN(new_n1443_));
  AOI21_X1   g01251(.A1(new_n1443_), .A2(new_n720_), .B(new_n1402_), .ZN(new_n1444_));
  OAI21_X1   g01252(.A1(new_n1429_), .A2(new_n1442_), .B(\asqrt[54] ), .ZN(new_n1445_));
  NAND2_X1   g01253(.A1(new_n1445_), .A2(new_n630_), .ZN(new_n1446_));
  OAI21_X1   g01254(.A1(new_n1444_), .A2(new_n1446_), .B(new_n1399_), .ZN(new_n1447_));
  INV_X1     g01255(.I(new_n1445_), .ZN(new_n1448_));
  OAI21_X1   g01256(.A1(new_n1444_), .A2(new_n1448_), .B(\asqrt[55] ), .ZN(new_n1449_));
  NAND3_X1   g01257(.A1(new_n1447_), .A2(new_n1449_), .A3(new_n545_), .ZN(new_n1450_));
  NAND2_X1   g01258(.A1(new_n1450_), .A2(new_n1396_), .ZN(new_n1451_));
  NAND2_X1   g01259(.A1(new_n1447_), .A2(new_n1449_), .ZN(new_n1452_));
  AOI21_X1   g01260(.A1(new_n1452_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1453_));
  AOI21_X1   g01261(.A1(new_n1453_), .A2(new_n1451_), .B(new_n1393_), .ZN(new_n1454_));
  INV_X1     g01262(.I(new_n1399_), .ZN(new_n1455_));
  NOR2_X1    g01263(.A1(new_n1439_), .A2(new_n1440_), .ZN(new_n1456_));
  INV_X1     g01264(.I(new_n1425_), .ZN(new_n1457_));
  AOI21_X1   g01265(.A1(new_n1456_), .A2(new_n962_), .B(new_n1457_), .ZN(new_n1458_));
  NAND2_X1   g01266(.A1(new_n1441_), .A2(new_n842_), .ZN(new_n1459_));
  OAI21_X1   g01267(.A1(new_n1458_), .A2(new_n1459_), .B(new_n1405_), .ZN(new_n1460_));
  INV_X1     g01268(.I(new_n1441_), .ZN(new_n1461_));
  OAI21_X1   g01269(.A1(new_n1458_), .A2(new_n1461_), .B(\asqrt[53] ), .ZN(new_n1462_));
  NAND3_X1   g01270(.A1(new_n1460_), .A2(new_n1462_), .A3(new_n720_), .ZN(new_n1463_));
  NAND2_X1   g01271(.A1(new_n1463_), .A2(new_n1401_), .ZN(new_n1464_));
  NAND2_X1   g01272(.A1(new_n1460_), .A2(new_n1462_), .ZN(new_n1465_));
  AOI21_X1   g01273(.A1(new_n1465_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1466_));
  AOI21_X1   g01274(.A1(new_n1466_), .A2(new_n1464_), .B(new_n1455_), .ZN(new_n1467_));
  AOI21_X1   g01275(.A1(new_n1464_), .A2(new_n1445_), .B(new_n630_), .ZN(new_n1468_));
  OAI21_X1   g01276(.A1(new_n1467_), .A2(new_n1468_), .B(\asqrt[56] ), .ZN(new_n1469_));
  AOI21_X1   g01277(.A1(new_n1451_), .A2(new_n1469_), .B(new_n450_), .ZN(new_n1470_));
  NOR2_X1    g01278(.A1(new_n1454_), .A2(new_n1470_), .ZN(new_n1471_));
  AOI21_X1   g01279(.A1(new_n1471_), .A2(new_n403_), .B(new_n1390_), .ZN(new_n1472_));
  OAI21_X1   g01280(.A1(new_n1454_), .A2(new_n1470_), .B(\asqrt[58] ), .ZN(new_n1473_));
  NAND2_X1   g01281(.A1(new_n1473_), .A2(new_n339_), .ZN(new_n1474_));
  OAI21_X1   g01282(.A1(new_n1472_), .A2(new_n1474_), .B(new_n1386_), .ZN(new_n1475_));
  INV_X1     g01283(.I(new_n1473_), .ZN(new_n1476_));
  OAI21_X1   g01284(.A1(new_n1472_), .A2(new_n1476_), .B(\asqrt[59] ), .ZN(new_n1477_));
  NAND3_X1   g01285(.A1(new_n1475_), .A2(new_n1477_), .A3(new_n288_), .ZN(new_n1478_));
  NAND2_X1   g01286(.A1(new_n1478_), .A2(new_n1384_), .ZN(new_n1479_));
  INV_X1     g01287(.I(new_n1386_), .ZN(new_n1480_));
  INV_X1     g01288(.I(new_n1396_), .ZN(new_n1481_));
  NOR2_X1    g01289(.A1(new_n1467_), .A2(new_n1468_), .ZN(new_n1482_));
  AOI21_X1   g01290(.A1(new_n1482_), .A2(new_n545_), .B(new_n1481_), .ZN(new_n1483_));
  NAND2_X1   g01291(.A1(new_n1469_), .A2(new_n450_), .ZN(new_n1484_));
  OAI21_X1   g01292(.A1(new_n1483_), .A2(new_n1484_), .B(new_n1392_), .ZN(new_n1485_));
  INV_X1     g01293(.I(new_n1469_), .ZN(new_n1486_));
  OAI21_X1   g01294(.A1(new_n1483_), .A2(new_n1486_), .B(\asqrt[57] ), .ZN(new_n1487_));
  NAND3_X1   g01295(.A1(new_n1485_), .A2(new_n1487_), .A3(new_n403_), .ZN(new_n1488_));
  NAND2_X1   g01296(.A1(new_n1488_), .A2(new_n1389_), .ZN(new_n1489_));
  NAND2_X1   g01297(.A1(new_n1485_), .A2(new_n1487_), .ZN(new_n1490_));
  AOI21_X1   g01298(.A1(new_n1490_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1491_));
  AOI21_X1   g01299(.A1(new_n1491_), .A2(new_n1489_), .B(new_n1480_), .ZN(new_n1492_));
  AOI21_X1   g01300(.A1(new_n1489_), .A2(new_n1473_), .B(new_n339_), .ZN(new_n1493_));
  OAI21_X1   g01301(.A1(new_n1492_), .A2(new_n1493_), .B(\asqrt[60] ), .ZN(new_n1494_));
  AOI21_X1   g01302(.A1(new_n1479_), .A2(new_n1494_), .B(new_n242_), .ZN(new_n1495_));
  NAND3_X1   g01303(.A1(\asqrt[49] ), .A2(new_n1313_), .A3(new_n1329_), .ZN(new_n1496_));
  XOR2_X1    g01304(.A1(new_n1496_), .A2(new_n1341_), .Z(new_n1497_));
  INV_X1     g01305(.I(new_n1497_), .ZN(new_n1498_));
  NAND2_X1   g01306(.A1(new_n1475_), .A2(new_n1477_), .ZN(new_n1499_));
  AOI21_X1   g01307(.A1(new_n1499_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1500_));
  AOI21_X1   g01308(.A1(new_n1500_), .A2(new_n1479_), .B(new_n1498_), .ZN(new_n1501_));
  OAI21_X1   g01309(.A1(new_n1501_), .A2(new_n1495_), .B(\asqrt[62] ), .ZN(new_n1502_));
  INV_X1     g01310(.I(new_n1502_), .ZN(new_n1503_));
  NOR2_X1    g01311(.A1(new_n1501_), .A2(new_n1495_), .ZN(new_n1504_));
  AOI21_X1   g01312(.A1(new_n1314_), .A2(new_n1335_), .B(new_n1330_), .ZN(new_n1505_));
  NAND2_X1   g01313(.A1(\asqrt[49] ), .A2(new_n1505_), .ZN(new_n1506_));
  XOR2_X1    g01314(.A1(new_n1506_), .A2(new_n1333_), .Z(new_n1507_));
  INV_X1     g01315(.I(new_n1507_), .ZN(new_n1508_));
  AOI21_X1   g01316(.A1(new_n1504_), .A2(new_n234_), .B(new_n1508_), .ZN(new_n1509_));
  OAI21_X1   g01317(.A1(new_n1509_), .A2(new_n1503_), .B(new_n1381_), .ZN(new_n1510_));
  OAI21_X1   g01318(.A1(new_n1510_), .A2(new_n1380_), .B(new_n193_), .ZN(new_n1511_));
  NOR2_X1    g01319(.A1(new_n1509_), .A2(new_n1503_), .ZN(new_n1512_));
  NAND2_X1   g01320(.A1(new_n1512_), .A2(new_n1380_), .ZN(new_n1513_));
  NOR2_X1    g01321(.A1(\asqrt[49] ), .A2(new_n1361_), .ZN(new_n1514_));
  INV_X1     g01322(.I(new_n1514_), .ZN(new_n1515_));
  NAND4_X1   g01323(.A1(new_n1511_), .A2(new_n1372_), .A3(new_n1513_), .A4(new_n1515_), .ZN(\asqrt[48] ));
  AOI21_X1   g01324(.A1(\asqrt[48] ), .A2(new_n197_), .B(new_n198_), .ZN(new_n1517_));
  INV_X1     g01325(.I(new_n1380_), .ZN(new_n1518_));
  INV_X1     g01326(.I(new_n1381_), .ZN(new_n1519_));
  INV_X1     g01327(.I(new_n1384_), .ZN(new_n1520_));
  NOR2_X1    g01328(.A1(new_n1492_), .A2(new_n1493_), .ZN(new_n1521_));
  AOI21_X1   g01329(.A1(new_n1521_), .A2(new_n288_), .B(new_n1520_), .ZN(new_n1522_));
  INV_X1     g01330(.I(new_n1494_), .ZN(new_n1523_));
  OAI21_X1   g01331(.A1(new_n1522_), .A2(new_n1523_), .B(\asqrt[61] ), .ZN(new_n1524_));
  NAND2_X1   g01332(.A1(new_n1494_), .A2(new_n242_), .ZN(new_n1525_));
  OAI21_X1   g01333(.A1(new_n1522_), .A2(new_n1525_), .B(new_n1497_), .ZN(new_n1526_));
  NAND3_X1   g01334(.A1(new_n1526_), .A2(new_n1524_), .A3(new_n234_), .ZN(new_n1527_));
  NAND2_X1   g01335(.A1(new_n1527_), .A2(new_n1507_), .ZN(new_n1528_));
  AOI21_X1   g01336(.A1(new_n1528_), .A2(new_n1502_), .B(new_n1519_), .ZN(new_n1529_));
  AOI21_X1   g01337(.A1(new_n1529_), .A2(new_n1518_), .B(\asqrt[63] ), .ZN(new_n1530_));
  NAND2_X1   g01338(.A1(new_n1528_), .A2(new_n1502_), .ZN(new_n1531_));
  NOR2_X1    g01339(.A1(new_n1531_), .A2(new_n1518_), .ZN(new_n1532_));
  NOR4_X1    g01340(.A1(new_n1530_), .A2(new_n1371_), .A3(new_n1532_), .A4(new_n1514_), .ZN(new_n1533_));
  NOR3_X1    g01341(.A1(new_n1533_), .A2(\a[96] ), .A3(\a[97] ), .ZN(new_n1534_));
  NOR2_X1    g01342(.A1(new_n1517_), .A2(new_n1534_), .ZN(new_n1535_));
  INV_X1     g01343(.I(\a[94] ), .ZN(new_n1536_));
  INV_X1     g01344(.I(\a[95] ), .ZN(new_n1537_));
  NAND3_X1   g01345(.A1(new_n1536_), .A2(new_n1537_), .A3(new_n197_), .ZN(new_n1538_));
  NAND2_X1   g01346(.A1(\asqrt[48] ), .A2(\a[96] ), .ZN(new_n1539_));
  AOI21_X1   g01347(.A1(new_n1539_), .A2(new_n1538_), .B(new_n1368_), .ZN(new_n1540_));
  OAI21_X1   g01348(.A1(new_n1533_), .A2(new_n197_), .B(new_n1538_), .ZN(new_n1541_));
  NOR2_X1    g01349(.A1(new_n1541_), .A2(\asqrt[49] ), .ZN(new_n1542_));
  NAND2_X1   g01350(.A1(new_n1531_), .A2(new_n1380_), .ZN(new_n1543_));
  NOR2_X1    g01351(.A1(new_n1533_), .A2(new_n1380_), .ZN(new_n1544_));
  NAND2_X1   g01352(.A1(new_n1544_), .A2(new_n1512_), .ZN(new_n1545_));
  AOI21_X1   g01353(.A1(new_n1545_), .A2(new_n1543_), .B(new_n193_), .ZN(new_n1546_));
  NAND3_X1   g01354(.A1(\asqrt[48] ), .A2(new_n1502_), .A3(new_n1527_), .ZN(new_n1547_));
  XOR2_X1    g01355(.A1(new_n1547_), .A2(new_n1507_), .Z(new_n1548_));
  INV_X1     g01356(.I(new_n1548_), .ZN(new_n1549_));
  AOI21_X1   g01357(.A1(new_n1544_), .A2(new_n1531_), .B(new_n1532_), .ZN(new_n1550_));
  INV_X1     g01358(.I(new_n1550_), .ZN(new_n1551_));
  OAI21_X1   g01359(.A1(new_n1472_), .A2(new_n1474_), .B(new_n1477_), .ZN(new_n1552_));
  NOR2_X1    g01360(.A1(new_n1533_), .A2(new_n1552_), .ZN(new_n1553_));
  XOR2_X1    g01361(.A1(new_n1553_), .A2(new_n1386_), .Z(new_n1554_));
  NAND3_X1   g01362(.A1(\asqrt[48] ), .A2(new_n1488_), .A3(new_n1473_), .ZN(new_n1555_));
  XOR2_X1    g01363(.A1(new_n1555_), .A2(new_n1390_), .Z(new_n1556_));
  OAI21_X1   g01364(.A1(new_n1483_), .A2(new_n1484_), .B(new_n1487_), .ZN(new_n1557_));
  NOR2_X1    g01365(.A1(new_n1533_), .A2(new_n1557_), .ZN(new_n1558_));
  XOR2_X1    g01366(.A1(new_n1558_), .A2(new_n1392_), .Z(new_n1559_));
  INV_X1     g01367(.I(new_n1559_), .ZN(new_n1560_));
  NAND3_X1   g01368(.A1(\asqrt[48] ), .A2(new_n1450_), .A3(new_n1469_), .ZN(new_n1561_));
  XOR2_X1    g01369(.A1(new_n1561_), .A2(new_n1481_), .Z(new_n1562_));
  INV_X1     g01370(.I(new_n1562_), .ZN(new_n1563_));
  OAI21_X1   g01371(.A1(new_n1444_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n1564_));
  NOR2_X1    g01372(.A1(new_n1533_), .A2(new_n1564_), .ZN(new_n1565_));
  XOR2_X1    g01373(.A1(new_n1565_), .A2(new_n1399_), .Z(new_n1566_));
  NAND3_X1   g01374(.A1(\asqrt[48] ), .A2(new_n1463_), .A3(new_n1445_), .ZN(new_n1567_));
  XOR2_X1    g01375(.A1(new_n1567_), .A2(new_n1402_), .Z(new_n1568_));
  OAI21_X1   g01376(.A1(new_n1458_), .A2(new_n1459_), .B(new_n1462_), .ZN(new_n1569_));
  NOR2_X1    g01377(.A1(new_n1533_), .A2(new_n1569_), .ZN(new_n1570_));
  XOR2_X1    g01378(.A1(new_n1570_), .A2(new_n1405_), .Z(new_n1571_));
  INV_X1     g01379(.I(new_n1571_), .ZN(new_n1572_));
  NAND3_X1   g01380(.A1(\asqrt[48] ), .A2(new_n1423_), .A3(new_n1441_), .ZN(new_n1573_));
  XOR2_X1    g01381(.A1(new_n1573_), .A2(new_n1457_), .Z(new_n1574_));
  INV_X1     g01382(.I(new_n1574_), .ZN(new_n1575_));
  NAND2_X1   g01383(.A1(new_n1438_), .A2(new_n1088_), .ZN(new_n1576_));
  NAND3_X1   g01384(.A1(\asqrt[48] ), .A2(new_n1576_), .A3(new_n1422_), .ZN(new_n1577_));
  XOR2_X1    g01385(.A1(new_n1577_), .A2(new_n1432_), .Z(new_n1578_));
  NOR4_X1    g01386(.A1(new_n1530_), .A2(new_n1368_), .A3(new_n1371_), .A4(new_n1532_), .ZN(new_n1579_));
  OAI21_X1   g01387(.A1(new_n1534_), .A2(new_n1579_), .B(new_n1257_), .ZN(new_n1580_));
  NAND3_X1   g01388(.A1(\asqrt[48] ), .A2(new_n197_), .A3(new_n198_), .ZN(new_n1581_));
  INV_X1     g01389(.I(new_n1579_), .ZN(new_n1582_));
  NAND3_X1   g01390(.A1(new_n1581_), .A2(\a[98] ), .A3(new_n1582_), .ZN(new_n1583_));
  NAND2_X1   g01391(.A1(new_n1580_), .A2(new_n1583_), .ZN(new_n1584_));
  NAND3_X1   g01392(.A1(new_n1539_), .A2(new_n1368_), .A3(new_n1538_), .ZN(new_n1585_));
  AOI21_X1   g01393(.A1(new_n1535_), .A2(new_n1585_), .B(new_n1540_), .ZN(new_n1586_));
  AOI21_X1   g01394(.A1(new_n1586_), .A2(new_n1228_), .B(new_n1584_), .ZN(new_n1587_));
  NOR2_X1    g01395(.A1(new_n1586_), .A2(new_n1228_), .ZN(new_n1588_));
  NOR3_X1    g01396(.A1(new_n1587_), .A2(\asqrt[51] ), .A3(new_n1588_), .ZN(new_n1589_));
  NOR3_X1    g01397(.A1(new_n1533_), .A2(new_n1434_), .A3(new_n1419_), .ZN(new_n1590_));
  XOR2_X1    g01398(.A1(new_n1590_), .A2(new_n1436_), .Z(new_n1591_));
  INV_X1     g01399(.I(new_n1591_), .ZN(new_n1592_));
  OAI21_X1   g01400(.A1(new_n1587_), .A2(new_n1588_), .B(\asqrt[51] ), .ZN(new_n1593_));
  OAI21_X1   g01401(.A1(new_n1589_), .A2(new_n1592_), .B(new_n1593_), .ZN(new_n1594_));
  OAI21_X1   g01402(.A1(new_n1594_), .A2(\asqrt[52] ), .B(new_n1578_), .ZN(new_n1595_));
  AOI21_X1   g01403(.A1(new_n1594_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n1596_));
  AOI21_X1   g01404(.A1(new_n1596_), .A2(new_n1595_), .B(new_n1575_), .ZN(new_n1597_));
  NAND2_X1   g01405(.A1(new_n1594_), .A2(\asqrt[52] ), .ZN(new_n1598_));
  AOI21_X1   g01406(.A1(new_n1595_), .A2(new_n1598_), .B(new_n842_), .ZN(new_n1599_));
  NOR2_X1    g01407(.A1(new_n1597_), .A2(new_n1599_), .ZN(new_n1600_));
  AOI21_X1   g01408(.A1(new_n1600_), .A2(new_n720_), .B(new_n1572_), .ZN(new_n1601_));
  OAI21_X1   g01409(.A1(new_n1597_), .A2(new_n1599_), .B(\asqrt[54] ), .ZN(new_n1602_));
  NAND2_X1   g01410(.A1(new_n1602_), .A2(new_n630_), .ZN(new_n1603_));
  OAI21_X1   g01411(.A1(new_n1601_), .A2(new_n1603_), .B(new_n1568_), .ZN(new_n1604_));
  INV_X1     g01412(.I(new_n1602_), .ZN(new_n1605_));
  OAI21_X1   g01413(.A1(new_n1601_), .A2(new_n1605_), .B(\asqrt[55] ), .ZN(new_n1606_));
  NAND3_X1   g01414(.A1(new_n1604_), .A2(new_n1606_), .A3(new_n545_), .ZN(new_n1607_));
  NAND2_X1   g01415(.A1(new_n1607_), .A2(new_n1566_), .ZN(new_n1608_));
  NAND2_X1   g01416(.A1(new_n1604_), .A2(new_n1606_), .ZN(new_n1609_));
  AOI21_X1   g01417(.A1(new_n1609_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1610_));
  AOI21_X1   g01418(.A1(new_n1610_), .A2(new_n1608_), .B(new_n1563_), .ZN(new_n1611_));
  INV_X1     g01419(.I(new_n1568_), .ZN(new_n1612_));
  INV_X1     g01420(.I(new_n1578_), .ZN(new_n1613_));
  AOI21_X1   g01421(.A1(new_n1581_), .A2(new_n1582_), .B(\a[98] ), .ZN(new_n1614_));
  NOR3_X1    g01422(.A1(new_n1534_), .A2(new_n1257_), .A3(new_n1579_), .ZN(new_n1615_));
  NOR2_X1    g01423(.A1(new_n1615_), .A2(new_n1614_), .ZN(new_n1616_));
  OAI21_X1   g01424(.A1(new_n1533_), .A2(\a[96] ), .B(\a[97] ), .ZN(new_n1617_));
  NAND2_X1   g01425(.A1(new_n1617_), .A2(new_n1581_), .ZN(new_n1618_));
  NAND2_X1   g01426(.A1(new_n1541_), .A2(\asqrt[49] ), .ZN(new_n1619_));
  OAI21_X1   g01427(.A1(new_n1618_), .A2(new_n1542_), .B(new_n1619_), .ZN(new_n1620_));
  OAI21_X1   g01428(.A1(\asqrt[50] ), .A2(new_n1620_), .B(new_n1616_), .ZN(new_n1621_));
  NAND2_X1   g01429(.A1(new_n1620_), .A2(\asqrt[50] ), .ZN(new_n1622_));
  NAND3_X1   g01430(.A1(new_n1621_), .A2(new_n1088_), .A3(new_n1622_), .ZN(new_n1623_));
  AOI21_X1   g01431(.A1(new_n1621_), .A2(new_n1622_), .B(new_n1088_), .ZN(new_n1624_));
  AOI21_X1   g01432(.A1(new_n1623_), .A2(new_n1591_), .B(new_n1624_), .ZN(new_n1625_));
  AOI21_X1   g01433(.A1(new_n1625_), .A2(new_n962_), .B(new_n1613_), .ZN(new_n1626_));
  OAI21_X1   g01434(.A1(new_n1625_), .A2(new_n962_), .B(new_n842_), .ZN(new_n1627_));
  OAI21_X1   g01435(.A1(new_n1626_), .A2(new_n1627_), .B(new_n1574_), .ZN(new_n1628_));
  NOR2_X1    g01436(.A1(new_n1625_), .A2(new_n962_), .ZN(new_n1629_));
  OAI21_X1   g01437(.A1(new_n1626_), .A2(new_n1629_), .B(\asqrt[53] ), .ZN(new_n1630_));
  NAND3_X1   g01438(.A1(new_n1628_), .A2(new_n1630_), .A3(new_n720_), .ZN(new_n1631_));
  NAND2_X1   g01439(.A1(new_n1631_), .A2(new_n1571_), .ZN(new_n1632_));
  NAND2_X1   g01440(.A1(new_n1628_), .A2(new_n1630_), .ZN(new_n1633_));
  AOI21_X1   g01441(.A1(new_n1633_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1634_));
  AOI21_X1   g01442(.A1(new_n1634_), .A2(new_n1632_), .B(new_n1612_), .ZN(new_n1635_));
  AOI21_X1   g01443(.A1(new_n1632_), .A2(new_n1602_), .B(new_n630_), .ZN(new_n1636_));
  OAI21_X1   g01444(.A1(new_n1635_), .A2(new_n1636_), .B(\asqrt[56] ), .ZN(new_n1637_));
  AOI21_X1   g01445(.A1(new_n1608_), .A2(new_n1637_), .B(new_n450_), .ZN(new_n1638_));
  NOR2_X1    g01446(.A1(new_n1611_), .A2(new_n1638_), .ZN(new_n1639_));
  AOI21_X1   g01447(.A1(new_n1639_), .A2(new_n403_), .B(new_n1560_), .ZN(new_n1640_));
  OAI21_X1   g01448(.A1(new_n1611_), .A2(new_n1638_), .B(\asqrt[58] ), .ZN(new_n1641_));
  NAND2_X1   g01449(.A1(new_n1641_), .A2(new_n339_), .ZN(new_n1642_));
  OAI21_X1   g01450(.A1(new_n1640_), .A2(new_n1642_), .B(new_n1556_), .ZN(new_n1643_));
  INV_X1     g01451(.I(new_n1641_), .ZN(new_n1644_));
  OAI21_X1   g01452(.A1(new_n1640_), .A2(new_n1644_), .B(\asqrt[59] ), .ZN(new_n1645_));
  NAND3_X1   g01453(.A1(new_n1643_), .A2(new_n1645_), .A3(new_n288_), .ZN(new_n1646_));
  NAND2_X1   g01454(.A1(new_n1646_), .A2(new_n1554_), .ZN(new_n1647_));
  INV_X1     g01455(.I(new_n1556_), .ZN(new_n1648_));
  INV_X1     g01456(.I(new_n1566_), .ZN(new_n1649_));
  NOR2_X1    g01457(.A1(new_n1635_), .A2(new_n1636_), .ZN(new_n1650_));
  AOI21_X1   g01458(.A1(new_n1650_), .A2(new_n545_), .B(new_n1649_), .ZN(new_n1651_));
  NAND2_X1   g01459(.A1(new_n1637_), .A2(new_n450_), .ZN(new_n1652_));
  OAI21_X1   g01460(.A1(new_n1651_), .A2(new_n1652_), .B(new_n1562_), .ZN(new_n1653_));
  INV_X1     g01461(.I(new_n1637_), .ZN(new_n1654_));
  OAI21_X1   g01462(.A1(new_n1651_), .A2(new_n1654_), .B(\asqrt[57] ), .ZN(new_n1655_));
  NAND3_X1   g01463(.A1(new_n1653_), .A2(new_n1655_), .A3(new_n403_), .ZN(new_n1656_));
  NAND2_X1   g01464(.A1(new_n1656_), .A2(new_n1559_), .ZN(new_n1657_));
  NAND2_X1   g01465(.A1(new_n1653_), .A2(new_n1655_), .ZN(new_n1658_));
  AOI21_X1   g01466(.A1(new_n1658_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1659_));
  AOI21_X1   g01467(.A1(new_n1659_), .A2(new_n1657_), .B(new_n1648_), .ZN(new_n1660_));
  AOI21_X1   g01468(.A1(new_n1657_), .A2(new_n1641_), .B(new_n339_), .ZN(new_n1661_));
  OAI21_X1   g01469(.A1(new_n1660_), .A2(new_n1661_), .B(\asqrt[60] ), .ZN(new_n1662_));
  AOI21_X1   g01470(.A1(new_n1647_), .A2(new_n1662_), .B(new_n242_), .ZN(new_n1663_));
  NAND3_X1   g01471(.A1(\asqrt[48] ), .A2(new_n1478_), .A3(new_n1494_), .ZN(new_n1664_));
  XOR2_X1    g01472(.A1(new_n1664_), .A2(new_n1520_), .Z(new_n1665_));
  INV_X1     g01473(.I(new_n1665_), .ZN(new_n1666_));
  NAND2_X1   g01474(.A1(new_n1643_), .A2(new_n1645_), .ZN(new_n1667_));
  AOI21_X1   g01475(.A1(new_n1667_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1668_));
  AOI21_X1   g01476(.A1(new_n1668_), .A2(new_n1647_), .B(new_n1666_), .ZN(new_n1669_));
  OAI21_X1   g01477(.A1(new_n1669_), .A2(new_n1663_), .B(\asqrt[62] ), .ZN(new_n1670_));
  AOI21_X1   g01478(.A1(new_n1479_), .A2(new_n1500_), .B(new_n1495_), .ZN(new_n1671_));
  NAND2_X1   g01479(.A1(\asqrt[48] ), .A2(new_n1671_), .ZN(new_n1672_));
  XOR2_X1    g01480(.A1(new_n1672_), .A2(new_n1498_), .Z(new_n1673_));
  INV_X1     g01481(.I(new_n1554_), .ZN(new_n1674_));
  NOR2_X1    g01482(.A1(new_n1660_), .A2(new_n1661_), .ZN(new_n1675_));
  AOI21_X1   g01483(.A1(new_n1675_), .A2(new_n288_), .B(new_n1674_), .ZN(new_n1676_));
  INV_X1     g01484(.I(new_n1662_), .ZN(new_n1677_));
  OAI21_X1   g01485(.A1(new_n1676_), .A2(new_n1677_), .B(\asqrt[61] ), .ZN(new_n1678_));
  NAND2_X1   g01486(.A1(new_n1662_), .A2(new_n242_), .ZN(new_n1679_));
  OAI21_X1   g01487(.A1(new_n1676_), .A2(new_n1679_), .B(new_n1665_), .ZN(new_n1680_));
  NAND3_X1   g01488(.A1(new_n1680_), .A2(new_n1678_), .A3(new_n234_), .ZN(new_n1681_));
  NAND2_X1   g01489(.A1(new_n1681_), .A2(new_n1673_), .ZN(new_n1682_));
  AOI21_X1   g01490(.A1(new_n1682_), .A2(new_n1670_), .B(new_n1551_), .ZN(new_n1683_));
  AOI21_X1   g01491(.A1(new_n1683_), .A2(new_n1549_), .B(\asqrt[63] ), .ZN(new_n1684_));
  NAND2_X1   g01492(.A1(new_n1682_), .A2(new_n1670_), .ZN(new_n1685_));
  NOR2_X1    g01493(.A1(new_n1685_), .A2(new_n1549_), .ZN(new_n1686_));
  NOR2_X1    g01494(.A1(\asqrt[48] ), .A2(new_n1518_), .ZN(new_n1687_));
  NOR4_X1    g01495(.A1(new_n1684_), .A2(new_n1546_), .A3(new_n1686_), .A4(new_n1687_), .ZN(new_n1688_));
  NOR3_X1    g01496(.A1(new_n1688_), .A2(new_n1540_), .A3(new_n1542_), .ZN(new_n1689_));
  XOR2_X1    g01497(.A1(new_n1689_), .A2(new_n1535_), .Z(new_n1690_));
  INV_X1     g01498(.I(new_n1690_), .ZN(new_n1691_));
  INV_X1     g01499(.I(new_n1546_), .ZN(new_n1692_));
  INV_X1     g01500(.I(new_n1670_), .ZN(new_n1693_));
  NOR2_X1    g01501(.A1(new_n1669_), .A2(new_n1663_), .ZN(new_n1694_));
  INV_X1     g01502(.I(new_n1673_), .ZN(new_n1695_));
  AOI21_X1   g01503(.A1(new_n1694_), .A2(new_n234_), .B(new_n1695_), .ZN(new_n1696_));
  OAI21_X1   g01504(.A1(new_n1696_), .A2(new_n1693_), .B(new_n1550_), .ZN(new_n1697_));
  OAI21_X1   g01505(.A1(new_n1697_), .A2(new_n1548_), .B(new_n193_), .ZN(new_n1698_));
  NOR2_X1    g01506(.A1(new_n1696_), .A2(new_n1693_), .ZN(new_n1699_));
  NAND2_X1   g01507(.A1(new_n1699_), .A2(new_n1548_), .ZN(new_n1700_));
  INV_X1     g01508(.I(new_n1687_), .ZN(new_n1701_));
  NAND4_X1   g01509(.A1(new_n1698_), .A2(new_n1692_), .A3(new_n1700_), .A4(new_n1701_), .ZN(\asqrt[47] ));
  NAND3_X1   g01510(.A1(\asqrt[47] ), .A2(new_n1536_), .A3(new_n1537_), .ZN(new_n1703_));
  NAND4_X1   g01511(.A1(new_n1698_), .A2(\asqrt[48] ), .A3(new_n1700_), .A4(new_n1692_), .ZN(new_n1704_));
  AOI21_X1   g01512(.A1(new_n1703_), .A2(new_n1704_), .B(\a[96] ), .ZN(new_n1705_));
  NOR3_X1    g01513(.A1(new_n1688_), .A2(\a[94] ), .A3(\a[95] ), .ZN(new_n1706_));
  INV_X1     g01514(.I(new_n1704_), .ZN(new_n1707_));
  NOR3_X1    g01515(.A1(new_n1706_), .A2(new_n197_), .A3(new_n1707_), .ZN(new_n1708_));
  NOR2_X1    g01516(.A1(new_n1708_), .A2(new_n1705_), .ZN(new_n1709_));
  INV_X1     g01517(.I(\a[92] ), .ZN(new_n1710_));
  INV_X1     g01518(.I(\a[93] ), .ZN(new_n1711_));
  NAND3_X1   g01519(.A1(new_n1710_), .A2(new_n1711_), .A3(new_n1536_), .ZN(new_n1712_));
  OAI21_X1   g01520(.A1(new_n1688_), .A2(new_n1536_), .B(new_n1712_), .ZN(new_n1713_));
  NAND2_X1   g01521(.A1(new_n1713_), .A2(\asqrt[48] ), .ZN(new_n1714_));
  OAI21_X1   g01522(.A1(new_n1688_), .A2(\a[94] ), .B(\a[95] ), .ZN(new_n1715_));
  NAND2_X1   g01523(.A1(new_n1715_), .A2(new_n1703_), .ZN(new_n1716_));
  NOR2_X1    g01524(.A1(new_n1713_), .A2(\asqrt[48] ), .ZN(new_n1717_));
  OAI21_X1   g01525(.A1(new_n1716_), .A2(new_n1717_), .B(new_n1714_), .ZN(new_n1718_));
  OAI21_X1   g01526(.A1(new_n1718_), .A2(\asqrt[49] ), .B(new_n1709_), .ZN(new_n1719_));
  NAND2_X1   g01527(.A1(new_n1718_), .A2(\asqrt[49] ), .ZN(new_n1720_));
  NAND3_X1   g01528(.A1(new_n1719_), .A2(new_n1228_), .A3(new_n1720_), .ZN(new_n1721_));
  OAI21_X1   g01529(.A1(new_n1706_), .A2(new_n1707_), .B(new_n197_), .ZN(new_n1722_));
  NAND3_X1   g01530(.A1(new_n1703_), .A2(\a[96] ), .A3(new_n1704_), .ZN(new_n1723_));
  NAND2_X1   g01531(.A1(new_n1722_), .A2(new_n1723_), .ZN(new_n1724_));
  NAND2_X1   g01532(.A1(\asqrt[47] ), .A2(\a[94] ), .ZN(new_n1725_));
  AOI21_X1   g01533(.A1(new_n1725_), .A2(new_n1712_), .B(new_n1533_), .ZN(new_n1726_));
  AOI21_X1   g01534(.A1(\asqrt[47] ), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n1727_));
  NOR2_X1    g01535(.A1(new_n1706_), .A2(new_n1727_), .ZN(new_n1728_));
  NAND3_X1   g01536(.A1(new_n1725_), .A2(new_n1533_), .A3(new_n1712_), .ZN(new_n1729_));
  AOI21_X1   g01537(.A1(new_n1728_), .A2(new_n1729_), .B(new_n1726_), .ZN(new_n1730_));
  AOI21_X1   g01538(.A1(new_n1730_), .A2(new_n1368_), .B(new_n1724_), .ZN(new_n1731_));
  NOR2_X1    g01539(.A1(new_n1730_), .A2(new_n1368_), .ZN(new_n1732_));
  OAI21_X1   g01540(.A1(new_n1731_), .A2(new_n1732_), .B(\asqrt[50] ), .ZN(new_n1733_));
  NAND2_X1   g01541(.A1(new_n1685_), .A2(new_n1548_), .ZN(new_n1734_));
  NOR2_X1    g01542(.A1(new_n1688_), .A2(new_n1548_), .ZN(new_n1735_));
  NAND2_X1   g01543(.A1(new_n1735_), .A2(new_n1699_), .ZN(new_n1736_));
  AOI21_X1   g01544(.A1(new_n1736_), .A2(new_n1734_), .B(new_n193_), .ZN(new_n1737_));
  INV_X1     g01545(.I(new_n1737_), .ZN(new_n1738_));
  NAND3_X1   g01546(.A1(\asqrt[47] ), .A2(new_n1670_), .A3(new_n1681_), .ZN(new_n1739_));
  XOR2_X1    g01547(.A1(new_n1739_), .A2(new_n1673_), .Z(new_n1740_));
  AOI21_X1   g01548(.A1(new_n1735_), .A2(new_n1685_), .B(new_n1686_), .ZN(new_n1741_));
  OAI21_X1   g01549(.A1(new_n1640_), .A2(new_n1642_), .B(new_n1645_), .ZN(new_n1742_));
  NOR2_X1    g01550(.A1(new_n1688_), .A2(new_n1742_), .ZN(new_n1743_));
  XOR2_X1    g01551(.A1(new_n1743_), .A2(new_n1556_), .Z(new_n1744_));
  NAND3_X1   g01552(.A1(\asqrt[47] ), .A2(new_n1656_), .A3(new_n1641_), .ZN(new_n1745_));
  XOR2_X1    g01553(.A1(new_n1745_), .A2(new_n1560_), .Z(new_n1746_));
  OAI21_X1   g01554(.A1(new_n1651_), .A2(new_n1652_), .B(new_n1655_), .ZN(new_n1747_));
  NOR2_X1    g01555(.A1(new_n1688_), .A2(new_n1747_), .ZN(new_n1748_));
  XOR2_X1    g01556(.A1(new_n1748_), .A2(new_n1562_), .Z(new_n1749_));
  INV_X1     g01557(.I(new_n1749_), .ZN(new_n1750_));
  NAND3_X1   g01558(.A1(\asqrt[47] ), .A2(new_n1607_), .A3(new_n1637_), .ZN(new_n1751_));
  XOR2_X1    g01559(.A1(new_n1751_), .A2(new_n1649_), .Z(new_n1752_));
  INV_X1     g01560(.I(new_n1752_), .ZN(new_n1753_));
  OAI21_X1   g01561(.A1(new_n1601_), .A2(new_n1603_), .B(new_n1606_), .ZN(new_n1754_));
  NOR2_X1    g01562(.A1(new_n1688_), .A2(new_n1754_), .ZN(new_n1755_));
  XOR2_X1    g01563(.A1(new_n1755_), .A2(new_n1568_), .Z(new_n1756_));
  NAND3_X1   g01564(.A1(\asqrt[47] ), .A2(new_n1631_), .A3(new_n1602_), .ZN(new_n1757_));
  XOR2_X1    g01565(.A1(new_n1757_), .A2(new_n1572_), .Z(new_n1758_));
  AOI21_X1   g01566(.A1(new_n1595_), .A2(new_n1596_), .B(new_n1599_), .ZN(new_n1759_));
  NAND2_X1   g01567(.A1(\asqrt[47] ), .A2(new_n1759_), .ZN(new_n1760_));
  XOR2_X1    g01568(.A1(new_n1760_), .A2(new_n1575_), .Z(new_n1761_));
  INV_X1     g01569(.I(new_n1761_), .ZN(new_n1762_));
  NOR2_X1    g01570(.A1(new_n1594_), .A2(\asqrt[52] ), .ZN(new_n1763_));
  NOR3_X1    g01571(.A1(new_n1688_), .A2(new_n1763_), .A3(new_n1629_), .ZN(new_n1764_));
  XOR2_X1    g01572(.A1(new_n1764_), .A2(new_n1578_), .Z(new_n1765_));
  INV_X1     g01573(.I(new_n1765_), .ZN(new_n1766_));
  NOR3_X1    g01574(.A1(new_n1688_), .A2(new_n1589_), .A3(new_n1624_), .ZN(new_n1767_));
  XOR2_X1    g01575(.A1(new_n1767_), .A2(new_n1591_), .Z(new_n1768_));
  NOR2_X1    g01576(.A1(new_n1620_), .A2(\asqrt[50] ), .ZN(new_n1769_));
  NOR3_X1    g01577(.A1(new_n1688_), .A2(new_n1769_), .A3(new_n1588_), .ZN(new_n1770_));
  XOR2_X1    g01578(.A1(new_n1770_), .A2(new_n1616_), .Z(new_n1771_));
  NOR2_X1    g01579(.A1(new_n1731_), .A2(new_n1732_), .ZN(new_n1772_));
  AOI21_X1   g01580(.A1(new_n1772_), .A2(new_n1228_), .B(new_n1691_), .ZN(new_n1773_));
  NAND2_X1   g01581(.A1(new_n1733_), .A2(new_n1088_), .ZN(new_n1774_));
  OAI21_X1   g01582(.A1(new_n1773_), .A2(new_n1774_), .B(new_n1771_), .ZN(new_n1775_));
  INV_X1     g01583(.I(new_n1733_), .ZN(new_n1776_));
  OAI21_X1   g01584(.A1(new_n1773_), .A2(new_n1776_), .B(\asqrt[51] ), .ZN(new_n1777_));
  NAND3_X1   g01585(.A1(new_n1775_), .A2(new_n1777_), .A3(new_n962_), .ZN(new_n1778_));
  NAND2_X1   g01586(.A1(new_n1778_), .A2(new_n1768_), .ZN(new_n1779_));
  NAND2_X1   g01587(.A1(new_n1775_), .A2(new_n1777_), .ZN(new_n1780_));
  AOI21_X1   g01588(.A1(new_n1780_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n1781_));
  AOI21_X1   g01589(.A1(new_n1781_), .A2(new_n1779_), .B(new_n1766_), .ZN(new_n1782_));
  INV_X1     g01590(.I(new_n1771_), .ZN(new_n1783_));
  NAND2_X1   g01591(.A1(new_n1721_), .A2(new_n1690_), .ZN(new_n1784_));
  NAND2_X1   g01592(.A1(new_n1719_), .A2(new_n1720_), .ZN(new_n1785_));
  AOI21_X1   g01593(.A1(new_n1785_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n1786_));
  AOI21_X1   g01594(.A1(new_n1786_), .A2(new_n1784_), .B(new_n1783_), .ZN(new_n1787_));
  AOI21_X1   g01595(.A1(new_n1784_), .A2(new_n1733_), .B(new_n1088_), .ZN(new_n1788_));
  OAI21_X1   g01596(.A1(new_n1787_), .A2(new_n1788_), .B(\asqrt[52] ), .ZN(new_n1789_));
  AOI21_X1   g01597(.A1(new_n1779_), .A2(new_n1789_), .B(new_n842_), .ZN(new_n1790_));
  NOR2_X1    g01598(.A1(new_n1782_), .A2(new_n1790_), .ZN(new_n1791_));
  AOI21_X1   g01599(.A1(new_n1791_), .A2(new_n720_), .B(new_n1762_), .ZN(new_n1792_));
  OAI21_X1   g01600(.A1(new_n1782_), .A2(new_n1790_), .B(\asqrt[54] ), .ZN(new_n1793_));
  NAND2_X1   g01601(.A1(new_n1793_), .A2(new_n630_), .ZN(new_n1794_));
  OAI21_X1   g01602(.A1(new_n1792_), .A2(new_n1794_), .B(new_n1758_), .ZN(new_n1795_));
  INV_X1     g01603(.I(new_n1793_), .ZN(new_n1796_));
  OAI21_X1   g01604(.A1(new_n1792_), .A2(new_n1796_), .B(\asqrt[55] ), .ZN(new_n1797_));
  NAND3_X1   g01605(.A1(new_n1795_), .A2(new_n1797_), .A3(new_n545_), .ZN(new_n1798_));
  NAND2_X1   g01606(.A1(new_n1798_), .A2(new_n1756_), .ZN(new_n1799_));
  NAND2_X1   g01607(.A1(new_n1795_), .A2(new_n1797_), .ZN(new_n1800_));
  AOI21_X1   g01608(.A1(new_n1800_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1801_));
  AOI21_X1   g01609(.A1(new_n1801_), .A2(new_n1799_), .B(new_n1753_), .ZN(new_n1802_));
  INV_X1     g01610(.I(new_n1758_), .ZN(new_n1803_));
  INV_X1     g01611(.I(new_n1768_), .ZN(new_n1804_));
  NOR2_X1    g01612(.A1(new_n1787_), .A2(new_n1788_), .ZN(new_n1805_));
  AOI21_X1   g01613(.A1(new_n1805_), .A2(new_n962_), .B(new_n1804_), .ZN(new_n1806_));
  NAND2_X1   g01614(.A1(new_n1789_), .A2(new_n842_), .ZN(new_n1807_));
  OAI21_X1   g01615(.A1(new_n1806_), .A2(new_n1807_), .B(new_n1765_), .ZN(new_n1808_));
  INV_X1     g01616(.I(new_n1789_), .ZN(new_n1809_));
  OAI21_X1   g01617(.A1(new_n1806_), .A2(new_n1809_), .B(\asqrt[53] ), .ZN(new_n1810_));
  NAND3_X1   g01618(.A1(new_n1808_), .A2(new_n1810_), .A3(new_n720_), .ZN(new_n1811_));
  NAND2_X1   g01619(.A1(new_n1811_), .A2(new_n1761_), .ZN(new_n1812_));
  NAND2_X1   g01620(.A1(new_n1808_), .A2(new_n1810_), .ZN(new_n1813_));
  AOI21_X1   g01621(.A1(new_n1813_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1814_));
  AOI21_X1   g01622(.A1(new_n1814_), .A2(new_n1812_), .B(new_n1803_), .ZN(new_n1815_));
  AOI21_X1   g01623(.A1(new_n1812_), .A2(new_n1793_), .B(new_n630_), .ZN(new_n1816_));
  OAI21_X1   g01624(.A1(new_n1815_), .A2(new_n1816_), .B(\asqrt[56] ), .ZN(new_n1817_));
  AOI21_X1   g01625(.A1(new_n1799_), .A2(new_n1817_), .B(new_n450_), .ZN(new_n1818_));
  NOR2_X1    g01626(.A1(new_n1802_), .A2(new_n1818_), .ZN(new_n1819_));
  AOI21_X1   g01627(.A1(new_n1819_), .A2(new_n403_), .B(new_n1750_), .ZN(new_n1820_));
  OAI21_X1   g01628(.A1(new_n1802_), .A2(new_n1818_), .B(\asqrt[58] ), .ZN(new_n1821_));
  NAND2_X1   g01629(.A1(new_n1821_), .A2(new_n339_), .ZN(new_n1822_));
  OAI21_X1   g01630(.A1(new_n1820_), .A2(new_n1822_), .B(new_n1746_), .ZN(new_n1823_));
  INV_X1     g01631(.I(new_n1821_), .ZN(new_n1824_));
  OAI21_X1   g01632(.A1(new_n1820_), .A2(new_n1824_), .B(\asqrt[59] ), .ZN(new_n1825_));
  NAND3_X1   g01633(.A1(new_n1823_), .A2(new_n1825_), .A3(new_n288_), .ZN(new_n1826_));
  NAND2_X1   g01634(.A1(new_n1826_), .A2(new_n1744_), .ZN(new_n1827_));
  INV_X1     g01635(.I(new_n1746_), .ZN(new_n1828_));
  INV_X1     g01636(.I(new_n1756_), .ZN(new_n1829_));
  NOR2_X1    g01637(.A1(new_n1815_), .A2(new_n1816_), .ZN(new_n1830_));
  AOI21_X1   g01638(.A1(new_n1830_), .A2(new_n545_), .B(new_n1829_), .ZN(new_n1831_));
  NAND2_X1   g01639(.A1(new_n1817_), .A2(new_n450_), .ZN(new_n1832_));
  OAI21_X1   g01640(.A1(new_n1831_), .A2(new_n1832_), .B(new_n1752_), .ZN(new_n1833_));
  INV_X1     g01641(.I(new_n1817_), .ZN(new_n1834_));
  OAI21_X1   g01642(.A1(new_n1831_), .A2(new_n1834_), .B(\asqrt[57] ), .ZN(new_n1835_));
  NAND3_X1   g01643(.A1(new_n1833_), .A2(new_n1835_), .A3(new_n403_), .ZN(new_n1836_));
  NAND2_X1   g01644(.A1(new_n1836_), .A2(new_n1749_), .ZN(new_n1837_));
  NAND2_X1   g01645(.A1(new_n1833_), .A2(new_n1835_), .ZN(new_n1838_));
  AOI21_X1   g01646(.A1(new_n1838_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1839_));
  AOI21_X1   g01647(.A1(new_n1839_), .A2(new_n1837_), .B(new_n1828_), .ZN(new_n1840_));
  AOI21_X1   g01648(.A1(new_n1837_), .A2(new_n1821_), .B(new_n339_), .ZN(new_n1841_));
  OAI21_X1   g01649(.A1(new_n1840_), .A2(new_n1841_), .B(\asqrt[60] ), .ZN(new_n1842_));
  AOI21_X1   g01650(.A1(new_n1827_), .A2(new_n1842_), .B(new_n242_), .ZN(new_n1843_));
  NAND3_X1   g01651(.A1(\asqrt[47] ), .A2(new_n1646_), .A3(new_n1662_), .ZN(new_n1844_));
  XOR2_X1    g01652(.A1(new_n1844_), .A2(new_n1674_), .Z(new_n1845_));
  INV_X1     g01653(.I(new_n1845_), .ZN(new_n1846_));
  NAND2_X1   g01654(.A1(new_n1823_), .A2(new_n1825_), .ZN(new_n1847_));
  AOI21_X1   g01655(.A1(new_n1847_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1848_));
  AOI21_X1   g01656(.A1(new_n1848_), .A2(new_n1827_), .B(new_n1846_), .ZN(new_n1849_));
  OAI21_X1   g01657(.A1(new_n1849_), .A2(new_n1843_), .B(\asqrt[62] ), .ZN(new_n1850_));
  INV_X1     g01658(.I(new_n1850_), .ZN(new_n1851_));
  NOR2_X1    g01659(.A1(new_n1849_), .A2(new_n1843_), .ZN(new_n1852_));
  AOI21_X1   g01660(.A1(new_n1647_), .A2(new_n1668_), .B(new_n1663_), .ZN(new_n1853_));
  NAND2_X1   g01661(.A1(\asqrt[47] ), .A2(new_n1853_), .ZN(new_n1854_));
  XOR2_X1    g01662(.A1(new_n1854_), .A2(new_n1666_), .Z(new_n1855_));
  INV_X1     g01663(.I(new_n1855_), .ZN(new_n1856_));
  AOI21_X1   g01664(.A1(new_n1852_), .A2(new_n234_), .B(new_n1856_), .ZN(new_n1857_));
  OAI21_X1   g01665(.A1(new_n1857_), .A2(new_n1851_), .B(new_n1741_), .ZN(new_n1858_));
  OAI21_X1   g01666(.A1(new_n1858_), .A2(new_n1740_), .B(new_n193_), .ZN(new_n1859_));
  NOR2_X1    g01667(.A1(new_n1857_), .A2(new_n1851_), .ZN(new_n1860_));
  NAND2_X1   g01668(.A1(new_n1860_), .A2(new_n1740_), .ZN(new_n1861_));
  NOR2_X1    g01669(.A1(\asqrt[47] ), .A2(new_n1549_), .ZN(new_n1862_));
  INV_X1     g01670(.I(new_n1862_), .ZN(new_n1863_));
  NAND4_X1   g01671(.A1(new_n1859_), .A2(new_n1738_), .A3(new_n1861_), .A4(new_n1863_), .ZN(\asqrt[46] ));
  NAND3_X1   g01672(.A1(\asqrt[46] ), .A2(new_n1721_), .A3(new_n1733_), .ZN(new_n1865_));
  XOR2_X1    g01673(.A1(new_n1865_), .A2(new_n1691_), .Z(new_n1866_));
  INV_X1     g01674(.I(new_n1866_), .ZN(new_n1867_));
  INV_X1     g01675(.I(new_n1744_), .ZN(new_n1868_));
  NOR2_X1    g01676(.A1(new_n1840_), .A2(new_n1841_), .ZN(new_n1869_));
  AOI21_X1   g01677(.A1(new_n1869_), .A2(new_n288_), .B(new_n1868_), .ZN(new_n1870_));
  INV_X1     g01678(.I(new_n1842_), .ZN(new_n1871_));
  OAI21_X1   g01679(.A1(new_n1870_), .A2(new_n1871_), .B(\asqrt[61] ), .ZN(new_n1872_));
  NAND2_X1   g01680(.A1(new_n1842_), .A2(new_n242_), .ZN(new_n1873_));
  OAI21_X1   g01681(.A1(new_n1870_), .A2(new_n1873_), .B(new_n1845_), .ZN(new_n1874_));
  NAND3_X1   g01682(.A1(new_n1874_), .A2(new_n1872_), .A3(new_n234_), .ZN(new_n1875_));
  NAND2_X1   g01683(.A1(new_n1875_), .A2(new_n1855_), .ZN(new_n1876_));
  NAND2_X1   g01684(.A1(new_n1876_), .A2(new_n1850_), .ZN(new_n1877_));
  NAND2_X1   g01685(.A1(new_n1877_), .A2(new_n1740_), .ZN(new_n1878_));
  INV_X1     g01686(.I(new_n1740_), .ZN(new_n1879_));
  INV_X1     g01687(.I(new_n1741_), .ZN(new_n1880_));
  AOI21_X1   g01688(.A1(new_n1876_), .A2(new_n1850_), .B(new_n1880_), .ZN(new_n1881_));
  AOI21_X1   g01689(.A1(new_n1881_), .A2(new_n1879_), .B(\asqrt[63] ), .ZN(new_n1882_));
  NOR2_X1    g01690(.A1(new_n1877_), .A2(new_n1879_), .ZN(new_n1883_));
  NOR4_X1    g01691(.A1(new_n1882_), .A2(new_n1737_), .A3(new_n1883_), .A4(new_n1862_), .ZN(new_n1884_));
  NOR2_X1    g01692(.A1(new_n1884_), .A2(new_n1740_), .ZN(new_n1885_));
  NAND2_X1   g01693(.A1(new_n1885_), .A2(new_n1860_), .ZN(new_n1886_));
  AOI21_X1   g01694(.A1(new_n1886_), .A2(new_n1878_), .B(new_n193_), .ZN(new_n1887_));
  INV_X1     g01695(.I(new_n1887_), .ZN(new_n1888_));
  NAND3_X1   g01696(.A1(\asqrt[46] ), .A2(new_n1850_), .A3(new_n1875_), .ZN(new_n1889_));
  XOR2_X1    g01697(.A1(new_n1889_), .A2(new_n1855_), .Z(new_n1890_));
  AOI21_X1   g01698(.A1(new_n1885_), .A2(new_n1877_), .B(new_n1883_), .ZN(new_n1891_));
  OAI21_X1   g01699(.A1(new_n1820_), .A2(new_n1822_), .B(new_n1825_), .ZN(new_n1892_));
  NOR2_X1    g01700(.A1(new_n1884_), .A2(new_n1892_), .ZN(new_n1893_));
  XOR2_X1    g01701(.A1(new_n1893_), .A2(new_n1746_), .Z(new_n1894_));
  NAND3_X1   g01702(.A1(\asqrt[46] ), .A2(new_n1836_), .A3(new_n1821_), .ZN(new_n1895_));
  XOR2_X1    g01703(.A1(new_n1895_), .A2(new_n1750_), .Z(new_n1896_));
  OAI21_X1   g01704(.A1(new_n1831_), .A2(new_n1832_), .B(new_n1835_), .ZN(new_n1897_));
  NOR2_X1    g01705(.A1(new_n1884_), .A2(new_n1897_), .ZN(new_n1898_));
  XOR2_X1    g01706(.A1(new_n1898_), .A2(new_n1752_), .Z(new_n1899_));
  INV_X1     g01707(.I(new_n1899_), .ZN(new_n1900_));
  NAND3_X1   g01708(.A1(\asqrt[46] ), .A2(new_n1798_), .A3(new_n1817_), .ZN(new_n1901_));
  XOR2_X1    g01709(.A1(new_n1901_), .A2(new_n1829_), .Z(new_n1902_));
  INV_X1     g01710(.I(new_n1902_), .ZN(new_n1903_));
  OAI21_X1   g01711(.A1(new_n1792_), .A2(new_n1794_), .B(new_n1797_), .ZN(new_n1904_));
  NOR2_X1    g01712(.A1(new_n1884_), .A2(new_n1904_), .ZN(new_n1905_));
  XOR2_X1    g01713(.A1(new_n1905_), .A2(new_n1758_), .Z(new_n1906_));
  NAND3_X1   g01714(.A1(\asqrt[46] ), .A2(new_n1811_), .A3(new_n1793_), .ZN(new_n1907_));
  XOR2_X1    g01715(.A1(new_n1907_), .A2(new_n1762_), .Z(new_n1908_));
  OAI21_X1   g01716(.A1(new_n1806_), .A2(new_n1807_), .B(new_n1810_), .ZN(new_n1909_));
  NOR2_X1    g01717(.A1(new_n1884_), .A2(new_n1909_), .ZN(new_n1910_));
  XOR2_X1    g01718(.A1(new_n1910_), .A2(new_n1765_), .Z(new_n1911_));
  INV_X1     g01719(.I(new_n1911_), .ZN(new_n1912_));
  NAND3_X1   g01720(.A1(\asqrt[46] ), .A2(new_n1778_), .A3(new_n1789_), .ZN(new_n1913_));
  XOR2_X1    g01721(.A1(new_n1913_), .A2(new_n1804_), .Z(new_n1914_));
  INV_X1     g01722(.I(new_n1914_), .ZN(new_n1915_));
  OAI21_X1   g01723(.A1(new_n1773_), .A2(new_n1774_), .B(new_n1777_), .ZN(new_n1916_));
  NOR2_X1    g01724(.A1(new_n1884_), .A2(new_n1916_), .ZN(new_n1917_));
  XOR2_X1    g01725(.A1(new_n1917_), .A2(new_n1771_), .Z(new_n1918_));
  NOR2_X1    g01726(.A1(new_n1718_), .A2(\asqrt[49] ), .ZN(new_n1919_));
  NOR3_X1    g01727(.A1(new_n1884_), .A2(new_n1919_), .A3(new_n1732_), .ZN(new_n1920_));
  XOR2_X1    g01728(.A1(new_n1920_), .A2(new_n1709_), .Z(new_n1921_));
  INV_X1     g01729(.I(new_n1921_), .ZN(new_n1922_));
  NAND3_X1   g01730(.A1(\asqrt[46] ), .A2(new_n1710_), .A3(new_n1711_), .ZN(new_n1923_));
  NOR4_X1    g01731(.A1(new_n1882_), .A2(new_n1688_), .A3(new_n1737_), .A4(new_n1883_), .ZN(new_n1924_));
  INV_X1     g01732(.I(new_n1924_), .ZN(new_n1925_));
  AOI21_X1   g01733(.A1(new_n1923_), .A2(new_n1925_), .B(\a[94] ), .ZN(new_n1926_));
  NOR3_X1    g01734(.A1(new_n1884_), .A2(\a[92] ), .A3(\a[93] ), .ZN(new_n1927_));
  NOR3_X1    g01735(.A1(new_n1927_), .A2(new_n1536_), .A3(new_n1924_), .ZN(new_n1928_));
  NOR2_X1    g01736(.A1(new_n1928_), .A2(new_n1926_), .ZN(new_n1929_));
  INV_X1     g01737(.I(\a[90] ), .ZN(new_n1930_));
  INV_X1     g01738(.I(\a[91] ), .ZN(new_n1931_));
  NAND3_X1   g01739(.A1(new_n1930_), .A2(new_n1931_), .A3(new_n1710_), .ZN(new_n1932_));
  OAI21_X1   g01740(.A1(new_n1884_), .A2(new_n1710_), .B(new_n1932_), .ZN(new_n1933_));
  NAND2_X1   g01741(.A1(new_n1933_), .A2(\asqrt[47] ), .ZN(new_n1934_));
  OAI21_X1   g01742(.A1(new_n1884_), .A2(\a[92] ), .B(\a[93] ), .ZN(new_n1935_));
  NAND2_X1   g01743(.A1(new_n1935_), .A2(new_n1923_), .ZN(new_n1936_));
  NOR2_X1    g01744(.A1(new_n1933_), .A2(\asqrt[47] ), .ZN(new_n1937_));
  OAI21_X1   g01745(.A1(new_n1936_), .A2(new_n1937_), .B(new_n1934_), .ZN(new_n1938_));
  OAI21_X1   g01746(.A1(new_n1938_), .A2(\asqrt[48] ), .B(new_n1929_), .ZN(new_n1939_));
  NAND2_X1   g01747(.A1(new_n1938_), .A2(\asqrt[48] ), .ZN(new_n1940_));
  NAND3_X1   g01748(.A1(new_n1939_), .A2(new_n1368_), .A3(new_n1940_), .ZN(new_n1941_));
  NOR3_X1    g01749(.A1(new_n1884_), .A2(new_n1726_), .A3(new_n1717_), .ZN(new_n1942_));
  XOR2_X1    g01750(.A1(new_n1942_), .A2(new_n1728_), .Z(new_n1943_));
  AOI21_X1   g01751(.A1(new_n1939_), .A2(new_n1940_), .B(new_n1368_), .ZN(new_n1944_));
  AOI21_X1   g01752(.A1(new_n1941_), .A2(new_n1943_), .B(new_n1944_), .ZN(new_n1945_));
  AOI21_X1   g01753(.A1(new_n1945_), .A2(new_n1228_), .B(new_n1922_), .ZN(new_n1946_));
  OAI21_X1   g01754(.A1(new_n1945_), .A2(new_n1228_), .B(new_n1088_), .ZN(new_n1947_));
  OAI21_X1   g01755(.A1(new_n1946_), .A2(new_n1947_), .B(new_n1866_), .ZN(new_n1948_));
  NOR2_X1    g01756(.A1(new_n1945_), .A2(new_n1228_), .ZN(new_n1949_));
  OAI21_X1   g01757(.A1(new_n1946_), .A2(new_n1949_), .B(\asqrt[51] ), .ZN(new_n1950_));
  NAND3_X1   g01758(.A1(new_n1948_), .A2(new_n1950_), .A3(new_n962_), .ZN(new_n1951_));
  NAND2_X1   g01759(.A1(new_n1951_), .A2(new_n1918_), .ZN(new_n1952_));
  NAND2_X1   g01760(.A1(new_n1948_), .A2(new_n1950_), .ZN(new_n1953_));
  AOI21_X1   g01761(.A1(new_n1953_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n1954_));
  AOI21_X1   g01762(.A1(new_n1954_), .A2(new_n1952_), .B(new_n1915_), .ZN(new_n1955_));
  OAI21_X1   g01763(.A1(new_n1927_), .A2(new_n1924_), .B(new_n1536_), .ZN(new_n1956_));
  NAND3_X1   g01764(.A1(new_n1923_), .A2(new_n1925_), .A3(\a[94] ), .ZN(new_n1957_));
  NAND2_X1   g01765(.A1(new_n1956_), .A2(new_n1957_), .ZN(new_n1958_));
  NAND2_X1   g01766(.A1(\asqrt[46] ), .A2(\a[92] ), .ZN(new_n1959_));
  AOI21_X1   g01767(.A1(new_n1959_), .A2(new_n1932_), .B(new_n1688_), .ZN(new_n1960_));
  AOI21_X1   g01768(.A1(\asqrt[46] ), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n1961_));
  NOR2_X1    g01769(.A1(new_n1927_), .A2(new_n1961_), .ZN(new_n1962_));
  NAND3_X1   g01770(.A1(new_n1959_), .A2(new_n1688_), .A3(new_n1932_), .ZN(new_n1963_));
  AOI21_X1   g01771(.A1(new_n1962_), .A2(new_n1963_), .B(new_n1960_), .ZN(new_n1964_));
  AOI21_X1   g01772(.A1(new_n1964_), .A2(new_n1533_), .B(new_n1958_), .ZN(new_n1965_));
  NOR2_X1    g01773(.A1(new_n1964_), .A2(new_n1533_), .ZN(new_n1966_));
  NOR3_X1    g01774(.A1(new_n1965_), .A2(\asqrt[49] ), .A3(new_n1966_), .ZN(new_n1967_));
  INV_X1     g01775(.I(new_n1943_), .ZN(new_n1968_));
  OAI21_X1   g01776(.A1(new_n1965_), .A2(new_n1966_), .B(\asqrt[49] ), .ZN(new_n1969_));
  OAI21_X1   g01777(.A1(new_n1967_), .A2(new_n1968_), .B(new_n1969_), .ZN(new_n1970_));
  OAI21_X1   g01778(.A1(new_n1970_), .A2(\asqrt[50] ), .B(new_n1921_), .ZN(new_n1971_));
  AOI21_X1   g01779(.A1(new_n1970_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n1972_));
  AOI21_X1   g01780(.A1(new_n1972_), .A2(new_n1971_), .B(new_n1867_), .ZN(new_n1973_));
  NAND2_X1   g01781(.A1(new_n1970_), .A2(\asqrt[50] ), .ZN(new_n1974_));
  AOI21_X1   g01782(.A1(new_n1971_), .A2(new_n1974_), .B(new_n1088_), .ZN(new_n1975_));
  OAI21_X1   g01783(.A1(new_n1973_), .A2(new_n1975_), .B(\asqrt[52] ), .ZN(new_n1976_));
  AOI21_X1   g01784(.A1(new_n1952_), .A2(new_n1976_), .B(new_n842_), .ZN(new_n1977_));
  NOR2_X1    g01785(.A1(new_n1955_), .A2(new_n1977_), .ZN(new_n1978_));
  AOI21_X1   g01786(.A1(new_n1978_), .A2(new_n720_), .B(new_n1912_), .ZN(new_n1979_));
  OAI21_X1   g01787(.A1(new_n1955_), .A2(new_n1977_), .B(\asqrt[54] ), .ZN(new_n1980_));
  NAND2_X1   g01788(.A1(new_n1980_), .A2(new_n630_), .ZN(new_n1981_));
  OAI21_X1   g01789(.A1(new_n1979_), .A2(new_n1981_), .B(new_n1908_), .ZN(new_n1982_));
  INV_X1     g01790(.I(new_n1980_), .ZN(new_n1983_));
  OAI21_X1   g01791(.A1(new_n1979_), .A2(new_n1983_), .B(\asqrt[55] ), .ZN(new_n1984_));
  NAND3_X1   g01792(.A1(new_n1982_), .A2(new_n1984_), .A3(new_n545_), .ZN(new_n1985_));
  NAND2_X1   g01793(.A1(new_n1985_), .A2(new_n1906_), .ZN(new_n1986_));
  NAND2_X1   g01794(.A1(new_n1982_), .A2(new_n1984_), .ZN(new_n1987_));
  AOI21_X1   g01795(.A1(new_n1987_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1988_));
  AOI21_X1   g01796(.A1(new_n1988_), .A2(new_n1986_), .B(new_n1903_), .ZN(new_n1989_));
  INV_X1     g01797(.I(new_n1908_), .ZN(new_n1990_));
  INV_X1     g01798(.I(new_n1918_), .ZN(new_n1991_));
  NOR2_X1    g01799(.A1(new_n1973_), .A2(new_n1975_), .ZN(new_n1992_));
  AOI21_X1   g01800(.A1(new_n1992_), .A2(new_n962_), .B(new_n1991_), .ZN(new_n1993_));
  NAND2_X1   g01801(.A1(new_n1976_), .A2(new_n842_), .ZN(new_n1994_));
  OAI21_X1   g01802(.A1(new_n1993_), .A2(new_n1994_), .B(new_n1914_), .ZN(new_n1995_));
  INV_X1     g01803(.I(new_n1976_), .ZN(new_n1996_));
  OAI21_X1   g01804(.A1(new_n1993_), .A2(new_n1996_), .B(\asqrt[53] ), .ZN(new_n1997_));
  NAND3_X1   g01805(.A1(new_n1995_), .A2(new_n1997_), .A3(new_n720_), .ZN(new_n1998_));
  NAND2_X1   g01806(.A1(new_n1998_), .A2(new_n1911_), .ZN(new_n1999_));
  NAND2_X1   g01807(.A1(new_n1995_), .A2(new_n1997_), .ZN(new_n2000_));
  AOI21_X1   g01808(.A1(new_n2000_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n2001_));
  AOI21_X1   g01809(.A1(new_n2001_), .A2(new_n1999_), .B(new_n1990_), .ZN(new_n2002_));
  AOI21_X1   g01810(.A1(new_n1999_), .A2(new_n1980_), .B(new_n630_), .ZN(new_n2003_));
  OAI21_X1   g01811(.A1(new_n2002_), .A2(new_n2003_), .B(\asqrt[56] ), .ZN(new_n2004_));
  AOI21_X1   g01812(.A1(new_n1986_), .A2(new_n2004_), .B(new_n450_), .ZN(new_n2005_));
  NOR2_X1    g01813(.A1(new_n1989_), .A2(new_n2005_), .ZN(new_n2006_));
  AOI21_X1   g01814(.A1(new_n2006_), .A2(new_n403_), .B(new_n1900_), .ZN(new_n2007_));
  OAI21_X1   g01815(.A1(new_n1989_), .A2(new_n2005_), .B(\asqrt[58] ), .ZN(new_n2008_));
  NAND2_X1   g01816(.A1(new_n2008_), .A2(new_n339_), .ZN(new_n2009_));
  OAI21_X1   g01817(.A1(new_n2007_), .A2(new_n2009_), .B(new_n1896_), .ZN(new_n2010_));
  INV_X1     g01818(.I(new_n2008_), .ZN(new_n2011_));
  OAI21_X1   g01819(.A1(new_n2007_), .A2(new_n2011_), .B(\asqrt[59] ), .ZN(new_n2012_));
  NAND3_X1   g01820(.A1(new_n2010_), .A2(new_n2012_), .A3(new_n288_), .ZN(new_n2013_));
  NAND2_X1   g01821(.A1(new_n2013_), .A2(new_n1894_), .ZN(new_n2014_));
  INV_X1     g01822(.I(new_n1896_), .ZN(new_n2015_));
  INV_X1     g01823(.I(new_n1906_), .ZN(new_n2016_));
  NOR2_X1    g01824(.A1(new_n2002_), .A2(new_n2003_), .ZN(new_n2017_));
  AOI21_X1   g01825(.A1(new_n2017_), .A2(new_n545_), .B(new_n2016_), .ZN(new_n2018_));
  NAND2_X1   g01826(.A1(new_n2004_), .A2(new_n450_), .ZN(new_n2019_));
  OAI21_X1   g01827(.A1(new_n2018_), .A2(new_n2019_), .B(new_n1902_), .ZN(new_n2020_));
  INV_X1     g01828(.I(new_n2004_), .ZN(new_n2021_));
  OAI21_X1   g01829(.A1(new_n2018_), .A2(new_n2021_), .B(\asqrt[57] ), .ZN(new_n2022_));
  NAND3_X1   g01830(.A1(new_n2020_), .A2(new_n2022_), .A3(new_n403_), .ZN(new_n2023_));
  NAND2_X1   g01831(.A1(new_n2023_), .A2(new_n1899_), .ZN(new_n2024_));
  NAND2_X1   g01832(.A1(new_n2020_), .A2(new_n2022_), .ZN(new_n2025_));
  AOI21_X1   g01833(.A1(new_n2025_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n2026_));
  AOI21_X1   g01834(.A1(new_n2026_), .A2(new_n2024_), .B(new_n2015_), .ZN(new_n2027_));
  AOI21_X1   g01835(.A1(new_n2024_), .A2(new_n2008_), .B(new_n339_), .ZN(new_n2028_));
  OAI21_X1   g01836(.A1(new_n2027_), .A2(new_n2028_), .B(\asqrt[60] ), .ZN(new_n2029_));
  AOI21_X1   g01837(.A1(new_n2014_), .A2(new_n2029_), .B(new_n242_), .ZN(new_n2030_));
  NAND3_X1   g01838(.A1(\asqrt[46] ), .A2(new_n1826_), .A3(new_n1842_), .ZN(new_n2031_));
  XOR2_X1    g01839(.A1(new_n2031_), .A2(new_n1868_), .Z(new_n2032_));
  INV_X1     g01840(.I(new_n2032_), .ZN(new_n2033_));
  NAND2_X1   g01841(.A1(new_n2010_), .A2(new_n2012_), .ZN(new_n2034_));
  AOI21_X1   g01842(.A1(new_n2034_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n2035_));
  AOI21_X1   g01843(.A1(new_n2035_), .A2(new_n2014_), .B(new_n2033_), .ZN(new_n2036_));
  OAI21_X1   g01844(.A1(new_n2036_), .A2(new_n2030_), .B(\asqrt[62] ), .ZN(new_n2037_));
  INV_X1     g01845(.I(new_n2037_), .ZN(new_n2038_));
  NOR2_X1    g01846(.A1(new_n2036_), .A2(new_n2030_), .ZN(new_n2039_));
  AOI21_X1   g01847(.A1(new_n1827_), .A2(new_n1848_), .B(new_n1843_), .ZN(new_n2040_));
  NAND2_X1   g01848(.A1(\asqrt[46] ), .A2(new_n2040_), .ZN(new_n2041_));
  XOR2_X1    g01849(.A1(new_n2041_), .A2(new_n1846_), .Z(new_n2042_));
  INV_X1     g01850(.I(new_n2042_), .ZN(new_n2043_));
  AOI21_X1   g01851(.A1(new_n2039_), .A2(new_n234_), .B(new_n2043_), .ZN(new_n2044_));
  OAI21_X1   g01852(.A1(new_n2044_), .A2(new_n2038_), .B(new_n1891_), .ZN(new_n2045_));
  OAI21_X1   g01853(.A1(new_n2045_), .A2(new_n1890_), .B(new_n193_), .ZN(new_n2046_));
  NOR2_X1    g01854(.A1(new_n2044_), .A2(new_n2038_), .ZN(new_n2047_));
  NAND2_X1   g01855(.A1(new_n2047_), .A2(new_n1890_), .ZN(new_n2048_));
  NOR2_X1    g01856(.A1(\asqrt[46] ), .A2(new_n1879_), .ZN(new_n2049_));
  INV_X1     g01857(.I(new_n2049_), .ZN(new_n2050_));
  NAND4_X1   g01858(.A1(new_n2046_), .A2(new_n1888_), .A3(new_n2048_), .A4(new_n2050_), .ZN(\asqrt[45] ));
  AOI21_X1   g01859(.A1(new_n1971_), .A2(new_n1972_), .B(new_n1975_), .ZN(new_n2052_));
  NAND2_X1   g01860(.A1(\asqrt[45] ), .A2(new_n2052_), .ZN(new_n2053_));
  XOR2_X1    g01861(.A1(new_n2053_), .A2(new_n1867_), .Z(new_n2054_));
  INV_X1     g01862(.I(new_n2054_), .ZN(new_n2055_));
  NOR2_X1    g01863(.A1(new_n1970_), .A2(\asqrt[50] ), .ZN(new_n2056_));
  INV_X1     g01864(.I(new_n1890_), .ZN(new_n2057_));
  INV_X1     g01865(.I(new_n1891_), .ZN(new_n2058_));
  INV_X1     g01866(.I(new_n1894_), .ZN(new_n2059_));
  NOR2_X1    g01867(.A1(new_n2027_), .A2(new_n2028_), .ZN(new_n2060_));
  AOI21_X1   g01868(.A1(new_n2060_), .A2(new_n288_), .B(new_n2059_), .ZN(new_n2061_));
  INV_X1     g01869(.I(new_n2029_), .ZN(new_n2062_));
  OAI21_X1   g01870(.A1(new_n2061_), .A2(new_n2062_), .B(\asqrt[61] ), .ZN(new_n2063_));
  NAND2_X1   g01871(.A1(new_n2029_), .A2(new_n242_), .ZN(new_n2064_));
  OAI21_X1   g01872(.A1(new_n2061_), .A2(new_n2064_), .B(new_n2032_), .ZN(new_n2065_));
  NAND3_X1   g01873(.A1(new_n2065_), .A2(new_n2063_), .A3(new_n234_), .ZN(new_n2066_));
  NAND2_X1   g01874(.A1(new_n2066_), .A2(new_n2042_), .ZN(new_n2067_));
  AOI21_X1   g01875(.A1(new_n2067_), .A2(new_n2037_), .B(new_n2058_), .ZN(new_n2068_));
  AOI21_X1   g01876(.A1(new_n2068_), .A2(new_n2057_), .B(\asqrt[63] ), .ZN(new_n2069_));
  NAND2_X1   g01877(.A1(new_n2067_), .A2(new_n2037_), .ZN(new_n2070_));
  NOR2_X1    g01878(.A1(new_n2070_), .A2(new_n2057_), .ZN(new_n2071_));
  NOR4_X1    g01879(.A1(new_n2069_), .A2(new_n1887_), .A3(new_n2071_), .A4(new_n2049_), .ZN(new_n2072_));
  NOR3_X1    g01880(.A1(new_n2072_), .A2(new_n2056_), .A3(new_n1949_), .ZN(new_n2073_));
  XOR2_X1    g01881(.A1(new_n2073_), .A2(new_n1921_), .Z(new_n2074_));
  NOR3_X1    g01882(.A1(new_n2072_), .A2(new_n1967_), .A3(new_n1944_), .ZN(new_n2075_));
  XOR2_X1    g01883(.A1(new_n2075_), .A2(new_n1943_), .Z(new_n2076_));
  INV_X1     g01884(.I(new_n2076_), .ZN(new_n2077_));
  NOR2_X1    g01885(.A1(new_n1938_), .A2(\asqrt[48] ), .ZN(new_n2078_));
  NOR3_X1    g01886(.A1(new_n2072_), .A2(new_n2078_), .A3(new_n1966_), .ZN(new_n2079_));
  XOR2_X1    g01887(.A1(new_n2079_), .A2(new_n1929_), .Z(new_n2080_));
  INV_X1     g01888(.I(new_n2080_), .ZN(new_n2081_));
  NAND3_X1   g01889(.A1(\asqrt[45] ), .A2(new_n1930_), .A3(new_n1931_), .ZN(new_n2082_));
  NOR4_X1    g01890(.A1(new_n2069_), .A2(new_n1884_), .A3(new_n1887_), .A4(new_n2071_), .ZN(new_n2083_));
  INV_X1     g01891(.I(new_n2083_), .ZN(new_n2084_));
  AOI21_X1   g01892(.A1(new_n2082_), .A2(new_n2084_), .B(\a[92] ), .ZN(new_n2085_));
  NOR3_X1    g01893(.A1(new_n2072_), .A2(\a[90] ), .A3(\a[91] ), .ZN(new_n2086_));
  NOR3_X1    g01894(.A1(new_n2086_), .A2(new_n1710_), .A3(new_n2083_), .ZN(new_n2087_));
  NOR2_X1    g01895(.A1(new_n2087_), .A2(new_n2085_), .ZN(new_n2088_));
  INV_X1     g01896(.I(\a[88] ), .ZN(new_n2089_));
  INV_X1     g01897(.I(\a[89] ), .ZN(new_n2090_));
  NAND3_X1   g01898(.A1(new_n2089_), .A2(new_n2090_), .A3(new_n1930_), .ZN(new_n2091_));
  OAI21_X1   g01899(.A1(new_n2072_), .A2(new_n1930_), .B(new_n2091_), .ZN(new_n2092_));
  NAND2_X1   g01900(.A1(new_n2092_), .A2(\asqrt[46] ), .ZN(new_n2093_));
  OAI21_X1   g01901(.A1(new_n2072_), .A2(\a[90] ), .B(\a[91] ), .ZN(new_n2094_));
  NAND2_X1   g01902(.A1(new_n2094_), .A2(new_n2082_), .ZN(new_n2095_));
  NOR2_X1    g01903(.A1(new_n2092_), .A2(\asqrt[46] ), .ZN(new_n2096_));
  OAI21_X1   g01904(.A1(new_n2095_), .A2(new_n2096_), .B(new_n2093_), .ZN(new_n2097_));
  OAI21_X1   g01905(.A1(\asqrt[47] ), .A2(new_n2097_), .B(new_n2088_), .ZN(new_n2098_));
  NAND2_X1   g01906(.A1(new_n2097_), .A2(\asqrt[47] ), .ZN(new_n2099_));
  NAND3_X1   g01907(.A1(new_n2098_), .A2(new_n1533_), .A3(new_n2099_), .ZN(new_n2100_));
  NOR3_X1    g01908(.A1(new_n2072_), .A2(new_n1960_), .A3(new_n1937_), .ZN(new_n2101_));
  XOR2_X1    g01909(.A1(new_n2101_), .A2(new_n1962_), .Z(new_n2102_));
  NAND2_X1   g01910(.A1(new_n2100_), .A2(new_n2102_), .ZN(new_n2103_));
  NAND2_X1   g01911(.A1(new_n2098_), .A2(new_n2099_), .ZN(new_n2104_));
  AOI21_X1   g01912(.A1(new_n2104_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n2105_));
  AOI21_X1   g01913(.A1(new_n2105_), .A2(new_n2103_), .B(new_n2081_), .ZN(new_n2106_));
  OAI21_X1   g01914(.A1(new_n2086_), .A2(new_n2083_), .B(new_n1710_), .ZN(new_n2107_));
  NAND3_X1   g01915(.A1(new_n2082_), .A2(\a[92] ), .A3(new_n2084_), .ZN(new_n2108_));
  NAND2_X1   g01916(.A1(new_n2107_), .A2(new_n2108_), .ZN(new_n2109_));
  NAND2_X1   g01917(.A1(\asqrt[45] ), .A2(\a[90] ), .ZN(new_n2110_));
  AOI21_X1   g01918(.A1(new_n2110_), .A2(new_n2091_), .B(new_n1884_), .ZN(new_n2111_));
  AOI21_X1   g01919(.A1(\asqrt[45] ), .A2(new_n1930_), .B(new_n1931_), .ZN(new_n2112_));
  NOR2_X1    g01920(.A1(new_n2112_), .A2(new_n2086_), .ZN(new_n2113_));
  NAND3_X1   g01921(.A1(new_n2110_), .A2(new_n1884_), .A3(new_n2091_), .ZN(new_n2114_));
  AOI21_X1   g01922(.A1(new_n2113_), .A2(new_n2114_), .B(new_n2111_), .ZN(new_n2115_));
  AOI21_X1   g01923(.A1(new_n2115_), .A2(new_n1688_), .B(new_n2109_), .ZN(new_n2116_));
  NOR2_X1    g01924(.A1(new_n2115_), .A2(new_n1688_), .ZN(new_n2117_));
  OAI21_X1   g01925(.A1(new_n2116_), .A2(new_n2117_), .B(\asqrt[48] ), .ZN(new_n2118_));
  AOI21_X1   g01926(.A1(new_n2103_), .A2(new_n2118_), .B(new_n1368_), .ZN(new_n2119_));
  NOR2_X1    g01927(.A1(new_n2106_), .A2(new_n2119_), .ZN(new_n2120_));
  AOI21_X1   g01928(.A1(new_n2120_), .A2(new_n1228_), .B(new_n2077_), .ZN(new_n2121_));
  OAI21_X1   g01929(.A1(new_n2106_), .A2(new_n2119_), .B(\asqrt[50] ), .ZN(new_n2122_));
  NAND2_X1   g01930(.A1(new_n2122_), .A2(new_n1088_), .ZN(new_n2123_));
  OAI21_X1   g01931(.A1(new_n2121_), .A2(new_n2123_), .B(new_n2074_), .ZN(new_n2124_));
  INV_X1     g01932(.I(new_n2122_), .ZN(new_n2125_));
  OAI21_X1   g01933(.A1(new_n2121_), .A2(new_n2125_), .B(\asqrt[51] ), .ZN(new_n2126_));
  NAND3_X1   g01934(.A1(new_n2124_), .A2(new_n2126_), .A3(new_n962_), .ZN(new_n2127_));
  INV_X1     g01935(.I(new_n2074_), .ZN(new_n2128_));
  NOR2_X1    g01936(.A1(new_n2116_), .A2(new_n2117_), .ZN(new_n2129_));
  INV_X1     g01937(.I(new_n2102_), .ZN(new_n2130_));
  AOI21_X1   g01938(.A1(new_n2129_), .A2(new_n1533_), .B(new_n2130_), .ZN(new_n2131_));
  NAND2_X1   g01939(.A1(new_n2118_), .A2(new_n1368_), .ZN(new_n2132_));
  OAI21_X1   g01940(.A1(new_n2131_), .A2(new_n2132_), .B(new_n2080_), .ZN(new_n2133_));
  INV_X1     g01941(.I(new_n2118_), .ZN(new_n2134_));
  OAI21_X1   g01942(.A1(new_n2131_), .A2(new_n2134_), .B(\asqrt[49] ), .ZN(new_n2135_));
  NAND3_X1   g01943(.A1(new_n2133_), .A2(new_n2135_), .A3(new_n1228_), .ZN(new_n2136_));
  NAND2_X1   g01944(.A1(new_n2136_), .A2(new_n2076_), .ZN(new_n2137_));
  NAND2_X1   g01945(.A1(new_n2133_), .A2(new_n2135_), .ZN(new_n2138_));
  AOI21_X1   g01946(.A1(new_n2138_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n2139_));
  AOI21_X1   g01947(.A1(new_n2139_), .A2(new_n2137_), .B(new_n2128_), .ZN(new_n2140_));
  AOI21_X1   g01948(.A1(new_n2137_), .A2(new_n2122_), .B(new_n1088_), .ZN(new_n2141_));
  OAI21_X1   g01949(.A1(new_n2140_), .A2(new_n2141_), .B(\asqrt[52] ), .ZN(new_n2142_));
  NAND2_X1   g01950(.A1(new_n2070_), .A2(new_n1890_), .ZN(new_n2143_));
  NOR2_X1    g01951(.A1(new_n2072_), .A2(new_n1890_), .ZN(new_n2144_));
  NAND2_X1   g01952(.A1(new_n2144_), .A2(new_n2047_), .ZN(new_n2145_));
  AOI21_X1   g01953(.A1(new_n2145_), .A2(new_n2143_), .B(new_n193_), .ZN(new_n2146_));
  INV_X1     g01954(.I(new_n2146_), .ZN(new_n2147_));
  NAND3_X1   g01955(.A1(\asqrt[45] ), .A2(new_n2037_), .A3(new_n2066_), .ZN(new_n2148_));
  XOR2_X1    g01956(.A1(new_n2148_), .A2(new_n2042_), .Z(new_n2149_));
  AOI21_X1   g01957(.A1(new_n2144_), .A2(new_n2070_), .B(new_n2071_), .ZN(new_n2150_));
  OAI21_X1   g01958(.A1(new_n2007_), .A2(new_n2009_), .B(new_n2012_), .ZN(new_n2151_));
  NOR2_X1    g01959(.A1(new_n2072_), .A2(new_n2151_), .ZN(new_n2152_));
  XOR2_X1    g01960(.A1(new_n2152_), .A2(new_n1896_), .Z(new_n2153_));
  NAND3_X1   g01961(.A1(\asqrt[45] ), .A2(new_n2023_), .A3(new_n2008_), .ZN(new_n2154_));
  XOR2_X1    g01962(.A1(new_n2154_), .A2(new_n1900_), .Z(new_n2155_));
  OAI21_X1   g01963(.A1(new_n2018_), .A2(new_n2019_), .B(new_n2022_), .ZN(new_n2156_));
  NOR2_X1    g01964(.A1(new_n2072_), .A2(new_n2156_), .ZN(new_n2157_));
  XOR2_X1    g01965(.A1(new_n2157_), .A2(new_n1902_), .Z(new_n2158_));
  INV_X1     g01966(.I(new_n2158_), .ZN(new_n2159_));
  NAND3_X1   g01967(.A1(\asqrt[45] ), .A2(new_n1985_), .A3(new_n2004_), .ZN(new_n2160_));
  XOR2_X1    g01968(.A1(new_n2160_), .A2(new_n2016_), .Z(new_n2161_));
  INV_X1     g01969(.I(new_n2161_), .ZN(new_n2162_));
  OAI21_X1   g01970(.A1(new_n1979_), .A2(new_n1981_), .B(new_n1984_), .ZN(new_n2163_));
  NOR2_X1    g01971(.A1(new_n2072_), .A2(new_n2163_), .ZN(new_n2164_));
  XOR2_X1    g01972(.A1(new_n2164_), .A2(new_n1908_), .Z(new_n2165_));
  NAND3_X1   g01973(.A1(\asqrt[45] ), .A2(new_n1998_), .A3(new_n1980_), .ZN(new_n2166_));
  XOR2_X1    g01974(.A1(new_n2166_), .A2(new_n1912_), .Z(new_n2167_));
  OAI21_X1   g01975(.A1(new_n1993_), .A2(new_n1994_), .B(new_n1997_), .ZN(new_n2168_));
  NOR2_X1    g01976(.A1(new_n2072_), .A2(new_n2168_), .ZN(new_n2169_));
  XOR2_X1    g01977(.A1(new_n2169_), .A2(new_n1914_), .Z(new_n2170_));
  INV_X1     g01978(.I(new_n2170_), .ZN(new_n2171_));
  NAND3_X1   g01979(.A1(\asqrt[45] ), .A2(new_n1951_), .A3(new_n1976_), .ZN(new_n2172_));
  XOR2_X1    g01980(.A1(new_n2172_), .A2(new_n1991_), .Z(new_n2173_));
  INV_X1     g01981(.I(new_n2173_), .ZN(new_n2174_));
  NAND2_X1   g01982(.A1(new_n2127_), .A2(new_n2054_), .ZN(new_n2175_));
  NAND2_X1   g01983(.A1(new_n2124_), .A2(new_n2126_), .ZN(new_n2176_));
  AOI21_X1   g01984(.A1(new_n2176_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n2177_));
  AOI21_X1   g01985(.A1(new_n2177_), .A2(new_n2175_), .B(new_n2174_), .ZN(new_n2178_));
  AOI21_X1   g01986(.A1(new_n2175_), .A2(new_n2142_), .B(new_n842_), .ZN(new_n2179_));
  NOR2_X1    g01987(.A1(new_n2178_), .A2(new_n2179_), .ZN(new_n2180_));
  AOI21_X1   g01988(.A1(new_n2180_), .A2(new_n720_), .B(new_n2171_), .ZN(new_n2181_));
  OAI21_X1   g01989(.A1(new_n2178_), .A2(new_n2179_), .B(\asqrt[54] ), .ZN(new_n2182_));
  NAND2_X1   g01990(.A1(new_n2182_), .A2(new_n630_), .ZN(new_n2183_));
  OAI21_X1   g01991(.A1(new_n2181_), .A2(new_n2183_), .B(new_n2167_), .ZN(new_n2184_));
  INV_X1     g01992(.I(new_n2182_), .ZN(new_n2185_));
  OAI21_X1   g01993(.A1(new_n2181_), .A2(new_n2185_), .B(\asqrt[55] ), .ZN(new_n2186_));
  NAND3_X1   g01994(.A1(new_n2184_), .A2(new_n2186_), .A3(new_n545_), .ZN(new_n2187_));
  NAND2_X1   g01995(.A1(new_n2187_), .A2(new_n2165_), .ZN(new_n2188_));
  NAND2_X1   g01996(.A1(new_n2184_), .A2(new_n2186_), .ZN(new_n2189_));
  AOI21_X1   g01997(.A1(new_n2189_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n2190_));
  AOI21_X1   g01998(.A1(new_n2190_), .A2(new_n2188_), .B(new_n2162_), .ZN(new_n2191_));
  INV_X1     g01999(.I(new_n2167_), .ZN(new_n2192_));
  NOR2_X1    g02000(.A1(new_n2140_), .A2(new_n2141_), .ZN(new_n2193_));
  AOI21_X1   g02001(.A1(new_n2193_), .A2(new_n962_), .B(new_n2055_), .ZN(new_n2194_));
  NAND2_X1   g02002(.A1(new_n2142_), .A2(new_n842_), .ZN(new_n2195_));
  OAI21_X1   g02003(.A1(new_n2194_), .A2(new_n2195_), .B(new_n2173_), .ZN(new_n2196_));
  INV_X1     g02004(.I(new_n2142_), .ZN(new_n2197_));
  OAI21_X1   g02005(.A1(new_n2194_), .A2(new_n2197_), .B(\asqrt[53] ), .ZN(new_n2198_));
  NAND3_X1   g02006(.A1(new_n2196_), .A2(new_n2198_), .A3(new_n720_), .ZN(new_n2199_));
  NAND2_X1   g02007(.A1(new_n2199_), .A2(new_n2170_), .ZN(new_n2200_));
  NAND2_X1   g02008(.A1(new_n2196_), .A2(new_n2198_), .ZN(new_n2201_));
  AOI21_X1   g02009(.A1(new_n2201_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n2202_));
  AOI21_X1   g02010(.A1(new_n2202_), .A2(new_n2200_), .B(new_n2192_), .ZN(new_n2203_));
  AOI21_X1   g02011(.A1(new_n2200_), .A2(new_n2182_), .B(new_n630_), .ZN(new_n2204_));
  OAI21_X1   g02012(.A1(new_n2203_), .A2(new_n2204_), .B(\asqrt[56] ), .ZN(new_n2205_));
  AOI21_X1   g02013(.A1(new_n2188_), .A2(new_n2205_), .B(new_n450_), .ZN(new_n2206_));
  NOR2_X1    g02014(.A1(new_n2191_), .A2(new_n2206_), .ZN(new_n2207_));
  AOI21_X1   g02015(.A1(new_n2207_), .A2(new_n403_), .B(new_n2159_), .ZN(new_n2208_));
  OAI21_X1   g02016(.A1(new_n2191_), .A2(new_n2206_), .B(\asqrt[58] ), .ZN(new_n2209_));
  NAND2_X1   g02017(.A1(new_n2209_), .A2(new_n339_), .ZN(new_n2210_));
  OAI21_X1   g02018(.A1(new_n2208_), .A2(new_n2210_), .B(new_n2155_), .ZN(new_n2211_));
  INV_X1     g02019(.I(new_n2209_), .ZN(new_n2212_));
  OAI21_X1   g02020(.A1(new_n2208_), .A2(new_n2212_), .B(\asqrt[59] ), .ZN(new_n2213_));
  NAND3_X1   g02021(.A1(new_n2211_), .A2(new_n2213_), .A3(new_n288_), .ZN(new_n2214_));
  NAND2_X1   g02022(.A1(new_n2214_), .A2(new_n2153_), .ZN(new_n2215_));
  INV_X1     g02023(.I(new_n2155_), .ZN(new_n2216_));
  INV_X1     g02024(.I(new_n2165_), .ZN(new_n2217_));
  NOR2_X1    g02025(.A1(new_n2203_), .A2(new_n2204_), .ZN(new_n2218_));
  AOI21_X1   g02026(.A1(new_n2218_), .A2(new_n545_), .B(new_n2217_), .ZN(new_n2219_));
  NAND2_X1   g02027(.A1(new_n2205_), .A2(new_n450_), .ZN(new_n2220_));
  OAI21_X1   g02028(.A1(new_n2219_), .A2(new_n2220_), .B(new_n2161_), .ZN(new_n2221_));
  INV_X1     g02029(.I(new_n2205_), .ZN(new_n2222_));
  OAI21_X1   g02030(.A1(new_n2219_), .A2(new_n2222_), .B(\asqrt[57] ), .ZN(new_n2223_));
  NAND3_X1   g02031(.A1(new_n2221_), .A2(new_n2223_), .A3(new_n403_), .ZN(new_n2224_));
  NAND2_X1   g02032(.A1(new_n2224_), .A2(new_n2158_), .ZN(new_n2225_));
  NAND2_X1   g02033(.A1(new_n2221_), .A2(new_n2223_), .ZN(new_n2226_));
  AOI21_X1   g02034(.A1(new_n2226_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n2227_));
  AOI21_X1   g02035(.A1(new_n2227_), .A2(new_n2225_), .B(new_n2216_), .ZN(new_n2228_));
  AOI21_X1   g02036(.A1(new_n2225_), .A2(new_n2209_), .B(new_n339_), .ZN(new_n2229_));
  OAI21_X1   g02037(.A1(new_n2228_), .A2(new_n2229_), .B(\asqrt[60] ), .ZN(new_n2230_));
  AOI21_X1   g02038(.A1(new_n2215_), .A2(new_n2230_), .B(new_n242_), .ZN(new_n2231_));
  NAND3_X1   g02039(.A1(\asqrt[45] ), .A2(new_n2013_), .A3(new_n2029_), .ZN(new_n2232_));
  XOR2_X1    g02040(.A1(new_n2232_), .A2(new_n2059_), .Z(new_n2233_));
  INV_X1     g02041(.I(new_n2233_), .ZN(new_n2234_));
  NAND2_X1   g02042(.A1(new_n2211_), .A2(new_n2213_), .ZN(new_n2235_));
  AOI21_X1   g02043(.A1(new_n2235_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n2236_));
  AOI21_X1   g02044(.A1(new_n2236_), .A2(new_n2215_), .B(new_n2234_), .ZN(new_n2237_));
  OAI21_X1   g02045(.A1(new_n2237_), .A2(new_n2231_), .B(\asqrt[62] ), .ZN(new_n2238_));
  INV_X1     g02046(.I(new_n2238_), .ZN(new_n2239_));
  NOR2_X1    g02047(.A1(new_n2237_), .A2(new_n2231_), .ZN(new_n2240_));
  AOI21_X1   g02048(.A1(new_n2014_), .A2(new_n2035_), .B(new_n2030_), .ZN(new_n2241_));
  NAND2_X1   g02049(.A1(\asqrt[45] ), .A2(new_n2241_), .ZN(new_n2242_));
  XOR2_X1    g02050(.A1(new_n2242_), .A2(new_n2033_), .Z(new_n2243_));
  INV_X1     g02051(.I(new_n2243_), .ZN(new_n2244_));
  AOI21_X1   g02052(.A1(new_n2240_), .A2(new_n234_), .B(new_n2244_), .ZN(new_n2245_));
  OAI21_X1   g02053(.A1(new_n2245_), .A2(new_n2239_), .B(new_n2150_), .ZN(new_n2246_));
  OAI21_X1   g02054(.A1(new_n2246_), .A2(new_n2149_), .B(new_n193_), .ZN(new_n2247_));
  NOR2_X1    g02055(.A1(new_n2245_), .A2(new_n2239_), .ZN(new_n2248_));
  NAND2_X1   g02056(.A1(new_n2248_), .A2(new_n2149_), .ZN(new_n2249_));
  NOR2_X1    g02057(.A1(\asqrt[45] ), .A2(new_n2057_), .ZN(new_n2250_));
  INV_X1     g02058(.I(new_n2250_), .ZN(new_n2251_));
  NAND4_X1   g02059(.A1(new_n2247_), .A2(new_n2147_), .A3(new_n2249_), .A4(new_n2251_), .ZN(\asqrt[44] ));
  NAND3_X1   g02060(.A1(\asqrt[44] ), .A2(new_n2127_), .A3(new_n2142_), .ZN(new_n2253_));
  XOR2_X1    g02061(.A1(new_n2253_), .A2(new_n2055_), .Z(new_n2254_));
  INV_X1     g02062(.I(new_n2153_), .ZN(new_n2255_));
  NOR2_X1    g02063(.A1(new_n2228_), .A2(new_n2229_), .ZN(new_n2256_));
  AOI21_X1   g02064(.A1(new_n2256_), .A2(new_n288_), .B(new_n2255_), .ZN(new_n2257_));
  INV_X1     g02065(.I(new_n2230_), .ZN(new_n2258_));
  OAI21_X1   g02066(.A1(new_n2257_), .A2(new_n2258_), .B(\asqrt[61] ), .ZN(new_n2259_));
  NAND2_X1   g02067(.A1(new_n2230_), .A2(new_n242_), .ZN(new_n2260_));
  OAI21_X1   g02068(.A1(new_n2257_), .A2(new_n2260_), .B(new_n2233_), .ZN(new_n2261_));
  NAND3_X1   g02069(.A1(new_n2261_), .A2(new_n2259_), .A3(new_n234_), .ZN(new_n2262_));
  NAND2_X1   g02070(.A1(new_n2262_), .A2(new_n2243_), .ZN(new_n2263_));
  NAND2_X1   g02071(.A1(new_n2263_), .A2(new_n2238_), .ZN(new_n2264_));
  NAND2_X1   g02072(.A1(new_n2264_), .A2(new_n2149_), .ZN(new_n2265_));
  INV_X1     g02073(.I(new_n2149_), .ZN(new_n2266_));
  INV_X1     g02074(.I(new_n2150_), .ZN(new_n2267_));
  AOI21_X1   g02075(.A1(new_n2263_), .A2(new_n2238_), .B(new_n2267_), .ZN(new_n2268_));
  AOI21_X1   g02076(.A1(new_n2268_), .A2(new_n2266_), .B(\asqrt[63] ), .ZN(new_n2269_));
  NOR2_X1    g02077(.A1(new_n2264_), .A2(new_n2266_), .ZN(new_n2270_));
  NOR4_X1    g02078(.A1(new_n2269_), .A2(new_n2146_), .A3(new_n2270_), .A4(new_n2250_), .ZN(new_n2271_));
  NOR2_X1    g02079(.A1(new_n2271_), .A2(new_n2149_), .ZN(new_n2272_));
  NAND2_X1   g02080(.A1(new_n2272_), .A2(new_n2248_), .ZN(new_n2273_));
  AOI21_X1   g02081(.A1(new_n2273_), .A2(new_n2265_), .B(new_n193_), .ZN(new_n2274_));
  NAND3_X1   g02082(.A1(\asqrt[44] ), .A2(new_n2238_), .A3(new_n2262_), .ZN(new_n2275_));
  XOR2_X1    g02083(.A1(new_n2275_), .A2(new_n2243_), .Z(new_n2276_));
  INV_X1     g02084(.I(new_n2276_), .ZN(new_n2277_));
  AOI21_X1   g02085(.A1(new_n2272_), .A2(new_n2264_), .B(new_n2270_), .ZN(new_n2278_));
  INV_X1     g02086(.I(new_n2278_), .ZN(new_n2279_));
  OAI21_X1   g02087(.A1(new_n2208_), .A2(new_n2210_), .B(new_n2213_), .ZN(new_n2280_));
  NOR2_X1    g02088(.A1(new_n2271_), .A2(new_n2280_), .ZN(new_n2281_));
  XOR2_X1    g02089(.A1(new_n2281_), .A2(new_n2155_), .Z(new_n2282_));
  NAND3_X1   g02090(.A1(\asqrt[44] ), .A2(new_n2224_), .A3(new_n2209_), .ZN(new_n2283_));
  XOR2_X1    g02091(.A1(new_n2283_), .A2(new_n2159_), .Z(new_n2284_));
  OAI21_X1   g02092(.A1(new_n2219_), .A2(new_n2220_), .B(new_n2223_), .ZN(new_n2285_));
  NOR2_X1    g02093(.A1(new_n2271_), .A2(new_n2285_), .ZN(new_n2286_));
  XOR2_X1    g02094(.A1(new_n2286_), .A2(new_n2161_), .Z(new_n2287_));
  INV_X1     g02095(.I(new_n2287_), .ZN(new_n2288_));
  NAND3_X1   g02096(.A1(\asqrt[44] ), .A2(new_n2187_), .A3(new_n2205_), .ZN(new_n2289_));
  XOR2_X1    g02097(.A1(new_n2289_), .A2(new_n2217_), .Z(new_n2290_));
  INV_X1     g02098(.I(new_n2290_), .ZN(new_n2291_));
  OAI21_X1   g02099(.A1(new_n2181_), .A2(new_n2183_), .B(new_n2186_), .ZN(new_n2292_));
  NOR2_X1    g02100(.A1(new_n2271_), .A2(new_n2292_), .ZN(new_n2293_));
  XOR2_X1    g02101(.A1(new_n2293_), .A2(new_n2167_), .Z(new_n2294_));
  NAND3_X1   g02102(.A1(\asqrt[44] ), .A2(new_n2199_), .A3(new_n2182_), .ZN(new_n2295_));
  XOR2_X1    g02103(.A1(new_n2295_), .A2(new_n2171_), .Z(new_n2296_));
  OAI21_X1   g02104(.A1(new_n2194_), .A2(new_n2195_), .B(new_n2198_), .ZN(new_n2297_));
  NOR2_X1    g02105(.A1(new_n2271_), .A2(new_n2297_), .ZN(new_n2298_));
  XOR2_X1    g02106(.A1(new_n2298_), .A2(new_n2173_), .Z(new_n2299_));
  INV_X1     g02107(.I(new_n2299_), .ZN(new_n2300_));
  INV_X1     g02108(.I(new_n2254_), .ZN(new_n2301_));
  OAI21_X1   g02109(.A1(new_n2121_), .A2(new_n2123_), .B(new_n2126_), .ZN(new_n2302_));
  NOR2_X1    g02110(.A1(new_n2271_), .A2(new_n2302_), .ZN(new_n2303_));
  XOR2_X1    g02111(.A1(new_n2303_), .A2(new_n2074_), .Z(new_n2304_));
  NAND3_X1   g02112(.A1(\asqrt[44] ), .A2(new_n2136_), .A3(new_n2122_), .ZN(new_n2305_));
  XOR2_X1    g02113(.A1(new_n2305_), .A2(new_n2077_), .Z(new_n2306_));
  OAI21_X1   g02114(.A1(new_n2131_), .A2(new_n2132_), .B(new_n2135_), .ZN(new_n2307_));
  NOR2_X1    g02115(.A1(new_n2271_), .A2(new_n2307_), .ZN(new_n2308_));
  XOR2_X1    g02116(.A1(new_n2308_), .A2(new_n2080_), .Z(new_n2309_));
  INV_X1     g02117(.I(new_n2309_), .ZN(new_n2310_));
  NAND3_X1   g02118(.A1(\asqrt[44] ), .A2(new_n2100_), .A3(new_n2118_), .ZN(new_n2311_));
  XOR2_X1    g02119(.A1(new_n2311_), .A2(new_n2130_), .Z(new_n2312_));
  INV_X1     g02120(.I(new_n2312_), .ZN(new_n2313_));
  NOR2_X1    g02121(.A1(new_n2097_), .A2(\asqrt[47] ), .ZN(new_n2314_));
  NOR3_X1    g02122(.A1(new_n2271_), .A2(new_n2314_), .A3(new_n2117_), .ZN(new_n2315_));
  XOR2_X1    g02123(.A1(new_n2315_), .A2(new_n2088_), .Z(new_n2316_));
  NOR3_X1    g02124(.A1(new_n2271_), .A2(\a[88] ), .A3(\a[89] ), .ZN(new_n2317_));
  NOR4_X1    g02125(.A1(new_n2269_), .A2(new_n2072_), .A3(new_n2146_), .A4(new_n2270_), .ZN(new_n2318_));
  OAI21_X1   g02126(.A1(new_n2317_), .A2(new_n2318_), .B(new_n1930_), .ZN(new_n2319_));
  NAND3_X1   g02127(.A1(\asqrt[44] ), .A2(new_n2089_), .A3(new_n2090_), .ZN(new_n2320_));
  INV_X1     g02128(.I(new_n2318_), .ZN(new_n2321_));
  NAND3_X1   g02129(.A1(new_n2320_), .A2(\a[90] ), .A3(new_n2321_), .ZN(new_n2322_));
  NAND2_X1   g02130(.A1(new_n2319_), .A2(new_n2322_), .ZN(new_n2323_));
  INV_X1     g02131(.I(\a[86] ), .ZN(new_n2324_));
  INV_X1     g02132(.I(\a[87] ), .ZN(new_n2325_));
  NAND3_X1   g02133(.A1(new_n2324_), .A2(new_n2325_), .A3(new_n2089_), .ZN(new_n2326_));
  NAND2_X1   g02134(.A1(\asqrt[44] ), .A2(\a[88] ), .ZN(new_n2327_));
  AOI21_X1   g02135(.A1(new_n2327_), .A2(new_n2326_), .B(new_n2072_), .ZN(new_n2328_));
  AOI21_X1   g02136(.A1(\asqrt[44] ), .A2(new_n2089_), .B(new_n2090_), .ZN(new_n2329_));
  NOR2_X1    g02137(.A1(new_n2317_), .A2(new_n2329_), .ZN(new_n2330_));
  NAND3_X1   g02138(.A1(new_n2327_), .A2(new_n2072_), .A3(new_n2326_), .ZN(new_n2331_));
  AOI21_X1   g02139(.A1(new_n2330_), .A2(new_n2331_), .B(new_n2328_), .ZN(new_n2332_));
  AOI21_X1   g02140(.A1(new_n2332_), .A2(new_n1884_), .B(new_n2323_), .ZN(new_n2333_));
  NOR2_X1    g02141(.A1(new_n2332_), .A2(new_n1884_), .ZN(new_n2334_));
  NOR3_X1    g02142(.A1(new_n2333_), .A2(\asqrt[47] ), .A3(new_n2334_), .ZN(new_n2335_));
  NOR3_X1    g02143(.A1(new_n2271_), .A2(new_n2111_), .A3(new_n2096_), .ZN(new_n2336_));
  XOR2_X1    g02144(.A1(new_n2336_), .A2(new_n2113_), .Z(new_n2337_));
  INV_X1     g02145(.I(new_n2337_), .ZN(new_n2338_));
  OAI21_X1   g02146(.A1(new_n2333_), .A2(new_n2334_), .B(\asqrt[47] ), .ZN(new_n2339_));
  OAI21_X1   g02147(.A1(new_n2335_), .A2(new_n2338_), .B(new_n2339_), .ZN(new_n2340_));
  OAI21_X1   g02148(.A1(new_n2340_), .A2(\asqrt[48] ), .B(new_n2316_), .ZN(new_n2341_));
  AOI21_X1   g02149(.A1(new_n2340_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n2342_));
  AOI21_X1   g02150(.A1(new_n2342_), .A2(new_n2341_), .B(new_n2313_), .ZN(new_n2343_));
  NAND2_X1   g02151(.A1(new_n2340_), .A2(\asqrt[48] ), .ZN(new_n2344_));
  AOI21_X1   g02152(.A1(new_n2341_), .A2(new_n2344_), .B(new_n1368_), .ZN(new_n2345_));
  NOR2_X1    g02153(.A1(new_n2343_), .A2(new_n2345_), .ZN(new_n2346_));
  AOI21_X1   g02154(.A1(new_n2346_), .A2(new_n1228_), .B(new_n2310_), .ZN(new_n2347_));
  OAI21_X1   g02155(.A1(new_n2343_), .A2(new_n2345_), .B(\asqrt[50] ), .ZN(new_n2348_));
  NAND2_X1   g02156(.A1(new_n2348_), .A2(new_n1088_), .ZN(new_n2349_));
  OAI21_X1   g02157(.A1(new_n2347_), .A2(new_n2349_), .B(new_n2306_), .ZN(new_n2350_));
  INV_X1     g02158(.I(new_n2348_), .ZN(new_n2351_));
  OAI21_X1   g02159(.A1(new_n2347_), .A2(new_n2351_), .B(\asqrt[51] ), .ZN(new_n2352_));
  NAND3_X1   g02160(.A1(new_n2350_), .A2(new_n2352_), .A3(new_n962_), .ZN(new_n2353_));
  NAND2_X1   g02161(.A1(new_n2353_), .A2(new_n2304_), .ZN(new_n2354_));
  NAND2_X1   g02162(.A1(new_n2350_), .A2(new_n2352_), .ZN(new_n2355_));
  AOI21_X1   g02163(.A1(new_n2355_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n2356_));
  AOI21_X1   g02164(.A1(new_n2356_), .A2(new_n2354_), .B(new_n2301_), .ZN(new_n2357_));
  INV_X1     g02165(.I(new_n2306_), .ZN(new_n2358_));
  INV_X1     g02166(.I(new_n2316_), .ZN(new_n2359_));
  AOI21_X1   g02167(.A1(new_n2320_), .A2(new_n2321_), .B(\a[90] ), .ZN(new_n2360_));
  NOR3_X1    g02168(.A1(new_n2317_), .A2(new_n1930_), .A3(new_n2318_), .ZN(new_n2361_));
  NOR2_X1    g02169(.A1(new_n2361_), .A2(new_n2360_), .ZN(new_n2362_));
  OAI21_X1   g02170(.A1(new_n2271_), .A2(new_n2089_), .B(new_n2326_), .ZN(new_n2363_));
  NAND2_X1   g02171(.A1(new_n2363_), .A2(\asqrt[45] ), .ZN(new_n2364_));
  OAI21_X1   g02172(.A1(new_n2271_), .A2(\a[88] ), .B(\a[89] ), .ZN(new_n2365_));
  NAND2_X1   g02173(.A1(new_n2365_), .A2(new_n2320_), .ZN(new_n2366_));
  NOR2_X1    g02174(.A1(new_n2363_), .A2(\asqrt[45] ), .ZN(new_n2367_));
  OAI21_X1   g02175(.A1(new_n2366_), .A2(new_n2367_), .B(new_n2364_), .ZN(new_n2368_));
  OAI21_X1   g02176(.A1(\asqrt[46] ), .A2(new_n2368_), .B(new_n2362_), .ZN(new_n2369_));
  NAND2_X1   g02177(.A1(new_n2368_), .A2(\asqrt[46] ), .ZN(new_n2370_));
  NAND3_X1   g02178(.A1(new_n2369_), .A2(new_n1688_), .A3(new_n2370_), .ZN(new_n2371_));
  AOI21_X1   g02179(.A1(new_n2369_), .A2(new_n2370_), .B(new_n1688_), .ZN(new_n2372_));
  AOI21_X1   g02180(.A1(new_n2371_), .A2(new_n2337_), .B(new_n2372_), .ZN(new_n2373_));
  AOI21_X1   g02181(.A1(new_n2373_), .A2(new_n1533_), .B(new_n2359_), .ZN(new_n2374_));
  OAI21_X1   g02182(.A1(new_n2373_), .A2(new_n1533_), .B(new_n1368_), .ZN(new_n2375_));
  OAI21_X1   g02183(.A1(new_n2374_), .A2(new_n2375_), .B(new_n2312_), .ZN(new_n2376_));
  NOR2_X1    g02184(.A1(new_n2373_), .A2(new_n1533_), .ZN(new_n2377_));
  OAI21_X1   g02185(.A1(new_n2374_), .A2(new_n2377_), .B(\asqrt[49] ), .ZN(new_n2378_));
  NAND3_X1   g02186(.A1(new_n2376_), .A2(new_n2378_), .A3(new_n1228_), .ZN(new_n2379_));
  NAND2_X1   g02187(.A1(new_n2379_), .A2(new_n2309_), .ZN(new_n2380_));
  NAND2_X1   g02188(.A1(new_n2376_), .A2(new_n2378_), .ZN(new_n2381_));
  AOI21_X1   g02189(.A1(new_n2381_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n2382_));
  AOI21_X1   g02190(.A1(new_n2382_), .A2(new_n2380_), .B(new_n2358_), .ZN(new_n2383_));
  AOI21_X1   g02191(.A1(new_n2380_), .A2(new_n2348_), .B(new_n1088_), .ZN(new_n2384_));
  OAI21_X1   g02192(.A1(new_n2383_), .A2(new_n2384_), .B(\asqrt[52] ), .ZN(new_n2385_));
  AOI21_X1   g02193(.A1(new_n2354_), .A2(new_n2385_), .B(new_n842_), .ZN(new_n2386_));
  NOR2_X1    g02194(.A1(new_n2357_), .A2(new_n2386_), .ZN(new_n2387_));
  AOI21_X1   g02195(.A1(new_n2387_), .A2(new_n720_), .B(new_n2300_), .ZN(new_n2388_));
  OAI21_X1   g02196(.A1(new_n2357_), .A2(new_n2386_), .B(\asqrt[54] ), .ZN(new_n2389_));
  NAND2_X1   g02197(.A1(new_n2389_), .A2(new_n630_), .ZN(new_n2390_));
  OAI21_X1   g02198(.A1(new_n2388_), .A2(new_n2390_), .B(new_n2296_), .ZN(new_n2391_));
  INV_X1     g02199(.I(new_n2389_), .ZN(new_n2392_));
  OAI21_X1   g02200(.A1(new_n2388_), .A2(new_n2392_), .B(\asqrt[55] ), .ZN(new_n2393_));
  NAND3_X1   g02201(.A1(new_n2391_), .A2(new_n2393_), .A3(new_n545_), .ZN(new_n2394_));
  NAND2_X1   g02202(.A1(new_n2394_), .A2(new_n2294_), .ZN(new_n2395_));
  NAND2_X1   g02203(.A1(new_n2391_), .A2(new_n2393_), .ZN(new_n2396_));
  AOI21_X1   g02204(.A1(new_n2396_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n2397_));
  AOI21_X1   g02205(.A1(new_n2397_), .A2(new_n2395_), .B(new_n2291_), .ZN(new_n2398_));
  INV_X1     g02206(.I(new_n2296_), .ZN(new_n2399_));
  INV_X1     g02207(.I(new_n2304_), .ZN(new_n2400_));
  NOR2_X1    g02208(.A1(new_n2383_), .A2(new_n2384_), .ZN(new_n2401_));
  AOI21_X1   g02209(.A1(new_n2401_), .A2(new_n962_), .B(new_n2400_), .ZN(new_n2402_));
  NAND2_X1   g02210(.A1(new_n2385_), .A2(new_n842_), .ZN(new_n2403_));
  OAI21_X1   g02211(.A1(new_n2402_), .A2(new_n2403_), .B(new_n2254_), .ZN(new_n2404_));
  INV_X1     g02212(.I(new_n2385_), .ZN(new_n2405_));
  OAI21_X1   g02213(.A1(new_n2402_), .A2(new_n2405_), .B(\asqrt[53] ), .ZN(new_n2406_));
  NAND3_X1   g02214(.A1(new_n2404_), .A2(new_n2406_), .A3(new_n720_), .ZN(new_n2407_));
  NAND2_X1   g02215(.A1(new_n2407_), .A2(new_n2299_), .ZN(new_n2408_));
  NAND2_X1   g02216(.A1(new_n2404_), .A2(new_n2406_), .ZN(new_n2409_));
  AOI21_X1   g02217(.A1(new_n2409_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n2410_));
  AOI21_X1   g02218(.A1(new_n2410_), .A2(new_n2408_), .B(new_n2399_), .ZN(new_n2411_));
  AOI21_X1   g02219(.A1(new_n2408_), .A2(new_n2389_), .B(new_n630_), .ZN(new_n2412_));
  OAI21_X1   g02220(.A1(new_n2411_), .A2(new_n2412_), .B(\asqrt[56] ), .ZN(new_n2413_));
  AOI21_X1   g02221(.A1(new_n2395_), .A2(new_n2413_), .B(new_n450_), .ZN(new_n2414_));
  NOR2_X1    g02222(.A1(new_n2398_), .A2(new_n2414_), .ZN(new_n2415_));
  AOI21_X1   g02223(.A1(new_n2415_), .A2(new_n403_), .B(new_n2288_), .ZN(new_n2416_));
  OAI21_X1   g02224(.A1(new_n2398_), .A2(new_n2414_), .B(\asqrt[58] ), .ZN(new_n2417_));
  NAND2_X1   g02225(.A1(new_n2417_), .A2(new_n339_), .ZN(new_n2418_));
  OAI21_X1   g02226(.A1(new_n2416_), .A2(new_n2418_), .B(new_n2284_), .ZN(new_n2419_));
  INV_X1     g02227(.I(new_n2417_), .ZN(new_n2420_));
  OAI21_X1   g02228(.A1(new_n2416_), .A2(new_n2420_), .B(\asqrt[59] ), .ZN(new_n2421_));
  NAND3_X1   g02229(.A1(new_n2419_), .A2(new_n2421_), .A3(new_n288_), .ZN(new_n2422_));
  NAND2_X1   g02230(.A1(new_n2422_), .A2(new_n2282_), .ZN(new_n2423_));
  INV_X1     g02231(.I(new_n2284_), .ZN(new_n2424_));
  INV_X1     g02232(.I(new_n2294_), .ZN(new_n2425_));
  NOR2_X1    g02233(.A1(new_n2411_), .A2(new_n2412_), .ZN(new_n2426_));
  AOI21_X1   g02234(.A1(new_n2426_), .A2(new_n545_), .B(new_n2425_), .ZN(new_n2427_));
  NAND2_X1   g02235(.A1(new_n2413_), .A2(new_n450_), .ZN(new_n2428_));
  OAI21_X1   g02236(.A1(new_n2427_), .A2(new_n2428_), .B(new_n2290_), .ZN(new_n2429_));
  INV_X1     g02237(.I(new_n2413_), .ZN(new_n2430_));
  OAI21_X1   g02238(.A1(new_n2427_), .A2(new_n2430_), .B(\asqrt[57] ), .ZN(new_n2431_));
  NAND3_X1   g02239(.A1(new_n2429_), .A2(new_n2431_), .A3(new_n403_), .ZN(new_n2432_));
  NAND2_X1   g02240(.A1(new_n2432_), .A2(new_n2287_), .ZN(new_n2433_));
  NAND2_X1   g02241(.A1(new_n2429_), .A2(new_n2431_), .ZN(new_n2434_));
  AOI21_X1   g02242(.A1(new_n2434_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n2435_));
  AOI21_X1   g02243(.A1(new_n2435_), .A2(new_n2433_), .B(new_n2424_), .ZN(new_n2436_));
  AOI21_X1   g02244(.A1(new_n2433_), .A2(new_n2417_), .B(new_n339_), .ZN(new_n2437_));
  OAI21_X1   g02245(.A1(new_n2436_), .A2(new_n2437_), .B(\asqrt[60] ), .ZN(new_n2438_));
  AOI21_X1   g02246(.A1(new_n2423_), .A2(new_n2438_), .B(new_n242_), .ZN(new_n2439_));
  NAND3_X1   g02247(.A1(\asqrt[44] ), .A2(new_n2214_), .A3(new_n2230_), .ZN(new_n2440_));
  XOR2_X1    g02248(.A1(new_n2440_), .A2(new_n2255_), .Z(new_n2441_));
  INV_X1     g02249(.I(new_n2441_), .ZN(new_n2442_));
  NAND2_X1   g02250(.A1(new_n2419_), .A2(new_n2421_), .ZN(new_n2443_));
  AOI21_X1   g02251(.A1(new_n2443_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n2444_));
  AOI21_X1   g02252(.A1(new_n2444_), .A2(new_n2423_), .B(new_n2442_), .ZN(new_n2445_));
  OAI21_X1   g02253(.A1(new_n2445_), .A2(new_n2439_), .B(\asqrt[62] ), .ZN(new_n2446_));
  AOI21_X1   g02254(.A1(new_n2215_), .A2(new_n2236_), .B(new_n2231_), .ZN(new_n2447_));
  NAND2_X1   g02255(.A1(\asqrt[44] ), .A2(new_n2447_), .ZN(new_n2448_));
  XOR2_X1    g02256(.A1(new_n2448_), .A2(new_n2234_), .Z(new_n2449_));
  INV_X1     g02257(.I(new_n2282_), .ZN(new_n2450_));
  NOR2_X1    g02258(.A1(new_n2436_), .A2(new_n2437_), .ZN(new_n2451_));
  AOI21_X1   g02259(.A1(new_n2451_), .A2(new_n288_), .B(new_n2450_), .ZN(new_n2452_));
  INV_X1     g02260(.I(new_n2438_), .ZN(new_n2453_));
  OAI21_X1   g02261(.A1(new_n2452_), .A2(new_n2453_), .B(\asqrt[61] ), .ZN(new_n2454_));
  NAND2_X1   g02262(.A1(new_n2438_), .A2(new_n242_), .ZN(new_n2455_));
  OAI21_X1   g02263(.A1(new_n2452_), .A2(new_n2455_), .B(new_n2441_), .ZN(new_n2456_));
  NAND3_X1   g02264(.A1(new_n2456_), .A2(new_n2454_), .A3(new_n234_), .ZN(new_n2457_));
  NAND2_X1   g02265(.A1(new_n2457_), .A2(new_n2449_), .ZN(new_n2458_));
  AOI21_X1   g02266(.A1(new_n2458_), .A2(new_n2446_), .B(new_n2279_), .ZN(new_n2459_));
  AOI21_X1   g02267(.A1(new_n2459_), .A2(new_n2277_), .B(\asqrt[63] ), .ZN(new_n2460_));
  NAND2_X1   g02268(.A1(new_n2458_), .A2(new_n2446_), .ZN(new_n2461_));
  NOR2_X1    g02269(.A1(new_n2461_), .A2(new_n2277_), .ZN(new_n2462_));
  NOR2_X1    g02270(.A1(\asqrt[44] ), .A2(new_n2266_), .ZN(new_n2463_));
  NOR4_X1    g02271(.A1(new_n2460_), .A2(new_n2274_), .A3(new_n2462_), .A4(new_n2463_), .ZN(new_n2464_));
  OAI21_X1   g02272(.A1(new_n2402_), .A2(new_n2403_), .B(new_n2406_), .ZN(new_n2465_));
  NOR2_X1    g02273(.A1(new_n2464_), .A2(new_n2465_), .ZN(new_n2466_));
  XOR2_X1    g02274(.A1(new_n2466_), .A2(new_n2254_), .Z(new_n2467_));
  INV_X1     g02275(.I(new_n2467_), .ZN(new_n2468_));
  INV_X1     g02276(.I(new_n2274_), .ZN(new_n2469_));
  INV_X1     g02277(.I(new_n2446_), .ZN(new_n2470_));
  NOR2_X1    g02278(.A1(new_n2445_), .A2(new_n2439_), .ZN(new_n2471_));
  INV_X1     g02279(.I(new_n2449_), .ZN(new_n2472_));
  AOI21_X1   g02280(.A1(new_n2471_), .A2(new_n234_), .B(new_n2472_), .ZN(new_n2473_));
  OAI21_X1   g02281(.A1(new_n2473_), .A2(new_n2470_), .B(new_n2278_), .ZN(new_n2474_));
  OAI21_X1   g02282(.A1(new_n2474_), .A2(new_n2276_), .B(new_n193_), .ZN(new_n2475_));
  NOR2_X1    g02283(.A1(new_n2473_), .A2(new_n2470_), .ZN(new_n2476_));
  NAND2_X1   g02284(.A1(new_n2476_), .A2(new_n2276_), .ZN(new_n2477_));
  INV_X1     g02285(.I(new_n2463_), .ZN(new_n2478_));
  NAND4_X1   g02286(.A1(new_n2475_), .A2(new_n2469_), .A3(new_n2477_), .A4(new_n2478_), .ZN(\asqrt[43] ));
  NAND3_X1   g02287(.A1(\asqrt[43] ), .A2(new_n2353_), .A3(new_n2385_), .ZN(new_n2480_));
  XOR2_X1    g02288(.A1(new_n2480_), .A2(new_n2400_), .Z(new_n2481_));
  OAI21_X1   g02289(.A1(new_n2347_), .A2(new_n2349_), .B(new_n2352_), .ZN(new_n2482_));
  NOR2_X1    g02290(.A1(new_n2464_), .A2(new_n2482_), .ZN(new_n2483_));
  XOR2_X1    g02291(.A1(new_n2483_), .A2(new_n2306_), .Z(new_n2484_));
  INV_X1     g02292(.I(new_n2484_), .ZN(new_n2485_));
  NAND3_X1   g02293(.A1(\asqrt[43] ), .A2(new_n2379_), .A3(new_n2348_), .ZN(new_n2486_));
  XOR2_X1    g02294(.A1(new_n2486_), .A2(new_n2310_), .Z(new_n2487_));
  INV_X1     g02295(.I(new_n2487_), .ZN(new_n2488_));
  AOI21_X1   g02296(.A1(new_n2341_), .A2(new_n2342_), .B(new_n2345_), .ZN(new_n2489_));
  NAND2_X1   g02297(.A1(\asqrt[43] ), .A2(new_n2489_), .ZN(new_n2490_));
  XOR2_X1    g02298(.A1(new_n2490_), .A2(new_n2313_), .Z(new_n2491_));
  NOR2_X1    g02299(.A1(new_n2340_), .A2(\asqrt[48] ), .ZN(new_n2492_));
  NOR3_X1    g02300(.A1(new_n2464_), .A2(new_n2492_), .A3(new_n2377_), .ZN(new_n2493_));
  XOR2_X1    g02301(.A1(new_n2493_), .A2(new_n2316_), .Z(new_n2494_));
  NOR3_X1    g02302(.A1(new_n2464_), .A2(new_n2335_), .A3(new_n2372_), .ZN(new_n2495_));
  XOR2_X1    g02303(.A1(new_n2495_), .A2(new_n2337_), .Z(new_n2496_));
  INV_X1     g02304(.I(new_n2496_), .ZN(new_n2497_));
  NOR2_X1    g02305(.A1(new_n2368_), .A2(\asqrt[46] ), .ZN(new_n2498_));
  NOR3_X1    g02306(.A1(new_n2464_), .A2(new_n2498_), .A3(new_n2334_), .ZN(new_n2499_));
  XOR2_X1    g02307(.A1(new_n2499_), .A2(new_n2362_), .Z(new_n2500_));
  INV_X1     g02308(.I(new_n2500_), .ZN(new_n2501_));
  NAND3_X1   g02309(.A1(\asqrt[43] ), .A2(new_n2324_), .A3(new_n2325_), .ZN(new_n2502_));
  NAND4_X1   g02310(.A1(new_n2475_), .A2(\asqrt[44] ), .A3(new_n2477_), .A4(new_n2469_), .ZN(new_n2503_));
  AOI21_X1   g02311(.A1(new_n2502_), .A2(new_n2503_), .B(\a[88] ), .ZN(new_n2504_));
  NOR3_X1    g02312(.A1(new_n2464_), .A2(\a[86] ), .A3(\a[87] ), .ZN(new_n2505_));
  INV_X1     g02313(.I(new_n2503_), .ZN(new_n2506_));
  NOR3_X1    g02314(.A1(new_n2505_), .A2(new_n2089_), .A3(new_n2506_), .ZN(new_n2507_));
  NOR2_X1    g02315(.A1(new_n2507_), .A2(new_n2504_), .ZN(new_n2508_));
  INV_X1     g02316(.I(\a[84] ), .ZN(new_n2509_));
  INV_X1     g02317(.I(\a[85] ), .ZN(new_n2510_));
  NAND3_X1   g02318(.A1(new_n2509_), .A2(new_n2510_), .A3(new_n2324_), .ZN(new_n2511_));
  OAI21_X1   g02319(.A1(new_n2464_), .A2(new_n2324_), .B(new_n2511_), .ZN(new_n2512_));
  NAND2_X1   g02320(.A1(new_n2512_), .A2(\asqrt[44] ), .ZN(new_n2513_));
  OAI21_X1   g02321(.A1(new_n2464_), .A2(\a[86] ), .B(\a[87] ), .ZN(new_n2514_));
  NAND2_X1   g02322(.A1(new_n2514_), .A2(new_n2502_), .ZN(new_n2515_));
  NOR2_X1    g02323(.A1(new_n2512_), .A2(\asqrt[44] ), .ZN(new_n2516_));
  OAI21_X1   g02324(.A1(new_n2515_), .A2(new_n2516_), .B(new_n2513_), .ZN(new_n2517_));
  OAI21_X1   g02325(.A1(new_n2517_), .A2(\asqrt[45] ), .B(new_n2508_), .ZN(new_n2518_));
  NAND2_X1   g02326(.A1(new_n2517_), .A2(\asqrt[45] ), .ZN(new_n2519_));
  NAND3_X1   g02327(.A1(new_n2518_), .A2(new_n1884_), .A3(new_n2519_), .ZN(new_n2520_));
  NOR3_X1    g02328(.A1(new_n2464_), .A2(new_n2328_), .A3(new_n2367_), .ZN(new_n2521_));
  XOR2_X1    g02329(.A1(new_n2521_), .A2(new_n2330_), .Z(new_n2522_));
  NAND2_X1   g02330(.A1(new_n2520_), .A2(new_n2522_), .ZN(new_n2523_));
  NAND2_X1   g02331(.A1(new_n2518_), .A2(new_n2519_), .ZN(new_n2524_));
  AOI21_X1   g02332(.A1(new_n2524_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n2525_));
  AOI21_X1   g02333(.A1(new_n2525_), .A2(new_n2523_), .B(new_n2501_), .ZN(new_n2526_));
  OAI21_X1   g02334(.A1(new_n2505_), .A2(new_n2506_), .B(new_n2089_), .ZN(new_n2527_));
  NAND3_X1   g02335(.A1(new_n2502_), .A2(\a[88] ), .A3(new_n2503_), .ZN(new_n2528_));
  NAND2_X1   g02336(.A1(new_n2527_), .A2(new_n2528_), .ZN(new_n2529_));
  NAND2_X1   g02337(.A1(\asqrt[43] ), .A2(\a[86] ), .ZN(new_n2530_));
  AOI21_X1   g02338(.A1(new_n2530_), .A2(new_n2511_), .B(new_n2271_), .ZN(new_n2531_));
  AOI21_X1   g02339(.A1(\asqrt[43] ), .A2(new_n2324_), .B(new_n2325_), .ZN(new_n2532_));
  NOR2_X1    g02340(.A1(new_n2505_), .A2(new_n2532_), .ZN(new_n2533_));
  NAND3_X1   g02341(.A1(new_n2530_), .A2(new_n2271_), .A3(new_n2511_), .ZN(new_n2534_));
  AOI21_X1   g02342(.A1(new_n2533_), .A2(new_n2534_), .B(new_n2531_), .ZN(new_n2535_));
  AOI21_X1   g02343(.A1(new_n2535_), .A2(new_n2072_), .B(new_n2529_), .ZN(new_n2536_));
  NOR2_X1    g02344(.A1(new_n2535_), .A2(new_n2072_), .ZN(new_n2537_));
  OAI21_X1   g02345(.A1(new_n2536_), .A2(new_n2537_), .B(\asqrt[46] ), .ZN(new_n2538_));
  AOI21_X1   g02346(.A1(new_n2523_), .A2(new_n2538_), .B(new_n1688_), .ZN(new_n2539_));
  NOR2_X1    g02347(.A1(new_n2526_), .A2(new_n2539_), .ZN(new_n2540_));
  AOI21_X1   g02348(.A1(new_n2540_), .A2(new_n1533_), .B(new_n2497_), .ZN(new_n2541_));
  OAI21_X1   g02349(.A1(new_n2526_), .A2(new_n2539_), .B(\asqrt[48] ), .ZN(new_n2542_));
  NAND2_X1   g02350(.A1(new_n2542_), .A2(new_n1368_), .ZN(new_n2543_));
  OAI21_X1   g02351(.A1(new_n2541_), .A2(new_n2543_), .B(new_n2494_), .ZN(new_n2544_));
  INV_X1     g02352(.I(new_n2542_), .ZN(new_n2545_));
  OAI21_X1   g02353(.A1(new_n2541_), .A2(new_n2545_), .B(\asqrt[49] ), .ZN(new_n2546_));
  NAND3_X1   g02354(.A1(new_n2544_), .A2(new_n2546_), .A3(new_n1228_), .ZN(new_n2547_));
  NAND2_X1   g02355(.A1(new_n2547_), .A2(new_n2491_), .ZN(new_n2548_));
  NAND2_X1   g02356(.A1(new_n2544_), .A2(new_n2546_), .ZN(new_n2549_));
  AOI21_X1   g02357(.A1(new_n2549_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n2550_));
  AOI21_X1   g02358(.A1(new_n2550_), .A2(new_n2548_), .B(new_n2488_), .ZN(new_n2551_));
  INV_X1     g02359(.I(new_n2494_), .ZN(new_n2552_));
  NOR2_X1    g02360(.A1(new_n2536_), .A2(new_n2537_), .ZN(new_n2553_));
  INV_X1     g02361(.I(new_n2522_), .ZN(new_n2554_));
  AOI21_X1   g02362(.A1(new_n2553_), .A2(new_n1884_), .B(new_n2554_), .ZN(new_n2555_));
  NAND2_X1   g02363(.A1(new_n2538_), .A2(new_n1688_), .ZN(new_n2556_));
  OAI21_X1   g02364(.A1(new_n2555_), .A2(new_n2556_), .B(new_n2500_), .ZN(new_n2557_));
  INV_X1     g02365(.I(new_n2538_), .ZN(new_n2558_));
  OAI21_X1   g02366(.A1(new_n2555_), .A2(new_n2558_), .B(\asqrt[47] ), .ZN(new_n2559_));
  NAND3_X1   g02367(.A1(new_n2557_), .A2(new_n2559_), .A3(new_n1533_), .ZN(new_n2560_));
  NAND2_X1   g02368(.A1(new_n2560_), .A2(new_n2496_), .ZN(new_n2561_));
  NAND2_X1   g02369(.A1(new_n2557_), .A2(new_n2559_), .ZN(new_n2562_));
  AOI21_X1   g02370(.A1(new_n2562_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n2563_));
  AOI21_X1   g02371(.A1(new_n2563_), .A2(new_n2561_), .B(new_n2552_), .ZN(new_n2564_));
  AOI21_X1   g02372(.A1(new_n2561_), .A2(new_n2542_), .B(new_n1368_), .ZN(new_n2565_));
  OAI21_X1   g02373(.A1(new_n2564_), .A2(new_n2565_), .B(\asqrt[50] ), .ZN(new_n2566_));
  AOI21_X1   g02374(.A1(new_n2548_), .A2(new_n2566_), .B(new_n1088_), .ZN(new_n2567_));
  NOR2_X1    g02375(.A1(new_n2551_), .A2(new_n2567_), .ZN(new_n2568_));
  AOI21_X1   g02376(.A1(new_n2568_), .A2(new_n962_), .B(new_n2485_), .ZN(new_n2569_));
  OAI21_X1   g02377(.A1(new_n2551_), .A2(new_n2567_), .B(\asqrt[52] ), .ZN(new_n2570_));
  NAND2_X1   g02378(.A1(new_n2570_), .A2(new_n842_), .ZN(new_n2571_));
  OAI21_X1   g02379(.A1(new_n2569_), .A2(new_n2571_), .B(new_n2481_), .ZN(new_n2572_));
  INV_X1     g02380(.I(new_n2570_), .ZN(new_n2573_));
  OAI21_X1   g02381(.A1(new_n2569_), .A2(new_n2573_), .B(\asqrt[53] ), .ZN(new_n2574_));
  NAND3_X1   g02382(.A1(new_n2572_), .A2(new_n2574_), .A3(new_n720_), .ZN(new_n2575_));
  INV_X1     g02383(.I(new_n2481_), .ZN(new_n2576_));
  INV_X1     g02384(.I(new_n2491_), .ZN(new_n2577_));
  NOR2_X1    g02385(.A1(new_n2564_), .A2(new_n2565_), .ZN(new_n2578_));
  AOI21_X1   g02386(.A1(new_n2578_), .A2(new_n1228_), .B(new_n2577_), .ZN(new_n2579_));
  NAND2_X1   g02387(.A1(new_n2566_), .A2(new_n1088_), .ZN(new_n2580_));
  OAI21_X1   g02388(.A1(new_n2579_), .A2(new_n2580_), .B(new_n2487_), .ZN(new_n2581_));
  INV_X1     g02389(.I(new_n2566_), .ZN(new_n2582_));
  OAI21_X1   g02390(.A1(new_n2579_), .A2(new_n2582_), .B(\asqrt[51] ), .ZN(new_n2583_));
  NAND3_X1   g02391(.A1(new_n2581_), .A2(new_n2583_), .A3(new_n962_), .ZN(new_n2584_));
  NAND2_X1   g02392(.A1(new_n2584_), .A2(new_n2484_), .ZN(new_n2585_));
  NAND2_X1   g02393(.A1(new_n2581_), .A2(new_n2583_), .ZN(new_n2586_));
  AOI21_X1   g02394(.A1(new_n2586_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n2587_));
  AOI21_X1   g02395(.A1(new_n2587_), .A2(new_n2585_), .B(new_n2576_), .ZN(new_n2588_));
  AOI21_X1   g02396(.A1(new_n2585_), .A2(new_n2570_), .B(new_n842_), .ZN(new_n2589_));
  OAI21_X1   g02397(.A1(new_n2588_), .A2(new_n2589_), .B(\asqrt[54] ), .ZN(new_n2590_));
  NAND2_X1   g02398(.A1(new_n2461_), .A2(new_n2276_), .ZN(new_n2591_));
  NOR2_X1    g02399(.A1(new_n2464_), .A2(new_n2276_), .ZN(new_n2592_));
  NAND2_X1   g02400(.A1(new_n2592_), .A2(new_n2476_), .ZN(new_n2593_));
  AOI21_X1   g02401(.A1(new_n2593_), .A2(new_n2591_), .B(new_n193_), .ZN(new_n2594_));
  INV_X1     g02402(.I(new_n2594_), .ZN(new_n2595_));
  NAND3_X1   g02403(.A1(\asqrt[43] ), .A2(new_n2446_), .A3(new_n2457_), .ZN(new_n2596_));
  XOR2_X1    g02404(.A1(new_n2596_), .A2(new_n2449_), .Z(new_n2597_));
  AOI21_X1   g02405(.A1(new_n2592_), .A2(new_n2461_), .B(new_n2462_), .ZN(new_n2598_));
  OAI21_X1   g02406(.A1(new_n2416_), .A2(new_n2418_), .B(new_n2421_), .ZN(new_n2599_));
  NOR2_X1    g02407(.A1(new_n2464_), .A2(new_n2599_), .ZN(new_n2600_));
  XOR2_X1    g02408(.A1(new_n2600_), .A2(new_n2284_), .Z(new_n2601_));
  NAND3_X1   g02409(.A1(\asqrt[43] ), .A2(new_n2432_), .A3(new_n2417_), .ZN(new_n2602_));
  XOR2_X1    g02410(.A1(new_n2602_), .A2(new_n2288_), .Z(new_n2603_));
  OAI21_X1   g02411(.A1(new_n2427_), .A2(new_n2428_), .B(new_n2431_), .ZN(new_n2604_));
  NOR2_X1    g02412(.A1(new_n2464_), .A2(new_n2604_), .ZN(new_n2605_));
  XOR2_X1    g02413(.A1(new_n2605_), .A2(new_n2290_), .Z(new_n2606_));
  INV_X1     g02414(.I(new_n2606_), .ZN(new_n2607_));
  NAND3_X1   g02415(.A1(\asqrt[43] ), .A2(new_n2394_), .A3(new_n2413_), .ZN(new_n2608_));
  XOR2_X1    g02416(.A1(new_n2608_), .A2(new_n2425_), .Z(new_n2609_));
  INV_X1     g02417(.I(new_n2609_), .ZN(new_n2610_));
  OAI21_X1   g02418(.A1(new_n2388_), .A2(new_n2390_), .B(new_n2393_), .ZN(new_n2611_));
  NOR2_X1    g02419(.A1(new_n2464_), .A2(new_n2611_), .ZN(new_n2612_));
  XOR2_X1    g02420(.A1(new_n2612_), .A2(new_n2296_), .Z(new_n2613_));
  NAND3_X1   g02421(.A1(\asqrt[43] ), .A2(new_n2407_), .A3(new_n2389_), .ZN(new_n2614_));
  XOR2_X1    g02422(.A1(new_n2614_), .A2(new_n2300_), .Z(new_n2615_));
  NOR2_X1    g02423(.A1(new_n2588_), .A2(new_n2589_), .ZN(new_n2616_));
  AOI21_X1   g02424(.A1(new_n2616_), .A2(new_n720_), .B(new_n2468_), .ZN(new_n2617_));
  NAND2_X1   g02425(.A1(new_n2590_), .A2(new_n630_), .ZN(new_n2618_));
  OAI21_X1   g02426(.A1(new_n2617_), .A2(new_n2618_), .B(new_n2615_), .ZN(new_n2619_));
  INV_X1     g02427(.I(new_n2590_), .ZN(new_n2620_));
  OAI21_X1   g02428(.A1(new_n2617_), .A2(new_n2620_), .B(\asqrt[55] ), .ZN(new_n2621_));
  NAND3_X1   g02429(.A1(new_n2619_), .A2(new_n2621_), .A3(new_n545_), .ZN(new_n2622_));
  NAND2_X1   g02430(.A1(new_n2622_), .A2(new_n2613_), .ZN(new_n2623_));
  NAND2_X1   g02431(.A1(new_n2619_), .A2(new_n2621_), .ZN(new_n2624_));
  AOI21_X1   g02432(.A1(new_n2624_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n2625_));
  AOI21_X1   g02433(.A1(new_n2625_), .A2(new_n2623_), .B(new_n2610_), .ZN(new_n2626_));
  INV_X1     g02434(.I(new_n2615_), .ZN(new_n2627_));
  NAND2_X1   g02435(.A1(new_n2575_), .A2(new_n2467_), .ZN(new_n2628_));
  NAND2_X1   g02436(.A1(new_n2572_), .A2(new_n2574_), .ZN(new_n2629_));
  AOI21_X1   g02437(.A1(new_n2629_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n2630_));
  AOI21_X1   g02438(.A1(new_n2630_), .A2(new_n2628_), .B(new_n2627_), .ZN(new_n2631_));
  AOI21_X1   g02439(.A1(new_n2628_), .A2(new_n2590_), .B(new_n630_), .ZN(new_n2632_));
  OAI21_X1   g02440(.A1(new_n2631_), .A2(new_n2632_), .B(\asqrt[56] ), .ZN(new_n2633_));
  AOI21_X1   g02441(.A1(new_n2623_), .A2(new_n2633_), .B(new_n450_), .ZN(new_n2634_));
  NOR2_X1    g02442(.A1(new_n2626_), .A2(new_n2634_), .ZN(new_n2635_));
  AOI21_X1   g02443(.A1(new_n2635_), .A2(new_n403_), .B(new_n2607_), .ZN(new_n2636_));
  OAI21_X1   g02444(.A1(new_n2626_), .A2(new_n2634_), .B(\asqrt[58] ), .ZN(new_n2637_));
  NAND2_X1   g02445(.A1(new_n2637_), .A2(new_n339_), .ZN(new_n2638_));
  OAI21_X1   g02446(.A1(new_n2636_), .A2(new_n2638_), .B(new_n2603_), .ZN(new_n2639_));
  INV_X1     g02447(.I(new_n2637_), .ZN(new_n2640_));
  OAI21_X1   g02448(.A1(new_n2636_), .A2(new_n2640_), .B(\asqrt[59] ), .ZN(new_n2641_));
  NAND3_X1   g02449(.A1(new_n2639_), .A2(new_n2641_), .A3(new_n288_), .ZN(new_n2642_));
  NAND2_X1   g02450(.A1(new_n2642_), .A2(new_n2601_), .ZN(new_n2643_));
  INV_X1     g02451(.I(new_n2603_), .ZN(new_n2644_));
  INV_X1     g02452(.I(new_n2613_), .ZN(new_n2645_));
  NOR2_X1    g02453(.A1(new_n2631_), .A2(new_n2632_), .ZN(new_n2646_));
  AOI21_X1   g02454(.A1(new_n2646_), .A2(new_n545_), .B(new_n2645_), .ZN(new_n2647_));
  NAND2_X1   g02455(.A1(new_n2633_), .A2(new_n450_), .ZN(new_n2648_));
  OAI21_X1   g02456(.A1(new_n2647_), .A2(new_n2648_), .B(new_n2609_), .ZN(new_n2649_));
  INV_X1     g02457(.I(new_n2633_), .ZN(new_n2650_));
  OAI21_X1   g02458(.A1(new_n2647_), .A2(new_n2650_), .B(\asqrt[57] ), .ZN(new_n2651_));
  NAND3_X1   g02459(.A1(new_n2649_), .A2(new_n2651_), .A3(new_n403_), .ZN(new_n2652_));
  NAND2_X1   g02460(.A1(new_n2652_), .A2(new_n2606_), .ZN(new_n2653_));
  NAND2_X1   g02461(.A1(new_n2649_), .A2(new_n2651_), .ZN(new_n2654_));
  AOI21_X1   g02462(.A1(new_n2654_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n2655_));
  AOI21_X1   g02463(.A1(new_n2655_), .A2(new_n2653_), .B(new_n2644_), .ZN(new_n2656_));
  AOI21_X1   g02464(.A1(new_n2653_), .A2(new_n2637_), .B(new_n339_), .ZN(new_n2657_));
  OAI21_X1   g02465(.A1(new_n2656_), .A2(new_n2657_), .B(\asqrt[60] ), .ZN(new_n2658_));
  AOI21_X1   g02466(.A1(new_n2643_), .A2(new_n2658_), .B(new_n242_), .ZN(new_n2659_));
  NAND3_X1   g02467(.A1(\asqrt[43] ), .A2(new_n2422_), .A3(new_n2438_), .ZN(new_n2660_));
  XOR2_X1    g02468(.A1(new_n2660_), .A2(new_n2450_), .Z(new_n2661_));
  INV_X1     g02469(.I(new_n2661_), .ZN(new_n2662_));
  NAND2_X1   g02470(.A1(new_n2639_), .A2(new_n2641_), .ZN(new_n2663_));
  AOI21_X1   g02471(.A1(new_n2663_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n2664_));
  AOI21_X1   g02472(.A1(new_n2664_), .A2(new_n2643_), .B(new_n2662_), .ZN(new_n2665_));
  OAI21_X1   g02473(.A1(new_n2665_), .A2(new_n2659_), .B(\asqrt[62] ), .ZN(new_n2666_));
  INV_X1     g02474(.I(new_n2666_), .ZN(new_n2667_));
  NOR2_X1    g02475(.A1(new_n2665_), .A2(new_n2659_), .ZN(new_n2668_));
  AOI21_X1   g02476(.A1(new_n2423_), .A2(new_n2444_), .B(new_n2439_), .ZN(new_n2669_));
  NAND2_X1   g02477(.A1(\asqrt[43] ), .A2(new_n2669_), .ZN(new_n2670_));
  XOR2_X1    g02478(.A1(new_n2670_), .A2(new_n2442_), .Z(new_n2671_));
  INV_X1     g02479(.I(new_n2671_), .ZN(new_n2672_));
  AOI21_X1   g02480(.A1(new_n2668_), .A2(new_n234_), .B(new_n2672_), .ZN(new_n2673_));
  OAI21_X1   g02481(.A1(new_n2673_), .A2(new_n2667_), .B(new_n2598_), .ZN(new_n2674_));
  OAI21_X1   g02482(.A1(new_n2674_), .A2(new_n2597_), .B(new_n193_), .ZN(new_n2675_));
  NOR2_X1    g02483(.A1(new_n2673_), .A2(new_n2667_), .ZN(new_n2676_));
  NAND2_X1   g02484(.A1(new_n2676_), .A2(new_n2597_), .ZN(new_n2677_));
  NOR2_X1    g02485(.A1(\asqrt[43] ), .A2(new_n2277_), .ZN(new_n2678_));
  INV_X1     g02486(.I(new_n2678_), .ZN(new_n2679_));
  NAND4_X1   g02487(.A1(new_n2675_), .A2(new_n2595_), .A3(new_n2677_), .A4(new_n2679_), .ZN(\asqrt[42] ));
  NAND3_X1   g02488(.A1(\asqrt[42] ), .A2(new_n2575_), .A3(new_n2590_), .ZN(new_n2681_));
  XOR2_X1    g02489(.A1(new_n2681_), .A2(new_n2468_), .Z(new_n2682_));
  INV_X1     g02490(.I(new_n2601_), .ZN(new_n2683_));
  NOR2_X1    g02491(.A1(new_n2656_), .A2(new_n2657_), .ZN(new_n2684_));
  AOI21_X1   g02492(.A1(new_n2684_), .A2(new_n288_), .B(new_n2683_), .ZN(new_n2685_));
  INV_X1     g02493(.I(new_n2658_), .ZN(new_n2686_));
  OAI21_X1   g02494(.A1(new_n2685_), .A2(new_n2686_), .B(\asqrt[61] ), .ZN(new_n2687_));
  NAND2_X1   g02495(.A1(new_n2658_), .A2(new_n242_), .ZN(new_n2688_));
  OAI21_X1   g02496(.A1(new_n2685_), .A2(new_n2688_), .B(new_n2661_), .ZN(new_n2689_));
  NAND3_X1   g02497(.A1(new_n2689_), .A2(new_n2687_), .A3(new_n234_), .ZN(new_n2690_));
  NAND2_X1   g02498(.A1(new_n2690_), .A2(new_n2671_), .ZN(new_n2691_));
  NAND2_X1   g02499(.A1(new_n2691_), .A2(new_n2666_), .ZN(new_n2692_));
  NAND2_X1   g02500(.A1(new_n2692_), .A2(new_n2597_), .ZN(new_n2693_));
  INV_X1     g02501(.I(new_n2597_), .ZN(new_n2694_));
  INV_X1     g02502(.I(new_n2598_), .ZN(new_n2695_));
  AOI21_X1   g02503(.A1(new_n2691_), .A2(new_n2666_), .B(new_n2695_), .ZN(new_n2696_));
  AOI21_X1   g02504(.A1(new_n2696_), .A2(new_n2694_), .B(\asqrt[63] ), .ZN(new_n2697_));
  NOR2_X1    g02505(.A1(new_n2692_), .A2(new_n2694_), .ZN(new_n2698_));
  NOR4_X1    g02506(.A1(new_n2697_), .A2(new_n2594_), .A3(new_n2698_), .A4(new_n2678_), .ZN(new_n2699_));
  NOR2_X1    g02507(.A1(new_n2699_), .A2(new_n2597_), .ZN(new_n2700_));
  NAND2_X1   g02508(.A1(new_n2700_), .A2(new_n2676_), .ZN(new_n2701_));
  AOI21_X1   g02509(.A1(new_n2701_), .A2(new_n2693_), .B(new_n193_), .ZN(new_n2702_));
  NAND3_X1   g02510(.A1(\asqrt[42] ), .A2(new_n2666_), .A3(new_n2690_), .ZN(new_n2703_));
  XOR2_X1    g02511(.A1(new_n2703_), .A2(new_n2671_), .Z(new_n2704_));
  INV_X1     g02512(.I(new_n2704_), .ZN(new_n2705_));
  AOI21_X1   g02513(.A1(new_n2700_), .A2(new_n2692_), .B(new_n2698_), .ZN(new_n2706_));
  INV_X1     g02514(.I(new_n2706_), .ZN(new_n2707_));
  OAI21_X1   g02515(.A1(new_n2636_), .A2(new_n2638_), .B(new_n2641_), .ZN(new_n2708_));
  NOR2_X1    g02516(.A1(new_n2699_), .A2(new_n2708_), .ZN(new_n2709_));
  XOR2_X1    g02517(.A1(new_n2709_), .A2(new_n2603_), .Z(new_n2710_));
  NAND3_X1   g02518(.A1(\asqrt[42] ), .A2(new_n2652_), .A3(new_n2637_), .ZN(new_n2711_));
  XOR2_X1    g02519(.A1(new_n2711_), .A2(new_n2607_), .Z(new_n2712_));
  OAI21_X1   g02520(.A1(new_n2647_), .A2(new_n2648_), .B(new_n2651_), .ZN(new_n2713_));
  NOR2_X1    g02521(.A1(new_n2699_), .A2(new_n2713_), .ZN(new_n2714_));
  XOR2_X1    g02522(.A1(new_n2714_), .A2(new_n2609_), .Z(new_n2715_));
  INV_X1     g02523(.I(new_n2715_), .ZN(new_n2716_));
  NAND3_X1   g02524(.A1(\asqrt[42] ), .A2(new_n2622_), .A3(new_n2633_), .ZN(new_n2717_));
  XOR2_X1    g02525(.A1(new_n2717_), .A2(new_n2645_), .Z(new_n2718_));
  INV_X1     g02526(.I(new_n2718_), .ZN(new_n2719_));
  OAI21_X1   g02527(.A1(new_n2617_), .A2(new_n2618_), .B(new_n2621_), .ZN(new_n2720_));
  NOR2_X1    g02528(.A1(new_n2699_), .A2(new_n2720_), .ZN(new_n2721_));
  XOR2_X1    g02529(.A1(new_n2721_), .A2(new_n2615_), .Z(new_n2722_));
  OAI21_X1   g02530(.A1(new_n2569_), .A2(new_n2571_), .B(new_n2574_), .ZN(new_n2723_));
  NOR2_X1    g02531(.A1(new_n2699_), .A2(new_n2723_), .ZN(new_n2724_));
  XOR2_X1    g02532(.A1(new_n2724_), .A2(new_n2481_), .Z(new_n2725_));
  INV_X1     g02533(.I(new_n2725_), .ZN(new_n2726_));
  NAND3_X1   g02534(.A1(\asqrt[42] ), .A2(new_n2584_), .A3(new_n2570_), .ZN(new_n2727_));
  XOR2_X1    g02535(.A1(new_n2727_), .A2(new_n2485_), .Z(new_n2728_));
  INV_X1     g02536(.I(new_n2728_), .ZN(new_n2729_));
  OAI21_X1   g02537(.A1(new_n2579_), .A2(new_n2580_), .B(new_n2583_), .ZN(new_n2730_));
  NOR2_X1    g02538(.A1(new_n2699_), .A2(new_n2730_), .ZN(new_n2731_));
  XOR2_X1    g02539(.A1(new_n2731_), .A2(new_n2487_), .Z(new_n2732_));
  NAND3_X1   g02540(.A1(\asqrt[42] ), .A2(new_n2547_), .A3(new_n2566_), .ZN(new_n2733_));
  XOR2_X1    g02541(.A1(new_n2733_), .A2(new_n2577_), .Z(new_n2734_));
  OAI21_X1   g02542(.A1(new_n2541_), .A2(new_n2543_), .B(new_n2546_), .ZN(new_n2735_));
  NOR2_X1    g02543(.A1(new_n2699_), .A2(new_n2735_), .ZN(new_n2736_));
  XOR2_X1    g02544(.A1(new_n2736_), .A2(new_n2494_), .Z(new_n2737_));
  INV_X1     g02545(.I(new_n2737_), .ZN(new_n2738_));
  NAND3_X1   g02546(.A1(\asqrt[42] ), .A2(new_n2560_), .A3(new_n2542_), .ZN(new_n2739_));
  XOR2_X1    g02547(.A1(new_n2739_), .A2(new_n2497_), .Z(new_n2740_));
  INV_X1     g02548(.I(new_n2740_), .ZN(new_n2741_));
  OAI21_X1   g02549(.A1(new_n2555_), .A2(new_n2556_), .B(new_n2559_), .ZN(new_n2742_));
  NOR2_X1    g02550(.A1(new_n2699_), .A2(new_n2742_), .ZN(new_n2743_));
  XOR2_X1    g02551(.A1(new_n2743_), .A2(new_n2500_), .Z(new_n2744_));
  NAND3_X1   g02552(.A1(\asqrt[42] ), .A2(new_n2520_), .A3(new_n2538_), .ZN(new_n2745_));
  XOR2_X1    g02553(.A1(new_n2745_), .A2(new_n2554_), .Z(new_n2746_));
  NOR2_X1    g02554(.A1(new_n2517_), .A2(\asqrt[45] ), .ZN(new_n2747_));
  NOR3_X1    g02555(.A1(new_n2699_), .A2(new_n2747_), .A3(new_n2537_), .ZN(new_n2748_));
  XOR2_X1    g02556(.A1(new_n2748_), .A2(new_n2508_), .Z(new_n2749_));
  INV_X1     g02557(.I(new_n2749_), .ZN(new_n2750_));
  NAND3_X1   g02558(.A1(\asqrt[42] ), .A2(new_n2509_), .A3(new_n2510_), .ZN(new_n2751_));
  NOR4_X1    g02559(.A1(new_n2697_), .A2(new_n2464_), .A3(new_n2594_), .A4(new_n2698_), .ZN(new_n2752_));
  INV_X1     g02560(.I(new_n2752_), .ZN(new_n2753_));
  AOI21_X1   g02561(.A1(new_n2751_), .A2(new_n2753_), .B(\a[86] ), .ZN(new_n2754_));
  NOR3_X1    g02562(.A1(new_n2699_), .A2(\a[84] ), .A3(\a[85] ), .ZN(new_n2755_));
  NOR3_X1    g02563(.A1(new_n2755_), .A2(new_n2324_), .A3(new_n2752_), .ZN(new_n2756_));
  NOR2_X1    g02564(.A1(new_n2756_), .A2(new_n2754_), .ZN(new_n2757_));
  INV_X1     g02565(.I(\a[82] ), .ZN(new_n2758_));
  INV_X1     g02566(.I(\a[83] ), .ZN(new_n2759_));
  NAND3_X1   g02567(.A1(new_n2758_), .A2(new_n2759_), .A3(new_n2509_), .ZN(new_n2760_));
  OAI21_X1   g02568(.A1(new_n2699_), .A2(new_n2509_), .B(new_n2760_), .ZN(new_n2761_));
  NAND2_X1   g02569(.A1(new_n2761_), .A2(\asqrt[43] ), .ZN(new_n2762_));
  OAI21_X1   g02570(.A1(new_n2699_), .A2(\a[84] ), .B(\a[85] ), .ZN(new_n2763_));
  NAND2_X1   g02571(.A1(new_n2763_), .A2(new_n2751_), .ZN(new_n2764_));
  NOR2_X1    g02572(.A1(new_n2761_), .A2(\asqrt[43] ), .ZN(new_n2765_));
  OAI21_X1   g02573(.A1(new_n2764_), .A2(new_n2765_), .B(new_n2762_), .ZN(new_n2766_));
  OAI21_X1   g02574(.A1(new_n2766_), .A2(\asqrt[44] ), .B(new_n2757_), .ZN(new_n2767_));
  NAND2_X1   g02575(.A1(new_n2766_), .A2(\asqrt[44] ), .ZN(new_n2768_));
  NAND3_X1   g02576(.A1(new_n2767_), .A2(new_n2072_), .A3(new_n2768_), .ZN(new_n2769_));
  NOR3_X1    g02577(.A1(new_n2699_), .A2(new_n2531_), .A3(new_n2516_), .ZN(new_n2770_));
  XOR2_X1    g02578(.A1(new_n2770_), .A2(new_n2533_), .Z(new_n2771_));
  AOI21_X1   g02579(.A1(new_n2767_), .A2(new_n2768_), .B(new_n2072_), .ZN(new_n2772_));
  AOI21_X1   g02580(.A1(new_n2769_), .A2(new_n2771_), .B(new_n2772_), .ZN(new_n2773_));
  AOI21_X1   g02581(.A1(new_n2773_), .A2(new_n1884_), .B(new_n2750_), .ZN(new_n2774_));
  OAI21_X1   g02582(.A1(new_n2773_), .A2(new_n1884_), .B(new_n1688_), .ZN(new_n2775_));
  OAI21_X1   g02583(.A1(new_n2774_), .A2(new_n2775_), .B(new_n2746_), .ZN(new_n2776_));
  NOR2_X1    g02584(.A1(new_n2773_), .A2(new_n1884_), .ZN(new_n2777_));
  OAI21_X1   g02585(.A1(new_n2774_), .A2(new_n2777_), .B(\asqrt[47] ), .ZN(new_n2778_));
  NAND3_X1   g02586(.A1(new_n2776_), .A2(new_n2778_), .A3(new_n1533_), .ZN(new_n2779_));
  NAND2_X1   g02587(.A1(new_n2779_), .A2(new_n2744_), .ZN(new_n2780_));
  NAND2_X1   g02588(.A1(new_n2776_), .A2(new_n2778_), .ZN(new_n2781_));
  AOI21_X1   g02589(.A1(new_n2781_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n2782_));
  AOI21_X1   g02590(.A1(new_n2782_), .A2(new_n2780_), .B(new_n2741_), .ZN(new_n2783_));
  INV_X1     g02591(.I(new_n2746_), .ZN(new_n2784_));
  OAI21_X1   g02592(.A1(new_n2755_), .A2(new_n2752_), .B(new_n2324_), .ZN(new_n2785_));
  NAND3_X1   g02593(.A1(new_n2751_), .A2(new_n2753_), .A3(\a[86] ), .ZN(new_n2786_));
  NAND2_X1   g02594(.A1(new_n2785_), .A2(new_n2786_), .ZN(new_n2787_));
  NAND2_X1   g02595(.A1(\asqrt[42] ), .A2(\a[84] ), .ZN(new_n2788_));
  AOI21_X1   g02596(.A1(new_n2788_), .A2(new_n2760_), .B(new_n2464_), .ZN(new_n2789_));
  AOI21_X1   g02597(.A1(\asqrt[42] ), .A2(new_n2509_), .B(new_n2510_), .ZN(new_n2790_));
  NOR2_X1    g02598(.A1(new_n2755_), .A2(new_n2790_), .ZN(new_n2791_));
  NAND3_X1   g02599(.A1(new_n2788_), .A2(new_n2464_), .A3(new_n2760_), .ZN(new_n2792_));
  AOI21_X1   g02600(.A1(new_n2791_), .A2(new_n2792_), .B(new_n2789_), .ZN(new_n2793_));
  AOI21_X1   g02601(.A1(new_n2793_), .A2(new_n2271_), .B(new_n2787_), .ZN(new_n2794_));
  NOR2_X1    g02602(.A1(new_n2793_), .A2(new_n2271_), .ZN(new_n2795_));
  NOR3_X1    g02603(.A1(new_n2794_), .A2(\asqrt[45] ), .A3(new_n2795_), .ZN(new_n2796_));
  INV_X1     g02604(.I(new_n2771_), .ZN(new_n2797_));
  OAI21_X1   g02605(.A1(new_n2794_), .A2(new_n2795_), .B(\asqrt[45] ), .ZN(new_n2798_));
  OAI21_X1   g02606(.A1(new_n2796_), .A2(new_n2797_), .B(new_n2798_), .ZN(new_n2799_));
  OAI21_X1   g02607(.A1(new_n2799_), .A2(\asqrt[46] ), .B(new_n2749_), .ZN(new_n2800_));
  AOI21_X1   g02608(.A1(new_n2799_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n2801_));
  AOI21_X1   g02609(.A1(new_n2801_), .A2(new_n2800_), .B(new_n2784_), .ZN(new_n2802_));
  NAND2_X1   g02610(.A1(new_n2799_), .A2(\asqrt[46] ), .ZN(new_n2803_));
  AOI21_X1   g02611(.A1(new_n2800_), .A2(new_n2803_), .B(new_n1688_), .ZN(new_n2804_));
  OAI21_X1   g02612(.A1(new_n2802_), .A2(new_n2804_), .B(\asqrt[48] ), .ZN(new_n2805_));
  AOI21_X1   g02613(.A1(new_n2780_), .A2(new_n2805_), .B(new_n1368_), .ZN(new_n2806_));
  NOR2_X1    g02614(.A1(new_n2783_), .A2(new_n2806_), .ZN(new_n2807_));
  AOI21_X1   g02615(.A1(new_n2807_), .A2(new_n1228_), .B(new_n2738_), .ZN(new_n2808_));
  OAI21_X1   g02616(.A1(new_n2783_), .A2(new_n2806_), .B(\asqrt[50] ), .ZN(new_n2809_));
  NAND2_X1   g02617(.A1(new_n2809_), .A2(new_n1088_), .ZN(new_n2810_));
  OAI21_X1   g02618(.A1(new_n2808_), .A2(new_n2810_), .B(new_n2734_), .ZN(new_n2811_));
  INV_X1     g02619(.I(new_n2809_), .ZN(new_n2812_));
  OAI21_X1   g02620(.A1(new_n2808_), .A2(new_n2812_), .B(\asqrt[51] ), .ZN(new_n2813_));
  NAND3_X1   g02621(.A1(new_n2811_), .A2(new_n2813_), .A3(new_n962_), .ZN(new_n2814_));
  NAND2_X1   g02622(.A1(new_n2814_), .A2(new_n2732_), .ZN(new_n2815_));
  NAND2_X1   g02623(.A1(new_n2811_), .A2(new_n2813_), .ZN(new_n2816_));
  AOI21_X1   g02624(.A1(new_n2816_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n2817_));
  AOI21_X1   g02625(.A1(new_n2817_), .A2(new_n2815_), .B(new_n2729_), .ZN(new_n2818_));
  INV_X1     g02626(.I(new_n2734_), .ZN(new_n2819_));
  INV_X1     g02627(.I(new_n2744_), .ZN(new_n2820_));
  NOR2_X1    g02628(.A1(new_n2802_), .A2(new_n2804_), .ZN(new_n2821_));
  AOI21_X1   g02629(.A1(new_n2821_), .A2(new_n1533_), .B(new_n2820_), .ZN(new_n2822_));
  NAND2_X1   g02630(.A1(new_n2805_), .A2(new_n1368_), .ZN(new_n2823_));
  OAI21_X1   g02631(.A1(new_n2822_), .A2(new_n2823_), .B(new_n2740_), .ZN(new_n2824_));
  INV_X1     g02632(.I(new_n2805_), .ZN(new_n2825_));
  OAI21_X1   g02633(.A1(new_n2822_), .A2(new_n2825_), .B(\asqrt[49] ), .ZN(new_n2826_));
  NAND3_X1   g02634(.A1(new_n2824_), .A2(new_n2826_), .A3(new_n1228_), .ZN(new_n2827_));
  NAND2_X1   g02635(.A1(new_n2827_), .A2(new_n2737_), .ZN(new_n2828_));
  NAND2_X1   g02636(.A1(new_n2824_), .A2(new_n2826_), .ZN(new_n2829_));
  AOI21_X1   g02637(.A1(new_n2829_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n2830_));
  AOI21_X1   g02638(.A1(new_n2830_), .A2(new_n2828_), .B(new_n2819_), .ZN(new_n2831_));
  AOI21_X1   g02639(.A1(new_n2828_), .A2(new_n2809_), .B(new_n1088_), .ZN(new_n2832_));
  OAI21_X1   g02640(.A1(new_n2831_), .A2(new_n2832_), .B(\asqrt[52] ), .ZN(new_n2833_));
  AOI21_X1   g02641(.A1(new_n2815_), .A2(new_n2833_), .B(new_n842_), .ZN(new_n2834_));
  NOR2_X1    g02642(.A1(new_n2818_), .A2(new_n2834_), .ZN(new_n2835_));
  AOI21_X1   g02643(.A1(new_n2835_), .A2(new_n720_), .B(new_n2726_), .ZN(new_n2836_));
  OAI21_X1   g02644(.A1(new_n2818_), .A2(new_n2834_), .B(\asqrt[54] ), .ZN(new_n2837_));
  NAND2_X1   g02645(.A1(new_n2837_), .A2(new_n630_), .ZN(new_n2838_));
  OAI21_X1   g02646(.A1(new_n2836_), .A2(new_n2838_), .B(new_n2682_), .ZN(new_n2839_));
  INV_X1     g02647(.I(new_n2837_), .ZN(new_n2840_));
  OAI21_X1   g02648(.A1(new_n2836_), .A2(new_n2840_), .B(\asqrt[55] ), .ZN(new_n2841_));
  NAND3_X1   g02649(.A1(new_n2839_), .A2(new_n2841_), .A3(new_n545_), .ZN(new_n2842_));
  NAND2_X1   g02650(.A1(new_n2842_), .A2(new_n2722_), .ZN(new_n2843_));
  NAND2_X1   g02651(.A1(new_n2839_), .A2(new_n2841_), .ZN(new_n2844_));
  AOI21_X1   g02652(.A1(new_n2844_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n2845_));
  AOI21_X1   g02653(.A1(new_n2845_), .A2(new_n2843_), .B(new_n2719_), .ZN(new_n2846_));
  INV_X1     g02654(.I(new_n2682_), .ZN(new_n2847_));
  INV_X1     g02655(.I(new_n2732_), .ZN(new_n2848_));
  NOR2_X1    g02656(.A1(new_n2831_), .A2(new_n2832_), .ZN(new_n2849_));
  AOI21_X1   g02657(.A1(new_n2849_), .A2(new_n962_), .B(new_n2848_), .ZN(new_n2850_));
  NAND2_X1   g02658(.A1(new_n2833_), .A2(new_n842_), .ZN(new_n2851_));
  OAI21_X1   g02659(.A1(new_n2850_), .A2(new_n2851_), .B(new_n2728_), .ZN(new_n2852_));
  INV_X1     g02660(.I(new_n2833_), .ZN(new_n2853_));
  OAI21_X1   g02661(.A1(new_n2850_), .A2(new_n2853_), .B(\asqrt[53] ), .ZN(new_n2854_));
  NAND3_X1   g02662(.A1(new_n2852_), .A2(new_n2854_), .A3(new_n720_), .ZN(new_n2855_));
  NAND2_X1   g02663(.A1(new_n2855_), .A2(new_n2725_), .ZN(new_n2856_));
  NAND2_X1   g02664(.A1(new_n2852_), .A2(new_n2854_), .ZN(new_n2857_));
  AOI21_X1   g02665(.A1(new_n2857_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n2858_));
  AOI21_X1   g02666(.A1(new_n2858_), .A2(new_n2856_), .B(new_n2847_), .ZN(new_n2859_));
  AOI21_X1   g02667(.A1(new_n2856_), .A2(new_n2837_), .B(new_n630_), .ZN(new_n2860_));
  OAI21_X1   g02668(.A1(new_n2859_), .A2(new_n2860_), .B(\asqrt[56] ), .ZN(new_n2861_));
  AOI21_X1   g02669(.A1(new_n2843_), .A2(new_n2861_), .B(new_n450_), .ZN(new_n2862_));
  NOR2_X1    g02670(.A1(new_n2846_), .A2(new_n2862_), .ZN(new_n2863_));
  AOI21_X1   g02671(.A1(new_n2863_), .A2(new_n403_), .B(new_n2716_), .ZN(new_n2864_));
  OAI21_X1   g02672(.A1(new_n2846_), .A2(new_n2862_), .B(\asqrt[58] ), .ZN(new_n2865_));
  NAND2_X1   g02673(.A1(new_n2865_), .A2(new_n339_), .ZN(new_n2866_));
  OAI21_X1   g02674(.A1(new_n2864_), .A2(new_n2866_), .B(new_n2712_), .ZN(new_n2867_));
  INV_X1     g02675(.I(new_n2865_), .ZN(new_n2868_));
  OAI21_X1   g02676(.A1(new_n2864_), .A2(new_n2868_), .B(\asqrt[59] ), .ZN(new_n2869_));
  NAND3_X1   g02677(.A1(new_n2867_), .A2(new_n2869_), .A3(new_n288_), .ZN(new_n2870_));
  NAND2_X1   g02678(.A1(new_n2870_), .A2(new_n2710_), .ZN(new_n2871_));
  INV_X1     g02679(.I(new_n2712_), .ZN(new_n2872_));
  INV_X1     g02680(.I(new_n2722_), .ZN(new_n2873_));
  NOR2_X1    g02681(.A1(new_n2859_), .A2(new_n2860_), .ZN(new_n2874_));
  AOI21_X1   g02682(.A1(new_n2874_), .A2(new_n545_), .B(new_n2873_), .ZN(new_n2875_));
  NAND2_X1   g02683(.A1(new_n2861_), .A2(new_n450_), .ZN(new_n2876_));
  OAI21_X1   g02684(.A1(new_n2875_), .A2(new_n2876_), .B(new_n2718_), .ZN(new_n2877_));
  INV_X1     g02685(.I(new_n2861_), .ZN(new_n2878_));
  OAI21_X1   g02686(.A1(new_n2875_), .A2(new_n2878_), .B(\asqrt[57] ), .ZN(new_n2879_));
  NAND3_X1   g02687(.A1(new_n2877_), .A2(new_n2879_), .A3(new_n403_), .ZN(new_n2880_));
  NAND2_X1   g02688(.A1(new_n2880_), .A2(new_n2715_), .ZN(new_n2881_));
  NAND2_X1   g02689(.A1(new_n2877_), .A2(new_n2879_), .ZN(new_n2882_));
  AOI21_X1   g02690(.A1(new_n2882_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n2883_));
  AOI21_X1   g02691(.A1(new_n2883_), .A2(new_n2881_), .B(new_n2872_), .ZN(new_n2884_));
  AOI21_X1   g02692(.A1(new_n2881_), .A2(new_n2865_), .B(new_n339_), .ZN(new_n2885_));
  OAI21_X1   g02693(.A1(new_n2884_), .A2(new_n2885_), .B(\asqrt[60] ), .ZN(new_n2886_));
  AOI21_X1   g02694(.A1(new_n2871_), .A2(new_n2886_), .B(new_n242_), .ZN(new_n2887_));
  NAND3_X1   g02695(.A1(\asqrt[42] ), .A2(new_n2642_), .A3(new_n2658_), .ZN(new_n2888_));
  XOR2_X1    g02696(.A1(new_n2888_), .A2(new_n2683_), .Z(new_n2889_));
  INV_X1     g02697(.I(new_n2889_), .ZN(new_n2890_));
  NAND2_X1   g02698(.A1(new_n2867_), .A2(new_n2869_), .ZN(new_n2891_));
  AOI21_X1   g02699(.A1(new_n2891_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n2892_));
  AOI21_X1   g02700(.A1(new_n2892_), .A2(new_n2871_), .B(new_n2890_), .ZN(new_n2893_));
  OAI21_X1   g02701(.A1(new_n2893_), .A2(new_n2887_), .B(\asqrt[62] ), .ZN(new_n2894_));
  AOI21_X1   g02702(.A1(new_n2643_), .A2(new_n2664_), .B(new_n2659_), .ZN(new_n2895_));
  NAND2_X1   g02703(.A1(\asqrt[42] ), .A2(new_n2895_), .ZN(new_n2896_));
  XOR2_X1    g02704(.A1(new_n2896_), .A2(new_n2662_), .Z(new_n2897_));
  INV_X1     g02705(.I(new_n2710_), .ZN(new_n2898_));
  NOR2_X1    g02706(.A1(new_n2884_), .A2(new_n2885_), .ZN(new_n2899_));
  AOI21_X1   g02707(.A1(new_n2899_), .A2(new_n288_), .B(new_n2898_), .ZN(new_n2900_));
  INV_X1     g02708(.I(new_n2886_), .ZN(new_n2901_));
  OAI21_X1   g02709(.A1(new_n2900_), .A2(new_n2901_), .B(\asqrt[61] ), .ZN(new_n2902_));
  NAND2_X1   g02710(.A1(new_n2886_), .A2(new_n242_), .ZN(new_n2903_));
  OAI21_X1   g02711(.A1(new_n2900_), .A2(new_n2903_), .B(new_n2889_), .ZN(new_n2904_));
  NAND3_X1   g02712(.A1(new_n2904_), .A2(new_n2902_), .A3(new_n234_), .ZN(new_n2905_));
  NAND2_X1   g02713(.A1(new_n2905_), .A2(new_n2897_), .ZN(new_n2906_));
  AOI21_X1   g02714(.A1(new_n2906_), .A2(new_n2894_), .B(new_n2707_), .ZN(new_n2907_));
  AOI21_X1   g02715(.A1(new_n2907_), .A2(new_n2705_), .B(\asqrt[63] ), .ZN(new_n2908_));
  NAND2_X1   g02716(.A1(new_n2906_), .A2(new_n2894_), .ZN(new_n2909_));
  NOR2_X1    g02717(.A1(new_n2909_), .A2(new_n2705_), .ZN(new_n2910_));
  NOR2_X1    g02718(.A1(\asqrt[42] ), .A2(new_n2694_), .ZN(new_n2911_));
  NOR4_X1    g02719(.A1(new_n2908_), .A2(new_n2702_), .A3(new_n2910_), .A4(new_n2911_), .ZN(new_n2912_));
  OAI21_X1   g02720(.A1(new_n2836_), .A2(new_n2838_), .B(new_n2841_), .ZN(new_n2913_));
  NOR2_X1    g02721(.A1(new_n2912_), .A2(new_n2913_), .ZN(new_n2914_));
  XOR2_X1    g02722(.A1(new_n2914_), .A2(new_n2682_), .Z(new_n2915_));
  INV_X1     g02723(.I(new_n2915_), .ZN(new_n2916_));
  INV_X1     g02724(.I(new_n2702_), .ZN(new_n2917_));
  INV_X1     g02725(.I(new_n2894_), .ZN(new_n2918_));
  NOR2_X1    g02726(.A1(new_n2893_), .A2(new_n2887_), .ZN(new_n2919_));
  INV_X1     g02727(.I(new_n2897_), .ZN(new_n2920_));
  AOI21_X1   g02728(.A1(new_n2919_), .A2(new_n234_), .B(new_n2920_), .ZN(new_n2921_));
  OAI21_X1   g02729(.A1(new_n2921_), .A2(new_n2918_), .B(new_n2706_), .ZN(new_n2922_));
  OAI21_X1   g02730(.A1(new_n2922_), .A2(new_n2704_), .B(new_n193_), .ZN(new_n2923_));
  NOR2_X1    g02731(.A1(new_n2921_), .A2(new_n2918_), .ZN(new_n2924_));
  NAND2_X1   g02732(.A1(new_n2924_), .A2(new_n2704_), .ZN(new_n2925_));
  INV_X1     g02733(.I(new_n2911_), .ZN(new_n2926_));
  NAND4_X1   g02734(.A1(new_n2923_), .A2(new_n2917_), .A3(new_n2925_), .A4(new_n2926_), .ZN(\asqrt[41] ));
  NAND3_X1   g02735(.A1(\asqrt[41] ), .A2(new_n2855_), .A3(new_n2837_), .ZN(new_n2928_));
  XOR2_X1    g02736(.A1(new_n2928_), .A2(new_n2726_), .Z(new_n2929_));
  OAI21_X1   g02737(.A1(new_n2850_), .A2(new_n2851_), .B(new_n2854_), .ZN(new_n2930_));
  NOR2_X1    g02738(.A1(new_n2912_), .A2(new_n2930_), .ZN(new_n2931_));
  XOR2_X1    g02739(.A1(new_n2931_), .A2(new_n2728_), .Z(new_n2932_));
  INV_X1     g02740(.I(new_n2932_), .ZN(new_n2933_));
  NAND3_X1   g02741(.A1(\asqrt[41] ), .A2(new_n2814_), .A3(new_n2833_), .ZN(new_n2934_));
  XOR2_X1    g02742(.A1(new_n2934_), .A2(new_n2848_), .Z(new_n2935_));
  INV_X1     g02743(.I(new_n2935_), .ZN(new_n2936_));
  OAI21_X1   g02744(.A1(new_n2808_), .A2(new_n2810_), .B(new_n2813_), .ZN(new_n2937_));
  NOR2_X1    g02745(.A1(new_n2912_), .A2(new_n2937_), .ZN(new_n2938_));
  XOR2_X1    g02746(.A1(new_n2938_), .A2(new_n2734_), .Z(new_n2939_));
  NAND3_X1   g02747(.A1(\asqrt[41] ), .A2(new_n2827_), .A3(new_n2809_), .ZN(new_n2940_));
  XOR2_X1    g02748(.A1(new_n2940_), .A2(new_n2738_), .Z(new_n2941_));
  OAI21_X1   g02749(.A1(new_n2822_), .A2(new_n2823_), .B(new_n2826_), .ZN(new_n2942_));
  NOR2_X1    g02750(.A1(new_n2912_), .A2(new_n2942_), .ZN(new_n2943_));
  XOR2_X1    g02751(.A1(new_n2943_), .A2(new_n2740_), .Z(new_n2944_));
  INV_X1     g02752(.I(new_n2944_), .ZN(new_n2945_));
  NAND3_X1   g02753(.A1(\asqrt[41] ), .A2(new_n2779_), .A3(new_n2805_), .ZN(new_n2946_));
  XOR2_X1    g02754(.A1(new_n2946_), .A2(new_n2820_), .Z(new_n2947_));
  INV_X1     g02755(.I(new_n2947_), .ZN(new_n2948_));
  AOI21_X1   g02756(.A1(new_n2800_), .A2(new_n2801_), .B(new_n2804_), .ZN(new_n2949_));
  NAND2_X1   g02757(.A1(\asqrt[41] ), .A2(new_n2949_), .ZN(new_n2950_));
  XOR2_X1    g02758(.A1(new_n2950_), .A2(new_n2784_), .Z(new_n2951_));
  NOR2_X1    g02759(.A1(new_n2799_), .A2(\asqrt[46] ), .ZN(new_n2952_));
  NOR3_X1    g02760(.A1(new_n2912_), .A2(new_n2952_), .A3(new_n2777_), .ZN(new_n2953_));
  XOR2_X1    g02761(.A1(new_n2953_), .A2(new_n2749_), .Z(new_n2954_));
  NOR3_X1    g02762(.A1(new_n2912_), .A2(new_n2796_), .A3(new_n2772_), .ZN(new_n2955_));
  XOR2_X1    g02763(.A1(new_n2955_), .A2(new_n2771_), .Z(new_n2956_));
  INV_X1     g02764(.I(new_n2956_), .ZN(new_n2957_));
  NOR2_X1    g02765(.A1(new_n2766_), .A2(\asqrt[44] ), .ZN(new_n2958_));
  NOR3_X1    g02766(.A1(new_n2912_), .A2(new_n2958_), .A3(new_n2795_), .ZN(new_n2959_));
  XOR2_X1    g02767(.A1(new_n2959_), .A2(new_n2757_), .Z(new_n2960_));
  INV_X1     g02768(.I(new_n2960_), .ZN(new_n2961_));
  NAND3_X1   g02769(.A1(\asqrt[41] ), .A2(new_n2758_), .A3(new_n2759_), .ZN(new_n2962_));
  NOR4_X1    g02770(.A1(new_n2908_), .A2(new_n2699_), .A3(new_n2702_), .A4(new_n2910_), .ZN(new_n2963_));
  INV_X1     g02771(.I(new_n2963_), .ZN(new_n2964_));
  AOI21_X1   g02772(.A1(new_n2962_), .A2(new_n2964_), .B(\a[84] ), .ZN(new_n2965_));
  NOR3_X1    g02773(.A1(new_n2912_), .A2(\a[82] ), .A3(\a[83] ), .ZN(new_n2966_));
  NOR3_X1    g02774(.A1(new_n2966_), .A2(new_n2509_), .A3(new_n2963_), .ZN(new_n2967_));
  NOR2_X1    g02775(.A1(new_n2967_), .A2(new_n2965_), .ZN(new_n2968_));
  INV_X1     g02776(.I(\a[80] ), .ZN(new_n2969_));
  INV_X1     g02777(.I(\a[81] ), .ZN(new_n2970_));
  NAND3_X1   g02778(.A1(new_n2969_), .A2(new_n2970_), .A3(new_n2758_), .ZN(new_n2971_));
  OAI21_X1   g02779(.A1(new_n2912_), .A2(new_n2758_), .B(new_n2971_), .ZN(new_n2972_));
  NAND2_X1   g02780(.A1(new_n2972_), .A2(\asqrt[42] ), .ZN(new_n2973_));
  OAI21_X1   g02781(.A1(new_n2912_), .A2(\a[82] ), .B(\a[83] ), .ZN(new_n2974_));
  NAND2_X1   g02782(.A1(new_n2974_), .A2(new_n2962_), .ZN(new_n2975_));
  NOR2_X1    g02783(.A1(new_n2972_), .A2(\asqrt[42] ), .ZN(new_n2976_));
  OAI21_X1   g02784(.A1(new_n2975_), .A2(new_n2976_), .B(new_n2973_), .ZN(new_n2977_));
  OAI21_X1   g02785(.A1(\asqrt[43] ), .A2(new_n2977_), .B(new_n2968_), .ZN(new_n2978_));
  NAND2_X1   g02786(.A1(new_n2977_), .A2(\asqrt[43] ), .ZN(new_n2979_));
  NAND3_X1   g02787(.A1(new_n2978_), .A2(new_n2271_), .A3(new_n2979_), .ZN(new_n2980_));
  NOR3_X1    g02788(.A1(new_n2912_), .A2(new_n2789_), .A3(new_n2765_), .ZN(new_n2981_));
  XOR2_X1    g02789(.A1(new_n2981_), .A2(new_n2791_), .Z(new_n2982_));
  NAND2_X1   g02790(.A1(new_n2980_), .A2(new_n2982_), .ZN(new_n2983_));
  NAND2_X1   g02791(.A1(new_n2978_), .A2(new_n2979_), .ZN(new_n2984_));
  AOI21_X1   g02792(.A1(new_n2984_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n2985_));
  AOI21_X1   g02793(.A1(new_n2985_), .A2(new_n2983_), .B(new_n2961_), .ZN(new_n2986_));
  OAI21_X1   g02794(.A1(new_n2966_), .A2(new_n2963_), .B(new_n2509_), .ZN(new_n2987_));
  NAND3_X1   g02795(.A1(new_n2962_), .A2(\a[84] ), .A3(new_n2964_), .ZN(new_n2988_));
  NAND2_X1   g02796(.A1(new_n2987_), .A2(new_n2988_), .ZN(new_n2989_));
  NAND2_X1   g02797(.A1(\asqrt[41] ), .A2(\a[82] ), .ZN(new_n2990_));
  AOI21_X1   g02798(.A1(new_n2990_), .A2(new_n2971_), .B(new_n2699_), .ZN(new_n2991_));
  AOI21_X1   g02799(.A1(\asqrt[41] ), .A2(new_n2758_), .B(new_n2759_), .ZN(new_n2992_));
  NOR2_X1    g02800(.A1(new_n2992_), .A2(new_n2966_), .ZN(new_n2993_));
  NAND3_X1   g02801(.A1(new_n2990_), .A2(new_n2699_), .A3(new_n2971_), .ZN(new_n2994_));
  AOI21_X1   g02802(.A1(new_n2993_), .A2(new_n2994_), .B(new_n2991_), .ZN(new_n2995_));
  AOI21_X1   g02803(.A1(new_n2995_), .A2(new_n2464_), .B(new_n2989_), .ZN(new_n2996_));
  NOR2_X1    g02804(.A1(new_n2995_), .A2(new_n2464_), .ZN(new_n2997_));
  OAI21_X1   g02805(.A1(new_n2996_), .A2(new_n2997_), .B(\asqrt[44] ), .ZN(new_n2998_));
  AOI21_X1   g02806(.A1(new_n2983_), .A2(new_n2998_), .B(new_n2072_), .ZN(new_n2999_));
  NOR2_X1    g02807(.A1(new_n2986_), .A2(new_n2999_), .ZN(new_n3000_));
  AOI21_X1   g02808(.A1(new_n3000_), .A2(new_n1884_), .B(new_n2957_), .ZN(new_n3001_));
  OAI21_X1   g02809(.A1(new_n2986_), .A2(new_n2999_), .B(\asqrt[46] ), .ZN(new_n3002_));
  NAND2_X1   g02810(.A1(new_n3002_), .A2(new_n1688_), .ZN(new_n3003_));
  OAI21_X1   g02811(.A1(new_n3001_), .A2(new_n3003_), .B(new_n2954_), .ZN(new_n3004_));
  INV_X1     g02812(.I(new_n3002_), .ZN(new_n3005_));
  OAI21_X1   g02813(.A1(new_n3001_), .A2(new_n3005_), .B(\asqrt[47] ), .ZN(new_n3006_));
  NAND3_X1   g02814(.A1(new_n3004_), .A2(new_n3006_), .A3(new_n1533_), .ZN(new_n3007_));
  NAND2_X1   g02815(.A1(new_n3007_), .A2(new_n2951_), .ZN(new_n3008_));
  NAND2_X1   g02816(.A1(new_n3004_), .A2(new_n3006_), .ZN(new_n3009_));
  AOI21_X1   g02817(.A1(new_n3009_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n3010_));
  AOI21_X1   g02818(.A1(new_n3010_), .A2(new_n3008_), .B(new_n2948_), .ZN(new_n3011_));
  INV_X1     g02819(.I(new_n2954_), .ZN(new_n3012_));
  NOR2_X1    g02820(.A1(new_n2996_), .A2(new_n2997_), .ZN(new_n3013_));
  INV_X1     g02821(.I(new_n2982_), .ZN(new_n3014_));
  AOI21_X1   g02822(.A1(new_n3013_), .A2(new_n2271_), .B(new_n3014_), .ZN(new_n3015_));
  NAND2_X1   g02823(.A1(new_n2998_), .A2(new_n2072_), .ZN(new_n3016_));
  OAI21_X1   g02824(.A1(new_n3015_), .A2(new_n3016_), .B(new_n2960_), .ZN(new_n3017_));
  INV_X1     g02825(.I(new_n2998_), .ZN(new_n3018_));
  OAI21_X1   g02826(.A1(new_n3015_), .A2(new_n3018_), .B(\asqrt[45] ), .ZN(new_n3019_));
  NAND3_X1   g02827(.A1(new_n3017_), .A2(new_n3019_), .A3(new_n1884_), .ZN(new_n3020_));
  NAND2_X1   g02828(.A1(new_n3020_), .A2(new_n2956_), .ZN(new_n3021_));
  NAND2_X1   g02829(.A1(new_n3017_), .A2(new_n3019_), .ZN(new_n3022_));
  AOI21_X1   g02830(.A1(new_n3022_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n3023_));
  AOI21_X1   g02831(.A1(new_n3023_), .A2(new_n3021_), .B(new_n3012_), .ZN(new_n3024_));
  AOI21_X1   g02832(.A1(new_n3021_), .A2(new_n3002_), .B(new_n1688_), .ZN(new_n3025_));
  OAI21_X1   g02833(.A1(new_n3024_), .A2(new_n3025_), .B(\asqrt[48] ), .ZN(new_n3026_));
  AOI21_X1   g02834(.A1(new_n3008_), .A2(new_n3026_), .B(new_n1368_), .ZN(new_n3027_));
  NOR2_X1    g02835(.A1(new_n3011_), .A2(new_n3027_), .ZN(new_n3028_));
  AOI21_X1   g02836(.A1(new_n3028_), .A2(new_n1228_), .B(new_n2945_), .ZN(new_n3029_));
  OAI21_X1   g02837(.A1(new_n3011_), .A2(new_n3027_), .B(\asqrt[50] ), .ZN(new_n3030_));
  NAND2_X1   g02838(.A1(new_n3030_), .A2(new_n1088_), .ZN(new_n3031_));
  OAI21_X1   g02839(.A1(new_n3029_), .A2(new_n3031_), .B(new_n2941_), .ZN(new_n3032_));
  INV_X1     g02840(.I(new_n3030_), .ZN(new_n3033_));
  OAI21_X1   g02841(.A1(new_n3029_), .A2(new_n3033_), .B(\asqrt[51] ), .ZN(new_n3034_));
  NAND3_X1   g02842(.A1(new_n3032_), .A2(new_n3034_), .A3(new_n962_), .ZN(new_n3035_));
  NAND2_X1   g02843(.A1(new_n3035_), .A2(new_n2939_), .ZN(new_n3036_));
  NAND2_X1   g02844(.A1(new_n3032_), .A2(new_n3034_), .ZN(new_n3037_));
  AOI21_X1   g02845(.A1(new_n3037_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n3038_));
  AOI21_X1   g02846(.A1(new_n3038_), .A2(new_n3036_), .B(new_n2936_), .ZN(new_n3039_));
  INV_X1     g02847(.I(new_n2941_), .ZN(new_n3040_));
  INV_X1     g02848(.I(new_n2951_), .ZN(new_n3041_));
  NOR2_X1    g02849(.A1(new_n3024_), .A2(new_n3025_), .ZN(new_n3042_));
  AOI21_X1   g02850(.A1(new_n3042_), .A2(new_n1533_), .B(new_n3041_), .ZN(new_n3043_));
  NAND2_X1   g02851(.A1(new_n3026_), .A2(new_n1368_), .ZN(new_n3044_));
  OAI21_X1   g02852(.A1(new_n3043_), .A2(new_n3044_), .B(new_n2947_), .ZN(new_n3045_));
  INV_X1     g02853(.I(new_n3026_), .ZN(new_n3046_));
  OAI21_X1   g02854(.A1(new_n3043_), .A2(new_n3046_), .B(\asqrt[49] ), .ZN(new_n3047_));
  NAND3_X1   g02855(.A1(new_n3045_), .A2(new_n3047_), .A3(new_n1228_), .ZN(new_n3048_));
  NAND2_X1   g02856(.A1(new_n3048_), .A2(new_n2944_), .ZN(new_n3049_));
  NAND2_X1   g02857(.A1(new_n3045_), .A2(new_n3047_), .ZN(new_n3050_));
  AOI21_X1   g02858(.A1(new_n3050_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n3051_));
  AOI21_X1   g02859(.A1(new_n3051_), .A2(new_n3049_), .B(new_n3040_), .ZN(new_n3052_));
  AOI21_X1   g02860(.A1(new_n3049_), .A2(new_n3030_), .B(new_n1088_), .ZN(new_n3053_));
  OAI21_X1   g02861(.A1(new_n3052_), .A2(new_n3053_), .B(\asqrt[52] ), .ZN(new_n3054_));
  AOI21_X1   g02862(.A1(new_n3036_), .A2(new_n3054_), .B(new_n842_), .ZN(new_n3055_));
  NOR2_X1    g02863(.A1(new_n3039_), .A2(new_n3055_), .ZN(new_n3056_));
  AOI21_X1   g02864(.A1(new_n3056_), .A2(new_n720_), .B(new_n2933_), .ZN(new_n3057_));
  OAI21_X1   g02865(.A1(new_n3039_), .A2(new_n3055_), .B(\asqrt[54] ), .ZN(new_n3058_));
  NAND2_X1   g02866(.A1(new_n3058_), .A2(new_n630_), .ZN(new_n3059_));
  OAI21_X1   g02867(.A1(new_n3057_), .A2(new_n3059_), .B(new_n2929_), .ZN(new_n3060_));
  INV_X1     g02868(.I(new_n3058_), .ZN(new_n3061_));
  OAI21_X1   g02869(.A1(new_n3057_), .A2(new_n3061_), .B(\asqrt[55] ), .ZN(new_n3062_));
  NAND3_X1   g02870(.A1(new_n3060_), .A2(new_n3062_), .A3(new_n545_), .ZN(new_n3063_));
  INV_X1     g02871(.I(new_n2929_), .ZN(new_n3064_));
  INV_X1     g02872(.I(new_n2939_), .ZN(new_n3065_));
  NOR2_X1    g02873(.A1(new_n3052_), .A2(new_n3053_), .ZN(new_n3066_));
  AOI21_X1   g02874(.A1(new_n3066_), .A2(new_n962_), .B(new_n3065_), .ZN(new_n3067_));
  NAND2_X1   g02875(.A1(new_n3054_), .A2(new_n842_), .ZN(new_n3068_));
  OAI21_X1   g02876(.A1(new_n3067_), .A2(new_n3068_), .B(new_n2935_), .ZN(new_n3069_));
  INV_X1     g02877(.I(new_n3054_), .ZN(new_n3070_));
  OAI21_X1   g02878(.A1(new_n3067_), .A2(new_n3070_), .B(\asqrt[53] ), .ZN(new_n3071_));
  NAND3_X1   g02879(.A1(new_n3069_), .A2(new_n3071_), .A3(new_n720_), .ZN(new_n3072_));
  NAND2_X1   g02880(.A1(new_n3072_), .A2(new_n2932_), .ZN(new_n3073_));
  NAND2_X1   g02881(.A1(new_n3069_), .A2(new_n3071_), .ZN(new_n3074_));
  AOI21_X1   g02882(.A1(new_n3074_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n3075_));
  AOI21_X1   g02883(.A1(new_n3075_), .A2(new_n3073_), .B(new_n3064_), .ZN(new_n3076_));
  AOI21_X1   g02884(.A1(new_n3073_), .A2(new_n3058_), .B(new_n630_), .ZN(new_n3077_));
  OAI21_X1   g02885(.A1(new_n3076_), .A2(new_n3077_), .B(\asqrt[56] ), .ZN(new_n3078_));
  NAND2_X1   g02886(.A1(new_n2909_), .A2(new_n2704_), .ZN(new_n3079_));
  NOR2_X1    g02887(.A1(new_n2912_), .A2(new_n2704_), .ZN(new_n3080_));
  NAND2_X1   g02888(.A1(new_n3080_), .A2(new_n2924_), .ZN(new_n3081_));
  AOI21_X1   g02889(.A1(new_n3081_), .A2(new_n3079_), .B(new_n193_), .ZN(new_n3082_));
  INV_X1     g02890(.I(new_n3082_), .ZN(new_n3083_));
  NAND3_X1   g02891(.A1(\asqrt[41] ), .A2(new_n2894_), .A3(new_n2905_), .ZN(new_n3084_));
  XOR2_X1    g02892(.A1(new_n3084_), .A2(new_n2897_), .Z(new_n3085_));
  AOI21_X1   g02893(.A1(new_n3080_), .A2(new_n2909_), .B(new_n2910_), .ZN(new_n3086_));
  OAI21_X1   g02894(.A1(new_n2864_), .A2(new_n2866_), .B(new_n2869_), .ZN(new_n3087_));
  NOR2_X1    g02895(.A1(new_n2912_), .A2(new_n3087_), .ZN(new_n3088_));
  XOR2_X1    g02896(.A1(new_n3088_), .A2(new_n2712_), .Z(new_n3089_));
  NAND3_X1   g02897(.A1(\asqrt[41] ), .A2(new_n2880_), .A3(new_n2865_), .ZN(new_n3090_));
  XOR2_X1    g02898(.A1(new_n3090_), .A2(new_n2716_), .Z(new_n3091_));
  OAI21_X1   g02899(.A1(new_n2875_), .A2(new_n2876_), .B(new_n2879_), .ZN(new_n3092_));
  NOR2_X1    g02900(.A1(new_n2912_), .A2(new_n3092_), .ZN(new_n3093_));
  XOR2_X1    g02901(.A1(new_n3093_), .A2(new_n2718_), .Z(new_n3094_));
  INV_X1     g02902(.I(new_n3094_), .ZN(new_n3095_));
  NAND3_X1   g02903(.A1(\asqrt[41] ), .A2(new_n2842_), .A3(new_n2861_), .ZN(new_n3096_));
  XOR2_X1    g02904(.A1(new_n3096_), .A2(new_n2873_), .Z(new_n3097_));
  INV_X1     g02905(.I(new_n3097_), .ZN(new_n3098_));
  NAND2_X1   g02906(.A1(new_n3063_), .A2(new_n2915_), .ZN(new_n3099_));
  NAND2_X1   g02907(.A1(new_n3060_), .A2(new_n3062_), .ZN(new_n3100_));
  AOI21_X1   g02908(.A1(new_n3100_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n3101_));
  AOI21_X1   g02909(.A1(new_n3101_), .A2(new_n3099_), .B(new_n3098_), .ZN(new_n3102_));
  AOI21_X1   g02910(.A1(new_n3099_), .A2(new_n3078_), .B(new_n450_), .ZN(new_n3103_));
  NOR2_X1    g02911(.A1(new_n3102_), .A2(new_n3103_), .ZN(new_n3104_));
  AOI21_X1   g02912(.A1(new_n3104_), .A2(new_n403_), .B(new_n3095_), .ZN(new_n3105_));
  OAI21_X1   g02913(.A1(new_n3102_), .A2(new_n3103_), .B(\asqrt[58] ), .ZN(new_n3106_));
  NAND2_X1   g02914(.A1(new_n3106_), .A2(new_n339_), .ZN(new_n3107_));
  OAI21_X1   g02915(.A1(new_n3105_), .A2(new_n3107_), .B(new_n3091_), .ZN(new_n3108_));
  INV_X1     g02916(.I(new_n3106_), .ZN(new_n3109_));
  OAI21_X1   g02917(.A1(new_n3105_), .A2(new_n3109_), .B(\asqrt[59] ), .ZN(new_n3110_));
  NAND3_X1   g02918(.A1(new_n3108_), .A2(new_n3110_), .A3(new_n288_), .ZN(new_n3111_));
  NAND2_X1   g02919(.A1(new_n3111_), .A2(new_n3089_), .ZN(new_n3112_));
  INV_X1     g02920(.I(new_n3091_), .ZN(new_n3113_));
  NOR2_X1    g02921(.A1(new_n3076_), .A2(new_n3077_), .ZN(new_n3114_));
  AOI21_X1   g02922(.A1(new_n3114_), .A2(new_n545_), .B(new_n2916_), .ZN(new_n3115_));
  NAND2_X1   g02923(.A1(new_n3078_), .A2(new_n450_), .ZN(new_n3116_));
  OAI21_X1   g02924(.A1(new_n3115_), .A2(new_n3116_), .B(new_n3097_), .ZN(new_n3117_));
  INV_X1     g02925(.I(new_n3078_), .ZN(new_n3118_));
  OAI21_X1   g02926(.A1(new_n3115_), .A2(new_n3118_), .B(\asqrt[57] ), .ZN(new_n3119_));
  NAND3_X1   g02927(.A1(new_n3117_), .A2(new_n3119_), .A3(new_n403_), .ZN(new_n3120_));
  NAND2_X1   g02928(.A1(new_n3120_), .A2(new_n3094_), .ZN(new_n3121_));
  NAND2_X1   g02929(.A1(new_n3117_), .A2(new_n3119_), .ZN(new_n3122_));
  AOI21_X1   g02930(.A1(new_n3122_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n3123_));
  AOI21_X1   g02931(.A1(new_n3123_), .A2(new_n3121_), .B(new_n3113_), .ZN(new_n3124_));
  AOI21_X1   g02932(.A1(new_n3121_), .A2(new_n3106_), .B(new_n339_), .ZN(new_n3125_));
  OAI21_X1   g02933(.A1(new_n3124_), .A2(new_n3125_), .B(\asqrt[60] ), .ZN(new_n3126_));
  AOI21_X1   g02934(.A1(new_n3112_), .A2(new_n3126_), .B(new_n242_), .ZN(new_n3127_));
  NAND3_X1   g02935(.A1(\asqrt[41] ), .A2(new_n2870_), .A3(new_n2886_), .ZN(new_n3128_));
  XOR2_X1    g02936(.A1(new_n3128_), .A2(new_n2898_), .Z(new_n3129_));
  INV_X1     g02937(.I(new_n3129_), .ZN(new_n3130_));
  NAND2_X1   g02938(.A1(new_n3108_), .A2(new_n3110_), .ZN(new_n3131_));
  AOI21_X1   g02939(.A1(new_n3131_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n3132_));
  AOI21_X1   g02940(.A1(new_n3132_), .A2(new_n3112_), .B(new_n3130_), .ZN(new_n3133_));
  OAI21_X1   g02941(.A1(new_n3133_), .A2(new_n3127_), .B(\asqrt[62] ), .ZN(new_n3134_));
  INV_X1     g02942(.I(new_n3134_), .ZN(new_n3135_));
  NOR2_X1    g02943(.A1(new_n3133_), .A2(new_n3127_), .ZN(new_n3136_));
  AOI21_X1   g02944(.A1(new_n2871_), .A2(new_n2892_), .B(new_n2887_), .ZN(new_n3137_));
  NAND2_X1   g02945(.A1(\asqrt[41] ), .A2(new_n3137_), .ZN(new_n3138_));
  XOR2_X1    g02946(.A1(new_n3138_), .A2(new_n2890_), .Z(new_n3139_));
  INV_X1     g02947(.I(new_n3139_), .ZN(new_n3140_));
  AOI21_X1   g02948(.A1(new_n3136_), .A2(new_n234_), .B(new_n3140_), .ZN(new_n3141_));
  OAI21_X1   g02949(.A1(new_n3141_), .A2(new_n3135_), .B(new_n3086_), .ZN(new_n3142_));
  OAI21_X1   g02950(.A1(new_n3142_), .A2(new_n3085_), .B(new_n193_), .ZN(new_n3143_));
  NOR2_X1    g02951(.A1(new_n3141_), .A2(new_n3135_), .ZN(new_n3144_));
  NAND2_X1   g02952(.A1(new_n3144_), .A2(new_n3085_), .ZN(new_n3145_));
  NOR2_X1    g02953(.A1(\asqrt[41] ), .A2(new_n2705_), .ZN(new_n3146_));
  INV_X1     g02954(.I(new_n3146_), .ZN(new_n3147_));
  NAND4_X1   g02955(.A1(new_n3143_), .A2(new_n3083_), .A3(new_n3145_), .A4(new_n3147_), .ZN(\asqrt[40] ));
  NAND3_X1   g02956(.A1(\asqrt[40] ), .A2(new_n3063_), .A3(new_n3078_), .ZN(new_n3149_));
  XOR2_X1    g02957(.A1(new_n3149_), .A2(new_n2916_), .Z(new_n3150_));
  INV_X1     g02958(.I(new_n3089_), .ZN(new_n3151_));
  NOR2_X1    g02959(.A1(new_n3124_), .A2(new_n3125_), .ZN(new_n3152_));
  AOI21_X1   g02960(.A1(new_n3152_), .A2(new_n288_), .B(new_n3151_), .ZN(new_n3153_));
  INV_X1     g02961(.I(new_n3126_), .ZN(new_n3154_));
  OAI21_X1   g02962(.A1(new_n3153_), .A2(new_n3154_), .B(\asqrt[61] ), .ZN(new_n3155_));
  NAND2_X1   g02963(.A1(new_n3126_), .A2(new_n242_), .ZN(new_n3156_));
  OAI21_X1   g02964(.A1(new_n3153_), .A2(new_n3156_), .B(new_n3129_), .ZN(new_n3157_));
  NAND3_X1   g02965(.A1(new_n3157_), .A2(new_n3155_), .A3(new_n234_), .ZN(new_n3158_));
  NAND2_X1   g02966(.A1(new_n3158_), .A2(new_n3139_), .ZN(new_n3159_));
  NAND2_X1   g02967(.A1(new_n3159_), .A2(new_n3134_), .ZN(new_n3160_));
  NAND2_X1   g02968(.A1(new_n3160_), .A2(new_n3085_), .ZN(new_n3161_));
  INV_X1     g02969(.I(new_n3085_), .ZN(new_n3162_));
  INV_X1     g02970(.I(new_n3086_), .ZN(new_n3163_));
  AOI21_X1   g02971(.A1(new_n3159_), .A2(new_n3134_), .B(new_n3163_), .ZN(new_n3164_));
  AOI21_X1   g02972(.A1(new_n3164_), .A2(new_n3162_), .B(\asqrt[63] ), .ZN(new_n3165_));
  NOR2_X1    g02973(.A1(new_n3160_), .A2(new_n3162_), .ZN(new_n3166_));
  NOR4_X1    g02974(.A1(new_n3165_), .A2(new_n3082_), .A3(new_n3166_), .A4(new_n3146_), .ZN(new_n3167_));
  NOR2_X1    g02975(.A1(new_n3167_), .A2(new_n3085_), .ZN(new_n3168_));
  NAND2_X1   g02976(.A1(new_n3168_), .A2(new_n3144_), .ZN(new_n3169_));
  AOI21_X1   g02977(.A1(new_n3169_), .A2(new_n3161_), .B(new_n193_), .ZN(new_n3170_));
  NAND3_X1   g02978(.A1(\asqrt[40] ), .A2(new_n3134_), .A3(new_n3158_), .ZN(new_n3171_));
  XOR2_X1    g02979(.A1(new_n3171_), .A2(new_n3139_), .Z(new_n3172_));
  INV_X1     g02980(.I(new_n3172_), .ZN(new_n3173_));
  AOI21_X1   g02981(.A1(new_n3168_), .A2(new_n3160_), .B(new_n3166_), .ZN(new_n3174_));
  INV_X1     g02982(.I(new_n3174_), .ZN(new_n3175_));
  OAI21_X1   g02983(.A1(new_n3105_), .A2(new_n3107_), .B(new_n3110_), .ZN(new_n3176_));
  NOR2_X1    g02984(.A1(new_n3167_), .A2(new_n3176_), .ZN(new_n3177_));
  XOR2_X1    g02985(.A1(new_n3177_), .A2(new_n3091_), .Z(new_n3178_));
  NAND3_X1   g02986(.A1(\asqrt[40] ), .A2(new_n3120_), .A3(new_n3106_), .ZN(new_n3179_));
  XOR2_X1    g02987(.A1(new_n3179_), .A2(new_n3095_), .Z(new_n3180_));
  OAI21_X1   g02988(.A1(new_n3115_), .A2(new_n3116_), .B(new_n3119_), .ZN(new_n3181_));
  NOR2_X1    g02989(.A1(new_n3167_), .A2(new_n3181_), .ZN(new_n3182_));
  XOR2_X1    g02990(.A1(new_n3182_), .A2(new_n3097_), .Z(new_n3183_));
  INV_X1     g02991(.I(new_n3183_), .ZN(new_n3184_));
  INV_X1     g02992(.I(new_n3150_), .ZN(new_n3185_));
  OAI21_X1   g02993(.A1(new_n3057_), .A2(new_n3059_), .B(new_n3062_), .ZN(new_n3186_));
  NOR2_X1    g02994(.A1(new_n3167_), .A2(new_n3186_), .ZN(new_n3187_));
  XOR2_X1    g02995(.A1(new_n3187_), .A2(new_n2929_), .Z(new_n3188_));
  NAND3_X1   g02996(.A1(\asqrt[40] ), .A2(new_n3072_), .A3(new_n3058_), .ZN(new_n3189_));
  XOR2_X1    g02997(.A1(new_n3189_), .A2(new_n2933_), .Z(new_n3190_));
  OAI21_X1   g02998(.A1(new_n3067_), .A2(new_n3068_), .B(new_n3071_), .ZN(new_n3191_));
  NOR2_X1    g02999(.A1(new_n3167_), .A2(new_n3191_), .ZN(new_n3192_));
  XOR2_X1    g03000(.A1(new_n3192_), .A2(new_n2935_), .Z(new_n3193_));
  INV_X1     g03001(.I(new_n3193_), .ZN(new_n3194_));
  NAND3_X1   g03002(.A1(\asqrt[40] ), .A2(new_n3035_), .A3(new_n3054_), .ZN(new_n3195_));
  XOR2_X1    g03003(.A1(new_n3195_), .A2(new_n3065_), .Z(new_n3196_));
  INV_X1     g03004(.I(new_n3196_), .ZN(new_n3197_));
  OAI21_X1   g03005(.A1(new_n3029_), .A2(new_n3031_), .B(new_n3034_), .ZN(new_n3198_));
  NOR2_X1    g03006(.A1(new_n3167_), .A2(new_n3198_), .ZN(new_n3199_));
  XOR2_X1    g03007(.A1(new_n3199_), .A2(new_n2941_), .Z(new_n3200_));
  NAND3_X1   g03008(.A1(\asqrt[40] ), .A2(new_n3048_), .A3(new_n3030_), .ZN(new_n3201_));
  XOR2_X1    g03009(.A1(new_n3201_), .A2(new_n2945_), .Z(new_n3202_));
  OAI21_X1   g03010(.A1(new_n3043_), .A2(new_n3044_), .B(new_n3047_), .ZN(new_n3203_));
  NOR2_X1    g03011(.A1(new_n3167_), .A2(new_n3203_), .ZN(new_n3204_));
  XOR2_X1    g03012(.A1(new_n3204_), .A2(new_n2947_), .Z(new_n3205_));
  INV_X1     g03013(.I(new_n3205_), .ZN(new_n3206_));
  NAND3_X1   g03014(.A1(\asqrt[40] ), .A2(new_n3007_), .A3(new_n3026_), .ZN(new_n3207_));
  XOR2_X1    g03015(.A1(new_n3207_), .A2(new_n3041_), .Z(new_n3208_));
  INV_X1     g03016(.I(new_n3208_), .ZN(new_n3209_));
  OAI21_X1   g03017(.A1(new_n3001_), .A2(new_n3003_), .B(new_n3006_), .ZN(new_n3210_));
  NOR2_X1    g03018(.A1(new_n3167_), .A2(new_n3210_), .ZN(new_n3211_));
  XOR2_X1    g03019(.A1(new_n3211_), .A2(new_n2954_), .Z(new_n3212_));
  NAND3_X1   g03020(.A1(\asqrt[40] ), .A2(new_n3020_), .A3(new_n3002_), .ZN(new_n3213_));
  XOR2_X1    g03021(.A1(new_n3213_), .A2(new_n2957_), .Z(new_n3214_));
  OAI21_X1   g03022(.A1(new_n3015_), .A2(new_n3016_), .B(new_n3019_), .ZN(new_n3215_));
  NOR2_X1    g03023(.A1(new_n3167_), .A2(new_n3215_), .ZN(new_n3216_));
  XOR2_X1    g03024(.A1(new_n3216_), .A2(new_n2960_), .Z(new_n3217_));
  INV_X1     g03025(.I(new_n3217_), .ZN(new_n3218_));
  NAND3_X1   g03026(.A1(\asqrt[40] ), .A2(new_n2980_), .A3(new_n2998_), .ZN(new_n3219_));
  XOR2_X1    g03027(.A1(new_n3219_), .A2(new_n3014_), .Z(new_n3220_));
  INV_X1     g03028(.I(new_n3220_), .ZN(new_n3221_));
  NOR2_X1    g03029(.A1(new_n2977_), .A2(\asqrt[43] ), .ZN(new_n3222_));
  NOR3_X1    g03030(.A1(new_n3167_), .A2(new_n3222_), .A3(new_n2997_), .ZN(new_n3223_));
  XOR2_X1    g03031(.A1(new_n3223_), .A2(new_n2968_), .Z(new_n3224_));
  NOR3_X1    g03032(.A1(new_n3167_), .A2(\a[80] ), .A3(\a[81] ), .ZN(new_n3225_));
  NOR4_X1    g03033(.A1(new_n3165_), .A2(new_n2912_), .A3(new_n3082_), .A4(new_n3166_), .ZN(new_n3226_));
  OAI21_X1   g03034(.A1(new_n3225_), .A2(new_n3226_), .B(new_n2758_), .ZN(new_n3227_));
  NAND3_X1   g03035(.A1(\asqrt[40] ), .A2(new_n2969_), .A3(new_n2970_), .ZN(new_n3228_));
  INV_X1     g03036(.I(new_n3226_), .ZN(new_n3229_));
  NAND3_X1   g03037(.A1(new_n3228_), .A2(\a[82] ), .A3(new_n3229_), .ZN(new_n3230_));
  NAND2_X1   g03038(.A1(new_n3227_), .A2(new_n3230_), .ZN(new_n3231_));
  INV_X1     g03039(.I(\a[78] ), .ZN(new_n3232_));
  INV_X1     g03040(.I(\a[79] ), .ZN(new_n3233_));
  NAND3_X1   g03041(.A1(new_n3232_), .A2(new_n3233_), .A3(new_n2969_), .ZN(new_n3234_));
  NAND2_X1   g03042(.A1(\asqrt[40] ), .A2(\a[80] ), .ZN(new_n3235_));
  AOI21_X1   g03043(.A1(new_n3235_), .A2(new_n3234_), .B(new_n2912_), .ZN(new_n3236_));
  AOI21_X1   g03044(.A1(\asqrt[40] ), .A2(new_n2969_), .B(new_n2970_), .ZN(new_n3237_));
  NOR2_X1    g03045(.A1(new_n3225_), .A2(new_n3237_), .ZN(new_n3238_));
  NAND3_X1   g03046(.A1(new_n3235_), .A2(new_n2912_), .A3(new_n3234_), .ZN(new_n3239_));
  AOI21_X1   g03047(.A1(new_n3238_), .A2(new_n3239_), .B(new_n3236_), .ZN(new_n3240_));
  AOI21_X1   g03048(.A1(new_n3240_), .A2(new_n2699_), .B(new_n3231_), .ZN(new_n3241_));
  NOR2_X1    g03049(.A1(new_n3240_), .A2(new_n2699_), .ZN(new_n3242_));
  NOR3_X1    g03050(.A1(new_n3241_), .A2(\asqrt[43] ), .A3(new_n3242_), .ZN(new_n3243_));
  NOR3_X1    g03051(.A1(new_n3167_), .A2(new_n2991_), .A3(new_n2976_), .ZN(new_n3244_));
  XOR2_X1    g03052(.A1(new_n3244_), .A2(new_n2993_), .Z(new_n3245_));
  INV_X1     g03053(.I(new_n3245_), .ZN(new_n3246_));
  OAI21_X1   g03054(.A1(new_n3241_), .A2(new_n3242_), .B(\asqrt[43] ), .ZN(new_n3247_));
  OAI21_X1   g03055(.A1(new_n3243_), .A2(new_n3246_), .B(new_n3247_), .ZN(new_n3248_));
  OAI21_X1   g03056(.A1(new_n3248_), .A2(\asqrt[44] ), .B(new_n3224_), .ZN(new_n3249_));
  AOI21_X1   g03057(.A1(new_n3248_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n3250_));
  AOI21_X1   g03058(.A1(new_n3250_), .A2(new_n3249_), .B(new_n3221_), .ZN(new_n3251_));
  NAND2_X1   g03059(.A1(new_n3248_), .A2(\asqrt[44] ), .ZN(new_n3252_));
  AOI21_X1   g03060(.A1(new_n3249_), .A2(new_n3252_), .B(new_n2072_), .ZN(new_n3253_));
  NOR2_X1    g03061(.A1(new_n3251_), .A2(new_n3253_), .ZN(new_n3254_));
  AOI21_X1   g03062(.A1(new_n3254_), .A2(new_n1884_), .B(new_n3218_), .ZN(new_n3255_));
  OAI21_X1   g03063(.A1(new_n3251_), .A2(new_n3253_), .B(\asqrt[46] ), .ZN(new_n3256_));
  NAND2_X1   g03064(.A1(new_n3256_), .A2(new_n1688_), .ZN(new_n3257_));
  OAI21_X1   g03065(.A1(new_n3255_), .A2(new_n3257_), .B(new_n3214_), .ZN(new_n3258_));
  INV_X1     g03066(.I(new_n3256_), .ZN(new_n3259_));
  OAI21_X1   g03067(.A1(new_n3255_), .A2(new_n3259_), .B(\asqrt[47] ), .ZN(new_n3260_));
  NAND3_X1   g03068(.A1(new_n3258_), .A2(new_n3260_), .A3(new_n1533_), .ZN(new_n3261_));
  NAND2_X1   g03069(.A1(new_n3261_), .A2(new_n3212_), .ZN(new_n3262_));
  NAND2_X1   g03070(.A1(new_n3258_), .A2(new_n3260_), .ZN(new_n3263_));
  AOI21_X1   g03071(.A1(new_n3263_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n3264_));
  AOI21_X1   g03072(.A1(new_n3264_), .A2(new_n3262_), .B(new_n3209_), .ZN(new_n3265_));
  INV_X1     g03073(.I(new_n3214_), .ZN(new_n3266_));
  INV_X1     g03074(.I(new_n3224_), .ZN(new_n3267_));
  AOI21_X1   g03075(.A1(new_n3228_), .A2(new_n3229_), .B(\a[82] ), .ZN(new_n3268_));
  NOR3_X1    g03076(.A1(new_n3225_), .A2(new_n2758_), .A3(new_n3226_), .ZN(new_n3269_));
  NOR2_X1    g03077(.A1(new_n3269_), .A2(new_n3268_), .ZN(new_n3270_));
  OAI21_X1   g03078(.A1(new_n3167_), .A2(new_n2969_), .B(new_n3234_), .ZN(new_n3271_));
  NAND2_X1   g03079(.A1(new_n3271_), .A2(\asqrt[41] ), .ZN(new_n3272_));
  OAI21_X1   g03080(.A1(new_n3167_), .A2(\a[80] ), .B(\a[81] ), .ZN(new_n3273_));
  NAND2_X1   g03081(.A1(new_n3273_), .A2(new_n3228_), .ZN(new_n3274_));
  NOR2_X1    g03082(.A1(new_n3271_), .A2(\asqrt[41] ), .ZN(new_n3275_));
  OAI21_X1   g03083(.A1(new_n3274_), .A2(new_n3275_), .B(new_n3272_), .ZN(new_n3276_));
  OAI21_X1   g03084(.A1(\asqrt[42] ), .A2(new_n3276_), .B(new_n3270_), .ZN(new_n3277_));
  NAND2_X1   g03085(.A1(new_n3276_), .A2(\asqrt[42] ), .ZN(new_n3278_));
  NAND3_X1   g03086(.A1(new_n3277_), .A2(new_n2464_), .A3(new_n3278_), .ZN(new_n3279_));
  AOI21_X1   g03087(.A1(new_n3277_), .A2(new_n3278_), .B(new_n2464_), .ZN(new_n3280_));
  AOI21_X1   g03088(.A1(new_n3279_), .A2(new_n3245_), .B(new_n3280_), .ZN(new_n3281_));
  AOI21_X1   g03089(.A1(new_n3281_), .A2(new_n2271_), .B(new_n3267_), .ZN(new_n3282_));
  OAI21_X1   g03090(.A1(new_n3281_), .A2(new_n2271_), .B(new_n2072_), .ZN(new_n3283_));
  OAI21_X1   g03091(.A1(new_n3282_), .A2(new_n3283_), .B(new_n3220_), .ZN(new_n3284_));
  NOR2_X1    g03092(.A1(new_n3281_), .A2(new_n2271_), .ZN(new_n3285_));
  OAI21_X1   g03093(.A1(new_n3282_), .A2(new_n3285_), .B(\asqrt[45] ), .ZN(new_n3286_));
  NAND3_X1   g03094(.A1(new_n3284_), .A2(new_n3286_), .A3(new_n1884_), .ZN(new_n3287_));
  NAND2_X1   g03095(.A1(new_n3287_), .A2(new_n3217_), .ZN(new_n3288_));
  NAND2_X1   g03096(.A1(new_n3284_), .A2(new_n3286_), .ZN(new_n3289_));
  AOI21_X1   g03097(.A1(new_n3289_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n3290_));
  AOI21_X1   g03098(.A1(new_n3290_), .A2(new_n3288_), .B(new_n3266_), .ZN(new_n3291_));
  AOI21_X1   g03099(.A1(new_n3288_), .A2(new_n3256_), .B(new_n1688_), .ZN(new_n3292_));
  OAI21_X1   g03100(.A1(new_n3291_), .A2(new_n3292_), .B(\asqrt[48] ), .ZN(new_n3293_));
  AOI21_X1   g03101(.A1(new_n3262_), .A2(new_n3293_), .B(new_n1368_), .ZN(new_n3294_));
  NOR2_X1    g03102(.A1(new_n3265_), .A2(new_n3294_), .ZN(new_n3295_));
  AOI21_X1   g03103(.A1(new_n3295_), .A2(new_n1228_), .B(new_n3206_), .ZN(new_n3296_));
  OAI21_X1   g03104(.A1(new_n3265_), .A2(new_n3294_), .B(\asqrt[50] ), .ZN(new_n3297_));
  NAND2_X1   g03105(.A1(new_n3297_), .A2(new_n1088_), .ZN(new_n3298_));
  OAI21_X1   g03106(.A1(new_n3296_), .A2(new_n3298_), .B(new_n3202_), .ZN(new_n3299_));
  INV_X1     g03107(.I(new_n3297_), .ZN(new_n3300_));
  OAI21_X1   g03108(.A1(new_n3296_), .A2(new_n3300_), .B(\asqrt[51] ), .ZN(new_n3301_));
  NAND3_X1   g03109(.A1(new_n3299_), .A2(new_n3301_), .A3(new_n962_), .ZN(new_n3302_));
  NAND2_X1   g03110(.A1(new_n3302_), .A2(new_n3200_), .ZN(new_n3303_));
  NAND2_X1   g03111(.A1(new_n3299_), .A2(new_n3301_), .ZN(new_n3304_));
  AOI21_X1   g03112(.A1(new_n3304_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n3305_));
  AOI21_X1   g03113(.A1(new_n3305_), .A2(new_n3303_), .B(new_n3197_), .ZN(new_n3306_));
  INV_X1     g03114(.I(new_n3202_), .ZN(new_n3307_));
  INV_X1     g03115(.I(new_n3212_), .ZN(new_n3308_));
  NOR2_X1    g03116(.A1(new_n3291_), .A2(new_n3292_), .ZN(new_n3309_));
  AOI21_X1   g03117(.A1(new_n3309_), .A2(new_n1533_), .B(new_n3308_), .ZN(new_n3310_));
  NAND2_X1   g03118(.A1(new_n3293_), .A2(new_n1368_), .ZN(new_n3311_));
  OAI21_X1   g03119(.A1(new_n3310_), .A2(new_n3311_), .B(new_n3208_), .ZN(new_n3312_));
  INV_X1     g03120(.I(new_n3293_), .ZN(new_n3313_));
  OAI21_X1   g03121(.A1(new_n3310_), .A2(new_n3313_), .B(\asqrt[49] ), .ZN(new_n3314_));
  NAND3_X1   g03122(.A1(new_n3312_), .A2(new_n3314_), .A3(new_n1228_), .ZN(new_n3315_));
  NAND2_X1   g03123(.A1(new_n3315_), .A2(new_n3205_), .ZN(new_n3316_));
  NAND2_X1   g03124(.A1(new_n3312_), .A2(new_n3314_), .ZN(new_n3317_));
  AOI21_X1   g03125(.A1(new_n3317_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n3318_));
  AOI21_X1   g03126(.A1(new_n3318_), .A2(new_n3316_), .B(new_n3307_), .ZN(new_n3319_));
  AOI21_X1   g03127(.A1(new_n3316_), .A2(new_n3297_), .B(new_n1088_), .ZN(new_n3320_));
  OAI21_X1   g03128(.A1(new_n3319_), .A2(new_n3320_), .B(\asqrt[52] ), .ZN(new_n3321_));
  AOI21_X1   g03129(.A1(new_n3303_), .A2(new_n3321_), .B(new_n842_), .ZN(new_n3322_));
  NOR2_X1    g03130(.A1(new_n3306_), .A2(new_n3322_), .ZN(new_n3323_));
  AOI21_X1   g03131(.A1(new_n3323_), .A2(new_n720_), .B(new_n3194_), .ZN(new_n3324_));
  OAI21_X1   g03132(.A1(new_n3306_), .A2(new_n3322_), .B(\asqrt[54] ), .ZN(new_n3325_));
  NAND2_X1   g03133(.A1(new_n3325_), .A2(new_n630_), .ZN(new_n3326_));
  OAI21_X1   g03134(.A1(new_n3324_), .A2(new_n3326_), .B(new_n3190_), .ZN(new_n3327_));
  INV_X1     g03135(.I(new_n3325_), .ZN(new_n3328_));
  OAI21_X1   g03136(.A1(new_n3324_), .A2(new_n3328_), .B(\asqrt[55] ), .ZN(new_n3329_));
  NAND3_X1   g03137(.A1(new_n3327_), .A2(new_n3329_), .A3(new_n545_), .ZN(new_n3330_));
  NAND2_X1   g03138(.A1(new_n3330_), .A2(new_n3188_), .ZN(new_n3331_));
  NAND2_X1   g03139(.A1(new_n3327_), .A2(new_n3329_), .ZN(new_n3332_));
  AOI21_X1   g03140(.A1(new_n3332_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n3333_));
  AOI21_X1   g03141(.A1(new_n3333_), .A2(new_n3331_), .B(new_n3185_), .ZN(new_n3334_));
  INV_X1     g03142(.I(new_n3190_), .ZN(new_n3335_));
  INV_X1     g03143(.I(new_n3200_), .ZN(new_n3336_));
  NOR2_X1    g03144(.A1(new_n3319_), .A2(new_n3320_), .ZN(new_n3337_));
  AOI21_X1   g03145(.A1(new_n3337_), .A2(new_n962_), .B(new_n3336_), .ZN(new_n3338_));
  NAND2_X1   g03146(.A1(new_n3321_), .A2(new_n842_), .ZN(new_n3339_));
  OAI21_X1   g03147(.A1(new_n3338_), .A2(new_n3339_), .B(new_n3196_), .ZN(new_n3340_));
  INV_X1     g03148(.I(new_n3321_), .ZN(new_n3341_));
  OAI21_X1   g03149(.A1(new_n3338_), .A2(new_n3341_), .B(\asqrt[53] ), .ZN(new_n3342_));
  NAND3_X1   g03150(.A1(new_n3340_), .A2(new_n3342_), .A3(new_n720_), .ZN(new_n3343_));
  NAND2_X1   g03151(.A1(new_n3343_), .A2(new_n3193_), .ZN(new_n3344_));
  NAND2_X1   g03152(.A1(new_n3340_), .A2(new_n3342_), .ZN(new_n3345_));
  AOI21_X1   g03153(.A1(new_n3345_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n3346_));
  AOI21_X1   g03154(.A1(new_n3346_), .A2(new_n3344_), .B(new_n3335_), .ZN(new_n3347_));
  AOI21_X1   g03155(.A1(new_n3344_), .A2(new_n3325_), .B(new_n630_), .ZN(new_n3348_));
  OAI21_X1   g03156(.A1(new_n3347_), .A2(new_n3348_), .B(\asqrt[56] ), .ZN(new_n3349_));
  AOI21_X1   g03157(.A1(new_n3331_), .A2(new_n3349_), .B(new_n450_), .ZN(new_n3350_));
  NOR2_X1    g03158(.A1(new_n3334_), .A2(new_n3350_), .ZN(new_n3351_));
  AOI21_X1   g03159(.A1(new_n3351_), .A2(new_n403_), .B(new_n3184_), .ZN(new_n3352_));
  OAI21_X1   g03160(.A1(new_n3334_), .A2(new_n3350_), .B(\asqrt[58] ), .ZN(new_n3353_));
  NAND2_X1   g03161(.A1(new_n3353_), .A2(new_n339_), .ZN(new_n3354_));
  OAI21_X1   g03162(.A1(new_n3352_), .A2(new_n3354_), .B(new_n3180_), .ZN(new_n3355_));
  INV_X1     g03163(.I(new_n3353_), .ZN(new_n3356_));
  OAI21_X1   g03164(.A1(new_n3352_), .A2(new_n3356_), .B(\asqrt[59] ), .ZN(new_n3357_));
  NAND3_X1   g03165(.A1(new_n3355_), .A2(new_n3357_), .A3(new_n288_), .ZN(new_n3358_));
  NAND2_X1   g03166(.A1(new_n3358_), .A2(new_n3178_), .ZN(new_n3359_));
  INV_X1     g03167(.I(new_n3180_), .ZN(new_n3360_));
  INV_X1     g03168(.I(new_n3188_), .ZN(new_n3361_));
  NOR2_X1    g03169(.A1(new_n3347_), .A2(new_n3348_), .ZN(new_n3362_));
  AOI21_X1   g03170(.A1(new_n3362_), .A2(new_n545_), .B(new_n3361_), .ZN(new_n3363_));
  NAND2_X1   g03171(.A1(new_n3349_), .A2(new_n450_), .ZN(new_n3364_));
  OAI21_X1   g03172(.A1(new_n3363_), .A2(new_n3364_), .B(new_n3150_), .ZN(new_n3365_));
  INV_X1     g03173(.I(new_n3349_), .ZN(new_n3366_));
  OAI21_X1   g03174(.A1(new_n3363_), .A2(new_n3366_), .B(\asqrt[57] ), .ZN(new_n3367_));
  NAND3_X1   g03175(.A1(new_n3365_), .A2(new_n3367_), .A3(new_n403_), .ZN(new_n3368_));
  NAND2_X1   g03176(.A1(new_n3368_), .A2(new_n3183_), .ZN(new_n3369_));
  NAND2_X1   g03177(.A1(new_n3365_), .A2(new_n3367_), .ZN(new_n3370_));
  AOI21_X1   g03178(.A1(new_n3370_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n3371_));
  AOI21_X1   g03179(.A1(new_n3371_), .A2(new_n3369_), .B(new_n3360_), .ZN(new_n3372_));
  AOI21_X1   g03180(.A1(new_n3369_), .A2(new_n3353_), .B(new_n339_), .ZN(new_n3373_));
  OAI21_X1   g03181(.A1(new_n3372_), .A2(new_n3373_), .B(\asqrt[60] ), .ZN(new_n3374_));
  AOI21_X1   g03182(.A1(new_n3359_), .A2(new_n3374_), .B(new_n242_), .ZN(new_n3375_));
  NAND3_X1   g03183(.A1(\asqrt[40] ), .A2(new_n3111_), .A3(new_n3126_), .ZN(new_n3376_));
  XOR2_X1    g03184(.A1(new_n3376_), .A2(new_n3151_), .Z(new_n3377_));
  INV_X1     g03185(.I(new_n3377_), .ZN(new_n3378_));
  NAND2_X1   g03186(.A1(new_n3355_), .A2(new_n3357_), .ZN(new_n3379_));
  AOI21_X1   g03187(.A1(new_n3379_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n3380_));
  AOI21_X1   g03188(.A1(new_n3380_), .A2(new_n3359_), .B(new_n3378_), .ZN(new_n3381_));
  OAI21_X1   g03189(.A1(new_n3381_), .A2(new_n3375_), .B(\asqrt[62] ), .ZN(new_n3382_));
  AOI21_X1   g03190(.A1(new_n3112_), .A2(new_n3132_), .B(new_n3127_), .ZN(new_n3383_));
  NAND2_X1   g03191(.A1(\asqrt[40] ), .A2(new_n3383_), .ZN(new_n3384_));
  XOR2_X1    g03192(.A1(new_n3384_), .A2(new_n3130_), .Z(new_n3385_));
  INV_X1     g03193(.I(new_n3178_), .ZN(new_n3386_));
  NOR2_X1    g03194(.A1(new_n3372_), .A2(new_n3373_), .ZN(new_n3387_));
  AOI21_X1   g03195(.A1(new_n3387_), .A2(new_n288_), .B(new_n3386_), .ZN(new_n3388_));
  INV_X1     g03196(.I(new_n3374_), .ZN(new_n3389_));
  OAI21_X1   g03197(.A1(new_n3388_), .A2(new_n3389_), .B(\asqrt[61] ), .ZN(new_n3390_));
  NAND2_X1   g03198(.A1(new_n3374_), .A2(new_n242_), .ZN(new_n3391_));
  OAI21_X1   g03199(.A1(new_n3388_), .A2(new_n3391_), .B(new_n3377_), .ZN(new_n3392_));
  NAND3_X1   g03200(.A1(new_n3392_), .A2(new_n3390_), .A3(new_n234_), .ZN(new_n3393_));
  NAND2_X1   g03201(.A1(new_n3393_), .A2(new_n3385_), .ZN(new_n3394_));
  AOI21_X1   g03202(.A1(new_n3394_), .A2(new_n3382_), .B(new_n3175_), .ZN(new_n3395_));
  AOI21_X1   g03203(.A1(new_n3395_), .A2(new_n3173_), .B(\asqrt[63] ), .ZN(new_n3396_));
  NAND2_X1   g03204(.A1(new_n3394_), .A2(new_n3382_), .ZN(new_n3397_));
  NOR2_X1    g03205(.A1(new_n3397_), .A2(new_n3173_), .ZN(new_n3398_));
  NOR2_X1    g03206(.A1(\asqrt[40] ), .A2(new_n3162_), .ZN(new_n3399_));
  NOR4_X1    g03207(.A1(new_n3396_), .A2(new_n3170_), .A3(new_n3398_), .A4(new_n3399_), .ZN(new_n3400_));
  OAI21_X1   g03208(.A1(new_n3363_), .A2(new_n3364_), .B(new_n3367_), .ZN(new_n3401_));
  NOR2_X1    g03209(.A1(new_n3400_), .A2(new_n3401_), .ZN(new_n3402_));
  XOR2_X1    g03210(.A1(new_n3402_), .A2(new_n3150_), .Z(new_n3403_));
  INV_X1     g03211(.I(new_n3403_), .ZN(new_n3404_));
  INV_X1     g03212(.I(new_n3170_), .ZN(new_n3405_));
  INV_X1     g03213(.I(new_n3382_), .ZN(new_n3406_));
  NOR2_X1    g03214(.A1(new_n3381_), .A2(new_n3375_), .ZN(new_n3407_));
  INV_X1     g03215(.I(new_n3385_), .ZN(new_n3408_));
  AOI21_X1   g03216(.A1(new_n3407_), .A2(new_n234_), .B(new_n3408_), .ZN(new_n3409_));
  OAI21_X1   g03217(.A1(new_n3409_), .A2(new_n3406_), .B(new_n3174_), .ZN(new_n3410_));
  OAI21_X1   g03218(.A1(new_n3410_), .A2(new_n3172_), .B(new_n193_), .ZN(new_n3411_));
  NOR2_X1    g03219(.A1(new_n3409_), .A2(new_n3406_), .ZN(new_n3412_));
  NAND2_X1   g03220(.A1(new_n3412_), .A2(new_n3172_), .ZN(new_n3413_));
  INV_X1     g03221(.I(new_n3399_), .ZN(new_n3414_));
  NAND4_X1   g03222(.A1(new_n3411_), .A2(new_n3405_), .A3(new_n3413_), .A4(new_n3414_), .ZN(\asqrt[39] ));
  NAND3_X1   g03223(.A1(\asqrt[39] ), .A2(new_n3330_), .A3(new_n3349_), .ZN(new_n3416_));
  XOR2_X1    g03224(.A1(new_n3416_), .A2(new_n3361_), .Z(new_n3417_));
  OAI21_X1   g03225(.A1(new_n3324_), .A2(new_n3326_), .B(new_n3329_), .ZN(new_n3418_));
  NOR2_X1    g03226(.A1(new_n3400_), .A2(new_n3418_), .ZN(new_n3419_));
  XOR2_X1    g03227(.A1(new_n3419_), .A2(new_n3190_), .Z(new_n3420_));
  INV_X1     g03228(.I(new_n3420_), .ZN(new_n3421_));
  NAND3_X1   g03229(.A1(\asqrt[39] ), .A2(new_n3343_), .A3(new_n3325_), .ZN(new_n3422_));
  XOR2_X1    g03230(.A1(new_n3422_), .A2(new_n3194_), .Z(new_n3423_));
  INV_X1     g03231(.I(new_n3423_), .ZN(new_n3424_));
  OAI21_X1   g03232(.A1(new_n3338_), .A2(new_n3339_), .B(new_n3342_), .ZN(new_n3425_));
  NOR2_X1    g03233(.A1(new_n3400_), .A2(new_n3425_), .ZN(new_n3426_));
  XOR2_X1    g03234(.A1(new_n3426_), .A2(new_n3196_), .Z(new_n3427_));
  NAND3_X1   g03235(.A1(\asqrt[39] ), .A2(new_n3302_), .A3(new_n3321_), .ZN(new_n3428_));
  XOR2_X1    g03236(.A1(new_n3428_), .A2(new_n3336_), .Z(new_n3429_));
  OAI21_X1   g03237(.A1(new_n3296_), .A2(new_n3298_), .B(new_n3301_), .ZN(new_n3430_));
  NOR2_X1    g03238(.A1(new_n3400_), .A2(new_n3430_), .ZN(new_n3431_));
  XOR2_X1    g03239(.A1(new_n3431_), .A2(new_n3202_), .Z(new_n3432_));
  INV_X1     g03240(.I(new_n3432_), .ZN(new_n3433_));
  NAND3_X1   g03241(.A1(\asqrt[39] ), .A2(new_n3315_), .A3(new_n3297_), .ZN(new_n3434_));
  XOR2_X1    g03242(.A1(new_n3434_), .A2(new_n3206_), .Z(new_n3435_));
  INV_X1     g03243(.I(new_n3435_), .ZN(new_n3436_));
  OAI21_X1   g03244(.A1(new_n3310_), .A2(new_n3311_), .B(new_n3314_), .ZN(new_n3437_));
  NOR2_X1    g03245(.A1(new_n3400_), .A2(new_n3437_), .ZN(new_n3438_));
  XOR2_X1    g03246(.A1(new_n3438_), .A2(new_n3208_), .Z(new_n3439_));
  NAND3_X1   g03247(.A1(\asqrt[39] ), .A2(new_n3261_), .A3(new_n3293_), .ZN(new_n3440_));
  XOR2_X1    g03248(.A1(new_n3440_), .A2(new_n3308_), .Z(new_n3441_));
  OAI21_X1   g03249(.A1(new_n3255_), .A2(new_n3257_), .B(new_n3260_), .ZN(new_n3442_));
  NOR2_X1    g03250(.A1(new_n3400_), .A2(new_n3442_), .ZN(new_n3443_));
  XOR2_X1    g03251(.A1(new_n3443_), .A2(new_n3214_), .Z(new_n3444_));
  INV_X1     g03252(.I(new_n3444_), .ZN(new_n3445_));
  NAND3_X1   g03253(.A1(\asqrt[39] ), .A2(new_n3287_), .A3(new_n3256_), .ZN(new_n3446_));
  XOR2_X1    g03254(.A1(new_n3446_), .A2(new_n3218_), .Z(new_n3447_));
  INV_X1     g03255(.I(new_n3447_), .ZN(new_n3448_));
  AOI21_X1   g03256(.A1(new_n3249_), .A2(new_n3250_), .B(new_n3253_), .ZN(new_n3449_));
  NAND2_X1   g03257(.A1(\asqrt[39] ), .A2(new_n3449_), .ZN(new_n3450_));
  XOR2_X1    g03258(.A1(new_n3450_), .A2(new_n3221_), .Z(new_n3451_));
  NOR2_X1    g03259(.A1(new_n3248_), .A2(\asqrt[44] ), .ZN(new_n3452_));
  NOR3_X1    g03260(.A1(new_n3400_), .A2(new_n3452_), .A3(new_n3285_), .ZN(new_n3453_));
  XOR2_X1    g03261(.A1(new_n3453_), .A2(new_n3224_), .Z(new_n3454_));
  NOR3_X1    g03262(.A1(new_n3400_), .A2(new_n3243_), .A3(new_n3280_), .ZN(new_n3455_));
  XOR2_X1    g03263(.A1(new_n3455_), .A2(new_n3245_), .Z(new_n3456_));
  INV_X1     g03264(.I(new_n3456_), .ZN(new_n3457_));
  NOR2_X1    g03265(.A1(new_n3276_), .A2(\asqrt[42] ), .ZN(new_n3458_));
  NOR3_X1    g03266(.A1(new_n3400_), .A2(new_n3458_), .A3(new_n3242_), .ZN(new_n3459_));
  XOR2_X1    g03267(.A1(new_n3459_), .A2(new_n3270_), .Z(new_n3460_));
  INV_X1     g03268(.I(new_n3460_), .ZN(new_n3461_));
  NAND3_X1   g03269(.A1(\asqrt[39] ), .A2(new_n3232_), .A3(new_n3233_), .ZN(new_n3462_));
  NAND4_X1   g03270(.A1(new_n3411_), .A2(\asqrt[40] ), .A3(new_n3413_), .A4(new_n3405_), .ZN(new_n3463_));
  AOI21_X1   g03271(.A1(new_n3462_), .A2(new_n3463_), .B(\a[80] ), .ZN(new_n3464_));
  NOR3_X1    g03272(.A1(new_n3400_), .A2(\a[78] ), .A3(\a[79] ), .ZN(new_n3465_));
  INV_X1     g03273(.I(new_n3463_), .ZN(new_n3466_));
  NOR3_X1    g03274(.A1(new_n3465_), .A2(new_n2969_), .A3(new_n3466_), .ZN(new_n3467_));
  NOR2_X1    g03275(.A1(new_n3467_), .A2(new_n3464_), .ZN(new_n3468_));
  INV_X1     g03276(.I(\a[76] ), .ZN(new_n3469_));
  INV_X1     g03277(.I(\a[77] ), .ZN(new_n3470_));
  NAND3_X1   g03278(.A1(new_n3469_), .A2(new_n3470_), .A3(new_n3232_), .ZN(new_n3471_));
  OAI21_X1   g03279(.A1(new_n3400_), .A2(new_n3232_), .B(new_n3471_), .ZN(new_n3472_));
  NAND2_X1   g03280(.A1(new_n3472_), .A2(\asqrt[40] ), .ZN(new_n3473_));
  OAI21_X1   g03281(.A1(new_n3400_), .A2(\a[78] ), .B(\a[79] ), .ZN(new_n3474_));
  NAND2_X1   g03282(.A1(new_n3474_), .A2(new_n3462_), .ZN(new_n3475_));
  NOR2_X1    g03283(.A1(new_n3472_), .A2(\asqrt[40] ), .ZN(new_n3476_));
  OAI21_X1   g03284(.A1(new_n3475_), .A2(new_n3476_), .B(new_n3473_), .ZN(new_n3477_));
  OAI21_X1   g03285(.A1(new_n3477_), .A2(\asqrt[41] ), .B(new_n3468_), .ZN(new_n3478_));
  NAND2_X1   g03286(.A1(new_n3477_), .A2(\asqrt[41] ), .ZN(new_n3479_));
  NAND3_X1   g03287(.A1(new_n3478_), .A2(new_n2699_), .A3(new_n3479_), .ZN(new_n3480_));
  NOR3_X1    g03288(.A1(new_n3400_), .A2(new_n3236_), .A3(new_n3275_), .ZN(new_n3481_));
  XOR2_X1    g03289(.A1(new_n3481_), .A2(new_n3238_), .Z(new_n3482_));
  NAND2_X1   g03290(.A1(new_n3480_), .A2(new_n3482_), .ZN(new_n3483_));
  NAND2_X1   g03291(.A1(new_n3478_), .A2(new_n3479_), .ZN(new_n3484_));
  AOI21_X1   g03292(.A1(new_n3484_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n3485_));
  AOI21_X1   g03293(.A1(new_n3485_), .A2(new_n3483_), .B(new_n3461_), .ZN(new_n3486_));
  OAI21_X1   g03294(.A1(new_n3465_), .A2(new_n3466_), .B(new_n2969_), .ZN(new_n3487_));
  NAND3_X1   g03295(.A1(new_n3462_), .A2(\a[80] ), .A3(new_n3463_), .ZN(new_n3488_));
  NAND2_X1   g03296(.A1(new_n3487_), .A2(new_n3488_), .ZN(new_n3489_));
  NAND2_X1   g03297(.A1(\asqrt[39] ), .A2(\a[78] ), .ZN(new_n3490_));
  AOI21_X1   g03298(.A1(new_n3490_), .A2(new_n3471_), .B(new_n3167_), .ZN(new_n3491_));
  AOI21_X1   g03299(.A1(\asqrt[39] ), .A2(new_n3232_), .B(new_n3233_), .ZN(new_n3492_));
  NOR2_X1    g03300(.A1(new_n3465_), .A2(new_n3492_), .ZN(new_n3493_));
  NAND3_X1   g03301(.A1(new_n3490_), .A2(new_n3167_), .A3(new_n3471_), .ZN(new_n3494_));
  AOI21_X1   g03302(.A1(new_n3493_), .A2(new_n3494_), .B(new_n3491_), .ZN(new_n3495_));
  AOI21_X1   g03303(.A1(new_n3495_), .A2(new_n2912_), .B(new_n3489_), .ZN(new_n3496_));
  NOR2_X1    g03304(.A1(new_n3495_), .A2(new_n2912_), .ZN(new_n3497_));
  OAI21_X1   g03305(.A1(new_n3496_), .A2(new_n3497_), .B(\asqrt[42] ), .ZN(new_n3498_));
  AOI21_X1   g03306(.A1(new_n3483_), .A2(new_n3498_), .B(new_n2464_), .ZN(new_n3499_));
  NOR2_X1    g03307(.A1(new_n3486_), .A2(new_n3499_), .ZN(new_n3500_));
  AOI21_X1   g03308(.A1(new_n3500_), .A2(new_n2271_), .B(new_n3457_), .ZN(new_n3501_));
  OAI21_X1   g03309(.A1(new_n3486_), .A2(new_n3499_), .B(\asqrt[44] ), .ZN(new_n3502_));
  NAND2_X1   g03310(.A1(new_n3502_), .A2(new_n2072_), .ZN(new_n3503_));
  OAI21_X1   g03311(.A1(new_n3501_), .A2(new_n3503_), .B(new_n3454_), .ZN(new_n3504_));
  INV_X1     g03312(.I(new_n3502_), .ZN(new_n3505_));
  OAI21_X1   g03313(.A1(new_n3501_), .A2(new_n3505_), .B(\asqrt[45] ), .ZN(new_n3506_));
  NAND3_X1   g03314(.A1(new_n3504_), .A2(new_n3506_), .A3(new_n1884_), .ZN(new_n3507_));
  NAND2_X1   g03315(.A1(new_n3507_), .A2(new_n3451_), .ZN(new_n3508_));
  NAND2_X1   g03316(.A1(new_n3504_), .A2(new_n3506_), .ZN(new_n3509_));
  AOI21_X1   g03317(.A1(new_n3509_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n3510_));
  AOI21_X1   g03318(.A1(new_n3510_), .A2(new_n3508_), .B(new_n3448_), .ZN(new_n3511_));
  INV_X1     g03319(.I(new_n3454_), .ZN(new_n3512_));
  NOR2_X1    g03320(.A1(new_n3496_), .A2(new_n3497_), .ZN(new_n3513_));
  INV_X1     g03321(.I(new_n3482_), .ZN(new_n3514_));
  AOI21_X1   g03322(.A1(new_n3513_), .A2(new_n2699_), .B(new_n3514_), .ZN(new_n3515_));
  NAND2_X1   g03323(.A1(new_n3498_), .A2(new_n2464_), .ZN(new_n3516_));
  OAI21_X1   g03324(.A1(new_n3515_), .A2(new_n3516_), .B(new_n3460_), .ZN(new_n3517_));
  INV_X1     g03325(.I(new_n3498_), .ZN(new_n3518_));
  OAI21_X1   g03326(.A1(new_n3515_), .A2(new_n3518_), .B(\asqrt[43] ), .ZN(new_n3519_));
  NAND3_X1   g03327(.A1(new_n3517_), .A2(new_n3519_), .A3(new_n2271_), .ZN(new_n3520_));
  NAND2_X1   g03328(.A1(new_n3520_), .A2(new_n3456_), .ZN(new_n3521_));
  NAND2_X1   g03329(.A1(new_n3517_), .A2(new_n3519_), .ZN(new_n3522_));
  AOI21_X1   g03330(.A1(new_n3522_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n3523_));
  AOI21_X1   g03331(.A1(new_n3523_), .A2(new_n3521_), .B(new_n3512_), .ZN(new_n3524_));
  AOI21_X1   g03332(.A1(new_n3521_), .A2(new_n3502_), .B(new_n2072_), .ZN(new_n3525_));
  OAI21_X1   g03333(.A1(new_n3524_), .A2(new_n3525_), .B(\asqrt[46] ), .ZN(new_n3526_));
  AOI21_X1   g03334(.A1(new_n3508_), .A2(new_n3526_), .B(new_n1688_), .ZN(new_n3527_));
  NOR2_X1    g03335(.A1(new_n3511_), .A2(new_n3527_), .ZN(new_n3528_));
  AOI21_X1   g03336(.A1(new_n3528_), .A2(new_n1533_), .B(new_n3445_), .ZN(new_n3529_));
  OAI21_X1   g03337(.A1(new_n3511_), .A2(new_n3527_), .B(\asqrt[48] ), .ZN(new_n3530_));
  NAND2_X1   g03338(.A1(new_n3530_), .A2(new_n1368_), .ZN(new_n3531_));
  OAI21_X1   g03339(.A1(new_n3529_), .A2(new_n3531_), .B(new_n3441_), .ZN(new_n3532_));
  INV_X1     g03340(.I(new_n3530_), .ZN(new_n3533_));
  OAI21_X1   g03341(.A1(new_n3529_), .A2(new_n3533_), .B(\asqrt[49] ), .ZN(new_n3534_));
  NAND3_X1   g03342(.A1(new_n3532_), .A2(new_n3534_), .A3(new_n1228_), .ZN(new_n3535_));
  NAND2_X1   g03343(.A1(new_n3535_), .A2(new_n3439_), .ZN(new_n3536_));
  NAND2_X1   g03344(.A1(new_n3532_), .A2(new_n3534_), .ZN(new_n3537_));
  AOI21_X1   g03345(.A1(new_n3537_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n3538_));
  AOI21_X1   g03346(.A1(new_n3538_), .A2(new_n3536_), .B(new_n3436_), .ZN(new_n3539_));
  INV_X1     g03347(.I(new_n3441_), .ZN(new_n3540_));
  INV_X1     g03348(.I(new_n3451_), .ZN(new_n3541_));
  NOR2_X1    g03349(.A1(new_n3524_), .A2(new_n3525_), .ZN(new_n3542_));
  AOI21_X1   g03350(.A1(new_n3542_), .A2(new_n1884_), .B(new_n3541_), .ZN(new_n3543_));
  NAND2_X1   g03351(.A1(new_n3526_), .A2(new_n1688_), .ZN(new_n3544_));
  OAI21_X1   g03352(.A1(new_n3543_), .A2(new_n3544_), .B(new_n3447_), .ZN(new_n3545_));
  INV_X1     g03353(.I(new_n3526_), .ZN(new_n3546_));
  OAI21_X1   g03354(.A1(new_n3543_), .A2(new_n3546_), .B(\asqrt[47] ), .ZN(new_n3547_));
  NAND3_X1   g03355(.A1(new_n3545_), .A2(new_n3547_), .A3(new_n1533_), .ZN(new_n3548_));
  NAND2_X1   g03356(.A1(new_n3548_), .A2(new_n3444_), .ZN(new_n3549_));
  NAND2_X1   g03357(.A1(new_n3545_), .A2(new_n3547_), .ZN(new_n3550_));
  AOI21_X1   g03358(.A1(new_n3550_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n3551_));
  AOI21_X1   g03359(.A1(new_n3551_), .A2(new_n3549_), .B(new_n3540_), .ZN(new_n3552_));
  AOI21_X1   g03360(.A1(new_n3549_), .A2(new_n3530_), .B(new_n1368_), .ZN(new_n3553_));
  OAI21_X1   g03361(.A1(new_n3552_), .A2(new_n3553_), .B(\asqrt[50] ), .ZN(new_n3554_));
  AOI21_X1   g03362(.A1(new_n3536_), .A2(new_n3554_), .B(new_n1088_), .ZN(new_n3555_));
  NOR2_X1    g03363(.A1(new_n3539_), .A2(new_n3555_), .ZN(new_n3556_));
  AOI21_X1   g03364(.A1(new_n3556_), .A2(new_n962_), .B(new_n3433_), .ZN(new_n3557_));
  OAI21_X1   g03365(.A1(new_n3539_), .A2(new_n3555_), .B(\asqrt[52] ), .ZN(new_n3558_));
  NAND2_X1   g03366(.A1(new_n3558_), .A2(new_n842_), .ZN(new_n3559_));
  OAI21_X1   g03367(.A1(new_n3557_), .A2(new_n3559_), .B(new_n3429_), .ZN(new_n3560_));
  INV_X1     g03368(.I(new_n3558_), .ZN(new_n3561_));
  OAI21_X1   g03369(.A1(new_n3557_), .A2(new_n3561_), .B(\asqrt[53] ), .ZN(new_n3562_));
  NAND3_X1   g03370(.A1(new_n3560_), .A2(new_n3562_), .A3(new_n720_), .ZN(new_n3563_));
  NAND2_X1   g03371(.A1(new_n3563_), .A2(new_n3427_), .ZN(new_n3564_));
  NAND2_X1   g03372(.A1(new_n3560_), .A2(new_n3562_), .ZN(new_n3565_));
  AOI21_X1   g03373(.A1(new_n3565_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n3566_));
  AOI21_X1   g03374(.A1(new_n3566_), .A2(new_n3564_), .B(new_n3424_), .ZN(new_n3567_));
  INV_X1     g03375(.I(new_n3429_), .ZN(new_n3568_));
  INV_X1     g03376(.I(new_n3439_), .ZN(new_n3569_));
  NOR2_X1    g03377(.A1(new_n3552_), .A2(new_n3553_), .ZN(new_n3570_));
  AOI21_X1   g03378(.A1(new_n3570_), .A2(new_n1228_), .B(new_n3569_), .ZN(new_n3571_));
  NAND2_X1   g03379(.A1(new_n3554_), .A2(new_n1088_), .ZN(new_n3572_));
  OAI21_X1   g03380(.A1(new_n3571_), .A2(new_n3572_), .B(new_n3435_), .ZN(new_n3573_));
  INV_X1     g03381(.I(new_n3554_), .ZN(new_n3574_));
  OAI21_X1   g03382(.A1(new_n3571_), .A2(new_n3574_), .B(\asqrt[51] ), .ZN(new_n3575_));
  NAND3_X1   g03383(.A1(new_n3573_), .A2(new_n3575_), .A3(new_n962_), .ZN(new_n3576_));
  NAND2_X1   g03384(.A1(new_n3576_), .A2(new_n3432_), .ZN(new_n3577_));
  NAND2_X1   g03385(.A1(new_n3573_), .A2(new_n3575_), .ZN(new_n3578_));
  AOI21_X1   g03386(.A1(new_n3578_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n3579_));
  AOI21_X1   g03387(.A1(new_n3579_), .A2(new_n3577_), .B(new_n3568_), .ZN(new_n3580_));
  AOI21_X1   g03388(.A1(new_n3577_), .A2(new_n3558_), .B(new_n842_), .ZN(new_n3581_));
  OAI21_X1   g03389(.A1(new_n3580_), .A2(new_n3581_), .B(\asqrt[54] ), .ZN(new_n3582_));
  AOI21_X1   g03390(.A1(new_n3564_), .A2(new_n3582_), .B(new_n630_), .ZN(new_n3583_));
  NOR2_X1    g03391(.A1(new_n3567_), .A2(new_n3583_), .ZN(new_n3584_));
  AOI21_X1   g03392(.A1(new_n3584_), .A2(new_n545_), .B(new_n3421_), .ZN(new_n3585_));
  OAI21_X1   g03393(.A1(new_n3567_), .A2(new_n3583_), .B(\asqrt[56] ), .ZN(new_n3586_));
  NAND2_X1   g03394(.A1(new_n3586_), .A2(new_n450_), .ZN(new_n3587_));
  OAI21_X1   g03395(.A1(new_n3585_), .A2(new_n3587_), .B(new_n3417_), .ZN(new_n3588_));
  INV_X1     g03396(.I(new_n3586_), .ZN(new_n3589_));
  OAI21_X1   g03397(.A1(new_n3585_), .A2(new_n3589_), .B(\asqrt[57] ), .ZN(new_n3590_));
  NAND3_X1   g03398(.A1(new_n3588_), .A2(new_n3590_), .A3(new_n403_), .ZN(new_n3591_));
  INV_X1     g03399(.I(new_n3417_), .ZN(new_n3592_));
  INV_X1     g03400(.I(new_n3427_), .ZN(new_n3593_));
  NOR2_X1    g03401(.A1(new_n3580_), .A2(new_n3581_), .ZN(new_n3594_));
  AOI21_X1   g03402(.A1(new_n3594_), .A2(new_n720_), .B(new_n3593_), .ZN(new_n3595_));
  NAND2_X1   g03403(.A1(new_n3582_), .A2(new_n630_), .ZN(new_n3596_));
  OAI21_X1   g03404(.A1(new_n3595_), .A2(new_n3596_), .B(new_n3423_), .ZN(new_n3597_));
  INV_X1     g03405(.I(new_n3582_), .ZN(new_n3598_));
  OAI21_X1   g03406(.A1(new_n3595_), .A2(new_n3598_), .B(\asqrt[55] ), .ZN(new_n3599_));
  NAND3_X1   g03407(.A1(new_n3597_), .A2(new_n3599_), .A3(new_n545_), .ZN(new_n3600_));
  NAND2_X1   g03408(.A1(new_n3600_), .A2(new_n3420_), .ZN(new_n3601_));
  NAND2_X1   g03409(.A1(new_n3597_), .A2(new_n3599_), .ZN(new_n3602_));
  AOI21_X1   g03410(.A1(new_n3602_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n3603_));
  AOI21_X1   g03411(.A1(new_n3603_), .A2(new_n3601_), .B(new_n3592_), .ZN(new_n3604_));
  AOI21_X1   g03412(.A1(new_n3601_), .A2(new_n3586_), .B(new_n450_), .ZN(new_n3605_));
  OAI21_X1   g03413(.A1(new_n3604_), .A2(new_n3605_), .B(\asqrt[58] ), .ZN(new_n3606_));
  NAND2_X1   g03414(.A1(new_n3397_), .A2(new_n3172_), .ZN(new_n3607_));
  NOR2_X1    g03415(.A1(new_n3400_), .A2(new_n3172_), .ZN(new_n3608_));
  NAND2_X1   g03416(.A1(new_n3608_), .A2(new_n3412_), .ZN(new_n3609_));
  AOI21_X1   g03417(.A1(new_n3609_), .A2(new_n3607_), .B(new_n193_), .ZN(new_n3610_));
  INV_X1     g03418(.I(new_n3610_), .ZN(new_n3611_));
  NAND3_X1   g03419(.A1(\asqrt[39] ), .A2(new_n3382_), .A3(new_n3393_), .ZN(new_n3612_));
  XOR2_X1    g03420(.A1(new_n3612_), .A2(new_n3385_), .Z(new_n3613_));
  AOI21_X1   g03421(.A1(new_n3608_), .A2(new_n3397_), .B(new_n3398_), .ZN(new_n3614_));
  OAI21_X1   g03422(.A1(new_n3352_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n3615_));
  NOR2_X1    g03423(.A1(new_n3400_), .A2(new_n3615_), .ZN(new_n3616_));
  XOR2_X1    g03424(.A1(new_n3616_), .A2(new_n3180_), .Z(new_n3617_));
  NAND3_X1   g03425(.A1(\asqrt[39] ), .A2(new_n3368_), .A3(new_n3353_), .ZN(new_n3618_));
  XOR2_X1    g03426(.A1(new_n3618_), .A2(new_n3184_), .Z(new_n3619_));
  NOR2_X1    g03427(.A1(new_n3604_), .A2(new_n3605_), .ZN(new_n3620_));
  AOI21_X1   g03428(.A1(new_n3620_), .A2(new_n403_), .B(new_n3404_), .ZN(new_n3621_));
  NAND2_X1   g03429(.A1(new_n3606_), .A2(new_n339_), .ZN(new_n3622_));
  OAI21_X1   g03430(.A1(new_n3621_), .A2(new_n3622_), .B(new_n3619_), .ZN(new_n3623_));
  INV_X1     g03431(.I(new_n3606_), .ZN(new_n3624_));
  OAI21_X1   g03432(.A1(new_n3621_), .A2(new_n3624_), .B(\asqrt[59] ), .ZN(new_n3625_));
  NAND3_X1   g03433(.A1(new_n3623_), .A2(new_n3625_), .A3(new_n288_), .ZN(new_n3626_));
  NAND2_X1   g03434(.A1(new_n3626_), .A2(new_n3617_), .ZN(new_n3627_));
  INV_X1     g03435(.I(new_n3619_), .ZN(new_n3628_));
  NAND2_X1   g03436(.A1(new_n3591_), .A2(new_n3403_), .ZN(new_n3629_));
  NAND2_X1   g03437(.A1(new_n3588_), .A2(new_n3590_), .ZN(new_n3630_));
  AOI21_X1   g03438(.A1(new_n3630_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n3631_));
  AOI21_X1   g03439(.A1(new_n3631_), .A2(new_n3629_), .B(new_n3628_), .ZN(new_n3632_));
  AOI21_X1   g03440(.A1(new_n3629_), .A2(new_n3606_), .B(new_n339_), .ZN(new_n3633_));
  OAI21_X1   g03441(.A1(new_n3632_), .A2(new_n3633_), .B(\asqrt[60] ), .ZN(new_n3634_));
  AOI21_X1   g03442(.A1(new_n3627_), .A2(new_n3634_), .B(new_n242_), .ZN(new_n3635_));
  NAND3_X1   g03443(.A1(\asqrt[39] ), .A2(new_n3358_), .A3(new_n3374_), .ZN(new_n3636_));
  XOR2_X1    g03444(.A1(new_n3636_), .A2(new_n3386_), .Z(new_n3637_));
  INV_X1     g03445(.I(new_n3637_), .ZN(new_n3638_));
  NAND2_X1   g03446(.A1(new_n3623_), .A2(new_n3625_), .ZN(new_n3639_));
  AOI21_X1   g03447(.A1(new_n3639_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n3640_));
  AOI21_X1   g03448(.A1(new_n3640_), .A2(new_n3627_), .B(new_n3638_), .ZN(new_n3641_));
  OAI21_X1   g03449(.A1(new_n3641_), .A2(new_n3635_), .B(\asqrt[62] ), .ZN(new_n3642_));
  INV_X1     g03450(.I(new_n3642_), .ZN(new_n3643_));
  NOR2_X1    g03451(.A1(new_n3641_), .A2(new_n3635_), .ZN(new_n3644_));
  AOI21_X1   g03452(.A1(new_n3359_), .A2(new_n3380_), .B(new_n3375_), .ZN(new_n3645_));
  NAND2_X1   g03453(.A1(\asqrt[39] ), .A2(new_n3645_), .ZN(new_n3646_));
  XOR2_X1    g03454(.A1(new_n3646_), .A2(new_n3378_), .Z(new_n3647_));
  INV_X1     g03455(.I(new_n3647_), .ZN(new_n3648_));
  AOI21_X1   g03456(.A1(new_n3644_), .A2(new_n234_), .B(new_n3648_), .ZN(new_n3649_));
  OAI21_X1   g03457(.A1(new_n3649_), .A2(new_n3643_), .B(new_n3614_), .ZN(new_n3650_));
  OAI21_X1   g03458(.A1(new_n3650_), .A2(new_n3613_), .B(new_n193_), .ZN(new_n3651_));
  NOR2_X1    g03459(.A1(new_n3649_), .A2(new_n3643_), .ZN(new_n3652_));
  NAND2_X1   g03460(.A1(new_n3652_), .A2(new_n3613_), .ZN(new_n3653_));
  NOR2_X1    g03461(.A1(\asqrt[39] ), .A2(new_n3173_), .ZN(new_n3654_));
  INV_X1     g03462(.I(new_n3654_), .ZN(new_n3655_));
  NAND4_X1   g03463(.A1(new_n3651_), .A2(new_n3611_), .A3(new_n3653_), .A4(new_n3655_), .ZN(\asqrt[38] ));
  NAND3_X1   g03464(.A1(\asqrt[38] ), .A2(new_n3591_), .A3(new_n3606_), .ZN(new_n3657_));
  XOR2_X1    g03465(.A1(new_n3657_), .A2(new_n3404_), .Z(new_n3658_));
  INV_X1     g03466(.I(new_n3617_), .ZN(new_n3659_));
  NOR2_X1    g03467(.A1(new_n3632_), .A2(new_n3633_), .ZN(new_n3660_));
  AOI21_X1   g03468(.A1(new_n3660_), .A2(new_n288_), .B(new_n3659_), .ZN(new_n3661_));
  INV_X1     g03469(.I(new_n3634_), .ZN(new_n3662_));
  OAI21_X1   g03470(.A1(new_n3661_), .A2(new_n3662_), .B(\asqrt[61] ), .ZN(new_n3663_));
  NAND2_X1   g03471(.A1(new_n3634_), .A2(new_n242_), .ZN(new_n3664_));
  OAI21_X1   g03472(.A1(new_n3661_), .A2(new_n3664_), .B(new_n3637_), .ZN(new_n3665_));
  NAND3_X1   g03473(.A1(new_n3665_), .A2(new_n3663_), .A3(new_n234_), .ZN(new_n3666_));
  NAND2_X1   g03474(.A1(new_n3666_), .A2(new_n3647_), .ZN(new_n3667_));
  NAND2_X1   g03475(.A1(new_n3667_), .A2(new_n3642_), .ZN(new_n3668_));
  NAND2_X1   g03476(.A1(new_n3668_), .A2(new_n3613_), .ZN(new_n3669_));
  INV_X1     g03477(.I(new_n3613_), .ZN(new_n3670_));
  INV_X1     g03478(.I(new_n3614_), .ZN(new_n3671_));
  AOI21_X1   g03479(.A1(new_n3667_), .A2(new_n3642_), .B(new_n3671_), .ZN(new_n3672_));
  AOI21_X1   g03480(.A1(new_n3672_), .A2(new_n3670_), .B(\asqrt[63] ), .ZN(new_n3673_));
  NOR2_X1    g03481(.A1(new_n3668_), .A2(new_n3670_), .ZN(new_n3674_));
  NOR4_X1    g03482(.A1(new_n3673_), .A2(new_n3610_), .A3(new_n3674_), .A4(new_n3654_), .ZN(new_n3675_));
  NOR2_X1    g03483(.A1(new_n3675_), .A2(new_n3613_), .ZN(new_n3676_));
  NAND2_X1   g03484(.A1(new_n3676_), .A2(new_n3652_), .ZN(new_n3677_));
  AOI21_X1   g03485(.A1(new_n3677_), .A2(new_n3669_), .B(new_n193_), .ZN(new_n3678_));
  NAND3_X1   g03486(.A1(\asqrt[38] ), .A2(new_n3642_), .A3(new_n3666_), .ZN(new_n3679_));
  XOR2_X1    g03487(.A1(new_n3679_), .A2(new_n3647_), .Z(new_n3680_));
  INV_X1     g03488(.I(new_n3680_), .ZN(new_n3681_));
  AOI21_X1   g03489(.A1(new_n3676_), .A2(new_n3668_), .B(new_n3674_), .ZN(new_n3682_));
  INV_X1     g03490(.I(new_n3682_), .ZN(new_n3683_));
  OAI21_X1   g03491(.A1(new_n3621_), .A2(new_n3622_), .B(new_n3625_), .ZN(new_n3684_));
  NOR2_X1    g03492(.A1(new_n3675_), .A2(new_n3684_), .ZN(new_n3685_));
  XOR2_X1    g03493(.A1(new_n3685_), .A2(new_n3619_), .Z(new_n3686_));
  OAI21_X1   g03494(.A1(new_n3585_), .A2(new_n3587_), .B(new_n3590_), .ZN(new_n3687_));
  NOR2_X1    g03495(.A1(new_n3675_), .A2(new_n3687_), .ZN(new_n3688_));
  XOR2_X1    g03496(.A1(new_n3688_), .A2(new_n3417_), .Z(new_n3689_));
  INV_X1     g03497(.I(new_n3689_), .ZN(new_n3690_));
  NAND3_X1   g03498(.A1(\asqrt[38] ), .A2(new_n3600_), .A3(new_n3586_), .ZN(new_n3691_));
  XOR2_X1    g03499(.A1(new_n3691_), .A2(new_n3421_), .Z(new_n3692_));
  INV_X1     g03500(.I(new_n3692_), .ZN(new_n3693_));
  OAI21_X1   g03501(.A1(new_n3595_), .A2(new_n3596_), .B(new_n3599_), .ZN(new_n3694_));
  NOR2_X1    g03502(.A1(new_n3675_), .A2(new_n3694_), .ZN(new_n3695_));
  XOR2_X1    g03503(.A1(new_n3695_), .A2(new_n3423_), .Z(new_n3696_));
  NAND3_X1   g03504(.A1(\asqrt[38] ), .A2(new_n3563_), .A3(new_n3582_), .ZN(new_n3697_));
  XOR2_X1    g03505(.A1(new_n3697_), .A2(new_n3593_), .Z(new_n3698_));
  OAI21_X1   g03506(.A1(new_n3557_), .A2(new_n3559_), .B(new_n3562_), .ZN(new_n3699_));
  NOR2_X1    g03507(.A1(new_n3675_), .A2(new_n3699_), .ZN(new_n3700_));
  XOR2_X1    g03508(.A1(new_n3700_), .A2(new_n3429_), .Z(new_n3701_));
  INV_X1     g03509(.I(new_n3701_), .ZN(new_n3702_));
  NAND3_X1   g03510(.A1(\asqrt[38] ), .A2(new_n3576_), .A3(new_n3558_), .ZN(new_n3703_));
  XOR2_X1    g03511(.A1(new_n3703_), .A2(new_n3433_), .Z(new_n3704_));
  INV_X1     g03512(.I(new_n3704_), .ZN(new_n3705_));
  OAI21_X1   g03513(.A1(new_n3571_), .A2(new_n3572_), .B(new_n3575_), .ZN(new_n3706_));
  NOR2_X1    g03514(.A1(new_n3675_), .A2(new_n3706_), .ZN(new_n3707_));
  XOR2_X1    g03515(.A1(new_n3707_), .A2(new_n3435_), .Z(new_n3708_));
  NAND3_X1   g03516(.A1(\asqrt[38] ), .A2(new_n3535_), .A3(new_n3554_), .ZN(new_n3709_));
  XOR2_X1    g03517(.A1(new_n3709_), .A2(new_n3569_), .Z(new_n3710_));
  OAI21_X1   g03518(.A1(new_n3529_), .A2(new_n3531_), .B(new_n3534_), .ZN(new_n3711_));
  NOR2_X1    g03519(.A1(new_n3675_), .A2(new_n3711_), .ZN(new_n3712_));
  XOR2_X1    g03520(.A1(new_n3712_), .A2(new_n3441_), .Z(new_n3713_));
  INV_X1     g03521(.I(new_n3713_), .ZN(new_n3714_));
  NAND3_X1   g03522(.A1(\asqrt[38] ), .A2(new_n3548_), .A3(new_n3530_), .ZN(new_n3715_));
  XOR2_X1    g03523(.A1(new_n3715_), .A2(new_n3445_), .Z(new_n3716_));
  INV_X1     g03524(.I(new_n3716_), .ZN(new_n3717_));
  OAI21_X1   g03525(.A1(new_n3543_), .A2(new_n3544_), .B(new_n3547_), .ZN(new_n3718_));
  NOR2_X1    g03526(.A1(new_n3675_), .A2(new_n3718_), .ZN(new_n3719_));
  XOR2_X1    g03527(.A1(new_n3719_), .A2(new_n3447_), .Z(new_n3720_));
  NAND3_X1   g03528(.A1(\asqrt[38] ), .A2(new_n3507_), .A3(new_n3526_), .ZN(new_n3721_));
  XOR2_X1    g03529(.A1(new_n3721_), .A2(new_n3541_), .Z(new_n3722_));
  OAI21_X1   g03530(.A1(new_n3501_), .A2(new_n3503_), .B(new_n3506_), .ZN(new_n3723_));
  NOR2_X1    g03531(.A1(new_n3675_), .A2(new_n3723_), .ZN(new_n3724_));
  XOR2_X1    g03532(.A1(new_n3724_), .A2(new_n3454_), .Z(new_n3725_));
  INV_X1     g03533(.I(new_n3725_), .ZN(new_n3726_));
  NAND3_X1   g03534(.A1(\asqrt[38] ), .A2(new_n3520_), .A3(new_n3502_), .ZN(new_n3727_));
  XOR2_X1    g03535(.A1(new_n3727_), .A2(new_n3457_), .Z(new_n3728_));
  INV_X1     g03536(.I(new_n3728_), .ZN(new_n3729_));
  OAI21_X1   g03537(.A1(new_n3515_), .A2(new_n3516_), .B(new_n3519_), .ZN(new_n3730_));
  NOR2_X1    g03538(.A1(new_n3675_), .A2(new_n3730_), .ZN(new_n3731_));
  XOR2_X1    g03539(.A1(new_n3731_), .A2(new_n3460_), .Z(new_n3732_));
  NAND3_X1   g03540(.A1(\asqrt[38] ), .A2(new_n3480_), .A3(new_n3498_), .ZN(new_n3733_));
  XOR2_X1    g03541(.A1(new_n3733_), .A2(new_n3514_), .Z(new_n3734_));
  NOR2_X1    g03542(.A1(new_n3477_), .A2(\asqrt[41] ), .ZN(new_n3735_));
  NOR3_X1    g03543(.A1(new_n3675_), .A2(new_n3735_), .A3(new_n3497_), .ZN(new_n3736_));
  XOR2_X1    g03544(.A1(new_n3736_), .A2(new_n3468_), .Z(new_n3737_));
  INV_X1     g03545(.I(new_n3737_), .ZN(new_n3738_));
  NAND3_X1   g03546(.A1(\asqrt[38] ), .A2(new_n3469_), .A3(new_n3470_), .ZN(new_n3739_));
  NOR4_X1    g03547(.A1(new_n3673_), .A2(new_n3400_), .A3(new_n3610_), .A4(new_n3674_), .ZN(new_n3740_));
  INV_X1     g03548(.I(new_n3740_), .ZN(new_n3741_));
  AOI21_X1   g03549(.A1(new_n3739_), .A2(new_n3741_), .B(\a[78] ), .ZN(new_n3742_));
  NOR3_X1    g03550(.A1(new_n3675_), .A2(\a[76] ), .A3(\a[77] ), .ZN(new_n3743_));
  NOR3_X1    g03551(.A1(new_n3743_), .A2(new_n3232_), .A3(new_n3740_), .ZN(new_n3744_));
  NOR2_X1    g03552(.A1(new_n3744_), .A2(new_n3742_), .ZN(new_n3745_));
  INV_X1     g03553(.I(\a[74] ), .ZN(new_n3746_));
  INV_X1     g03554(.I(\a[75] ), .ZN(new_n3747_));
  NAND3_X1   g03555(.A1(new_n3746_), .A2(new_n3747_), .A3(new_n3469_), .ZN(new_n3748_));
  OAI21_X1   g03556(.A1(new_n3675_), .A2(new_n3469_), .B(new_n3748_), .ZN(new_n3749_));
  NAND2_X1   g03557(.A1(new_n3749_), .A2(\asqrt[39] ), .ZN(new_n3750_));
  OAI21_X1   g03558(.A1(new_n3675_), .A2(\a[76] ), .B(\a[77] ), .ZN(new_n3751_));
  NAND2_X1   g03559(.A1(new_n3751_), .A2(new_n3739_), .ZN(new_n3752_));
  NOR2_X1    g03560(.A1(new_n3749_), .A2(\asqrt[39] ), .ZN(new_n3753_));
  OAI21_X1   g03561(.A1(new_n3752_), .A2(new_n3753_), .B(new_n3750_), .ZN(new_n3754_));
  OAI21_X1   g03562(.A1(new_n3754_), .A2(\asqrt[40] ), .B(new_n3745_), .ZN(new_n3755_));
  NAND2_X1   g03563(.A1(new_n3754_), .A2(\asqrt[40] ), .ZN(new_n3756_));
  NAND3_X1   g03564(.A1(new_n3755_), .A2(new_n2912_), .A3(new_n3756_), .ZN(new_n3757_));
  NOR3_X1    g03565(.A1(new_n3675_), .A2(new_n3491_), .A3(new_n3476_), .ZN(new_n3758_));
  XOR2_X1    g03566(.A1(new_n3758_), .A2(new_n3493_), .Z(new_n3759_));
  AOI21_X1   g03567(.A1(new_n3755_), .A2(new_n3756_), .B(new_n2912_), .ZN(new_n3760_));
  AOI21_X1   g03568(.A1(new_n3757_), .A2(new_n3759_), .B(new_n3760_), .ZN(new_n3761_));
  AOI21_X1   g03569(.A1(new_n3761_), .A2(new_n2699_), .B(new_n3738_), .ZN(new_n3762_));
  OAI21_X1   g03570(.A1(new_n3761_), .A2(new_n2699_), .B(new_n2464_), .ZN(new_n3763_));
  OAI21_X1   g03571(.A1(new_n3762_), .A2(new_n3763_), .B(new_n3734_), .ZN(new_n3764_));
  NOR2_X1    g03572(.A1(new_n3761_), .A2(new_n2699_), .ZN(new_n3765_));
  OAI21_X1   g03573(.A1(new_n3762_), .A2(new_n3765_), .B(\asqrt[43] ), .ZN(new_n3766_));
  NAND3_X1   g03574(.A1(new_n3764_), .A2(new_n3766_), .A3(new_n2271_), .ZN(new_n3767_));
  NAND2_X1   g03575(.A1(new_n3767_), .A2(new_n3732_), .ZN(new_n3768_));
  NAND2_X1   g03576(.A1(new_n3764_), .A2(new_n3766_), .ZN(new_n3769_));
  AOI21_X1   g03577(.A1(new_n3769_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n3770_));
  AOI21_X1   g03578(.A1(new_n3770_), .A2(new_n3768_), .B(new_n3729_), .ZN(new_n3771_));
  INV_X1     g03579(.I(new_n3734_), .ZN(new_n3772_));
  OAI21_X1   g03580(.A1(new_n3743_), .A2(new_n3740_), .B(new_n3232_), .ZN(new_n3773_));
  NAND3_X1   g03581(.A1(new_n3739_), .A2(new_n3741_), .A3(\a[78] ), .ZN(new_n3774_));
  NAND2_X1   g03582(.A1(new_n3773_), .A2(new_n3774_), .ZN(new_n3775_));
  NAND2_X1   g03583(.A1(\asqrt[38] ), .A2(\a[76] ), .ZN(new_n3776_));
  AOI21_X1   g03584(.A1(new_n3776_), .A2(new_n3748_), .B(new_n3400_), .ZN(new_n3777_));
  AOI21_X1   g03585(.A1(\asqrt[38] ), .A2(new_n3469_), .B(new_n3470_), .ZN(new_n3778_));
  NOR2_X1    g03586(.A1(new_n3743_), .A2(new_n3778_), .ZN(new_n3779_));
  NAND3_X1   g03587(.A1(new_n3776_), .A2(new_n3400_), .A3(new_n3748_), .ZN(new_n3780_));
  AOI21_X1   g03588(.A1(new_n3779_), .A2(new_n3780_), .B(new_n3777_), .ZN(new_n3781_));
  AOI21_X1   g03589(.A1(new_n3781_), .A2(new_n3167_), .B(new_n3775_), .ZN(new_n3782_));
  NOR2_X1    g03590(.A1(new_n3781_), .A2(new_n3167_), .ZN(new_n3783_));
  NOR3_X1    g03591(.A1(new_n3782_), .A2(\asqrt[41] ), .A3(new_n3783_), .ZN(new_n3784_));
  INV_X1     g03592(.I(new_n3759_), .ZN(new_n3785_));
  OAI21_X1   g03593(.A1(new_n3782_), .A2(new_n3783_), .B(\asqrt[41] ), .ZN(new_n3786_));
  OAI21_X1   g03594(.A1(new_n3784_), .A2(new_n3785_), .B(new_n3786_), .ZN(new_n3787_));
  OAI21_X1   g03595(.A1(new_n3787_), .A2(\asqrt[42] ), .B(new_n3737_), .ZN(new_n3788_));
  AOI21_X1   g03596(.A1(new_n3787_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n3789_));
  AOI21_X1   g03597(.A1(new_n3789_), .A2(new_n3788_), .B(new_n3772_), .ZN(new_n3790_));
  NAND2_X1   g03598(.A1(new_n3787_), .A2(\asqrt[42] ), .ZN(new_n3791_));
  AOI21_X1   g03599(.A1(new_n3788_), .A2(new_n3791_), .B(new_n2464_), .ZN(new_n3792_));
  OAI21_X1   g03600(.A1(new_n3790_), .A2(new_n3792_), .B(\asqrt[44] ), .ZN(new_n3793_));
  AOI21_X1   g03601(.A1(new_n3768_), .A2(new_n3793_), .B(new_n2072_), .ZN(new_n3794_));
  NOR2_X1    g03602(.A1(new_n3771_), .A2(new_n3794_), .ZN(new_n3795_));
  AOI21_X1   g03603(.A1(new_n3795_), .A2(new_n1884_), .B(new_n3726_), .ZN(new_n3796_));
  OAI21_X1   g03604(.A1(new_n3771_), .A2(new_n3794_), .B(\asqrt[46] ), .ZN(new_n3797_));
  NAND2_X1   g03605(.A1(new_n3797_), .A2(new_n1688_), .ZN(new_n3798_));
  OAI21_X1   g03606(.A1(new_n3796_), .A2(new_n3798_), .B(new_n3722_), .ZN(new_n3799_));
  INV_X1     g03607(.I(new_n3797_), .ZN(new_n3800_));
  OAI21_X1   g03608(.A1(new_n3796_), .A2(new_n3800_), .B(\asqrt[47] ), .ZN(new_n3801_));
  NAND3_X1   g03609(.A1(new_n3799_), .A2(new_n3801_), .A3(new_n1533_), .ZN(new_n3802_));
  NAND2_X1   g03610(.A1(new_n3802_), .A2(new_n3720_), .ZN(new_n3803_));
  NAND2_X1   g03611(.A1(new_n3799_), .A2(new_n3801_), .ZN(new_n3804_));
  AOI21_X1   g03612(.A1(new_n3804_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n3805_));
  AOI21_X1   g03613(.A1(new_n3805_), .A2(new_n3803_), .B(new_n3717_), .ZN(new_n3806_));
  INV_X1     g03614(.I(new_n3722_), .ZN(new_n3807_));
  INV_X1     g03615(.I(new_n3732_), .ZN(new_n3808_));
  NOR2_X1    g03616(.A1(new_n3790_), .A2(new_n3792_), .ZN(new_n3809_));
  AOI21_X1   g03617(.A1(new_n3809_), .A2(new_n2271_), .B(new_n3808_), .ZN(new_n3810_));
  NAND2_X1   g03618(.A1(new_n3793_), .A2(new_n2072_), .ZN(new_n3811_));
  OAI21_X1   g03619(.A1(new_n3810_), .A2(new_n3811_), .B(new_n3728_), .ZN(new_n3812_));
  INV_X1     g03620(.I(new_n3793_), .ZN(new_n3813_));
  OAI21_X1   g03621(.A1(new_n3810_), .A2(new_n3813_), .B(\asqrt[45] ), .ZN(new_n3814_));
  NAND3_X1   g03622(.A1(new_n3812_), .A2(new_n3814_), .A3(new_n1884_), .ZN(new_n3815_));
  NAND2_X1   g03623(.A1(new_n3815_), .A2(new_n3725_), .ZN(new_n3816_));
  NAND2_X1   g03624(.A1(new_n3812_), .A2(new_n3814_), .ZN(new_n3817_));
  AOI21_X1   g03625(.A1(new_n3817_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n3818_));
  AOI21_X1   g03626(.A1(new_n3818_), .A2(new_n3816_), .B(new_n3807_), .ZN(new_n3819_));
  AOI21_X1   g03627(.A1(new_n3816_), .A2(new_n3797_), .B(new_n1688_), .ZN(new_n3820_));
  OAI21_X1   g03628(.A1(new_n3819_), .A2(new_n3820_), .B(\asqrt[48] ), .ZN(new_n3821_));
  AOI21_X1   g03629(.A1(new_n3803_), .A2(new_n3821_), .B(new_n1368_), .ZN(new_n3822_));
  NOR2_X1    g03630(.A1(new_n3806_), .A2(new_n3822_), .ZN(new_n3823_));
  AOI21_X1   g03631(.A1(new_n3823_), .A2(new_n1228_), .B(new_n3714_), .ZN(new_n3824_));
  OAI21_X1   g03632(.A1(new_n3806_), .A2(new_n3822_), .B(\asqrt[50] ), .ZN(new_n3825_));
  NAND2_X1   g03633(.A1(new_n3825_), .A2(new_n1088_), .ZN(new_n3826_));
  OAI21_X1   g03634(.A1(new_n3824_), .A2(new_n3826_), .B(new_n3710_), .ZN(new_n3827_));
  INV_X1     g03635(.I(new_n3825_), .ZN(new_n3828_));
  OAI21_X1   g03636(.A1(new_n3824_), .A2(new_n3828_), .B(\asqrt[51] ), .ZN(new_n3829_));
  NAND3_X1   g03637(.A1(new_n3827_), .A2(new_n3829_), .A3(new_n962_), .ZN(new_n3830_));
  NAND2_X1   g03638(.A1(new_n3830_), .A2(new_n3708_), .ZN(new_n3831_));
  NAND2_X1   g03639(.A1(new_n3827_), .A2(new_n3829_), .ZN(new_n3832_));
  AOI21_X1   g03640(.A1(new_n3832_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n3833_));
  AOI21_X1   g03641(.A1(new_n3833_), .A2(new_n3831_), .B(new_n3705_), .ZN(new_n3834_));
  INV_X1     g03642(.I(new_n3710_), .ZN(new_n3835_));
  INV_X1     g03643(.I(new_n3720_), .ZN(new_n3836_));
  NOR2_X1    g03644(.A1(new_n3819_), .A2(new_n3820_), .ZN(new_n3837_));
  AOI21_X1   g03645(.A1(new_n3837_), .A2(new_n1533_), .B(new_n3836_), .ZN(new_n3838_));
  NAND2_X1   g03646(.A1(new_n3821_), .A2(new_n1368_), .ZN(new_n3839_));
  OAI21_X1   g03647(.A1(new_n3838_), .A2(new_n3839_), .B(new_n3716_), .ZN(new_n3840_));
  INV_X1     g03648(.I(new_n3821_), .ZN(new_n3841_));
  OAI21_X1   g03649(.A1(new_n3838_), .A2(new_n3841_), .B(\asqrt[49] ), .ZN(new_n3842_));
  NAND3_X1   g03650(.A1(new_n3840_), .A2(new_n3842_), .A3(new_n1228_), .ZN(new_n3843_));
  NAND2_X1   g03651(.A1(new_n3843_), .A2(new_n3713_), .ZN(new_n3844_));
  NAND2_X1   g03652(.A1(new_n3840_), .A2(new_n3842_), .ZN(new_n3845_));
  AOI21_X1   g03653(.A1(new_n3845_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n3846_));
  AOI21_X1   g03654(.A1(new_n3846_), .A2(new_n3844_), .B(new_n3835_), .ZN(new_n3847_));
  AOI21_X1   g03655(.A1(new_n3844_), .A2(new_n3825_), .B(new_n1088_), .ZN(new_n3848_));
  OAI21_X1   g03656(.A1(new_n3847_), .A2(new_n3848_), .B(\asqrt[52] ), .ZN(new_n3849_));
  AOI21_X1   g03657(.A1(new_n3831_), .A2(new_n3849_), .B(new_n842_), .ZN(new_n3850_));
  NOR2_X1    g03658(.A1(new_n3834_), .A2(new_n3850_), .ZN(new_n3851_));
  AOI21_X1   g03659(.A1(new_n3851_), .A2(new_n720_), .B(new_n3702_), .ZN(new_n3852_));
  OAI21_X1   g03660(.A1(new_n3834_), .A2(new_n3850_), .B(\asqrt[54] ), .ZN(new_n3853_));
  NAND2_X1   g03661(.A1(new_n3853_), .A2(new_n630_), .ZN(new_n3854_));
  OAI21_X1   g03662(.A1(new_n3852_), .A2(new_n3854_), .B(new_n3698_), .ZN(new_n3855_));
  INV_X1     g03663(.I(new_n3853_), .ZN(new_n3856_));
  OAI21_X1   g03664(.A1(new_n3852_), .A2(new_n3856_), .B(\asqrt[55] ), .ZN(new_n3857_));
  NAND3_X1   g03665(.A1(new_n3855_), .A2(new_n3857_), .A3(new_n545_), .ZN(new_n3858_));
  NAND2_X1   g03666(.A1(new_n3858_), .A2(new_n3696_), .ZN(new_n3859_));
  NAND2_X1   g03667(.A1(new_n3855_), .A2(new_n3857_), .ZN(new_n3860_));
  AOI21_X1   g03668(.A1(new_n3860_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n3861_));
  AOI21_X1   g03669(.A1(new_n3861_), .A2(new_n3859_), .B(new_n3693_), .ZN(new_n3862_));
  INV_X1     g03670(.I(new_n3698_), .ZN(new_n3863_));
  INV_X1     g03671(.I(new_n3708_), .ZN(new_n3864_));
  NOR2_X1    g03672(.A1(new_n3847_), .A2(new_n3848_), .ZN(new_n3865_));
  AOI21_X1   g03673(.A1(new_n3865_), .A2(new_n962_), .B(new_n3864_), .ZN(new_n3866_));
  NAND2_X1   g03674(.A1(new_n3849_), .A2(new_n842_), .ZN(new_n3867_));
  OAI21_X1   g03675(.A1(new_n3866_), .A2(new_n3867_), .B(new_n3704_), .ZN(new_n3868_));
  INV_X1     g03676(.I(new_n3849_), .ZN(new_n3869_));
  OAI21_X1   g03677(.A1(new_n3866_), .A2(new_n3869_), .B(\asqrt[53] ), .ZN(new_n3870_));
  NAND3_X1   g03678(.A1(new_n3868_), .A2(new_n3870_), .A3(new_n720_), .ZN(new_n3871_));
  NAND2_X1   g03679(.A1(new_n3871_), .A2(new_n3701_), .ZN(new_n3872_));
  NAND2_X1   g03680(.A1(new_n3868_), .A2(new_n3870_), .ZN(new_n3873_));
  AOI21_X1   g03681(.A1(new_n3873_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n3874_));
  AOI21_X1   g03682(.A1(new_n3874_), .A2(new_n3872_), .B(new_n3863_), .ZN(new_n3875_));
  AOI21_X1   g03683(.A1(new_n3872_), .A2(new_n3853_), .B(new_n630_), .ZN(new_n3876_));
  OAI21_X1   g03684(.A1(new_n3875_), .A2(new_n3876_), .B(\asqrt[56] ), .ZN(new_n3877_));
  AOI21_X1   g03685(.A1(new_n3859_), .A2(new_n3877_), .B(new_n450_), .ZN(new_n3878_));
  NOR2_X1    g03686(.A1(new_n3862_), .A2(new_n3878_), .ZN(new_n3879_));
  AOI21_X1   g03687(.A1(new_n3879_), .A2(new_n403_), .B(new_n3690_), .ZN(new_n3880_));
  OAI21_X1   g03688(.A1(new_n3862_), .A2(new_n3878_), .B(\asqrt[58] ), .ZN(new_n3881_));
  NAND2_X1   g03689(.A1(new_n3881_), .A2(new_n339_), .ZN(new_n3882_));
  OAI21_X1   g03690(.A1(new_n3880_), .A2(new_n3882_), .B(new_n3658_), .ZN(new_n3883_));
  INV_X1     g03691(.I(new_n3881_), .ZN(new_n3884_));
  OAI21_X1   g03692(.A1(new_n3880_), .A2(new_n3884_), .B(\asqrt[59] ), .ZN(new_n3885_));
  NAND3_X1   g03693(.A1(new_n3883_), .A2(new_n3885_), .A3(new_n288_), .ZN(new_n3886_));
  NAND2_X1   g03694(.A1(new_n3886_), .A2(new_n3686_), .ZN(new_n3887_));
  INV_X1     g03695(.I(new_n3658_), .ZN(new_n3888_));
  INV_X1     g03696(.I(new_n3696_), .ZN(new_n3889_));
  NOR2_X1    g03697(.A1(new_n3875_), .A2(new_n3876_), .ZN(new_n3890_));
  AOI21_X1   g03698(.A1(new_n3890_), .A2(new_n545_), .B(new_n3889_), .ZN(new_n3891_));
  NAND2_X1   g03699(.A1(new_n3877_), .A2(new_n450_), .ZN(new_n3892_));
  OAI21_X1   g03700(.A1(new_n3891_), .A2(new_n3892_), .B(new_n3692_), .ZN(new_n3893_));
  INV_X1     g03701(.I(new_n3877_), .ZN(new_n3894_));
  OAI21_X1   g03702(.A1(new_n3891_), .A2(new_n3894_), .B(\asqrt[57] ), .ZN(new_n3895_));
  NAND3_X1   g03703(.A1(new_n3893_), .A2(new_n3895_), .A3(new_n403_), .ZN(new_n3896_));
  NAND2_X1   g03704(.A1(new_n3896_), .A2(new_n3689_), .ZN(new_n3897_));
  NAND2_X1   g03705(.A1(new_n3893_), .A2(new_n3895_), .ZN(new_n3898_));
  AOI21_X1   g03706(.A1(new_n3898_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n3899_));
  AOI21_X1   g03707(.A1(new_n3899_), .A2(new_n3897_), .B(new_n3888_), .ZN(new_n3900_));
  AOI21_X1   g03708(.A1(new_n3897_), .A2(new_n3881_), .B(new_n339_), .ZN(new_n3901_));
  OAI21_X1   g03709(.A1(new_n3900_), .A2(new_n3901_), .B(\asqrt[60] ), .ZN(new_n3902_));
  AOI21_X1   g03710(.A1(new_n3887_), .A2(new_n3902_), .B(new_n242_), .ZN(new_n3903_));
  NAND3_X1   g03711(.A1(\asqrt[38] ), .A2(new_n3626_), .A3(new_n3634_), .ZN(new_n3904_));
  XOR2_X1    g03712(.A1(new_n3904_), .A2(new_n3659_), .Z(new_n3905_));
  INV_X1     g03713(.I(new_n3905_), .ZN(new_n3906_));
  NAND2_X1   g03714(.A1(new_n3883_), .A2(new_n3885_), .ZN(new_n3907_));
  AOI21_X1   g03715(.A1(new_n3907_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n3908_));
  AOI21_X1   g03716(.A1(new_n3908_), .A2(new_n3887_), .B(new_n3906_), .ZN(new_n3909_));
  OAI21_X1   g03717(.A1(new_n3909_), .A2(new_n3903_), .B(\asqrt[62] ), .ZN(new_n3910_));
  AOI21_X1   g03718(.A1(new_n3627_), .A2(new_n3640_), .B(new_n3635_), .ZN(new_n3911_));
  NAND2_X1   g03719(.A1(\asqrt[38] ), .A2(new_n3911_), .ZN(new_n3912_));
  XOR2_X1    g03720(.A1(new_n3912_), .A2(new_n3638_), .Z(new_n3913_));
  INV_X1     g03721(.I(new_n3686_), .ZN(new_n3914_));
  NOR2_X1    g03722(.A1(new_n3900_), .A2(new_n3901_), .ZN(new_n3915_));
  AOI21_X1   g03723(.A1(new_n3915_), .A2(new_n288_), .B(new_n3914_), .ZN(new_n3916_));
  INV_X1     g03724(.I(new_n3902_), .ZN(new_n3917_));
  OAI21_X1   g03725(.A1(new_n3916_), .A2(new_n3917_), .B(\asqrt[61] ), .ZN(new_n3918_));
  NAND2_X1   g03726(.A1(new_n3902_), .A2(new_n242_), .ZN(new_n3919_));
  OAI21_X1   g03727(.A1(new_n3916_), .A2(new_n3919_), .B(new_n3905_), .ZN(new_n3920_));
  NAND3_X1   g03728(.A1(new_n3920_), .A2(new_n3918_), .A3(new_n234_), .ZN(new_n3921_));
  NAND2_X1   g03729(.A1(new_n3921_), .A2(new_n3913_), .ZN(new_n3922_));
  AOI21_X1   g03730(.A1(new_n3922_), .A2(new_n3910_), .B(new_n3683_), .ZN(new_n3923_));
  AOI21_X1   g03731(.A1(new_n3923_), .A2(new_n3681_), .B(\asqrt[63] ), .ZN(new_n3924_));
  NAND2_X1   g03732(.A1(new_n3922_), .A2(new_n3910_), .ZN(new_n3925_));
  NOR2_X1    g03733(.A1(new_n3925_), .A2(new_n3681_), .ZN(new_n3926_));
  NOR2_X1    g03734(.A1(\asqrt[38] ), .A2(new_n3670_), .ZN(new_n3927_));
  NOR4_X1    g03735(.A1(new_n3924_), .A2(new_n3678_), .A3(new_n3926_), .A4(new_n3927_), .ZN(new_n3928_));
  OAI21_X1   g03736(.A1(new_n3880_), .A2(new_n3882_), .B(new_n3885_), .ZN(new_n3929_));
  NOR2_X1    g03737(.A1(new_n3928_), .A2(new_n3929_), .ZN(new_n3930_));
  XOR2_X1    g03738(.A1(new_n3930_), .A2(new_n3658_), .Z(new_n3931_));
  INV_X1     g03739(.I(new_n3931_), .ZN(new_n3932_));
  INV_X1     g03740(.I(new_n3678_), .ZN(new_n3933_));
  INV_X1     g03741(.I(new_n3910_), .ZN(new_n3934_));
  NOR2_X1    g03742(.A1(new_n3909_), .A2(new_n3903_), .ZN(new_n3935_));
  INV_X1     g03743(.I(new_n3913_), .ZN(new_n3936_));
  AOI21_X1   g03744(.A1(new_n3935_), .A2(new_n234_), .B(new_n3936_), .ZN(new_n3937_));
  OAI21_X1   g03745(.A1(new_n3937_), .A2(new_n3934_), .B(new_n3682_), .ZN(new_n3938_));
  OAI21_X1   g03746(.A1(new_n3938_), .A2(new_n3680_), .B(new_n193_), .ZN(new_n3939_));
  NOR2_X1    g03747(.A1(new_n3937_), .A2(new_n3934_), .ZN(new_n3940_));
  NAND2_X1   g03748(.A1(new_n3940_), .A2(new_n3680_), .ZN(new_n3941_));
  INV_X1     g03749(.I(new_n3927_), .ZN(new_n3942_));
  NAND4_X1   g03750(.A1(new_n3939_), .A2(new_n3933_), .A3(new_n3941_), .A4(new_n3942_), .ZN(\asqrt[37] ));
  NAND3_X1   g03751(.A1(\asqrt[37] ), .A2(new_n3896_), .A3(new_n3881_), .ZN(new_n3944_));
  XOR2_X1    g03752(.A1(new_n3944_), .A2(new_n3690_), .Z(new_n3945_));
  OAI21_X1   g03753(.A1(new_n3891_), .A2(new_n3892_), .B(new_n3895_), .ZN(new_n3946_));
  NOR2_X1    g03754(.A1(new_n3928_), .A2(new_n3946_), .ZN(new_n3947_));
  XOR2_X1    g03755(.A1(new_n3947_), .A2(new_n3692_), .Z(new_n3948_));
  INV_X1     g03756(.I(new_n3948_), .ZN(new_n3949_));
  NAND3_X1   g03757(.A1(\asqrt[37] ), .A2(new_n3858_), .A3(new_n3877_), .ZN(new_n3950_));
  XOR2_X1    g03758(.A1(new_n3950_), .A2(new_n3889_), .Z(new_n3951_));
  INV_X1     g03759(.I(new_n3951_), .ZN(new_n3952_));
  OAI21_X1   g03760(.A1(new_n3852_), .A2(new_n3854_), .B(new_n3857_), .ZN(new_n3953_));
  NOR2_X1    g03761(.A1(new_n3928_), .A2(new_n3953_), .ZN(new_n3954_));
  XOR2_X1    g03762(.A1(new_n3954_), .A2(new_n3698_), .Z(new_n3955_));
  NAND3_X1   g03763(.A1(\asqrt[37] ), .A2(new_n3871_), .A3(new_n3853_), .ZN(new_n3956_));
  XOR2_X1    g03764(.A1(new_n3956_), .A2(new_n3702_), .Z(new_n3957_));
  OAI21_X1   g03765(.A1(new_n3866_), .A2(new_n3867_), .B(new_n3870_), .ZN(new_n3958_));
  NOR2_X1    g03766(.A1(new_n3928_), .A2(new_n3958_), .ZN(new_n3959_));
  XOR2_X1    g03767(.A1(new_n3959_), .A2(new_n3704_), .Z(new_n3960_));
  INV_X1     g03768(.I(new_n3960_), .ZN(new_n3961_));
  NAND3_X1   g03769(.A1(\asqrt[37] ), .A2(new_n3830_), .A3(new_n3849_), .ZN(new_n3962_));
  XOR2_X1    g03770(.A1(new_n3962_), .A2(new_n3864_), .Z(new_n3963_));
  INV_X1     g03771(.I(new_n3963_), .ZN(new_n3964_));
  OAI21_X1   g03772(.A1(new_n3824_), .A2(new_n3826_), .B(new_n3829_), .ZN(new_n3965_));
  NOR2_X1    g03773(.A1(new_n3928_), .A2(new_n3965_), .ZN(new_n3966_));
  XOR2_X1    g03774(.A1(new_n3966_), .A2(new_n3710_), .Z(new_n3967_));
  NAND3_X1   g03775(.A1(\asqrt[37] ), .A2(new_n3843_), .A3(new_n3825_), .ZN(new_n3968_));
  XOR2_X1    g03776(.A1(new_n3968_), .A2(new_n3714_), .Z(new_n3969_));
  OAI21_X1   g03777(.A1(new_n3838_), .A2(new_n3839_), .B(new_n3842_), .ZN(new_n3970_));
  NOR2_X1    g03778(.A1(new_n3928_), .A2(new_n3970_), .ZN(new_n3971_));
  XOR2_X1    g03779(.A1(new_n3971_), .A2(new_n3716_), .Z(new_n3972_));
  INV_X1     g03780(.I(new_n3972_), .ZN(new_n3973_));
  NAND3_X1   g03781(.A1(\asqrt[37] ), .A2(new_n3802_), .A3(new_n3821_), .ZN(new_n3974_));
  XOR2_X1    g03782(.A1(new_n3974_), .A2(new_n3836_), .Z(new_n3975_));
  INV_X1     g03783(.I(new_n3975_), .ZN(new_n3976_));
  OAI21_X1   g03784(.A1(new_n3796_), .A2(new_n3798_), .B(new_n3801_), .ZN(new_n3977_));
  NOR2_X1    g03785(.A1(new_n3928_), .A2(new_n3977_), .ZN(new_n3978_));
  XOR2_X1    g03786(.A1(new_n3978_), .A2(new_n3722_), .Z(new_n3979_));
  NAND3_X1   g03787(.A1(\asqrt[37] ), .A2(new_n3815_), .A3(new_n3797_), .ZN(new_n3980_));
  XOR2_X1    g03788(.A1(new_n3980_), .A2(new_n3726_), .Z(new_n3981_));
  OAI21_X1   g03789(.A1(new_n3810_), .A2(new_n3811_), .B(new_n3814_), .ZN(new_n3982_));
  NOR2_X1    g03790(.A1(new_n3928_), .A2(new_n3982_), .ZN(new_n3983_));
  XOR2_X1    g03791(.A1(new_n3983_), .A2(new_n3728_), .Z(new_n3984_));
  INV_X1     g03792(.I(new_n3984_), .ZN(new_n3985_));
  NAND3_X1   g03793(.A1(\asqrt[37] ), .A2(new_n3767_), .A3(new_n3793_), .ZN(new_n3986_));
  XOR2_X1    g03794(.A1(new_n3986_), .A2(new_n3808_), .Z(new_n3987_));
  INV_X1     g03795(.I(new_n3987_), .ZN(new_n3988_));
  AOI21_X1   g03796(.A1(new_n3788_), .A2(new_n3789_), .B(new_n3792_), .ZN(new_n3989_));
  NAND2_X1   g03797(.A1(\asqrt[37] ), .A2(new_n3989_), .ZN(new_n3990_));
  XOR2_X1    g03798(.A1(new_n3990_), .A2(new_n3772_), .Z(new_n3991_));
  NOR2_X1    g03799(.A1(new_n3787_), .A2(\asqrt[42] ), .ZN(new_n3992_));
  NOR3_X1    g03800(.A1(new_n3928_), .A2(new_n3992_), .A3(new_n3765_), .ZN(new_n3993_));
  XOR2_X1    g03801(.A1(new_n3993_), .A2(new_n3737_), .Z(new_n3994_));
  NOR3_X1    g03802(.A1(new_n3928_), .A2(new_n3784_), .A3(new_n3760_), .ZN(new_n3995_));
  XOR2_X1    g03803(.A1(new_n3995_), .A2(new_n3759_), .Z(new_n3996_));
  INV_X1     g03804(.I(new_n3996_), .ZN(new_n3997_));
  NOR2_X1    g03805(.A1(new_n3754_), .A2(\asqrt[40] ), .ZN(new_n3998_));
  NOR3_X1    g03806(.A1(new_n3928_), .A2(new_n3998_), .A3(new_n3783_), .ZN(new_n3999_));
  XOR2_X1    g03807(.A1(new_n3999_), .A2(new_n3745_), .Z(new_n4000_));
  INV_X1     g03808(.I(new_n4000_), .ZN(new_n4001_));
  NAND3_X1   g03809(.A1(\asqrt[37] ), .A2(new_n3746_), .A3(new_n3747_), .ZN(new_n4002_));
  NOR4_X1    g03810(.A1(new_n3924_), .A2(new_n3675_), .A3(new_n3678_), .A4(new_n3926_), .ZN(new_n4003_));
  INV_X1     g03811(.I(new_n4003_), .ZN(new_n4004_));
  AOI21_X1   g03812(.A1(new_n4002_), .A2(new_n4004_), .B(\a[76] ), .ZN(new_n4005_));
  NOR3_X1    g03813(.A1(new_n3928_), .A2(\a[74] ), .A3(\a[75] ), .ZN(new_n4006_));
  NOR3_X1    g03814(.A1(new_n4006_), .A2(new_n3469_), .A3(new_n4003_), .ZN(new_n4007_));
  NOR2_X1    g03815(.A1(new_n4007_), .A2(new_n4005_), .ZN(new_n4008_));
  INV_X1     g03816(.I(\a[72] ), .ZN(new_n4009_));
  INV_X1     g03817(.I(\a[73] ), .ZN(new_n4010_));
  NAND3_X1   g03818(.A1(new_n4009_), .A2(new_n4010_), .A3(new_n3746_), .ZN(new_n4011_));
  OAI21_X1   g03819(.A1(new_n3928_), .A2(new_n3746_), .B(new_n4011_), .ZN(new_n4012_));
  NAND2_X1   g03820(.A1(new_n4012_), .A2(\asqrt[38] ), .ZN(new_n4013_));
  OAI21_X1   g03821(.A1(new_n3928_), .A2(\a[74] ), .B(\a[75] ), .ZN(new_n4014_));
  NAND2_X1   g03822(.A1(new_n4014_), .A2(new_n4002_), .ZN(new_n4015_));
  NOR2_X1    g03823(.A1(new_n4012_), .A2(\asqrt[38] ), .ZN(new_n4016_));
  OAI21_X1   g03824(.A1(new_n4015_), .A2(new_n4016_), .B(new_n4013_), .ZN(new_n4017_));
  OAI21_X1   g03825(.A1(\asqrt[39] ), .A2(new_n4017_), .B(new_n4008_), .ZN(new_n4018_));
  NAND2_X1   g03826(.A1(new_n4017_), .A2(\asqrt[39] ), .ZN(new_n4019_));
  NAND3_X1   g03827(.A1(new_n4018_), .A2(new_n3167_), .A3(new_n4019_), .ZN(new_n4020_));
  NOR3_X1    g03828(.A1(new_n3928_), .A2(new_n3777_), .A3(new_n3753_), .ZN(new_n4021_));
  XOR2_X1    g03829(.A1(new_n4021_), .A2(new_n3779_), .Z(new_n4022_));
  NAND2_X1   g03830(.A1(new_n4020_), .A2(new_n4022_), .ZN(new_n4023_));
  NAND2_X1   g03831(.A1(new_n4018_), .A2(new_n4019_), .ZN(new_n4024_));
  AOI21_X1   g03832(.A1(new_n4024_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n4025_));
  AOI21_X1   g03833(.A1(new_n4025_), .A2(new_n4023_), .B(new_n4001_), .ZN(new_n4026_));
  OAI21_X1   g03834(.A1(new_n4006_), .A2(new_n4003_), .B(new_n3469_), .ZN(new_n4027_));
  NAND3_X1   g03835(.A1(new_n4002_), .A2(\a[76] ), .A3(new_n4004_), .ZN(new_n4028_));
  NAND2_X1   g03836(.A1(new_n4027_), .A2(new_n4028_), .ZN(new_n4029_));
  NAND2_X1   g03837(.A1(\asqrt[37] ), .A2(\a[74] ), .ZN(new_n4030_));
  AOI21_X1   g03838(.A1(new_n4030_), .A2(new_n4011_), .B(new_n3675_), .ZN(new_n4031_));
  AOI21_X1   g03839(.A1(\asqrt[37] ), .A2(new_n3746_), .B(new_n3747_), .ZN(new_n4032_));
  NOR2_X1    g03840(.A1(new_n4032_), .A2(new_n4006_), .ZN(new_n4033_));
  NAND3_X1   g03841(.A1(new_n4030_), .A2(new_n3675_), .A3(new_n4011_), .ZN(new_n4034_));
  AOI21_X1   g03842(.A1(new_n4033_), .A2(new_n4034_), .B(new_n4031_), .ZN(new_n4035_));
  AOI21_X1   g03843(.A1(new_n4035_), .A2(new_n3400_), .B(new_n4029_), .ZN(new_n4036_));
  NOR2_X1    g03844(.A1(new_n4035_), .A2(new_n3400_), .ZN(new_n4037_));
  OAI21_X1   g03845(.A1(new_n4036_), .A2(new_n4037_), .B(\asqrt[40] ), .ZN(new_n4038_));
  AOI21_X1   g03846(.A1(new_n4023_), .A2(new_n4038_), .B(new_n2912_), .ZN(new_n4039_));
  NOR2_X1    g03847(.A1(new_n4026_), .A2(new_n4039_), .ZN(new_n4040_));
  AOI21_X1   g03848(.A1(new_n4040_), .A2(new_n2699_), .B(new_n3997_), .ZN(new_n4041_));
  OAI21_X1   g03849(.A1(new_n4026_), .A2(new_n4039_), .B(\asqrt[42] ), .ZN(new_n4042_));
  NAND2_X1   g03850(.A1(new_n4042_), .A2(new_n2464_), .ZN(new_n4043_));
  OAI21_X1   g03851(.A1(new_n4041_), .A2(new_n4043_), .B(new_n3994_), .ZN(new_n4044_));
  INV_X1     g03852(.I(new_n4042_), .ZN(new_n4045_));
  OAI21_X1   g03853(.A1(new_n4041_), .A2(new_n4045_), .B(\asqrt[43] ), .ZN(new_n4046_));
  NAND3_X1   g03854(.A1(new_n4044_), .A2(new_n4046_), .A3(new_n2271_), .ZN(new_n4047_));
  NAND2_X1   g03855(.A1(new_n4047_), .A2(new_n3991_), .ZN(new_n4048_));
  NAND2_X1   g03856(.A1(new_n4044_), .A2(new_n4046_), .ZN(new_n4049_));
  AOI21_X1   g03857(.A1(new_n4049_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n4050_));
  AOI21_X1   g03858(.A1(new_n4050_), .A2(new_n4048_), .B(new_n3988_), .ZN(new_n4051_));
  INV_X1     g03859(.I(new_n3994_), .ZN(new_n4052_));
  NOR2_X1    g03860(.A1(new_n4036_), .A2(new_n4037_), .ZN(new_n4053_));
  INV_X1     g03861(.I(new_n4022_), .ZN(new_n4054_));
  AOI21_X1   g03862(.A1(new_n4053_), .A2(new_n3167_), .B(new_n4054_), .ZN(new_n4055_));
  NAND2_X1   g03863(.A1(new_n4038_), .A2(new_n2912_), .ZN(new_n4056_));
  OAI21_X1   g03864(.A1(new_n4055_), .A2(new_n4056_), .B(new_n4000_), .ZN(new_n4057_));
  INV_X1     g03865(.I(new_n4038_), .ZN(new_n4058_));
  OAI21_X1   g03866(.A1(new_n4055_), .A2(new_n4058_), .B(\asqrt[41] ), .ZN(new_n4059_));
  NAND3_X1   g03867(.A1(new_n4057_), .A2(new_n4059_), .A3(new_n2699_), .ZN(new_n4060_));
  NAND2_X1   g03868(.A1(new_n4060_), .A2(new_n3996_), .ZN(new_n4061_));
  NAND2_X1   g03869(.A1(new_n4057_), .A2(new_n4059_), .ZN(new_n4062_));
  AOI21_X1   g03870(.A1(new_n4062_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n4063_));
  AOI21_X1   g03871(.A1(new_n4063_), .A2(new_n4061_), .B(new_n4052_), .ZN(new_n4064_));
  AOI21_X1   g03872(.A1(new_n4061_), .A2(new_n4042_), .B(new_n2464_), .ZN(new_n4065_));
  OAI21_X1   g03873(.A1(new_n4064_), .A2(new_n4065_), .B(\asqrt[44] ), .ZN(new_n4066_));
  AOI21_X1   g03874(.A1(new_n4048_), .A2(new_n4066_), .B(new_n2072_), .ZN(new_n4067_));
  NOR2_X1    g03875(.A1(new_n4051_), .A2(new_n4067_), .ZN(new_n4068_));
  AOI21_X1   g03876(.A1(new_n4068_), .A2(new_n1884_), .B(new_n3985_), .ZN(new_n4069_));
  OAI21_X1   g03877(.A1(new_n4051_), .A2(new_n4067_), .B(\asqrt[46] ), .ZN(new_n4070_));
  NAND2_X1   g03878(.A1(new_n4070_), .A2(new_n1688_), .ZN(new_n4071_));
  OAI21_X1   g03879(.A1(new_n4069_), .A2(new_n4071_), .B(new_n3981_), .ZN(new_n4072_));
  INV_X1     g03880(.I(new_n4070_), .ZN(new_n4073_));
  OAI21_X1   g03881(.A1(new_n4069_), .A2(new_n4073_), .B(\asqrt[47] ), .ZN(new_n4074_));
  NAND3_X1   g03882(.A1(new_n4072_), .A2(new_n4074_), .A3(new_n1533_), .ZN(new_n4075_));
  NAND2_X1   g03883(.A1(new_n4075_), .A2(new_n3979_), .ZN(new_n4076_));
  NAND2_X1   g03884(.A1(new_n4072_), .A2(new_n4074_), .ZN(new_n4077_));
  AOI21_X1   g03885(.A1(new_n4077_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n4078_));
  AOI21_X1   g03886(.A1(new_n4078_), .A2(new_n4076_), .B(new_n3976_), .ZN(new_n4079_));
  INV_X1     g03887(.I(new_n3981_), .ZN(new_n4080_));
  INV_X1     g03888(.I(new_n3991_), .ZN(new_n4081_));
  NOR2_X1    g03889(.A1(new_n4064_), .A2(new_n4065_), .ZN(new_n4082_));
  AOI21_X1   g03890(.A1(new_n4082_), .A2(new_n2271_), .B(new_n4081_), .ZN(new_n4083_));
  NAND2_X1   g03891(.A1(new_n4066_), .A2(new_n2072_), .ZN(new_n4084_));
  OAI21_X1   g03892(.A1(new_n4083_), .A2(new_n4084_), .B(new_n3987_), .ZN(new_n4085_));
  INV_X1     g03893(.I(new_n4066_), .ZN(new_n4086_));
  OAI21_X1   g03894(.A1(new_n4083_), .A2(new_n4086_), .B(\asqrt[45] ), .ZN(new_n4087_));
  NAND3_X1   g03895(.A1(new_n4085_), .A2(new_n4087_), .A3(new_n1884_), .ZN(new_n4088_));
  NAND2_X1   g03896(.A1(new_n4088_), .A2(new_n3984_), .ZN(new_n4089_));
  NAND2_X1   g03897(.A1(new_n4085_), .A2(new_n4087_), .ZN(new_n4090_));
  AOI21_X1   g03898(.A1(new_n4090_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n4091_));
  AOI21_X1   g03899(.A1(new_n4091_), .A2(new_n4089_), .B(new_n4080_), .ZN(new_n4092_));
  AOI21_X1   g03900(.A1(new_n4089_), .A2(new_n4070_), .B(new_n1688_), .ZN(new_n4093_));
  OAI21_X1   g03901(.A1(new_n4092_), .A2(new_n4093_), .B(\asqrt[48] ), .ZN(new_n4094_));
  AOI21_X1   g03902(.A1(new_n4076_), .A2(new_n4094_), .B(new_n1368_), .ZN(new_n4095_));
  NOR2_X1    g03903(.A1(new_n4079_), .A2(new_n4095_), .ZN(new_n4096_));
  AOI21_X1   g03904(.A1(new_n4096_), .A2(new_n1228_), .B(new_n3973_), .ZN(new_n4097_));
  OAI21_X1   g03905(.A1(new_n4079_), .A2(new_n4095_), .B(\asqrt[50] ), .ZN(new_n4098_));
  NAND2_X1   g03906(.A1(new_n4098_), .A2(new_n1088_), .ZN(new_n4099_));
  OAI21_X1   g03907(.A1(new_n4097_), .A2(new_n4099_), .B(new_n3969_), .ZN(new_n4100_));
  INV_X1     g03908(.I(new_n4098_), .ZN(new_n4101_));
  OAI21_X1   g03909(.A1(new_n4097_), .A2(new_n4101_), .B(\asqrt[51] ), .ZN(new_n4102_));
  NAND3_X1   g03910(.A1(new_n4100_), .A2(new_n4102_), .A3(new_n962_), .ZN(new_n4103_));
  NAND2_X1   g03911(.A1(new_n4103_), .A2(new_n3967_), .ZN(new_n4104_));
  NAND2_X1   g03912(.A1(new_n4100_), .A2(new_n4102_), .ZN(new_n4105_));
  AOI21_X1   g03913(.A1(new_n4105_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n4106_));
  AOI21_X1   g03914(.A1(new_n4106_), .A2(new_n4104_), .B(new_n3964_), .ZN(new_n4107_));
  INV_X1     g03915(.I(new_n3969_), .ZN(new_n4108_));
  INV_X1     g03916(.I(new_n3979_), .ZN(new_n4109_));
  NOR2_X1    g03917(.A1(new_n4092_), .A2(new_n4093_), .ZN(new_n4110_));
  AOI21_X1   g03918(.A1(new_n4110_), .A2(new_n1533_), .B(new_n4109_), .ZN(new_n4111_));
  NAND2_X1   g03919(.A1(new_n4094_), .A2(new_n1368_), .ZN(new_n4112_));
  OAI21_X1   g03920(.A1(new_n4111_), .A2(new_n4112_), .B(new_n3975_), .ZN(new_n4113_));
  INV_X1     g03921(.I(new_n4094_), .ZN(new_n4114_));
  OAI21_X1   g03922(.A1(new_n4111_), .A2(new_n4114_), .B(\asqrt[49] ), .ZN(new_n4115_));
  NAND3_X1   g03923(.A1(new_n4113_), .A2(new_n4115_), .A3(new_n1228_), .ZN(new_n4116_));
  NAND2_X1   g03924(.A1(new_n4116_), .A2(new_n3972_), .ZN(new_n4117_));
  NAND2_X1   g03925(.A1(new_n4113_), .A2(new_n4115_), .ZN(new_n4118_));
  AOI21_X1   g03926(.A1(new_n4118_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n4119_));
  AOI21_X1   g03927(.A1(new_n4119_), .A2(new_n4117_), .B(new_n4108_), .ZN(new_n4120_));
  AOI21_X1   g03928(.A1(new_n4117_), .A2(new_n4098_), .B(new_n1088_), .ZN(new_n4121_));
  OAI21_X1   g03929(.A1(new_n4120_), .A2(new_n4121_), .B(\asqrt[52] ), .ZN(new_n4122_));
  AOI21_X1   g03930(.A1(new_n4104_), .A2(new_n4122_), .B(new_n842_), .ZN(new_n4123_));
  NOR2_X1    g03931(.A1(new_n4107_), .A2(new_n4123_), .ZN(new_n4124_));
  AOI21_X1   g03932(.A1(new_n4124_), .A2(new_n720_), .B(new_n3961_), .ZN(new_n4125_));
  OAI21_X1   g03933(.A1(new_n4107_), .A2(new_n4123_), .B(\asqrt[54] ), .ZN(new_n4126_));
  NAND2_X1   g03934(.A1(new_n4126_), .A2(new_n630_), .ZN(new_n4127_));
  OAI21_X1   g03935(.A1(new_n4125_), .A2(new_n4127_), .B(new_n3957_), .ZN(new_n4128_));
  INV_X1     g03936(.I(new_n4126_), .ZN(new_n4129_));
  OAI21_X1   g03937(.A1(new_n4125_), .A2(new_n4129_), .B(\asqrt[55] ), .ZN(new_n4130_));
  NAND3_X1   g03938(.A1(new_n4128_), .A2(new_n4130_), .A3(new_n545_), .ZN(new_n4131_));
  NAND2_X1   g03939(.A1(new_n4131_), .A2(new_n3955_), .ZN(new_n4132_));
  NAND2_X1   g03940(.A1(new_n4128_), .A2(new_n4130_), .ZN(new_n4133_));
  AOI21_X1   g03941(.A1(new_n4133_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n4134_));
  AOI21_X1   g03942(.A1(new_n4134_), .A2(new_n4132_), .B(new_n3952_), .ZN(new_n4135_));
  INV_X1     g03943(.I(new_n3957_), .ZN(new_n4136_));
  INV_X1     g03944(.I(new_n3967_), .ZN(new_n4137_));
  NOR2_X1    g03945(.A1(new_n4120_), .A2(new_n4121_), .ZN(new_n4138_));
  AOI21_X1   g03946(.A1(new_n4138_), .A2(new_n962_), .B(new_n4137_), .ZN(new_n4139_));
  NAND2_X1   g03947(.A1(new_n4122_), .A2(new_n842_), .ZN(new_n4140_));
  OAI21_X1   g03948(.A1(new_n4139_), .A2(new_n4140_), .B(new_n3963_), .ZN(new_n4141_));
  INV_X1     g03949(.I(new_n4122_), .ZN(new_n4142_));
  OAI21_X1   g03950(.A1(new_n4139_), .A2(new_n4142_), .B(\asqrt[53] ), .ZN(new_n4143_));
  NAND3_X1   g03951(.A1(new_n4141_), .A2(new_n4143_), .A3(new_n720_), .ZN(new_n4144_));
  NAND2_X1   g03952(.A1(new_n4144_), .A2(new_n3960_), .ZN(new_n4145_));
  NAND2_X1   g03953(.A1(new_n4141_), .A2(new_n4143_), .ZN(new_n4146_));
  AOI21_X1   g03954(.A1(new_n4146_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n4147_));
  AOI21_X1   g03955(.A1(new_n4147_), .A2(new_n4145_), .B(new_n4136_), .ZN(new_n4148_));
  AOI21_X1   g03956(.A1(new_n4145_), .A2(new_n4126_), .B(new_n630_), .ZN(new_n4149_));
  OAI21_X1   g03957(.A1(new_n4148_), .A2(new_n4149_), .B(\asqrt[56] ), .ZN(new_n4150_));
  AOI21_X1   g03958(.A1(new_n4132_), .A2(new_n4150_), .B(new_n450_), .ZN(new_n4151_));
  NOR2_X1    g03959(.A1(new_n4135_), .A2(new_n4151_), .ZN(new_n4152_));
  AOI21_X1   g03960(.A1(new_n4152_), .A2(new_n403_), .B(new_n3949_), .ZN(new_n4153_));
  OAI21_X1   g03961(.A1(new_n4135_), .A2(new_n4151_), .B(\asqrt[58] ), .ZN(new_n4154_));
  NAND2_X1   g03962(.A1(new_n4154_), .A2(new_n339_), .ZN(new_n4155_));
  OAI21_X1   g03963(.A1(new_n4153_), .A2(new_n4155_), .B(new_n3945_), .ZN(new_n4156_));
  INV_X1     g03964(.I(new_n4154_), .ZN(new_n4157_));
  OAI21_X1   g03965(.A1(new_n4153_), .A2(new_n4157_), .B(\asqrt[59] ), .ZN(new_n4158_));
  NAND3_X1   g03966(.A1(new_n4156_), .A2(new_n4158_), .A3(new_n288_), .ZN(new_n4159_));
  INV_X1     g03967(.I(new_n3945_), .ZN(new_n4160_));
  INV_X1     g03968(.I(new_n3955_), .ZN(new_n4161_));
  NOR2_X1    g03969(.A1(new_n4148_), .A2(new_n4149_), .ZN(new_n4162_));
  AOI21_X1   g03970(.A1(new_n4162_), .A2(new_n545_), .B(new_n4161_), .ZN(new_n4163_));
  NAND2_X1   g03971(.A1(new_n4150_), .A2(new_n450_), .ZN(new_n4164_));
  OAI21_X1   g03972(.A1(new_n4163_), .A2(new_n4164_), .B(new_n3951_), .ZN(new_n4165_));
  INV_X1     g03973(.I(new_n4150_), .ZN(new_n4166_));
  OAI21_X1   g03974(.A1(new_n4163_), .A2(new_n4166_), .B(\asqrt[57] ), .ZN(new_n4167_));
  NAND3_X1   g03975(.A1(new_n4165_), .A2(new_n4167_), .A3(new_n403_), .ZN(new_n4168_));
  NAND2_X1   g03976(.A1(new_n4168_), .A2(new_n3948_), .ZN(new_n4169_));
  NAND2_X1   g03977(.A1(new_n4165_), .A2(new_n4167_), .ZN(new_n4170_));
  AOI21_X1   g03978(.A1(new_n4170_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n4171_));
  AOI21_X1   g03979(.A1(new_n4171_), .A2(new_n4169_), .B(new_n4160_), .ZN(new_n4172_));
  AOI21_X1   g03980(.A1(new_n4169_), .A2(new_n4154_), .B(new_n339_), .ZN(new_n4173_));
  OAI21_X1   g03981(.A1(new_n4172_), .A2(new_n4173_), .B(\asqrt[60] ), .ZN(new_n4174_));
  NAND2_X1   g03982(.A1(new_n3925_), .A2(new_n3680_), .ZN(new_n4175_));
  NOR2_X1    g03983(.A1(new_n3928_), .A2(new_n3680_), .ZN(new_n4176_));
  NAND2_X1   g03984(.A1(new_n4176_), .A2(new_n3940_), .ZN(new_n4177_));
  AOI21_X1   g03985(.A1(new_n4177_), .A2(new_n4175_), .B(new_n193_), .ZN(new_n4178_));
  INV_X1     g03986(.I(new_n4178_), .ZN(new_n4179_));
  NAND3_X1   g03987(.A1(\asqrt[37] ), .A2(new_n3910_), .A3(new_n3921_), .ZN(new_n4180_));
  XOR2_X1    g03988(.A1(new_n4180_), .A2(new_n3913_), .Z(new_n4181_));
  AOI21_X1   g03989(.A1(new_n4176_), .A2(new_n3925_), .B(new_n3926_), .ZN(new_n4182_));
  NAND2_X1   g03990(.A1(new_n4159_), .A2(new_n3931_), .ZN(new_n4183_));
  AOI21_X1   g03991(.A1(new_n4183_), .A2(new_n4174_), .B(new_n242_), .ZN(new_n4184_));
  NAND3_X1   g03992(.A1(\asqrt[37] ), .A2(new_n3886_), .A3(new_n3902_), .ZN(new_n4185_));
  XOR2_X1    g03993(.A1(new_n4185_), .A2(new_n3914_), .Z(new_n4186_));
  INV_X1     g03994(.I(new_n4186_), .ZN(new_n4187_));
  NAND2_X1   g03995(.A1(new_n4156_), .A2(new_n4158_), .ZN(new_n4188_));
  AOI21_X1   g03996(.A1(new_n4188_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n4189_));
  AOI21_X1   g03997(.A1(new_n4189_), .A2(new_n4183_), .B(new_n4187_), .ZN(new_n4190_));
  OAI21_X1   g03998(.A1(new_n4190_), .A2(new_n4184_), .B(\asqrt[62] ), .ZN(new_n4191_));
  INV_X1     g03999(.I(new_n4191_), .ZN(new_n4192_));
  NOR2_X1    g04000(.A1(new_n4190_), .A2(new_n4184_), .ZN(new_n4193_));
  AOI21_X1   g04001(.A1(new_n3887_), .A2(new_n3908_), .B(new_n3903_), .ZN(new_n4194_));
  NAND2_X1   g04002(.A1(\asqrt[37] ), .A2(new_n4194_), .ZN(new_n4195_));
  XOR2_X1    g04003(.A1(new_n4195_), .A2(new_n3906_), .Z(new_n4196_));
  INV_X1     g04004(.I(new_n4196_), .ZN(new_n4197_));
  AOI21_X1   g04005(.A1(new_n4193_), .A2(new_n234_), .B(new_n4197_), .ZN(new_n4198_));
  OAI21_X1   g04006(.A1(new_n4198_), .A2(new_n4192_), .B(new_n4182_), .ZN(new_n4199_));
  OAI21_X1   g04007(.A1(new_n4199_), .A2(new_n4181_), .B(new_n193_), .ZN(new_n4200_));
  NOR2_X1    g04008(.A1(new_n4198_), .A2(new_n4192_), .ZN(new_n4201_));
  NAND2_X1   g04009(.A1(new_n4201_), .A2(new_n4181_), .ZN(new_n4202_));
  NOR2_X1    g04010(.A1(\asqrt[37] ), .A2(new_n3681_), .ZN(new_n4203_));
  INV_X1     g04011(.I(new_n4203_), .ZN(new_n4204_));
  NAND4_X1   g04012(.A1(new_n4200_), .A2(new_n4179_), .A3(new_n4202_), .A4(new_n4204_), .ZN(\asqrt[36] ));
  NAND3_X1   g04013(.A1(\asqrt[36] ), .A2(new_n4159_), .A3(new_n4174_), .ZN(new_n4206_));
  XOR2_X1    g04014(.A1(new_n4206_), .A2(new_n3932_), .Z(new_n4207_));
  INV_X1     g04015(.I(new_n4207_), .ZN(new_n4208_));
  NOR2_X1    g04016(.A1(new_n4172_), .A2(new_n4173_), .ZN(new_n4209_));
  AOI21_X1   g04017(.A1(new_n4209_), .A2(new_n288_), .B(new_n3932_), .ZN(new_n4210_));
  INV_X1     g04018(.I(new_n4174_), .ZN(new_n4211_));
  OAI21_X1   g04019(.A1(new_n4210_), .A2(new_n4211_), .B(\asqrt[61] ), .ZN(new_n4212_));
  NAND2_X1   g04020(.A1(new_n4174_), .A2(new_n242_), .ZN(new_n4213_));
  OAI21_X1   g04021(.A1(new_n4210_), .A2(new_n4213_), .B(new_n4186_), .ZN(new_n4214_));
  NAND3_X1   g04022(.A1(new_n4214_), .A2(new_n4212_), .A3(new_n234_), .ZN(new_n4215_));
  NAND2_X1   g04023(.A1(new_n4215_), .A2(new_n4196_), .ZN(new_n4216_));
  NAND2_X1   g04024(.A1(new_n4216_), .A2(new_n4191_), .ZN(new_n4217_));
  NAND2_X1   g04025(.A1(new_n4217_), .A2(new_n4181_), .ZN(new_n4218_));
  INV_X1     g04026(.I(new_n4181_), .ZN(new_n4219_));
  INV_X1     g04027(.I(new_n4182_), .ZN(new_n4220_));
  AOI21_X1   g04028(.A1(new_n4216_), .A2(new_n4191_), .B(new_n4220_), .ZN(new_n4221_));
  AOI21_X1   g04029(.A1(new_n4221_), .A2(new_n4219_), .B(\asqrt[63] ), .ZN(new_n4222_));
  NOR2_X1    g04030(.A1(new_n4217_), .A2(new_n4219_), .ZN(new_n4223_));
  NOR4_X1    g04031(.A1(new_n4222_), .A2(new_n4178_), .A3(new_n4223_), .A4(new_n4203_), .ZN(new_n4224_));
  NOR2_X1    g04032(.A1(new_n4224_), .A2(new_n4181_), .ZN(new_n4225_));
  NAND2_X1   g04033(.A1(new_n4225_), .A2(new_n4201_), .ZN(new_n4226_));
  AOI21_X1   g04034(.A1(new_n4226_), .A2(new_n4218_), .B(new_n193_), .ZN(new_n4227_));
  INV_X1     g04035(.I(new_n4227_), .ZN(new_n4228_));
  NAND3_X1   g04036(.A1(\asqrt[36] ), .A2(new_n4191_), .A3(new_n4215_), .ZN(new_n4229_));
  XOR2_X1    g04037(.A1(new_n4229_), .A2(new_n4196_), .Z(new_n4230_));
  AOI21_X1   g04038(.A1(new_n4225_), .A2(new_n4217_), .B(new_n4223_), .ZN(new_n4231_));
  OAI21_X1   g04039(.A1(new_n4153_), .A2(new_n4155_), .B(new_n4158_), .ZN(new_n4232_));
  NOR2_X1    g04040(.A1(new_n4224_), .A2(new_n4232_), .ZN(new_n4233_));
  XOR2_X1    g04041(.A1(new_n4233_), .A2(new_n3945_), .Z(new_n4234_));
  NAND3_X1   g04042(.A1(\asqrt[36] ), .A2(new_n4168_), .A3(new_n4154_), .ZN(new_n4235_));
  XOR2_X1    g04043(.A1(new_n4235_), .A2(new_n3949_), .Z(new_n4236_));
  OAI21_X1   g04044(.A1(new_n4163_), .A2(new_n4164_), .B(new_n4167_), .ZN(new_n4237_));
  NOR2_X1    g04045(.A1(new_n4224_), .A2(new_n4237_), .ZN(new_n4238_));
  XOR2_X1    g04046(.A1(new_n4238_), .A2(new_n3951_), .Z(new_n4239_));
  INV_X1     g04047(.I(new_n4239_), .ZN(new_n4240_));
  NAND3_X1   g04048(.A1(\asqrt[36] ), .A2(new_n4131_), .A3(new_n4150_), .ZN(new_n4241_));
  XOR2_X1    g04049(.A1(new_n4241_), .A2(new_n4161_), .Z(new_n4242_));
  INV_X1     g04050(.I(new_n4242_), .ZN(new_n4243_));
  OAI21_X1   g04051(.A1(new_n4125_), .A2(new_n4127_), .B(new_n4130_), .ZN(new_n4244_));
  NOR2_X1    g04052(.A1(new_n4224_), .A2(new_n4244_), .ZN(new_n4245_));
  XOR2_X1    g04053(.A1(new_n4245_), .A2(new_n3957_), .Z(new_n4246_));
  NAND3_X1   g04054(.A1(\asqrt[36] ), .A2(new_n4144_), .A3(new_n4126_), .ZN(new_n4247_));
  XOR2_X1    g04055(.A1(new_n4247_), .A2(new_n3961_), .Z(new_n4248_));
  OAI21_X1   g04056(.A1(new_n4139_), .A2(new_n4140_), .B(new_n4143_), .ZN(new_n4249_));
  NOR2_X1    g04057(.A1(new_n4224_), .A2(new_n4249_), .ZN(new_n4250_));
  XOR2_X1    g04058(.A1(new_n4250_), .A2(new_n3963_), .Z(new_n4251_));
  INV_X1     g04059(.I(new_n4251_), .ZN(new_n4252_));
  NAND3_X1   g04060(.A1(\asqrt[36] ), .A2(new_n4103_), .A3(new_n4122_), .ZN(new_n4253_));
  XOR2_X1    g04061(.A1(new_n4253_), .A2(new_n4137_), .Z(new_n4254_));
  INV_X1     g04062(.I(new_n4254_), .ZN(new_n4255_));
  OAI21_X1   g04063(.A1(new_n4097_), .A2(new_n4099_), .B(new_n4102_), .ZN(new_n4256_));
  NOR2_X1    g04064(.A1(new_n4224_), .A2(new_n4256_), .ZN(new_n4257_));
  XOR2_X1    g04065(.A1(new_n4257_), .A2(new_n3969_), .Z(new_n4258_));
  NAND3_X1   g04066(.A1(\asqrt[36] ), .A2(new_n4116_), .A3(new_n4098_), .ZN(new_n4259_));
  XOR2_X1    g04067(.A1(new_n4259_), .A2(new_n3973_), .Z(new_n4260_));
  OAI21_X1   g04068(.A1(new_n4111_), .A2(new_n4112_), .B(new_n4115_), .ZN(new_n4261_));
  NOR2_X1    g04069(.A1(new_n4224_), .A2(new_n4261_), .ZN(new_n4262_));
  XOR2_X1    g04070(.A1(new_n4262_), .A2(new_n3975_), .Z(new_n4263_));
  INV_X1     g04071(.I(new_n4263_), .ZN(new_n4264_));
  NAND3_X1   g04072(.A1(\asqrt[36] ), .A2(new_n4075_), .A3(new_n4094_), .ZN(new_n4265_));
  XOR2_X1    g04073(.A1(new_n4265_), .A2(new_n4109_), .Z(new_n4266_));
  INV_X1     g04074(.I(new_n4266_), .ZN(new_n4267_));
  OAI21_X1   g04075(.A1(new_n4069_), .A2(new_n4071_), .B(new_n4074_), .ZN(new_n4268_));
  NOR2_X1    g04076(.A1(new_n4224_), .A2(new_n4268_), .ZN(new_n4269_));
  XOR2_X1    g04077(.A1(new_n4269_), .A2(new_n3981_), .Z(new_n4270_));
  NAND3_X1   g04078(.A1(\asqrt[36] ), .A2(new_n4088_), .A3(new_n4070_), .ZN(new_n4271_));
  XOR2_X1    g04079(.A1(new_n4271_), .A2(new_n3985_), .Z(new_n4272_));
  OAI21_X1   g04080(.A1(new_n4083_), .A2(new_n4084_), .B(new_n4087_), .ZN(new_n4273_));
  NOR2_X1    g04081(.A1(new_n4224_), .A2(new_n4273_), .ZN(new_n4274_));
  XOR2_X1    g04082(.A1(new_n4274_), .A2(new_n3987_), .Z(new_n4275_));
  INV_X1     g04083(.I(new_n4275_), .ZN(new_n4276_));
  NAND3_X1   g04084(.A1(\asqrt[36] ), .A2(new_n4047_), .A3(new_n4066_), .ZN(new_n4277_));
  XOR2_X1    g04085(.A1(new_n4277_), .A2(new_n4081_), .Z(new_n4278_));
  INV_X1     g04086(.I(new_n4278_), .ZN(new_n4279_));
  OAI21_X1   g04087(.A1(new_n4041_), .A2(new_n4043_), .B(new_n4046_), .ZN(new_n4280_));
  NOR2_X1    g04088(.A1(new_n4224_), .A2(new_n4280_), .ZN(new_n4281_));
  XOR2_X1    g04089(.A1(new_n4281_), .A2(new_n3994_), .Z(new_n4282_));
  NAND3_X1   g04090(.A1(\asqrt[36] ), .A2(new_n4060_), .A3(new_n4042_), .ZN(new_n4283_));
  XOR2_X1    g04091(.A1(new_n4283_), .A2(new_n3997_), .Z(new_n4284_));
  OAI21_X1   g04092(.A1(new_n4055_), .A2(new_n4056_), .B(new_n4059_), .ZN(new_n4285_));
  NOR2_X1    g04093(.A1(new_n4224_), .A2(new_n4285_), .ZN(new_n4286_));
  XOR2_X1    g04094(.A1(new_n4286_), .A2(new_n4000_), .Z(new_n4287_));
  INV_X1     g04095(.I(new_n4287_), .ZN(new_n4288_));
  NAND3_X1   g04096(.A1(\asqrt[36] ), .A2(new_n4020_), .A3(new_n4038_), .ZN(new_n4289_));
  XOR2_X1    g04097(.A1(new_n4289_), .A2(new_n4054_), .Z(new_n4290_));
  INV_X1     g04098(.I(new_n4290_), .ZN(new_n4291_));
  NOR2_X1    g04099(.A1(new_n4017_), .A2(\asqrt[39] ), .ZN(new_n4292_));
  NOR3_X1    g04100(.A1(new_n4224_), .A2(new_n4292_), .A3(new_n4037_), .ZN(new_n4293_));
  XOR2_X1    g04101(.A1(new_n4293_), .A2(new_n4008_), .Z(new_n4294_));
  NOR3_X1    g04102(.A1(new_n4224_), .A2(\a[72] ), .A3(\a[73] ), .ZN(new_n4295_));
  NOR4_X1    g04103(.A1(new_n4222_), .A2(new_n3928_), .A3(new_n4178_), .A4(new_n4223_), .ZN(new_n4296_));
  OAI21_X1   g04104(.A1(new_n4295_), .A2(new_n4296_), .B(new_n3746_), .ZN(new_n4297_));
  NAND3_X1   g04105(.A1(\asqrt[36] ), .A2(new_n4009_), .A3(new_n4010_), .ZN(new_n4298_));
  INV_X1     g04106(.I(new_n4296_), .ZN(new_n4299_));
  NAND3_X1   g04107(.A1(new_n4298_), .A2(\a[74] ), .A3(new_n4299_), .ZN(new_n4300_));
  NAND2_X1   g04108(.A1(new_n4297_), .A2(new_n4300_), .ZN(new_n4301_));
  INV_X1     g04109(.I(\a[70] ), .ZN(new_n4302_));
  INV_X1     g04110(.I(\a[71] ), .ZN(new_n4303_));
  NAND3_X1   g04111(.A1(new_n4302_), .A2(new_n4303_), .A3(new_n4009_), .ZN(new_n4304_));
  NAND2_X1   g04112(.A1(\asqrt[36] ), .A2(\a[72] ), .ZN(new_n4305_));
  AOI21_X1   g04113(.A1(new_n4305_), .A2(new_n4304_), .B(new_n3928_), .ZN(new_n4306_));
  AOI21_X1   g04114(.A1(\asqrt[36] ), .A2(new_n4009_), .B(new_n4010_), .ZN(new_n4307_));
  NOR2_X1    g04115(.A1(new_n4295_), .A2(new_n4307_), .ZN(new_n4308_));
  NAND3_X1   g04116(.A1(new_n4305_), .A2(new_n3928_), .A3(new_n4304_), .ZN(new_n4309_));
  AOI21_X1   g04117(.A1(new_n4308_), .A2(new_n4309_), .B(new_n4306_), .ZN(new_n4310_));
  AOI21_X1   g04118(.A1(new_n4310_), .A2(new_n3675_), .B(new_n4301_), .ZN(new_n4311_));
  NOR2_X1    g04119(.A1(new_n4310_), .A2(new_n3675_), .ZN(new_n4312_));
  NOR3_X1    g04120(.A1(new_n4311_), .A2(\asqrt[39] ), .A3(new_n4312_), .ZN(new_n4313_));
  NOR3_X1    g04121(.A1(new_n4224_), .A2(new_n4031_), .A3(new_n4016_), .ZN(new_n4314_));
  XOR2_X1    g04122(.A1(new_n4314_), .A2(new_n4033_), .Z(new_n4315_));
  INV_X1     g04123(.I(new_n4315_), .ZN(new_n4316_));
  OAI21_X1   g04124(.A1(new_n4311_), .A2(new_n4312_), .B(\asqrt[39] ), .ZN(new_n4317_));
  OAI21_X1   g04125(.A1(new_n4313_), .A2(new_n4316_), .B(new_n4317_), .ZN(new_n4318_));
  OAI21_X1   g04126(.A1(new_n4318_), .A2(\asqrt[40] ), .B(new_n4294_), .ZN(new_n4319_));
  AOI21_X1   g04127(.A1(new_n4318_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n4320_));
  AOI21_X1   g04128(.A1(new_n4320_), .A2(new_n4319_), .B(new_n4291_), .ZN(new_n4321_));
  NAND2_X1   g04129(.A1(new_n4318_), .A2(\asqrt[40] ), .ZN(new_n4322_));
  AOI21_X1   g04130(.A1(new_n4319_), .A2(new_n4322_), .B(new_n2912_), .ZN(new_n4323_));
  NOR2_X1    g04131(.A1(new_n4321_), .A2(new_n4323_), .ZN(new_n4324_));
  AOI21_X1   g04132(.A1(new_n4324_), .A2(new_n2699_), .B(new_n4288_), .ZN(new_n4325_));
  OAI21_X1   g04133(.A1(new_n4321_), .A2(new_n4323_), .B(\asqrt[42] ), .ZN(new_n4326_));
  NAND2_X1   g04134(.A1(new_n4326_), .A2(new_n2464_), .ZN(new_n4327_));
  OAI21_X1   g04135(.A1(new_n4325_), .A2(new_n4327_), .B(new_n4284_), .ZN(new_n4328_));
  INV_X1     g04136(.I(new_n4326_), .ZN(new_n4329_));
  OAI21_X1   g04137(.A1(new_n4325_), .A2(new_n4329_), .B(\asqrt[43] ), .ZN(new_n4330_));
  NAND3_X1   g04138(.A1(new_n4328_), .A2(new_n4330_), .A3(new_n2271_), .ZN(new_n4331_));
  NAND2_X1   g04139(.A1(new_n4331_), .A2(new_n4282_), .ZN(new_n4332_));
  NAND2_X1   g04140(.A1(new_n4328_), .A2(new_n4330_), .ZN(new_n4333_));
  AOI21_X1   g04141(.A1(new_n4333_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n4334_));
  AOI21_X1   g04142(.A1(new_n4334_), .A2(new_n4332_), .B(new_n4279_), .ZN(new_n4335_));
  INV_X1     g04143(.I(new_n4284_), .ZN(new_n4336_));
  INV_X1     g04144(.I(new_n4294_), .ZN(new_n4337_));
  AOI21_X1   g04145(.A1(new_n4298_), .A2(new_n4299_), .B(\a[74] ), .ZN(new_n4338_));
  NOR3_X1    g04146(.A1(new_n4295_), .A2(new_n3746_), .A3(new_n4296_), .ZN(new_n4339_));
  NOR2_X1    g04147(.A1(new_n4339_), .A2(new_n4338_), .ZN(new_n4340_));
  OAI21_X1   g04148(.A1(new_n4224_), .A2(new_n4009_), .B(new_n4304_), .ZN(new_n4341_));
  NAND2_X1   g04149(.A1(new_n4341_), .A2(\asqrt[37] ), .ZN(new_n4342_));
  OAI21_X1   g04150(.A1(new_n4224_), .A2(\a[72] ), .B(\a[73] ), .ZN(new_n4343_));
  NAND2_X1   g04151(.A1(new_n4343_), .A2(new_n4298_), .ZN(new_n4344_));
  NOR2_X1    g04152(.A1(new_n4341_), .A2(\asqrt[37] ), .ZN(new_n4345_));
  OAI21_X1   g04153(.A1(new_n4344_), .A2(new_n4345_), .B(new_n4342_), .ZN(new_n4346_));
  OAI21_X1   g04154(.A1(\asqrt[38] ), .A2(new_n4346_), .B(new_n4340_), .ZN(new_n4347_));
  NAND2_X1   g04155(.A1(new_n4346_), .A2(\asqrt[38] ), .ZN(new_n4348_));
  NAND3_X1   g04156(.A1(new_n4347_), .A2(new_n3400_), .A3(new_n4348_), .ZN(new_n4349_));
  AOI21_X1   g04157(.A1(new_n4347_), .A2(new_n4348_), .B(new_n3400_), .ZN(new_n4350_));
  AOI21_X1   g04158(.A1(new_n4349_), .A2(new_n4315_), .B(new_n4350_), .ZN(new_n4351_));
  AOI21_X1   g04159(.A1(new_n4351_), .A2(new_n3167_), .B(new_n4337_), .ZN(new_n4352_));
  OAI21_X1   g04160(.A1(new_n4351_), .A2(new_n3167_), .B(new_n2912_), .ZN(new_n4353_));
  OAI21_X1   g04161(.A1(new_n4352_), .A2(new_n4353_), .B(new_n4290_), .ZN(new_n4354_));
  NOR2_X1    g04162(.A1(new_n4351_), .A2(new_n3167_), .ZN(new_n4355_));
  OAI21_X1   g04163(.A1(new_n4352_), .A2(new_n4355_), .B(\asqrt[41] ), .ZN(new_n4356_));
  NAND3_X1   g04164(.A1(new_n4354_), .A2(new_n4356_), .A3(new_n2699_), .ZN(new_n4357_));
  NAND2_X1   g04165(.A1(new_n4357_), .A2(new_n4287_), .ZN(new_n4358_));
  NAND2_X1   g04166(.A1(new_n4354_), .A2(new_n4356_), .ZN(new_n4359_));
  AOI21_X1   g04167(.A1(new_n4359_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n4360_));
  AOI21_X1   g04168(.A1(new_n4360_), .A2(new_n4358_), .B(new_n4336_), .ZN(new_n4361_));
  AOI21_X1   g04169(.A1(new_n4358_), .A2(new_n4326_), .B(new_n2464_), .ZN(new_n4362_));
  OAI21_X1   g04170(.A1(new_n4361_), .A2(new_n4362_), .B(\asqrt[44] ), .ZN(new_n4363_));
  AOI21_X1   g04171(.A1(new_n4332_), .A2(new_n4363_), .B(new_n2072_), .ZN(new_n4364_));
  NOR2_X1    g04172(.A1(new_n4335_), .A2(new_n4364_), .ZN(new_n4365_));
  AOI21_X1   g04173(.A1(new_n4365_), .A2(new_n1884_), .B(new_n4276_), .ZN(new_n4366_));
  OAI21_X1   g04174(.A1(new_n4335_), .A2(new_n4364_), .B(\asqrt[46] ), .ZN(new_n4367_));
  NAND2_X1   g04175(.A1(new_n4367_), .A2(new_n1688_), .ZN(new_n4368_));
  OAI21_X1   g04176(.A1(new_n4366_), .A2(new_n4368_), .B(new_n4272_), .ZN(new_n4369_));
  INV_X1     g04177(.I(new_n4367_), .ZN(new_n4370_));
  OAI21_X1   g04178(.A1(new_n4366_), .A2(new_n4370_), .B(\asqrt[47] ), .ZN(new_n4371_));
  NAND3_X1   g04179(.A1(new_n4369_), .A2(new_n4371_), .A3(new_n1533_), .ZN(new_n4372_));
  NAND2_X1   g04180(.A1(new_n4372_), .A2(new_n4270_), .ZN(new_n4373_));
  NAND2_X1   g04181(.A1(new_n4369_), .A2(new_n4371_), .ZN(new_n4374_));
  AOI21_X1   g04182(.A1(new_n4374_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n4375_));
  AOI21_X1   g04183(.A1(new_n4375_), .A2(new_n4373_), .B(new_n4267_), .ZN(new_n4376_));
  INV_X1     g04184(.I(new_n4272_), .ZN(new_n4377_));
  INV_X1     g04185(.I(new_n4282_), .ZN(new_n4378_));
  NOR2_X1    g04186(.A1(new_n4361_), .A2(new_n4362_), .ZN(new_n4379_));
  AOI21_X1   g04187(.A1(new_n4379_), .A2(new_n2271_), .B(new_n4378_), .ZN(new_n4380_));
  NAND2_X1   g04188(.A1(new_n4363_), .A2(new_n2072_), .ZN(new_n4381_));
  OAI21_X1   g04189(.A1(new_n4380_), .A2(new_n4381_), .B(new_n4278_), .ZN(new_n4382_));
  INV_X1     g04190(.I(new_n4363_), .ZN(new_n4383_));
  OAI21_X1   g04191(.A1(new_n4380_), .A2(new_n4383_), .B(\asqrt[45] ), .ZN(new_n4384_));
  NAND3_X1   g04192(.A1(new_n4382_), .A2(new_n4384_), .A3(new_n1884_), .ZN(new_n4385_));
  NAND2_X1   g04193(.A1(new_n4385_), .A2(new_n4275_), .ZN(new_n4386_));
  NAND2_X1   g04194(.A1(new_n4382_), .A2(new_n4384_), .ZN(new_n4387_));
  AOI21_X1   g04195(.A1(new_n4387_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n4388_));
  AOI21_X1   g04196(.A1(new_n4388_), .A2(new_n4386_), .B(new_n4377_), .ZN(new_n4389_));
  AOI21_X1   g04197(.A1(new_n4386_), .A2(new_n4367_), .B(new_n1688_), .ZN(new_n4390_));
  OAI21_X1   g04198(.A1(new_n4389_), .A2(new_n4390_), .B(\asqrt[48] ), .ZN(new_n4391_));
  AOI21_X1   g04199(.A1(new_n4373_), .A2(new_n4391_), .B(new_n1368_), .ZN(new_n4392_));
  NOR2_X1    g04200(.A1(new_n4376_), .A2(new_n4392_), .ZN(new_n4393_));
  AOI21_X1   g04201(.A1(new_n4393_), .A2(new_n1228_), .B(new_n4264_), .ZN(new_n4394_));
  OAI21_X1   g04202(.A1(new_n4376_), .A2(new_n4392_), .B(\asqrt[50] ), .ZN(new_n4395_));
  NAND2_X1   g04203(.A1(new_n4395_), .A2(new_n1088_), .ZN(new_n4396_));
  OAI21_X1   g04204(.A1(new_n4394_), .A2(new_n4396_), .B(new_n4260_), .ZN(new_n4397_));
  INV_X1     g04205(.I(new_n4395_), .ZN(new_n4398_));
  OAI21_X1   g04206(.A1(new_n4394_), .A2(new_n4398_), .B(\asqrt[51] ), .ZN(new_n4399_));
  NAND3_X1   g04207(.A1(new_n4397_), .A2(new_n4399_), .A3(new_n962_), .ZN(new_n4400_));
  NAND2_X1   g04208(.A1(new_n4400_), .A2(new_n4258_), .ZN(new_n4401_));
  NAND2_X1   g04209(.A1(new_n4397_), .A2(new_n4399_), .ZN(new_n4402_));
  AOI21_X1   g04210(.A1(new_n4402_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n4403_));
  AOI21_X1   g04211(.A1(new_n4403_), .A2(new_n4401_), .B(new_n4255_), .ZN(new_n4404_));
  INV_X1     g04212(.I(new_n4260_), .ZN(new_n4405_));
  INV_X1     g04213(.I(new_n4270_), .ZN(new_n4406_));
  NOR2_X1    g04214(.A1(new_n4389_), .A2(new_n4390_), .ZN(new_n4407_));
  AOI21_X1   g04215(.A1(new_n4407_), .A2(new_n1533_), .B(new_n4406_), .ZN(new_n4408_));
  NAND2_X1   g04216(.A1(new_n4391_), .A2(new_n1368_), .ZN(new_n4409_));
  OAI21_X1   g04217(.A1(new_n4408_), .A2(new_n4409_), .B(new_n4266_), .ZN(new_n4410_));
  INV_X1     g04218(.I(new_n4391_), .ZN(new_n4411_));
  OAI21_X1   g04219(.A1(new_n4408_), .A2(new_n4411_), .B(\asqrt[49] ), .ZN(new_n4412_));
  NAND3_X1   g04220(.A1(new_n4410_), .A2(new_n4412_), .A3(new_n1228_), .ZN(new_n4413_));
  NAND2_X1   g04221(.A1(new_n4413_), .A2(new_n4263_), .ZN(new_n4414_));
  NAND2_X1   g04222(.A1(new_n4410_), .A2(new_n4412_), .ZN(new_n4415_));
  AOI21_X1   g04223(.A1(new_n4415_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n4416_));
  AOI21_X1   g04224(.A1(new_n4416_), .A2(new_n4414_), .B(new_n4405_), .ZN(new_n4417_));
  AOI21_X1   g04225(.A1(new_n4414_), .A2(new_n4395_), .B(new_n1088_), .ZN(new_n4418_));
  OAI21_X1   g04226(.A1(new_n4417_), .A2(new_n4418_), .B(\asqrt[52] ), .ZN(new_n4419_));
  AOI21_X1   g04227(.A1(new_n4401_), .A2(new_n4419_), .B(new_n842_), .ZN(new_n4420_));
  NOR2_X1    g04228(.A1(new_n4404_), .A2(new_n4420_), .ZN(new_n4421_));
  AOI21_X1   g04229(.A1(new_n4421_), .A2(new_n720_), .B(new_n4252_), .ZN(new_n4422_));
  OAI21_X1   g04230(.A1(new_n4404_), .A2(new_n4420_), .B(\asqrt[54] ), .ZN(new_n4423_));
  NAND2_X1   g04231(.A1(new_n4423_), .A2(new_n630_), .ZN(new_n4424_));
  OAI21_X1   g04232(.A1(new_n4422_), .A2(new_n4424_), .B(new_n4248_), .ZN(new_n4425_));
  INV_X1     g04233(.I(new_n4423_), .ZN(new_n4426_));
  OAI21_X1   g04234(.A1(new_n4422_), .A2(new_n4426_), .B(\asqrt[55] ), .ZN(new_n4427_));
  NAND3_X1   g04235(.A1(new_n4425_), .A2(new_n4427_), .A3(new_n545_), .ZN(new_n4428_));
  NAND2_X1   g04236(.A1(new_n4428_), .A2(new_n4246_), .ZN(new_n4429_));
  NAND2_X1   g04237(.A1(new_n4425_), .A2(new_n4427_), .ZN(new_n4430_));
  AOI21_X1   g04238(.A1(new_n4430_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n4431_));
  AOI21_X1   g04239(.A1(new_n4431_), .A2(new_n4429_), .B(new_n4243_), .ZN(new_n4432_));
  INV_X1     g04240(.I(new_n4248_), .ZN(new_n4433_));
  INV_X1     g04241(.I(new_n4258_), .ZN(new_n4434_));
  NOR2_X1    g04242(.A1(new_n4417_), .A2(new_n4418_), .ZN(new_n4435_));
  AOI21_X1   g04243(.A1(new_n4435_), .A2(new_n962_), .B(new_n4434_), .ZN(new_n4436_));
  NAND2_X1   g04244(.A1(new_n4419_), .A2(new_n842_), .ZN(new_n4437_));
  OAI21_X1   g04245(.A1(new_n4436_), .A2(new_n4437_), .B(new_n4254_), .ZN(new_n4438_));
  INV_X1     g04246(.I(new_n4419_), .ZN(new_n4439_));
  OAI21_X1   g04247(.A1(new_n4436_), .A2(new_n4439_), .B(\asqrt[53] ), .ZN(new_n4440_));
  NAND3_X1   g04248(.A1(new_n4438_), .A2(new_n4440_), .A3(new_n720_), .ZN(new_n4441_));
  NAND2_X1   g04249(.A1(new_n4441_), .A2(new_n4251_), .ZN(new_n4442_));
  NAND2_X1   g04250(.A1(new_n4438_), .A2(new_n4440_), .ZN(new_n4443_));
  AOI21_X1   g04251(.A1(new_n4443_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n4444_));
  AOI21_X1   g04252(.A1(new_n4444_), .A2(new_n4442_), .B(new_n4433_), .ZN(new_n4445_));
  AOI21_X1   g04253(.A1(new_n4442_), .A2(new_n4423_), .B(new_n630_), .ZN(new_n4446_));
  OAI21_X1   g04254(.A1(new_n4445_), .A2(new_n4446_), .B(\asqrt[56] ), .ZN(new_n4447_));
  AOI21_X1   g04255(.A1(new_n4429_), .A2(new_n4447_), .B(new_n450_), .ZN(new_n4448_));
  NOR2_X1    g04256(.A1(new_n4432_), .A2(new_n4448_), .ZN(new_n4449_));
  AOI21_X1   g04257(.A1(new_n4449_), .A2(new_n403_), .B(new_n4240_), .ZN(new_n4450_));
  OAI21_X1   g04258(.A1(new_n4432_), .A2(new_n4448_), .B(\asqrt[58] ), .ZN(new_n4451_));
  NAND2_X1   g04259(.A1(new_n4451_), .A2(new_n339_), .ZN(new_n4452_));
  OAI21_X1   g04260(.A1(new_n4450_), .A2(new_n4452_), .B(new_n4236_), .ZN(new_n4453_));
  INV_X1     g04261(.I(new_n4451_), .ZN(new_n4454_));
  OAI21_X1   g04262(.A1(new_n4450_), .A2(new_n4454_), .B(\asqrt[59] ), .ZN(new_n4455_));
  NAND3_X1   g04263(.A1(new_n4453_), .A2(new_n4455_), .A3(new_n288_), .ZN(new_n4456_));
  NAND2_X1   g04264(.A1(new_n4456_), .A2(new_n4234_), .ZN(new_n4457_));
  INV_X1     g04265(.I(new_n4236_), .ZN(new_n4458_));
  INV_X1     g04266(.I(new_n4246_), .ZN(new_n4459_));
  NOR2_X1    g04267(.A1(new_n4445_), .A2(new_n4446_), .ZN(new_n4460_));
  AOI21_X1   g04268(.A1(new_n4460_), .A2(new_n545_), .B(new_n4459_), .ZN(new_n4461_));
  NAND2_X1   g04269(.A1(new_n4447_), .A2(new_n450_), .ZN(new_n4462_));
  OAI21_X1   g04270(.A1(new_n4461_), .A2(new_n4462_), .B(new_n4242_), .ZN(new_n4463_));
  INV_X1     g04271(.I(new_n4447_), .ZN(new_n4464_));
  OAI21_X1   g04272(.A1(new_n4461_), .A2(new_n4464_), .B(\asqrt[57] ), .ZN(new_n4465_));
  NAND3_X1   g04273(.A1(new_n4463_), .A2(new_n4465_), .A3(new_n403_), .ZN(new_n4466_));
  NAND2_X1   g04274(.A1(new_n4466_), .A2(new_n4239_), .ZN(new_n4467_));
  NAND2_X1   g04275(.A1(new_n4463_), .A2(new_n4465_), .ZN(new_n4468_));
  AOI21_X1   g04276(.A1(new_n4468_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n4469_));
  AOI21_X1   g04277(.A1(new_n4469_), .A2(new_n4467_), .B(new_n4458_), .ZN(new_n4470_));
  AOI21_X1   g04278(.A1(new_n4467_), .A2(new_n4451_), .B(new_n339_), .ZN(new_n4471_));
  OAI21_X1   g04279(.A1(new_n4470_), .A2(new_n4471_), .B(\asqrt[60] ), .ZN(new_n4472_));
  AOI21_X1   g04280(.A1(new_n4457_), .A2(new_n4472_), .B(new_n242_), .ZN(new_n4473_));
  NAND2_X1   g04281(.A1(new_n4453_), .A2(new_n4455_), .ZN(new_n4474_));
  AOI21_X1   g04282(.A1(new_n4474_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n4475_));
  AOI21_X1   g04283(.A1(new_n4475_), .A2(new_n4457_), .B(new_n4208_), .ZN(new_n4476_));
  OAI21_X1   g04284(.A1(new_n4476_), .A2(new_n4473_), .B(\asqrt[62] ), .ZN(new_n4477_));
  INV_X1     g04285(.I(new_n4477_), .ZN(new_n4478_));
  NOR2_X1    g04286(.A1(new_n4476_), .A2(new_n4473_), .ZN(new_n4479_));
  AOI21_X1   g04287(.A1(new_n4183_), .A2(new_n4189_), .B(new_n4184_), .ZN(new_n4480_));
  NAND2_X1   g04288(.A1(\asqrt[36] ), .A2(new_n4480_), .ZN(new_n4481_));
  XOR2_X1    g04289(.A1(new_n4481_), .A2(new_n4187_), .Z(new_n4482_));
  INV_X1     g04290(.I(new_n4482_), .ZN(new_n4483_));
  AOI21_X1   g04291(.A1(new_n4479_), .A2(new_n234_), .B(new_n4483_), .ZN(new_n4484_));
  OAI21_X1   g04292(.A1(new_n4484_), .A2(new_n4478_), .B(new_n4231_), .ZN(new_n4485_));
  OAI21_X1   g04293(.A1(new_n4485_), .A2(new_n4230_), .B(new_n193_), .ZN(new_n4486_));
  NOR2_X1    g04294(.A1(new_n4484_), .A2(new_n4478_), .ZN(new_n4487_));
  NAND2_X1   g04295(.A1(new_n4487_), .A2(new_n4230_), .ZN(new_n4488_));
  NOR2_X1    g04296(.A1(\asqrt[36] ), .A2(new_n4219_), .ZN(new_n4489_));
  INV_X1     g04297(.I(new_n4489_), .ZN(new_n4490_));
  NAND4_X1   g04298(.A1(new_n4486_), .A2(new_n4228_), .A3(new_n4488_), .A4(new_n4490_), .ZN(\asqrt[35] ));
  AOI21_X1   g04299(.A1(new_n4457_), .A2(new_n4475_), .B(new_n4473_), .ZN(new_n4492_));
  NAND2_X1   g04300(.A1(\asqrt[35] ), .A2(new_n4492_), .ZN(new_n4493_));
  XOR2_X1    g04301(.A1(new_n4493_), .A2(new_n4208_), .Z(new_n4494_));
  INV_X1     g04302(.I(new_n4230_), .ZN(new_n4495_));
  INV_X1     g04303(.I(new_n4231_), .ZN(new_n4496_));
  INV_X1     g04304(.I(new_n4234_), .ZN(new_n4497_));
  NOR2_X1    g04305(.A1(new_n4470_), .A2(new_n4471_), .ZN(new_n4498_));
  AOI21_X1   g04306(.A1(new_n4498_), .A2(new_n288_), .B(new_n4497_), .ZN(new_n4499_));
  INV_X1     g04307(.I(new_n4472_), .ZN(new_n4500_));
  OAI21_X1   g04308(.A1(new_n4499_), .A2(new_n4500_), .B(\asqrt[61] ), .ZN(new_n4501_));
  NAND2_X1   g04309(.A1(new_n4472_), .A2(new_n242_), .ZN(new_n4502_));
  OAI21_X1   g04310(.A1(new_n4499_), .A2(new_n4502_), .B(new_n4207_), .ZN(new_n4503_));
  NAND3_X1   g04311(.A1(new_n4503_), .A2(new_n4501_), .A3(new_n234_), .ZN(new_n4504_));
  NAND2_X1   g04312(.A1(new_n4504_), .A2(new_n4482_), .ZN(new_n4505_));
  AOI21_X1   g04313(.A1(new_n4505_), .A2(new_n4477_), .B(new_n4496_), .ZN(new_n4506_));
  AOI21_X1   g04314(.A1(new_n4506_), .A2(new_n4495_), .B(\asqrt[63] ), .ZN(new_n4507_));
  NAND2_X1   g04315(.A1(new_n4505_), .A2(new_n4477_), .ZN(new_n4508_));
  NOR2_X1    g04316(.A1(new_n4508_), .A2(new_n4495_), .ZN(new_n4509_));
  NOR4_X1    g04317(.A1(new_n4507_), .A2(new_n4227_), .A3(new_n4509_), .A4(new_n4489_), .ZN(new_n4510_));
  OAI21_X1   g04318(.A1(new_n4450_), .A2(new_n4452_), .B(new_n4455_), .ZN(new_n4511_));
  NOR2_X1    g04319(.A1(new_n4510_), .A2(new_n4511_), .ZN(new_n4512_));
  XOR2_X1    g04320(.A1(new_n4512_), .A2(new_n4236_), .Z(new_n4513_));
  NAND3_X1   g04321(.A1(\asqrt[35] ), .A2(new_n4466_), .A3(new_n4451_), .ZN(new_n4514_));
  XOR2_X1    g04322(.A1(new_n4514_), .A2(new_n4240_), .Z(new_n4515_));
  OAI21_X1   g04323(.A1(new_n4461_), .A2(new_n4462_), .B(new_n4465_), .ZN(new_n4516_));
  NOR2_X1    g04324(.A1(new_n4510_), .A2(new_n4516_), .ZN(new_n4517_));
  XOR2_X1    g04325(.A1(new_n4517_), .A2(new_n4242_), .Z(new_n4518_));
  INV_X1     g04326(.I(new_n4518_), .ZN(new_n4519_));
  NAND3_X1   g04327(.A1(\asqrt[35] ), .A2(new_n4428_), .A3(new_n4447_), .ZN(new_n4520_));
  XOR2_X1    g04328(.A1(new_n4520_), .A2(new_n4459_), .Z(new_n4521_));
  INV_X1     g04329(.I(new_n4521_), .ZN(new_n4522_));
  OAI21_X1   g04330(.A1(new_n4422_), .A2(new_n4424_), .B(new_n4427_), .ZN(new_n4523_));
  NOR2_X1    g04331(.A1(new_n4510_), .A2(new_n4523_), .ZN(new_n4524_));
  XOR2_X1    g04332(.A1(new_n4524_), .A2(new_n4248_), .Z(new_n4525_));
  NAND3_X1   g04333(.A1(\asqrt[35] ), .A2(new_n4441_), .A3(new_n4423_), .ZN(new_n4526_));
  XOR2_X1    g04334(.A1(new_n4526_), .A2(new_n4252_), .Z(new_n4527_));
  OAI21_X1   g04335(.A1(new_n4436_), .A2(new_n4437_), .B(new_n4440_), .ZN(new_n4528_));
  NOR2_X1    g04336(.A1(new_n4510_), .A2(new_n4528_), .ZN(new_n4529_));
  XOR2_X1    g04337(.A1(new_n4529_), .A2(new_n4254_), .Z(new_n4530_));
  INV_X1     g04338(.I(new_n4530_), .ZN(new_n4531_));
  NAND3_X1   g04339(.A1(\asqrt[35] ), .A2(new_n4400_), .A3(new_n4419_), .ZN(new_n4532_));
  XOR2_X1    g04340(.A1(new_n4532_), .A2(new_n4434_), .Z(new_n4533_));
  INV_X1     g04341(.I(new_n4533_), .ZN(new_n4534_));
  OAI21_X1   g04342(.A1(new_n4394_), .A2(new_n4396_), .B(new_n4399_), .ZN(new_n4535_));
  NOR2_X1    g04343(.A1(new_n4510_), .A2(new_n4535_), .ZN(new_n4536_));
  XOR2_X1    g04344(.A1(new_n4536_), .A2(new_n4260_), .Z(new_n4537_));
  NAND3_X1   g04345(.A1(\asqrt[35] ), .A2(new_n4413_), .A3(new_n4395_), .ZN(new_n4538_));
  XOR2_X1    g04346(.A1(new_n4538_), .A2(new_n4264_), .Z(new_n4539_));
  OAI21_X1   g04347(.A1(new_n4408_), .A2(new_n4409_), .B(new_n4412_), .ZN(new_n4540_));
  NOR2_X1    g04348(.A1(new_n4510_), .A2(new_n4540_), .ZN(new_n4541_));
  XOR2_X1    g04349(.A1(new_n4541_), .A2(new_n4266_), .Z(new_n4542_));
  INV_X1     g04350(.I(new_n4542_), .ZN(new_n4543_));
  NAND3_X1   g04351(.A1(\asqrt[35] ), .A2(new_n4372_), .A3(new_n4391_), .ZN(new_n4544_));
  XOR2_X1    g04352(.A1(new_n4544_), .A2(new_n4406_), .Z(new_n4545_));
  INV_X1     g04353(.I(new_n4545_), .ZN(new_n4546_));
  OAI21_X1   g04354(.A1(new_n4366_), .A2(new_n4368_), .B(new_n4371_), .ZN(new_n4547_));
  NOR2_X1    g04355(.A1(new_n4510_), .A2(new_n4547_), .ZN(new_n4548_));
  XOR2_X1    g04356(.A1(new_n4548_), .A2(new_n4272_), .Z(new_n4549_));
  NAND3_X1   g04357(.A1(\asqrt[35] ), .A2(new_n4385_), .A3(new_n4367_), .ZN(new_n4550_));
  XOR2_X1    g04358(.A1(new_n4550_), .A2(new_n4276_), .Z(new_n4551_));
  OAI21_X1   g04359(.A1(new_n4380_), .A2(new_n4381_), .B(new_n4384_), .ZN(new_n4552_));
  NOR2_X1    g04360(.A1(new_n4510_), .A2(new_n4552_), .ZN(new_n4553_));
  XOR2_X1    g04361(.A1(new_n4553_), .A2(new_n4278_), .Z(new_n4554_));
  INV_X1     g04362(.I(new_n4554_), .ZN(new_n4555_));
  NAND3_X1   g04363(.A1(\asqrt[35] ), .A2(new_n4331_), .A3(new_n4363_), .ZN(new_n4556_));
  XOR2_X1    g04364(.A1(new_n4556_), .A2(new_n4378_), .Z(new_n4557_));
  INV_X1     g04365(.I(new_n4557_), .ZN(new_n4558_));
  OAI21_X1   g04366(.A1(new_n4325_), .A2(new_n4327_), .B(new_n4330_), .ZN(new_n4559_));
  NOR2_X1    g04367(.A1(new_n4510_), .A2(new_n4559_), .ZN(new_n4560_));
  XOR2_X1    g04368(.A1(new_n4560_), .A2(new_n4284_), .Z(new_n4561_));
  NAND3_X1   g04369(.A1(\asqrt[35] ), .A2(new_n4357_), .A3(new_n4326_), .ZN(new_n4562_));
  XOR2_X1    g04370(.A1(new_n4562_), .A2(new_n4288_), .Z(new_n4563_));
  AOI21_X1   g04371(.A1(new_n4319_), .A2(new_n4320_), .B(new_n4323_), .ZN(new_n4564_));
  NAND2_X1   g04372(.A1(\asqrt[35] ), .A2(new_n4564_), .ZN(new_n4565_));
  XOR2_X1    g04373(.A1(new_n4565_), .A2(new_n4291_), .Z(new_n4566_));
  INV_X1     g04374(.I(new_n4566_), .ZN(new_n4567_));
  NOR2_X1    g04375(.A1(new_n4318_), .A2(\asqrt[40] ), .ZN(new_n4568_));
  NOR3_X1    g04376(.A1(new_n4510_), .A2(new_n4568_), .A3(new_n4355_), .ZN(new_n4569_));
  XOR2_X1    g04377(.A1(new_n4569_), .A2(new_n4294_), .Z(new_n4570_));
  INV_X1     g04378(.I(new_n4570_), .ZN(new_n4571_));
  NOR3_X1    g04379(.A1(new_n4510_), .A2(new_n4313_), .A3(new_n4350_), .ZN(new_n4572_));
  XOR2_X1    g04380(.A1(new_n4572_), .A2(new_n4315_), .Z(new_n4573_));
  NOR2_X1    g04381(.A1(new_n4346_), .A2(\asqrt[38] ), .ZN(new_n4574_));
  NOR3_X1    g04382(.A1(new_n4510_), .A2(new_n4574_), .A3(new_n4312_), .ZN(new_n4575_));
  XOR2_X1    g04383(.A1(new_n4575_), .A2(new_n4340_), .Z(new_n4576_));
  NOR3_X1    g04384(.A1(new_n4510_), .A2(\a[70] ), .A3(\a[71] ), .ZN(new_n4577_));
  NAND4_X1   g04385(.A1(new_n4486_), .A2(\asqrt[36] ), .A3(new_n4488_), .A4(new_n4228_), .ZN(new_n4578_));
  INV_X1     g04386(.I(new_n4578_), .ZN(new_n4579_));
  OAI21_X1   g04387(.A1(new_n4577_), .A2(new_n4579_), .B(new_n4009_), .ZN(new_n4580_));
  NAND3_X1   g04388(.A1(\asqrt[35] ), .A2(new_n4302_), .A3(new_n4303_), .ZN(new_n4581_));
  NAND3_X1   g04389(.A1(new_n4581_), .A2(\a[72] ), .A3(new_n4578_), .ZN(new_n4582_));
  NAND2_X1   g04390(.A1(new_n4580_), .A2(new_n4582_), .ZN(new_n4583_));
  INV_X1     g04391(.I(\a[68] ), .ZN(new_n4584_));
  INV_X1     g04392(.I(\a[69] ), .ZN(new_n4585_));
  NAND3_X1   g04393(.A1(new_n4584_), .A2(new_n4585_), .A3(new_n4302_), .ZN(new_n4586_));
  NAND2_X1   g04394(.A1(\asqrt[35] ), .A2(\a[70] ), .ZN(new_n4587_));
  AOI21_X1   g04395(.A1(new_n4587_), .A2(new_n4586_), .B(new_n4224_), .ZN(new_n4588_));
  AOI21_X1   g04396(.A1(\asqrt[35] ), .A2(new_n4302_), .B(new_n4303_), .ZN(new_n4589_));
  NOR2_X1    g04397(.A1(new_n4577_), .A2(new_n4589_), .ZN(new_n4590_));
  NAND3_X1   g04398(.A1(new_n4587_), .A2(new_n4224_), .A3(new_n4586_), .ZN(new_n4591_));
  AOI21_X1   g04399(.A1(new_n4590_), .A2(new_n4591_), .B(new_n4588_), .ZN(new_n4592_));
  AOI21_X1   g04400(.A1(new_n4592_), .A2(new_n3928_), .B(new_n4583_), .ZN(new_n4593_));
  NOR2_X1    g04401(.A1(new_n4592_), .A2(new_n3928_), .ZN(new_n4594_));
  NOR2_X1    g04402(.A1(new_n4593_), .A2(new_n4594_), .ZN(new_n4595_));
  NOR3_X1    g04403(.A1(new_n4510_), .A2(new_n4306_), .A3(new_n4345_), .ZN(new_n4596_));
  XOR2_X1    g04404(.A1(new_n4596_), .A2(new_n4308_), .Z(new_n4597_));
  INV_X1     g04405(.I(new_n4597_), .ZN(new_n4598_));
  AOI21_X1   g04406(.A1(new_n4595_), .A2(new_n3675_), .B(new_n4598_), .ZN(new_n4599_));
  OAI21_X1   g04407(.A1(new_n4593_), .A2(new_n4594_), .B(\asqrt[38] ), .ZN(new_n4600_));
  NAND2_X1   g04408(.A1(new_n4600_), .A2(new_n3400_), .ZN(new_n4601_));
  OAI21_X1   g04409(.A1(new_n4599_), .A2(new_n4601_), .B(new_n4576_), .ZN(new_n4602_));
  INV_X1     g04410(.I(new_n4600_), .ZN(new_n4603_));
  OAI21_X1   g04411(.A1(new_n4599_), .A2(new_n4603_), .B(\asqrt[39] ), .ZN(new_n4604_));
  NAND3_X1   g04412(.A1(new_n4602_), .A2(new_n4604_), .A3(new_n3167_), .ZN(new_n4605_));
  NAND2_X1   g04413(.A1(new_n4605_), .A2(new_n4573_), .ZN(new_n4606_));
  NAND2_X1   g04414(.A1(new_n4602_), .A2(new_n4604_), .ZN(new_n4607_));
  AOI21_X1   g04415(.A1(new_n4607_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n4608_));
  AOI21_X1   g04416(.A1(new_n4608_), .A2(new_n4606_), .B(new_n4571_), .ZN(new_n4609_));
  INV_X1     g04417(.I(new_n4576_), .ZN(new_n4610_));
  AOI21_X1   g04418(.A1(new_n4581_), .A2(new_n4578_), .B(\a[72] ), .ZN(new_n4611_));
  NOR3_X1    g04419(.A1(new_n4577_), .A2(new_n4009_), .A3(new_n4579_), .ZN(new_n4612_));
  NOR2_X1    g04420(.A1(new_n4612_), .A2(new_n4611_), .ZN(new_n4613_));
  OAI21_X1   g04421(.A1(new_n4510_), .A2(new_n4302_), .B(new_n4586_), .ZN(new_n4614_));
  NAND2_X1   g04422(.A1(new_n4614_), .A2(\asqrt[36] ), .ZN(new_n4615_));
  OAI21_X1   g04423(.A1(new_n4510_), .A2(\a[70] ), .B(\a[71] ), .ZN(new_n4616_));
  NAND2_X1   g04424(.A1(new_n4616_), .A2(new_n4581_), .ZN(new_n4617_));
  NOR2_X1    g04425(.A1(new_n4614_), .A2(\asqrt[36] ), .ZN(new_n4618_));
  OAI21_X1   g04426(.A1(new_n4617_), .A2(new_n4618_), .B(new_n4615_), .ZN(new_n4619_));
  OAI21_X1   g04427(.A1(new_n4619_), .A2(\asqrt[37] ), .B(new_n4613_), .ZN(new_n4620_));
  NAND2_X1   g04428(.A1(new_n4619_), .A2(\asqrt[37] ), .ZN(new_n4621_));
  NAND3_X1   g04429(.A1(new_n4620_), .A2(new_n3675_), .A3(new_n4621_), .ZN(new_n4622_));
  NAND2_X1   g04430(.A1(new_n4622_), .A2(new_n4597_), .ZN(new_n4623_));
  NAND2_X1   g04431(.A1(new_n4620_), .A2(new_n4621_), .ZN(new_n4624_));
  AOI21_X1   g04432(.A1(new_n4624_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n4625_));
  AOI21_X1   g04433(.A1(new_n4625_), .A2(new_n4623_), .B(new_n4610_), .ZN(new_n4626_));
  AOI21_X1   g04434(.A1(new_n4623_), .A2(new_n4600_), .B(new_n3400_), .ZN(new_n4627_));
  OAI21_X1   g04435(.A1(new_n4626_), .A2(new_n4627_), .B(\asqrt[40] ), .ZN(new_n4628_));
  AOI21_X1   g04436(.A1(new_n4606_), .A2(new_n4628_), .B(new_n2912_), .ZN(new_n4629_));
  NOR2_X1    g04437(.A1(new_n4609_), .A2(new_n4629_), .ZN(new_n4630_));
  AOI21_X1   g04438(.A1(new_n4630_), .A2(new_n2699_), .B(new_n4567_), .ZN(new_n4631_));
  OAI21_X1   g04439(.A1(new_n4609_), .A2(new_n4629_), .B(\asqrt[42] ), .ZN(new_n4632_));
  NAND2_X1   g04440(.A1(new_n4632_), .A2(new_n2464_), .ZN(new_n4633_));
  OAI21_X1   g04441(.A1(new_n4631_), .A2(new_n4633_), .B(new_n4563_), .ZN(new_n4634_));
  INV_X1     g04442(.I(new_n4632_), .ZN(new_n4635_));
  OAI21_X1   g04443(.A1(new_n4631_), .A2(new_n4635_), .B(\asqrt[43] ), .ZN(new_n4636_));
  NAND3_X1   g04444(.A1(new_n4634_), .A2(new_n4636_), .A3(new_n2271_), .ZN(new_n4637_));
  NAND2_X1   g04445(.A1(new_n4637_), .A2(new_n4561_), .ZN(new_n4638_));
  NAND2_X1   g04446(.A1(new_n4634_), .A2(new_n4636_), .ZN(new_n4639_));
  AOI21_X1   g04447(.A1(new_n4639_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n4640_));
  AOI21_X1   g04448(.A1(new_n4640_), .A2(new_n4638_), .B(new_n4558_), .ZN(new_n4641_));
  INV_X1     g04449(.I(new_n4563_), .ZN(new_n4642_));
  INV_X1     g04450(.I(new_n4573_), .ZN(new_n4643_));
  NOR2_X1    g04451(.A1(new_n4626_), .A2(new_n4627_), .ZN(new_n4644_));
  AOI21_X1   g04452(.A1(new_n4644_), .A2(new_n3167_), .B(new_n4643_), .ZN(new_n4645_));
  NAND2_X1   g04453(.A1(new_n4628_), .A2(new_n2912_), .ZN(new_n4646_));
  OAI21_X1   g04454(.A1(new_n4645_), .A2(new_n4646_), .B(new_n4570_), .ZN(new_n4647_));
  INV_X1     g04455(.I(new_n4628_), .ZN(new_n4648_));
  OAI21_X1   g04456(.A1(new_n4645_), .A2(new_n4648_), .B(\asqrt[41] ), .ZN(new_n4649_));
  NAND3_X1   g04457(.A1(new_n4647_), .A2(new_n4649_), .A3(new_n2699_), .ZN(new_n4650_));
  NAND2_X1   g04458(.A1(new_n4650_), .A2(new_n4566_), .ZN(new_n4651_));
  NAND2_X1   g04459(.A1(new_n4647_), .A2(new_n4649_), .ZN(new_n4652_));
  AOI21_X1   g04460(.A1(new_n4652_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n4653_));
  AOI21_X1   g04461(.A1(new_n4653_), .A2(new_n4651_), .B(new_n4642_), .ZN(new_n4654_));
  AOI21_X1   g04462(.A1(new_n4651_), .A2(new_n4632_), .B(new_n2464_), .ZN(new_n4655_));
  OAI21_X1   g04463(.A1(new_n4654_), .A2(new_n4655_), .B(\asqrt[44] ), .ZN(new_n4656_));
  AOI21_X1   g04464(.A1(new_n4638_), .A2(new_n4656_), .B(new_n2072_), .ZN(new_n4657_));
  NOR2_X1    g04465(.A1(new_n4641_), .A2(new_n4657_), .ZN(new_n4658_));
  AOI21_X1   g04466(.A1(new_n4658_), .A2(new_n1884_), .B(new_n4555_), .ZN(new_n4659_));
  OAI21_X1   g04467(.A1(new_n4641_), .A2(new_n4657_), .B(\asqrt[46] ), .ZN(new_n4660_));
  NAND2_X1   g04468(.A1(new_n4660_), .A2(new_n1688_), .ZN(new_n4661_));
  OAI21_X1   g04469(.A1(new_n4659_), .A2(new_n4661_), .B(new_n4551_), .ZN(new_n4662_));
  INV_X1     g04470(.I(new_n4660_), .ZN(new_n4663_));
  OAI21_X1   g04471(.A1(new_n4659_), .A2(new_n4663_), .B(\asqrt[47] ), .ZN(new_n4664_));
  NAND3_X1   g04472(.A1(new_n4662_), .A2(new_n4664_), .A3(new_n1533_), .ZN(new_n4665_));
  NAND2_X1   g04473(.A1(new_n4665_), .A2(new_n4549_), .ZN(new_n4666_));
  NAND2_X1   g04474(.A1(new_n4662_), .A2(new_n4664_), .ZN(new_n4667_));
  AOI21_X1   g04475(.A1(new_n4667_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n4668_));
  AOI21_X1   g04476(.A1(new_n4668_), .A2(new_n4666_), .B(new_n4546_), .ZN(new_n4669_));
  INV_X1     g04477(.I(new_n4551_), .ZN(new_n4670_));
  INV_X1     g04478(.I(new_n4561_), .ZN(new_n4671_));
  NOR2_X1    g04479(.A1(new_n4654_), .A2(new_n4655_), .ZN(new_n4672_));
  AOI21_X1   g04480(.A1(new_n4672_), .A2(new_n2271_), .B(new_n4671_), .ZN(new_n4673_));
  NAND2_X1   g04481(.A1(new_n4656_), .A2(new_n2072_), .ZN(new_n4674_));
  OAI21_X1   g04482(.A1(new_n4673_), .A2(new_n4674_), .B(new_n4557_), .ZN(new_n4675_));
  INV_X1     g04483(.I(new_n4656_), .ZN(new_n4676_));
  OAI21_X1   g04484(.A1(new_n4673_), .A2(new_n4676_), .B(\asqrt[45] ), .ZN(new_n4677_));
  NAND3_X1   g04485(.A1(new_n4675_), .A2(new_n4677_), .A3(new_n1884_), .ZN(new_n4678_));
  NAND2_X1   g04486(.A1(new_n4678_), .A2(new_n4554_), .ZN(new_n4679_));
  NAND2_X1   g04487(.A1(new_n4675_), .A2(new_n4677_), .ZN(new_n4680_));
  AOI21_X1   g04488(.A1(new_n4680_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n4681_));
  AOI21_X1   g04489(.A1(new_n4681_), .A2(new_n4679_), .B(new_n4670_), .ZN(new_n4682_));
  AOI21_X1   g04490(.A1(new_n4679_), .A2(new_n4660_), .B(new_n1688_), .ZN(new_n4683_));
  OAI21_X1   g04491(.A1(new_n4682_), .A2(new_n4683_), .B(\asqrt[48] ), .ZN(new_n4684_));
  AOI21_X1   g04492(.A1(new_n4666_), .A2(new_n4684_), .B(new_n1368_), .ZN(new_n4685_));
  NOR2_X1    g04493(.A1(new_n4669_), .A2(new_n4685_), .ZN(new_n4686_));
  AOI21_X1   g04494(.A1(new_n4686_), .A2(new_n1228_), .B(new_n4543_), .ZN(new_n4687_));
  OAI21_X1   g04495(.A1(new_n4669_), .A2(new_n4685_), .B(\asqrt[50] ), .ZN(new_n4688_));
  NAND2_X1   g04496(.A1(new_n4688_), .A2(new_n1088_), .ZN(new_n4689_));
  OAI21_X1   g04497(.A1(new_n4687_), .A2(new_n4689_), .B(new_n4539_), .ZN(new_n4690_));
  INV_X1     g04498(.I(new_n4688_), .ZN(new_n4691_));
  OAI21_X1   g04499(.A1(new_n4687_), .A2(new_n4691_), .B(\asqrt[51] ), .ZN(new_n4692_));
  NAND3_X1   g04500(.A1(new_n4690_), .A2(new_n4692_), .A3(new_n962_), .ZN(new_n4693_));
  NAND2_X1   g04501(.A1(new_n4693_), .A2(new_n4537_), .ZN(new_n4694_));
  NAND2_X1   g04502(.A1(new_n4690_), .A2(new_n4692_), .ZN(new_n4695_));
  AOI21_X1   g04503(.A1(new_n4695_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n4696_));
  AOI21_X1   g04504(.A1(new_n4696_), .A2(new_n4694_), .B(new_n4534_), .ZN(new_n4697_));
  INV_X1     g04505(.I(new_n4539_), .ZN(new_n4698_));
  INV_X1     g04506(.I(new_n4549_), .ZN(new_n4699_));
  NOR2_X1    g04507(.A1(new_n4682_), .A2(new_n4683_), .ZN(new_n4700_));
  AOI21_X1   g04508(.A1(new_n4700_), .A2(new_n1533_), .B(new_n4699_), .ZN(new_n4701_));
  NAND2_X1   g04509(.A1(new_n4684_), .A2(new_n1368_), .ZN(new_n4702_));
  OAI21_X1   g04510(.A1(new_n4701_), .A2(new_n4702_), .B(new_n4545_), .ZN(new_n4703_));
  INV_X1     g04511(.I(new_n4684_), .ZN(new_n4704_));
  OAI21_X1   g04512(.A1(new_n4701_), .A2(new_n4704_), .B(\asqrt[49] ), .ZN(new_n4705_));
  NAND3_X1   g04513(.A1(new_n4703_), .A2(new_n4705_), .A3(new_n1228_), .ZN(new_n4706_));
  NAND2_X1   g04514(.A1(new_n4706_), .A2(new_n4542_), .ZN(new_n4707_));
  NAND2_X1   g04515(.A1(new_n4703_), .A2(new_n4705_), .ZN(new_n4708_));
  AOI21_X1   g04516(.A1(new_n4708_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n4709_));
  AOI21_X1   g04517(.A1(new_n4709_), .A2(new_n4707_), .B(new_n4698_), .ZN(new_n4710_));
  AOI21_X1   g04518(.A1(new_n4707_), .A2(new_n4688_), .B(new_n1088_), .ZN(new_n4711_));
  OAI21_X1   g04519(.A1(new_n4710_), .A2(new_n4711_), .B(\asqrt[52] ), .ZN(new_n4712_));
  AOI21_X1   g04520(.A1(new_n4694_), .A2(new_n4712_), .B(new_n842_), .ZN(new_n4713_));
  NOR2_X1    g04521(.A1(new_n4697_), .A2(new_n4713_), .ZN(new_n4714_));
  AOI21_X1   g04522(.A1(new_n4714_), .A2(new_n720_), .B(new_n4531_), .ZN(new_n4715_));
  OAI21_X1   g04523(.A1(new_n4697_), .A2(new_n4713_), .B(\asqrt[54] ), .ZN(new_n4716_));
  NAND2_X1   g04524(.A1(new_n4716_), .A2(new_n630_), .ZN(new_n4717_));
  OAI21_X1   g04525(.A1(new_n4715_), .A2(new_n4717_), .B(new_n4527_), .ZN(new_n4718_));
  INV_X1     g04526(.I(new_n4716_), .ZN(new_n4719_));
  OAI21_X1   g04527(.A1(new_n4715_), .A2(new_n4719_), .B(\asqrt[55] ), .ZN(new_n4720_));
  NAND3_X1   g04528(.A1(new_n4718_), .A2(new_n4720_), .A3(new_n545_), .ZN(new_n4721_));
  NAND2_X1   g04529(.A1(new_n4721_), .A2(new_n4525_), .ZN(new_n4722_));
  NAND2_X1   g04530(.A1(new_n4718_), .A2(new_n4720_), .ZN(new_n4723_));
  AOI21_X1   g04531(.A1(new_n4723_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n4724_));
  AOI21_X1   g04532(.A1(new_n4724_), .A2(new_n4722_), .B(new_n4522_), .ZN(new_n4725_));
  INV_X1     g04533(.I(new_n4527_), .ZN(new_n4726_));
  INV_X1     g04534(.I(new_n4537_), .ZN(new_n4727_));
  NOR2_X1    g04535(.A1(new_n4710_), .A2(new_n4711_), .ZN(new_n4728_));
  AOI21_X1   g04536(.A1(new_n4728_), .A2(new_n962_), .B(new_n4727_), .ZN(new_n4729_));
  NAND2_X1   g04537(.A1(new_n4712_), .A2(new_n842_), .ZN(new_n4730_));
  OAI21_X1   g04538(.A1(new_n4729_), .A2(new_n4730_), .B(new_n4533_), .ZN(new_n4731_));
  INV_X1     g04539(.I(new_n4712_), .ZN(new_n4732_));
  OAI21_X1   g04540(.A1(new_n4729_), .A2(new_n4732_), .B(\asqrt[53] ), .ZN(new_n4733_));
  NAND3_X1   g04541(.A1(new_n4731_), .A2(new_n4733_), .A3(new_n720_), .ZN(new_n4734_));
  NAND2_X1   g04542(.A1(new_n4734_), .A2(new_n4530_), .ZN(new_n4735_));
  NAND2_X1   g04543(.A1(new_n4731_), .A2(new_n4733_), .ZN(new_n4736_));
  AOI21_X1   g04544(.A1(new_n4736_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n4737_));
  AOI21_X1   g04545(.A1(new_n4737_), .A2(new_n4735_), .B(new_n4726_), .ZN(new_n4738_));
  AOI21_X1   g04546(.A1(new_n4735_), .A2(new_n4716_), .B(new_n630_), .ZN(new_n4739_));
  OAI21_X1   g04547(.A1(new_n4738_), .A2(new_n4739_), .B(\asqrt[56] ), .ZN(new_n4740_));
  AOI21_X1   g04548(.A1(new_n4722_), .A2(new_n4740_), .B(new_n450_), .ZN(new_n4741_));
  NOR2_X1    g04549(.A1(new_n4725_), .A2(new_n4741_), .ZN(new_n4742_));
  AOI21_X1   g04550(.A1(new_n4742_), .A2(new_n403_), .B(new_n4519_), .ZN(new_n4743_));
  OAI21_X1   g04551(.A1(new_n4725_), .A2(new_n4741_), .B(\asqrt[58] ), .ZN(new_n4744_));
  NAND2_X1   g04552(.A1(new_n4744_), .A2(new_n339_), .ZN(new_n4745_));
  OAI21_X1   g04553(.A1(new_n4743_), .A2(new_n4745_), .B(new_n4515_), .ZN(new_n4746_));
  INV_X1     g04554(.I(new_n4744_), .ZN(new_n4747_));
  OAI21_X1   g04555(.A1(new_n4743_), .A2(new_n4747_), .B(\asqrt[59] ), .ZN(new_n4748_));
  NAND3_X1   g04556(.A1(new_n4746_), .A2(new_n4748_), .A3(new_n288_), .ZN(new_n4749_));
  NAND2_X1   g04557(.A1(new_n4749_), .A2(new_n4513_), .ZN(new_n4750_));
  INV_X1     g04558(.I(new_n4515_), .ZN(new_n4751_));
  INV_X1     g04559(.I(new_n4525_), .ZN(new_n4752_));
  NOR2_X1    g04560(.A1(new_n4738_), .A2(new_n4739_), .ZN(new_n4753_));
  AOI21_X1   g04561(.A1(new_n4753_), .A2(new_n545_), .B(new_n4752_), .ZN(new_n4754_));
  NAND2_X1   g04562(.A1(new_n4740_), .A2(new_n450_), .ZN(new_n4755_));
  OAI21_X1   g04563(.A1(new_n4754_), .A2(new_n4755_), .B(new_n4521_), .ZN(new_n4756_));
  INV_X1     g04564(.I(new_n4740_), .ZN(new_n4757_));
  OAI21_X1   g04565(.A1(new_n4754_), .A2(new_n4757_), .B(\asqrt[57] ), .ZN(new_n4758_));
  NAND3_X1   g04566(.A1(new_n4756_), .A2(new_n4758_), .A3(new_n403_), .ZN(new_n4759_));
  NAND2_X1   g04567(.A1(new_n4759_), .A2(new_n4518_), .ZN(new_n4760_));
  NAND2_X1   g04568(.A1(new_n4756_), .A2(new_n4758_), .ZN(new_n4761_));
  AOI21_X1   g04569(.A1(new_n4761_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n4762_));
  AOI21_X1   g04570(.A1(new_n4762_), .A2(new_n4760_), .B(new_n4751_), .ZN(new_n4763_));
  AOI21_X1   g04571(.A1(new_n4760_), .A2(new_n4744_), .B(new_n339_), .ZN(new_n4764_));
  OAI21_X1   g04572(.A1(new_n4763_), .A2(new_n4764_), .B(\asqrt[60] ), .ZN(new_n4765_));
  AOI21_X1   g04573(.A1(new_n4750_), .A2(new_n4765_), .B(new_n242_), .ZN(new_n4766_));
  NAND3_X1   g04574(.A1(\asqrt[35] ), .A2(new_n4456_), .A3(new_n4472_), .ZN(new_n4767_));
  XOR2_X1    g04575(.A1(new_n4767_), .A2(new_n4497_), .Z(new_n4768_));
  INV_X1     g04576(.I(new_n4768_), .ZN(new_n4769_));
  NAND2_X1   g04577(.A1(new_n4746_), .A2(new_n4748_), .ZN(new_n4770_));
  AOI21_X1   g04578(.A1(new_n4770_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n4771_));
  AOI21_X1   g04579(.A1(new_n4771_), .A2(new_n4750_), .B(new_n4769_), .ZN(new_n4772_));
  OAI21_X1   g04580(.A1(new_n4772_), .A2(new_n4766_), .B(\asqrt[62] ), .ZN(new_n4773_));
  INV_X1     g04581(.I(new_n4513_), .ZN(new_n4774_));
  NOR2_X1    g04582(.A1(new_n4763_), .A2(new_n4764_), .ZN(new_n4775_));
  AOI21_X1   g04583(.A1(new_n4775_), .A2(new_n288_), .B(new_n4774_), .ZN(new_n4776_));
  INV_X1     g04584(.I(new_n4765_), .ZN(new_n4777_));
  OAI21_X1   g04585(.A1(new_n4776_), .A2(new_n4777_), .B(\asqrt[61] ), .ZN(new_n4778_));
  NAND2_X1   g04586(.A1(new_n4765_), .A2(new_n242_), .ZN(new_n4779_));
  OAI21_X1   g04587(.A1(new_n4776_), .A2(new_n4779_), .B(new_n4768_), .ZN(new_n4780_));
  NAND3_X1   g04588(.A1(new_n4780_), .A2(new_n4778_), .A3(new_n234_), .ZN(new_n4781_));
  NAND2_X1   g04589(.A1(new_n4508_), .A2(new_n4230_), .ZN(new_n4782_));
  NOR2_X1    g04590(.A1(new_n4510_), .A2(new_n4230_), .ZN(new_n4783_));
  NAND2_X1   g04591(.A1(new_n4783_), .A2(new_n4487_), .ZN(new_n4784_));
  AOI21_X1   g04592(.A1(new_n4784_), .A2(new_n4782_), .B(new_n193_), .ZN(new_n4785_));
  INV_X1     g04593(.I(new_n4785_), .ZN(new_n4786_));
  NAND3_X1   g04594(.A1(\asqrt[35] ), .A2(new_n4477_), .A3(new_n4504_), .ZN(new_n4787_));
  XOR2_X1    g04595(.A1(new_n4787_), .A2(new_n4482_), .Z(new_n4788_));
  INV_X1     g04596(.I(new_n4773_), .ZN(new_n4789_));
  AOI21_X1   g04597(.A1(new_n4783_), .A2(new_n4508_), .B(new_n4509_), .ZN(new_n4790_));
  INV_X1     g04598(.I(new_n4494_), .ZN(new_n4791_));
  NOR2_X1    g04599(.A1(new_n4772_), .A2(new_n4766_), .ZN(new_n4792_));
  AOI21_X1   g04600(.A1(new_n4792_), .A2(new_n234_), .B(new_n4791_), .ZN(new_n4793_));
  OAI21_X1   g04601(.A1(new_n4793_), .A2(new_n4789_), .B(new_n4790_), .ZN(new_n4794_));
  OAI21_X1   g04602(.A1(new_n4794_), .A2(new_n4788_), .B(new_n193_), .ZN(new_n4795_));
  NOR2_X1    g04603(.A1(new_n4793_), .A2(new_n4789_), .ZN(new_n4796_));
  NAND2_X1   g04604(.A1(new_n4796_), .A2(new_n4788_), .ZN(new_n4797_));
  NOR2_X1    g04605(.A1(\asqrt[35] ), .A2(new_n4495_), .ZN(new_n4798_));
  INV_X1     g04606(.I(new_n4798_), .ZN(new_n4799_));
  NAND4_X1   g04607(.A1(new_n4795_), .A2(new_n4786_), .A3(new_n4797_), .A4(new_n4799_), .ZN(\asqrt[34] ));
  NAND3_X1   g04608(.A1(\asqrt[34] ), .A2(new_n4773_), .A3(new_n4781_), .ZN(new_n4801_));
  XOR2_X1    g04609(.A1(new_n4801_), .A2(new_n4494_), .Z(new_n4802_));
  INV_X1     g04610(.I(new_n4788_), .ZN(new_n4803_));
  INV_X1     g04611(.I(new_n4790_), .ZN(new_n4804_));
  NAND2_X1   g04612(.A1(new_n4781_), .A2(new_n4494_), .ZN(new_n4805_));
  AOI21_X1   g04613(.A1(new_n4805_), .A2(new_n4773_), .B(new_n4804_), .ZN(new_n4806_));
  AOI21_X1   g04614(.A1(new_n4806_), .A2(new_n4803_), .B(\asqrt[63] ), .ZN(new_n4807_));
  NAND2_X1   g04615(.A1(new_n4805_), .A2(new_n4773_), .ZN(new_n4808_));
  NOR2_X1    g04616(.A1(new_n4808_), .A2(new_n4803_), .ZN(new_n4809_));
  NOR4_X1    g04617(.A1(new_n4807_), .A2(new_n4785_), .A3(new_n4809_), .A4(new_n4798_), .ZN(new_n4810_));
  OAI21_X1   g04618(.A1(new_n4743_), .A2(new_n4745_), .B(new_n4748_), .ZN(new_n4811_));
  NOR2_X1    g04619(.A1(new_n4810_), .A2(new_n4811_), .ZN(new_n4812_));
  XOR2_X1    g04620(.A1(new_n4812_), .A2(new_n4515_), .Z(new_n4813_));
  NAND3_X1   g04621(.A1(\asqrt[34] ), .A2(new_n4759_), .A3(new_n4744_), .ZN(new_n4814_));
  XOR2_X1    g04622(.A1(new_n4814_), .A2(new_n4519_), .Z(new_n4815_));
  OAI21_X1   g04623(.A1(new_n4754_), .A2(new_n4755_), .B(new_n4758_), .ZN(new_n4816_));
  NOR2_X1    g04624(.A1(new_n4810_), .A2(new_n4816_), .ZN(new_n4817_));
  XOR2_X1    g04625(.A1(new_n4817_), .A2(new_n4521_), .Z(new_n4818_));
  INV_X1     g04626(.I(new_n4818_), .ZN(new_n4819_));
  NAND3_X1   g04627(.A1(\asqrt[34] ), .A2(new_n4721_), .A3(new_n4740_), .ZN(new_n4820_));
  XOR2_X1    g04628(.A1(new_n4820_), .A2(new_n4752_), .Z(new_n4821_));
  INV_X1     g04629(.I(new_n4821_), .ZN(new_n4822_));
  OAI21_X1   g04630(.A1(new_n4715_), .A2(new_n4717_), .B(new_n4720_), .ZN(new_n4823_));
  NOR2_X1    g04631(.A1(new_n4810_), .A2(new_n4823_), .ZN(new_n4824_));
  XOR2_X1    g04632(.A1(new_n4824_), .A2(new_n4527_), .Z(new_n4825_));
  NAND3_X1   g04633(.A1(\asqrt[34] ), .A2(new_n4734_), .A3(new_n4716_), .ZN(new_n4826_));
  XOR2_X1    g04634(.A1(new_n4826_), .A2(new_n4531_), .Z(new_n4827_));
  OAI21_X1   g04635(.A1(new_n4729_), .A2(new_n4730_), .B(new_n4733_), .ZN(new_n4828_));
  NOR2_X1    g04636(.A1(new_n4810_), .A2(new_n4828_), .ZN(new_n4829_));
  XOR2_X1    g04637(.A1(new_n4829_), .A2(new_n4533_), .Z(new_n4830_));
  INV_X1     g04638(.I(new_n4830_), .ZN(new_n4831_));
  NAND3_X1   g04639(.A1(\asqrt[34] ), .A2(new_n4693_), .A3(new_n4712_), .ZN(new_n4832_));
  XOR2_X1    g04640(.A1(new_n4832_), .A2(new_n4727_), .Z(new_n4833_));
  INV_X1     g04641(.I(new_n4833_), .ZN(new_n4834_));
  OAI21_X1   g04642(.A1(new_n4687_), .A2(new_n4689_), .B(new_n4692_), .ZN(new_n4835_));
  NOR2_X1    g04643(.A1(new_n4810_), .A2(new_n4835_), .ZN(new_n4836_));
  XOR2_X1    g04644(.A1(new_n4836_), .A2(new_n4539_), .Z(new_n4837_));
  NAND3_X1   g04645(.A1(\asqrt[34] ), .A2(new_n4706_), .A3(new_n4688_), .ZN(new_n4838_));
  XOR2_X1    g04646(.A1(new_n4838_), .A2(new_n4543_), .Z(new_n4839_));
  OAI21_X1   g04647(.A1(new_n4701_), .A2(new_n4702_), .B(new_n4705_), .ZN(new_n4840_));
  NOR2_X1    g04648(.A1(new_n4810_), .A2(new_n4840_), .ZN(new_n4841_));
  XOR2_X1    g04649(.A1(new_n4841_), .A2(new_n4545_), .Z(new_n4842_));
  INV_X1     g04650(.I(new_n4842_), .ZN(new_n4843_));
  NAND3_X1   g04651(.A1(\asqrt[34] ), .A2(new_n4665_), .A3(new_n4684_), .ZN(new_n4844_));
  XOR2_X1    g04652(.A1(new_n4844_), .A2(new_n4699_), .Z(new_n4845_));
  INV_X1     g04653(.I(new_n4845_), .ZN(new_n4846_));
  OAI21_X1   g04654(.A1(new_n4659_), .A2(new_n4661_), .B(new_n4664_), .ZN(new_n4847_));
  NOR2_X1    g04655(.A1(new_n4810_), .A2(new_n4847_), .ZN(new_n4848_));
  XOR2_X1    g04656(.A1(new_n4848_), .A2(new_n4551_), .Z(new_n4849_));
  NAND3_X1   g04657(.A1(\asqrt[34] ), .A2(new_n4678_), .A3(new_n4660_), .ZN(new_n4850_));
  XOR2_X1    g04658(.A1(new_n4850_), .A2(new_n4555_), .Z(new_n4851_));
  OAI21_X1   g04659(.A1(new_n4673_), .A2(new_n4674_), .B(new_n4677_), .ZN(new_n4852_));
  NOR2_X1    g04660(.A1(new_n4810_), .A2(new_n4852_), .ZN(new_n4853_));
  XOR2_X1    g04661(.A1(new_n4853_), .A2(new_n4557_), .Z(new_n4854_));
  INV_X1     g04662(.I(new_n4854_), .ZN(new_n4855_));
  NAND3_X1   g04663(.A1(\asqrt[34] ), .A2(new_n4637_), .A3(new_n4656_), .ZN(new_n4856_));
  XOR2_X1    g04664(.A1(new_n4856_), .A2(new_n4671_), .Z(new_n4857_));
  INV_X1     g04665(.I(new_n4857_), .ZN(new_n4858_));
  OAI21_X1   g04666(.A1(new_n4631_), .A2(new_n4633_), .B(new_n4636_), .ZN(new_n4859_));
  NOR2_X1    g04667(.A1(new_n4810_), .A2(new_n4859_), .ZN(new_n4860_));
  XOR2_X1    g04668(.A1(new_n4860_), .A2(new_n4563_), .Z(new_n4861_));
  NAND3_X1   g04669(.A1(\asqrt[34] ), .A2(new_n4650_), .A3(new_n4632_), .ZN(new_n4862_));
  XOR2_X1    g04670(.A1(new_n4862_), .A2(new_n4567_), .Z(new_n4863_));
  OAI21_X1   g04671(.A1(new_n4645_), .A2(new_n4646_), .B(new_n4649_), .ZN(new_n4864_));
  NOR2_X1    g04672(.A1(new_n4810_), .A2(new_n4864_), .ZN(new_n4865_));
  XOR2_X1    g04673(.A1(new_n4865_), .A2(new_n4570_), .Z(new_n4866_));
  INV_X1     g04674(.I(new_n4866_), .ZN(new_n4867_));
  NAND3_X1   g04675(.A1(\asqrt[34] ), .A2(new_n4605_), .A3(new_n4628_), .ZN(new_n4868_));
  XOR2_X1    g04676(.A1(new_n4868_), .A2(new_n4643_), .Z(new_n4869_));
  INV_X1     g04677(.I(new_n4869_), .ZN(new_n4870_));
  OAI21_X1   g04678(.A1(new_n4599_), .A2(new_n4601_), .B(new_n4604_), .ZN(new_n4871_));
  NOR2_X1    g04679(.A1(new_n4810_), .A2(new_n4871_), .ZN(new_n4872_));
  XOR2_X1    g04680(.A1(new_n4872_), .A2(new_n4576_), .Z(new_n4873_));
  NAND3_X1   g04681(.A1(\asqrt[34] ), .A2(new_n4622_), .A3(new_n4600_), .ZN(new_n4874_));
  XOR2_X1    g04682(.A1(new_n4874_), .A2(new_n4598_), .Z(new_n4875_));
  NOR2_X1    g04683(.A1(new_n4619_), .A2(\asqrt[37] ), .ZN(new_n4876_));
  NOR3_X1    g04684(.A1(new_n4810_), .A2(new_n4876_), .A3(new_n4594_), .ZN(new_n4877_));
  XOR2_X1    g04685(.A1(new_n4877_), .A2(new_n4613_), .Z(new_n4878_));
  INV_X1     g04686(.I(new_n4878_), .ZN(new_n4879_));
  NAND3_X1   g04687(.A1(\asqrt[34] ), .A2(new_n4584_), .A3(new_n4585_), .ZN(new_n4880_));
  NOR4_X1    g04688(.A1(new_n4807_), .A2(new_n4510_), .A3(new_n4785_), .A4(new_n4809_), .ZN(new_n4881_));
  INV_X1     g04689(.I(new_n4881_), .ZN(new_n4882_));
  AOI21_X1   g04690(.A1(new_n4880_), .A2(new_n4882_), .B(\a[70] ), .ZN(new_n4883_));
  NOR3_X1    g04691(.A1(new_n4810_), .A2(\a[68] ), .A3(\a[69] ), .ZN(new_n4884_));
  NOR3_X1    g04692(.A1(new_n4884_), .A2(new_n4302_), .A3(new_n4881_), .ZN(new_n4885_));
  NOR2_X1    g04693(.A1(new_n4885_), .A2(new_n4883_), .ZN(new_n4886_));
  INV_X1     g04694(.I(\a[66] ), .ZN(new_n4887_));
  INV_X1     g04695(.I(\a[67] ), .ZN(new_n4888_));
  NAND3_X1   g04696(.A1(new_n4887_), .A2(new_n4888_), .A3(new_n4584_), .ZN(new_n4889_));
  OAI21_X1   g04697(.A1(new_n4810_), .A2(new_n4584_), .B(new_n4889_), .ZN(new_n4890_));
  NAND2_X1   g04698(.A1(new_n4890_), .A2(\asqrt[35] ), .ZN(new_n4891_));
  OAI21_X1   g04699(.A1(new_n4810_), .A2(\a[68] ), .B(\a[69] ), .ZN(new_n4892_));
  NAND2_X1   g04700(.A1(new_n4892_), .A2(new_n4880_), .ZN(new_n4893_));
  NOR2_X1    g04701(.A1(new_n4890_), .A2(\asqrt[35] ), .ZN(new_n4894_));
  OAI21_X1   g04702(.A1(new_n4893_), .A2(new_n4894_), .B(new_n4891_), .ZN(new_n4895_));
  OAI21_X1   g04703(.A1(new_n4895_), .A2(\asqrt[36] ), .B(new_n4886_), .ZN(new_n4896_));
  NAND2_X1   g04704(.A1(new_n4895_), .A2(\asqrt[36] ), .ZN(new_n4897_));
  NAND3_X1   g04705(.A1(new_n4896_), .A2(new_n3928_), .A3(new_n4897_), .ZN(new_n4898_));
  NOR3_X1    g04706(.A1(new_n4810_), .A2(new_n4588_), .A3(new_n4618_), .ZN(new_n4899_));
  XOR2_X1    g04707(.A1(new_n4899_), .A2(new_n4590_), .Z(new_n4900_));
  AOI21_X1   g04708(.A1(new_n4896_), .A2(new_n4897_), .B(new_n3928_), .ZN(new_n4901_));
  AOI21_X1   g04709(.A1(new_n4898_), .A2(new_n4900_), .B(new_n4901_), .ZN(new_n4902_));
  AOI21_X1   g04710(.A1(new_n4902_), .A2(new_n3675_), .B(new_n4879_), .ZN(new_n4903_));
  OAI21_X1   g04711(.A1(new_n4902_), .A2(new_n3675_), .B(new_n3400_), .ZN(new_n4904_));
  OAI21_X1   g04712(.A1(new_n4903_), .A2(new_n4904_), .B(new_n4875_), .ZN(new_n4905_));
  NOR2_X1    g04713(.A1(new_n4902_), .A2(new_n3675_), .ZN(new_n4906_));
  OAI21_X1   g04714(.A1(new_n4903_), .A2(new_n4906_), .B(\asqrt[39] ), .ZN(new_n4907_));
  NAND3_X1   g04715(.A1(new_n4905_), .A2(new_n4907_), .A3(new_n3167_), .ZN(new_n4908_));
  NAND2_X1   g04716(.A1(new_n4908_), .A2(new_n4873_), .ZN(new_n4909_));
  NAND2_X1   g04717(.A1(new_n4905_), .A2(new_n4907_), .ZN(new_n4910_));
  AOI21_X1   g04718(.A1(new_n4910_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n4911_));
  AOI21_X1   g04719(.A1(new_n4911_), .A2(new_n4909_), .B(new_n4870_), .ZN(new_n4912_));
  INV_X1     g04720(.I(new_n4875_), .ZN(new_n4913_));
  OAI21_X1   g04721(.A1(new_n4884_), .A2(new_n4881_), .B(new_n4302_), .ZN(new_n4914_));
  NAND3_X1   g04722(.A1(new_n4880_), .A2(new_n4882_), .A3(\a[70] ), .ZN(new_n4915_));
  NAND2_X1   g04723(.A1(new_n4914_), .A2(new_n4915_), .ZN(new_n4916_));
  NAND2_X1   g04724(.A1(\asqrt[34] ), .A2(\a[68] ), .ZN(new_n4917_));
  AOI21_X1   g04725(.A1(new_n4917_), .A2(new_n4889_), .B(new_n4510_), .ZN(new_n4918_));
  AOI21_X1   g04726(.A1(\asqrt[34] ), .A2(new_n4584_), .B(new_n4585_), .ZN(new_n4919_));
  NOR2_X1    g04727(.A1(new_n4884_), .A2(new_n4919_), .ZN(new_n4920_));
  NAND3_X1   g04728(.A1(new_n4917_), .A2(new_n4510_), .A3(new_n4889_), .ZN(new_n4921_));
  AOI21_X1   g04729(.A1(new_n4920_), .A2(new_n4921_), .B(new_n4918_), .ZN(new_n4922_));
  AOI21_X1   g04730(.A1(new_n4922_), .A2(new_n4224_), .B(new_n4916_), .ZN(new_n4923_));
  NOR2_X1    g04731(.A1(new_n4922_), .A2(new_n4224_), .ZN(new_n4924_));
  NOR3_X1    g04732(.A1(new_n4923_), .A2(\asqrt[37] ), .A3(new_n4924_), .ZN(new_n4925_));
  INV_X1     g04733(.I(new_n4900_), .ZN(new_n4926_));
  OAI21_X1   g04734(.A1(new_n4923_), .A2(new_n4924_), .B(\asqrt[37] ), .ZN(new_n4927_));
  OAI21_X1   g04735(.A1(new_n4925_), .A2(new_n4926_), .B(new_n4927_), .ZN(new_n4928_));
  OAI21_X1   g04736(.A1(new_n4928_), .A2(\asqrt[38] ), .B(new_n4878_), .ZN(new_n4929_));
  AOI21_X1   g04737(.A1(new_n4928_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n4930_));
  AOI21_X1   g04738(.A1(new_n4930_), .A2(new_n4929_), .B(new_n4913_), .ZN(new_n4931_));
  NAND2_X1   g04739(.A1(new_n4928_), .A2(\asqrt[38] ), .ZN(new_n4932_));
  AOI21_X1   g04740(.A1(new_n4929_), .A2(new_n4932_), .B(new_n3400_), .ZN(new_n4933_));
  OAI21_X1   g04741(.A1(new_n4931_), .A2(new_n4933_), .B(\asqrt[40] ), .ZN(new_n4934_));
  AOI21_X1   g04742(.A1(new_n4909_), .A2(new_n4934_), .B(new_n2912_), .ZN(new_n4935_));
  NOR2_X1    g04743(.A1(new_n4912_), .A2(new_n4935_), .ZN(new_n4936_));
  AOI21_X1   g04744(.A1(new_n4936_), .A2(new_n2699_), .B(new_n4867_), .ZN(new_n4937_));
  OAI21_X1   g04745(.A1(new_n4912_), .A2(new_n4935_), .B(\asqrt[42] ), .ZN(new_n4938_));
  NAND2_X1   g04746(.A1(new_n4938_), .A2(new_n2464_), .ZN(new_n4939_));
  OAI21_X1   g04747(.A1(new_n4937_), .A2(new_n4939_), .B(new_n4863_), .ZN(new_n4940_));
  INV_X1     g04748(.I(new_n4938_), .ZN(new_n4941_));
  OAI21_X1   g04749(.A1(new_n4937_), .A2(new_n4941_), .B(\asqrt[43] ), .ZN(new_n4942_));
  NAND3_X1   g04750(.A1(new_n4940_), .A2(new_n4942_), .A3(new_n2271_), .ZN(new_n4943_));
  NAND2_X1   g04751(.A1(new_n4943_), .A2(new_n4861_), .ZN(new_n4944_));
  NAND2_X1   g04752(.A1(new_n4940_), .A2(new_n4942_), .ZN(new_n4945_));
  AOI21_X1   g04753(.A1(new_n4945_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n4946_));
  AOI21_X1   g04754(.A1(new_n4946_), .A2(new_n4944_), .B(new_n4858_), .ZN(new_n4947_));
  INV_X1     g04755(.I(new_n4863_), .ZN(new_n4948_));
  INV_X1     g04756(.I(new_n4873_), .ZN(new_n4949_));
  NOR2_X1    g04757(.A1(new_n4931_), .A2(new_n4933_), .ZN(new_n4950_));
  AOI21_X1   g04758(.A1(new_n4950_), .A2(new_n3167_), .B(new_n4949_), .ZN(new_n4951_));
  NAND2_X1   g04759(.A1(new_n4934_), .A2(new_n2912_), .ZN(new_n4952_));
  OAI21_X1   g04760(.A1(new_n4951_), .A2(new_n4952_), .B(new_n4869_), .ZN(new_n4953_));
  INV_X1     g04761(.I(new_n4934_), .ZN(new_n4954_));
  OAI21_X1   g04762(.A1(new_n4951_), .A2(new_n4954_), .B(\asqrt[41] ), .ZN(new_n4955_));
  NAND3_X1   g04763(.A1(new_n4953_), .A2(new_n4955_), .A3(new_n2699_), .ZN(new_n4956_));
  NAND2_X1   g04764(.A1(new_n4956_), .A2(new_n4866_), .ZN(new_n4957_));
  NAND2_X1   g04765(.A1(new_n4953_), .A2(new_n4955_), .ZN(new_n4958_));
  AOI21_X1   g04766(.A1(new_n4958_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n4959_));
  AOI21_X1   g04767(.A1(new_n4959_), .A2(new_n4957_), .B(new_n4948_), .ZN(new_n4960_));
  AOI21_X1   g04768(.A1(new_n4957_), .A2(new_n4938_), .B(new_n2464_), .ZN(new_n4961_));
  OAI21_X1   g04769(.A1(new_n4960_), .A2(new_n4961_), .B(\asqrt[44] ), .ZN(new_n4962_));
  AOI21_X1   g04770(.A1(new_n4944_), .A2(new_n4962_), .B(new_n2072_), .ZN(new_n4963_));
  NOR2_X1    g04771(.A1(new_n4947_), .A2(new_n4963_), .ZN(new_n4964_));
  AOI21_X1   g04772(.A1(new_n4964_), .A2(new_n1884_), .B(new_n4855_), .ZN(new_n4965_));
  OAI21_X1   g04773(.A1(new_n4947_), .A2(new_n4963_), .B(\asqrt[46] ), .ZN(new_n4966_));
  NAND2_X1   g04774(.A1(new_n4966_), .A2(new_n1688_), .ZN(new_n4967_));
  OAI21_X1   g04775(.A1(new_n4965_), .A2(new_n4967_), .B(new_n4851_), .ZN(new_n4968_));
  INV_X1     g04776(.I(new_n4966_), .ZN(new_n4969_));
  OAI21_X1   g04777(.A1(new_n4965_), .A2(new_n4969_), .B(\asqrt[47] ), .ZN(new_n4970_));
  NAND3_X1   g04778(.A1(new_n4968_), .A2(new_n4970_), .A3(new_n1533_), .ZN(new_n4971_));
  NAND2_X1   g04779(.A1(new_n4971_), .A2(new_n4849_), .ZN(new_n4972_));
  NAND2_X1   g04780(.A1(new_n4968_), .A2(new_n4970_), .ZN(new_n4973_));
  AOI21_X1   g04781(.A1(new_n4973_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n4974_));
  AOI21_X1   g04782(.A1(new_n4974_), .A2(new_n4972_), .B(new_n4846_), .ZN(new_n4975_));
  INV_X1     g04783(.I(new_n4851_), .ZN(new_n4976_));
  INV_X1     g04784(.I(new_n4861_), .ZN(new_n4977_));
  NOR2_X1    g04785(.A1(new_n4960_), .A2(new_n4961_), .ZN(new_n4978_));
  AOI21_X1   g04786(.A1(new_n4978_), .A2(new_n2271_), .B(new_n4977_), .ZN(new_n4979_));
  NAND2_X1   g04787(.A1(new_n4962_), .A2(new_n2072_), .ZN(new_n4980_));
  OAI21_X1   g04788(.A1(new_n4979_), .A2(new_n4980_), .B(new_n4857_), .ZN(new_n4981_));
  INV_X1     g04789(.I(new_n4962_), .ZN(new_n4982_));
  OAI21_X1   g04790(.A1(new_n4979_), .A2(new_n4982_), .B(\asqrt[45] ), .ZN(new_n4983_));
  NAND3_X1   g04791(.A1(new_n4981_), .A2(new_n4983_), .A3(new_n1884_), .ZN(new_n4984_));
  NAND2_X1   g04792(.A1(new_n4984_), .A2(new_n4854_), .ZN(new_n4985_));
  NAND2_X1   g04793(.A1(new_n4981_), .A2(new_n4983_), .ZN(new_n4986_));
  AOI21_X1   g04794(.A1(new_n4986_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n4987_));
  AOI21_X1   g04795(.A1(new_n4987_), .A2(new_n4985_), .B(new_n4976_), .ZN(new_n4988_));
  AOI21_X1   g04796(.A1(new_n4985_), .A2(new_n4966_), .B(new_n1688_), .ZN(new_n4989_));
  OAI21_X1   g04797(.A1(new_n4988_), .A2(new_n4989_), .B(\asqrt[48] ), .ZN(new_n4990_));
  AOI21_X1   g04798(.A1(new_n4972_), .A2(new_n4990_), .B(new_n1368_), .ZN(new_n4991_));
  NOR2_X1    g04799(.A1(new_n4975_), .A2(new_n4991_), .ZN(new_n4992_));
  AOI21_X1   g04800(.A1(new_n4992_), .A2(new_n1228_), .B(new_n4843_), .ZN(new_n4993_));
  OAI21_X1   g04801(.A1(new_n4975_), .A2(new_n4991_), .B(\asqrt[50] ), .ZN(new_n4994_));
  NAND2_X1   g04802(.A1(new_n4994_), .A2(new_n1088_), .ZN(new_n4995_));
  OAI21_X1   g04803(.A1(new_n4993_), .A2(new_n4995_), .B(new_n4839_), .ZN(new_n4996_));
  INV_X1     g04804(.I(new_n4994_), .ZN(new_n4997_));
  OAI21_X1   g04805(.A1(new_n4993_), .A2(new_n4997_), .B(\asqrt[51] ), .ZN(new_n4998_));
  NAND3_X1   g04806(.A1(new_n4996_), .A2(new_n4998_), .A3(new_n962_), .ZN(new_n4999_));
  NAND2_X1   g04807(.A1(new_n4999_), .A2(new_n4837_), .ZN(new_n5000_));
  NAND2_X1   g04808(.A1(new_n4996_), .A2(new_n4998_), .ZN(new_n5001_));
  AOI21_X1   g04809(.A1(new_n5001_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n5002_));
  AOI21_X1   g04810(.A1(new_n5002_), .A2(new_n5000_), .B(new_n4834_), .ZN(new_n5003_));
  INV_X1     g04811(.I(new_n4839_), .ZN(new_n5004_));
  INV_X1     g04812(.I(new_n4849_), .ZN(new_n5005_));
  NOR2_X1    g04813(.A1(new_n4988_), .A2(new_n4989_), .ZN(new_n5006_));
  AOI21_X1   g04814(.A1(new_n5006_), .A2(new_n1533_), .B(new_n5005_), .ZN(new_n5007_));
  NAND2_X1   g04815(.A1(new_n4990_), .A2(new_n1368_), .ZN(new_n5008_));
  OAI21_X1   g04816(.A1(new_n5007_), .A2(new_n5008_), .B(new_n4845_), .ZN(new_n5009_));
  INV_X1     g04817(.I(new_n4990_), .ZN(new_n5010_));
  OAI21_X1   g04818(.A1(new_n5007_), .A2(new_n5010_), .B(\asqrt[49] ), .ZN(new_n5011_));
  NAND3_X1   g04819(.A1(new_n5009_), .A2(new_n5011_), .A3(new_n1228_), .ZN(new_n5012_));
  NAND2_X1   g04820(.A1(new_n5012_), .A2(new_n4842_), .ZN(new_n5013_));
  NAND2_X1   g04821(.A1(new_n5009_), .A2(new_n5011_), .ZN(new_n5014_));
  AOI21_X1   g04822(.A1(new_n5014_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n5015_));
  AOI21_X1   g04823(.A1(new_n5015_), .A2(new_n5013_), .B(new_n5004_), .ZN(new_n5016_));
  AOI21_X1   g04824(.A1(new_n5013_), .A2(new_n4994_), .B(new_n1088_), .ZN(new_n5017_));
  OAI21_X1   g04825(.A1(new_n5016_), .A2(new_n5017_), .B(\asqrt[52] ), .ZN(new_n5018_));
  AOI21_X1   g04826(.A1(new_n5000_), .A2(new_n5018_), .B(new_n842_), .ZN(new_n5019_));
  NOR2_X1    g04827(.A1(new_n5003_), .A2(new_n5019_), .ZN(new_n5020_));
  AOI21_X1   g04828(.A1(new_n5020_), .A2(new_n720_), .B(new_n4831_), .ZN(new_n5021_));
  OAI21_X1   g04829(.A1(new_n5003_), .A2(new_n5019_), .B(\asqrt[54] ), .ZN(new_n5022_));
  NAND2_X1   g04830(.A1(new_n5022_), .A2(new_n630_), .ZN(new_n5023_));
  OAI21_X1   g04831(.A1(new_n5021_), .A2(new_n5023_), .B(new_n4827_), .ZN(new_n5024_));
  INV_X1     g04832(.I(new_n5022_), .ZN(new_n5025_));
  OAI21_X1   g04833(.A1(new_n5021_), .A2(new_n5025_), .B(\asqrt[55] ), .ZN(new_n5026_));
  NAND3_X1   g04834(.A1(new_n5024_), .A2(new_n5026_), .A3(new_n545_), .ZN(new_n5027_));
  NAND2_X1   g04835(.A1(new_n5027_), .A2(new_n4825_), .ZN(new_n5028_));
  NAND2_X1   g04836(.A1(new_n5024_), .A2(new_n5026_), .ZN(new_n5029_));
  AOI21_X1   g04837(.A1(new_n5029_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n5030_));
  AOI21_X1   g04838(.A1(new_n5030_), .A2(new_n5028_), .B(new_n4822_), .ZN(new_n5031_));
  INV_X1     g04839(.I(new_n4827_), .ZN(new_n5032_));
  INV_X1     g04840(.I(new_n4837_), .ZN(new_n5033_));
  NOR2_X1    g04841(.A1(new_n5016_), .A2(new_n5017_), .ZN(new_n5034_));
  AOI21_X1   g04842(.A1(new_n5034_), .A2(new_n962_), .B(new_n5033_), .ZN(new_n5035_));
  NAND2_X1   g04843(.A1(new_n5018_), .A2(new_n842_), .ZN(new_n5036_));
  OAI21_X1   g04844(.A1(new_n5035_), .A2(new_n5036_), .B(new_n4833_), .ZN(new_n5037_));
  INV_X1     g04845(.I(new_n5018_), .ZN(new_n5038_));
  OAI21_X1   g04846(.A1(new_n5035_), .A2(new_n5038_), .B(\asqrt[53] ), .ZN(new_n5039_));
  NAND3_X1   g04847(.A1(new_n5037_), .A2(new_n5039_), .A3(new_n720_), .ZN(new_n5040_));
  NAND2_X1   g04848(.A1(new_n5040_), .A2(new_n4830_), .ZN(new_n5041_));
  NAND2_X1   g04849(.A1(new_n5037_), .A2(new_n5039_), .ZN(new_n5042_));
  AOI21_X1   g04850(.A1(new_n5042_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n5043_));
  AOI21_X1   g04851(.A1(new_n5043_), .A2(new_n5041_), .B(new_n5032_), .ZN(new_n5044_));
  AOI21_X1   g04852(.A1(new_n5041_), .A2(new_n5022_), .B(new_n630_), .ZN(new_n5045_));
  OAI21_X1   g04853(.A1(new_n5044_), .A2(new_n5045_), .B(\asqrt[56] ), .ZN(new_n5046_));
  AOI21_X1   g04854(.A1(new_n5028_), .A2(new_n5046_), .B(new_n450_), .ZN(new_n5047_));
  NOR2_X1    g04855(.A1(new_n5031_), .A2(new_n5047_), .ZN(new_n5048_));
  AOI21_X1   g04856(.A1(new_n5048_), .A2(new_n403_), .B(new_n4819_), .ZN(new_n5049_));
  OAI21_X1   g04857(.A1(new_n5031_), .A2(new_n5047_), .B(\asqrt[58] ), .ZN(new_n5050_));
  NAND2_X1   g04858(.A1(new_n5050_), .A2(new_n339_), .ZN(new_n5051_));
  OAI21_X1   g04859(.A1(new_n5049_), .A2(new_n5051_), .B(new_n4815_), .ZN(new_n5052_));
  INV_X1     g04860(.I(new_n5050_), .ZN(new_n5053_));
  OAI21_X1   g04861(.A1(new_n5049_), .A2(new_n5053_), .B(\asqrt[59] ), .ZN(new_n5054_));
  NAND3_X1   g04862(.A1(new_n5052_), .A2(new_n5054_), .A3(new_n288_), .ZN(new_n5055_));
  NAND2_X1   g04863(.A1(new_n5055_), .A2(new_n4813_), .ZN(new_n5056_));
  INV_X1     g04864(.I(new_n4815_), .ZN(new_n5057_));
  INV_X1     g04865(.I(new_n4825_), .ZN(new_n5058_));
  NOR2_X1    g04866(.A1(new_n5044_), .A2(new_n5045_), .ZN(new_n5059_));
  AOI21_X1   g04867(.A1(new_n5059_), .A2(new_n545_), .B(new_n5058_), .ZN(new_n5060_));
  NAND2_X1   g04868(.A1(new_n5046_), .A2(new_n450_), .ZN(new_n5061_));
  OAI21_X1   g04869(.A1(new_n5060_), .A2(new_n5061_), .B(new_n4821_), .ZN(new_n5062_));
  INV_X1     g04870(.I(new_n5046_), .ZN(new_n5063_));
  OAI21_X1   g04871(.A1(new_n5060_), .A2(new_n5063_), .B(\asqrt[57] ), .ZN(new_n5064_));
  NAND3_X1   g04872(.A1(new_n5062_), .A2(new_n5064_), .A3(new_n403_), .ZN(new_n5065_));
  NAND2_X1   g04873(.A1(new_n5065_), .A2(new_n4818_), .ZN(new_n5066_));
  NAND2_X1   g04874(.A1(new_n5062_), .A2(new_n5064_), .ZN(new_n5067_));
  AOI21_X1   g04875(.A1(new_n5067_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n5068_));
  AOI21_X1   g04876(.A1(new_n5068_), .A2(new_n5066_), .B(new_n5057_), .ZN(new_n5069_));
  AOI21_X1   g04877(.A1(new_n5066_), .A2(new_n5050_), .B(new_n339_), .ZN(new_n5070_));
  OAI21_X1   g04878(.A1(new_n5069_), .A2(new_n5070_), .B(\asqrt[60] ), .ZN(new_n5071_));
  AOI21_X1   g04879(.A1(new_n5056_), .A2(new_n5071_), .B(new_n242_), .ZN(new_n5072_));
  NAND3_X1   g04880(.A1(\asqrt[34] ), .A2(new_n4749_), .A3(new_n4765_), .ZN(new_n5073_));
  XOR2_X1    g04881(.A1(new_n5073_), .A2(new_n4774_), .Z(new_n5074_));
  INV_X1     g04882(.I(new_n5074_), .ZN(new_n5075_));
  NAND2_X1   g04883(.A1(new_n5052_), .A2(new_n5054_), .ZN(new_n5076_));
  AOI21_X1   g04884(.A1(new_n5076_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n5077_));
  AOI21_X1   g04885(.A1(new_n5077_), .A2(new_n5056_), .B(new_n5075_), .ZN(new_n5078_));
  OAI21_X1   g04886(.A1(new_n5078_), .A2(new_n5072_), .B(\asqrt[62] ), .ZN(new_n5079_));
  AOI21_X1   g04887(.A1(new_n4750_), .A2(new_n4771_), .B(new_n4766_), .ZN(new_n5080_));
  NAND2_X1   g04888(.A1(\asqrt[34] ), .A2(new_n5080_), .ZN(new_n5081_));
  XOR2_X1    g04889(.A1(new_n5081_), .A2(new_n4769_), .Z(new_n5082_));
  INV_X1     g04890(.I(new_n4813_), .ZN(new_n5083_));
  NOR2_X1    g04891(.A1(new_n5069_), .A2(new_n5070_), .ZN(new_n5084_));
  AOI21_X1   g04892(.A1(new_n5084_), .A2(new_n288_), .B(new_n5083_), .ZN(new_n5085_));
  INV_X1     g04893(.I(new_n5071_), .ZN(new_n5086_));
  OAI21_X1   g04894(.A1(new_n5085_), .A2(new_n5086_), .B(\asqrt[61] ), .ZN(new_n5087_));
  NAND2_X1   g04895(.A1(new_n5071_), .A2(new_n242_), .ZN(new_n5088_));
  OAI21_X1   g04896(.A1(new_n5085_), .A2(new_n5088_), .B(new_n5074_), .ZN(new_n5089_));
  NAND3_X1   g04897(.A1(new_n5089_), .A2(new_n5087_), .A3(new_n234_), .ZN(new_n5090_));
  NAND2_X1   g04898(.A1(new_n5090_), .A2(new_n5082_), .ZN(new_n5091_));
  NAND2_X1   g04899(.A1(new_n5091_), .A2(new_n5079_), .ZN(new_n5092_));
  NAND2_X1   g04900(.A1(new_n5092_), .A2(new_n4802_), .ZN(new_n5093_));
  INV_X1     g04901(.I(new_n5079_), .ZN(new_n5094_));
  NOR2_X1    g04902(.A1(new_n5078_), .A2(new_n5072_), .ZN(new_n5095_));
  INV_X1     g04903(.I(new_n5082_), .ZN(new_n5096_));
  AOI21_X1   g04904(.A1(new_n5095_), .A2(new_n234_), .B(new_n5096_), .ZN(new_n5097_));
  NOR2_X1    g04905(.A1(new_n5097_), .A2(new_n5094_), .ZN(new_n5098_));
  NAND2_X1   g04906(.A1(new_n4808_), .A2(new_n4788_), .ZN(new_n5099_));
  NOR2_X1    g04907(.A1(new_n4810_), .A2(new_n4788_), .ZN(new_n5100_));
  NAND2_X1   g04908(.A1(new_n5100_), .A2(new_n4796_), .ZN(new_n5101_));
  AOI21_X1   g04909(.A1(new_n5101_), .A2(new_n5099_), .B(new_n193_), .ZN(new_n5102_));
  INV_X1     g04910(.I(new_n4802_), .ZN(new_n5103_));
  AOI21_X1   g04911(.A1(new_n5100_), .A2(new_n4808_), .B(new_n4809_), .ZN(new_n5104_));
  INV_X1     g04912(.I(new_n5104_), .ZN(new_n5105_));
  AOI21_X1   g04913(.A1(new_n5091_), .A2(new_n5079_), .B(new_n5105_), .ZN(new_n5106_));
  AOI21_X1   g04914(.A1(new_n5106_), .A2(new_n5103_), .B(\asqrt[63] ), .ZN(new_n5107_));
  NOR2_X1    g04915(.A1(new_n5092_), .A2(new_n5103_), .ZN(new_n5108_));
  NOR2_X1    g04916(.A1(\asqrt[34] ), .A2(new_n4803_), .ZN(new_n5109_));
  NOR4_X1    g04917(.A1(new_n5107_), .A2(new_n5102_), .A3(new_n5108_), .A4(new_n5109_), .ZN(new_n5110_));
  NOR2_X1    g04918(.A1(new_n5110_), .A2(new_n4802_), .ZN(new_n5111_));
  NAND2_X1   g04919(.A1(new_n5111_), .A2(new_n5098_), .ZN(new_n5112_));
  AOI21_X1   g04920(.A1(new_n5112_), .A2(new_n5093_), .B(new_n193_), .ZN(new_n5113_));
  INV_X1     g04921(.I(new_n5113_), .ZN(new_n5114_));
  INV_X1     g04922(.I(new_n5102_), .ZN(new_n5115_));
  OAI21_X1   g04923(.A1(new_n5097_), .A2(new_n5094_), .B(new_n5104_), .ZN(new_n5116_));
  OAI21_X1   g04924(.A1(new_n5116_), .A2(new_n4802_), .B(new_n193_), .ZN(new_n5117_));
  NAND2_X1   g04925(.A1(new_n5098_), .A2(new_n4802_), .ZN(new_n5118_));
  INV_X1     g04926(.I(new_n5109_), .ZN(new_n5119_));
  NAND4_X1   g04927(.A1(new_n5117_), .A2(new_n5115_), .A3(new_n5118_), .A4(new_n5119_), .ZN(\asqrt[33] ));
  NAND3_X1   g04928(.A1(\asqrt[33] ), .A2(new_n5079_), .A3(new_n5090_), .ZN(new_n5121_));
  XOR2_X1    g04929(.A1(new_n5121_), .A2(new_n5082_), .Z(new_n5122_));
  AOI21_X1   g04930(.A1(new_n5111_), .A2(new_n5092_), .B(new_n5108_), .ZN(new_n5123_));
  OAI21_X1   g04931(.A1(new_n5049_), .A2(new_n5051_), .B(new_n5054_), .ZN(new_n5124_));
  NOR2_X1    g04932(.A1(new_n5110_), .A2(new_n5124_), .ZN(new_n5125_));
  XOR2_X1    g04933(.A1(new_n5125_), .A2(new_n4815_), .Z(new_n5126_));
  NAND3_X1   g04934(.A1(\asqrt[33] ), .A2(new_n5065_), .A3(new_n5050_), .ZN(new_n5127_));
  XOR2_X1    g04935(.A1(new_n5127_), .A2(new_n4819_), .Z(new_n5128_));
  OAI21_X1   g04936(.A1(new_n5060_), .A2(new_n5061_), .B(new_n5064_), .ZN(new_n5129_));
  NOR2_X1    g04937(.A1(new_n5110_), .A2(new_n5129_), .ZN(new_n5130_));
  XOR2_X1    g04938(.A1(new_n5130_), .A2(new_n4821_), .Z(new_n5131_));
  INV_X1     g04939(.I(new_n5131_), .ZN(new_n5132_));
  NAND3_X1   g04940(.A1(\asqrt[33] ), .A2(new_n5027_), .A3(new_n5046_), .ZN(new_n5133_));
  XOR2_X1    g04941(.A1(new_n5133_), .A2(new_n5058_), .Z(new_n5134_));
  INV_X1     g04942(.I(new_n5134_), .ZN(new_n5135_));
  OAI21_X1   g04943(.A1(new_n5021_), .A2(new_n5023_), .B(new_n5026_), .ZN(new_n5136_));
  NOR2_X1    g04944(.A1(new_n5110_), .A2(new_n5136_), .ZN(new_n5137_));
  XOR2_X1    g04945(.A1(new_n5137_), .A2(new_n4827_), .Z(new_n5138_));
  NAND3_X1   g04946(.A1(\asqrt[33] ), .A2(new_n5040_), .A3(new_n5022_), .ZN(new_n5139_));
  XOR2_X1    g04947(.A1(new_n5139_), .A2(new_n4831_), .Z(new_n5140_));
  OAI21_X1   g04948(.A1(new_n5035_), .A2(new_n5036_), .B(new_n5039_), .ZN(new_n5141_));
  NOR2_X1    g04949(.A1(new_n5110_), .A2(new_n5141_), .ZN(new_n5142_));
  XOR2_X1    g04950(.A1(new_n5142_), .A2(new_n4833_), .Z(new_n5143_));
  INV_X1     g04951(.I(new_n5143_), .ZN(new_n5144_));
  NAND3_X1   g04952(.A1(\asqrt[33] ), .A2(new_n4999_), .A3(new_n5018_), .ZN(new_n5145_));
  XOR2_X1    g04953(.A1(new_n5145_), .A2(new_n5033_), .Z(new_n5146_));
  INV_X1     g04954(.I(new_n5146_), .ZN(new_n5147_));
  OAI21_X1   g04955(.A1(new_n4993_), .A2(new_n4995_), .B(new_n4998_), .ZN(new_n5148_));
  NOR2_X1    g04956(.A1(new_n5110_), .A2(new_n5148_), .ZN(new_n5149_));
  XOR2_X1    g04957(.A1(new_n5149_), .A2(new_n4839_), .Z(new_n5150_));
  NAND3_X1   g04958(.A1(\asqrt[33] ), .A2(new_n5012_), .A3(new_n4994_), .ZN(new_n5151_));
  XOR2_X1    g04959(.A1(new_n5151_), .A2(new_n4843_), .Z(new_n5152_));
  OAI21_X1   g04960(.A1(new_n5007_), .A2(new_n5008_), .B(new_n5011_), .ZN(new_n5153_));
  NOR2_X1    g04961(.A1(new_n5110_), .A2(new_n5153_), .ZN(new_n5154_));
  XOR2_X1    g04962(.A1(new_n5154_), .A2(new_n4845_), .Z(new_n5155_));
  INV_X1     g04963(.I(new_n5155_), .ZN(new_n5156_));
  NAND3_X1   g04964(.A1(\asqrt[33] ), .A2(new_n4971_), .A3(new_n4990_), .ZN(new_n5157_));
  XOR2_X1    g04965(.A1(new_n5157_), .A2(new_n5005_), .Z(new_n5158_));
  INV_X1     g04966(.I(new_n5158_), .ZN(new_n5159_));
  OAI21_X1   g04967(.A1(new_n4965_), .A2(new_n4967_), .B(new_n4970_), .ZN(new_n5160_));
  NOR2_X1    g04968(.A1(new_n5110_), .A2(new_n5160_), .ZN(new_n5161_));
  XOR2_X1    g04969(.A1(new_n5161_), .A2(new_n4851_), .Z(new_n5162_));
  NAND3_X1   g04970(.A1(\asqrt[33] ), .A2(new_n4984_), .A3(new_n4966_), .ZN(new_n5163_));
  XOR2_X1    g04971(.A1(new_n5163_), .A2(new_n4855_), .Z(new_n5164_));
  OAI21_X1   g04972(.A1(new_n4979_), .A2(new_n4980_), .B(new_n4983_), .ZN(new_n5165_));
  NOR2_X1    g04973(.A1(new_n5110_), .A2(new_n5165_), .ZN(new_n5166_));
  XOR2_X1    g04974(.A1(new_n5166_), .A2(new_n4857_), .Z(new_n5167_));
  INV_X1     g04975(.I(new_n5167_), .ZN(new_n5168_));
  NAND3_X1   g04976(.A1(\asqrt[33] ), .A2(new_n4943_), .A3(new_n4962_), .ZN(new_n5169_));
  XOR2_X1    g04977(.A1(new_n5169_), .A2(new_n4977_), .Z(new_n5170_));
  INV_X1     g04978(.I(new_n5170_), .ZN(new_n5171_));
  OAI21_X1   g04979(.A1(new_n4937_), .A2(new_n4939_), .B(new_n4942_), .ZN(new_n5172_));
  NOR2_X1    g04980(.A1(new_n5110_), .A2(new_n5172_), .ZN(new_n5173_));
  XOR2_X1    g04981(.A1(new_n5173_), .A2(new_n4863_), .Z(new_n5174_));
  NAND3_X1   g04982(.A1(\asqrt[33] ), .A2(new_n4956_), .A3(new_n4938_), .ZN(new_n5175_));
  XOR2_X1    g04983(.A1(new_n5175_), .A2(new_n4867_), .Z(new_n5176_));
  OAI21_X1   g04984(.A1(new_n4951_), .A2(new_n4952_), .B(new_n4955_), .ZN(new_n5177_));
  NOR2_X1    g04985(.A1(new_n5110_), .A2(new_n5177_), .ZN(new_n5178_));
  XOR2_X1    g04986(.A1(new_n5178_), .A2(new_n4869_), .Z(new_n5179_));
  INV_X1     g04987(.I(new_n5179_), .ZN(new_n5180_));
  NAND3_X1   g04988(.A1(\asqrt[33] ), .A2(new_n4908_), .A3(new_n4934_), .ZN(new_n5181_));
  XOR2_X1    g04989(.A1(new_n5181_), .A2(new_n4949_), .Z(new_n5182_));
  INV_X1     g04990(.I(new_n5182_), .ZN(new_n5183_));
  AOI21_X1   g04991(.A1(new_n4929_), .A2(new_n4930_), .B(new_n4933_), .ZN(new_n5184_));
  NAND2_X1   g04992(.A1(\asqrt[33] ), .A2(new_n5184_), .ZN(new_n5185_));
  XOR2_X1    g04993(.A1(new_n5185_), .A2(new_n4913_), .Z(new_n5186_));
  NOR2_X1    g04994(.A1(new_n4928_), .A2(\asqrt[38] ), .ZN(new_n5187_));
  NOR3_X1    g04995(.A1(new_n5110_), .A2(new_n5187_), .A3(new_n4906_), .ZN(new_n5188_));
  XOR2_X1    g04996(.A1(new_n5188_), .A2(new_n4878_), .Z(new_n5189_));
  NOR3_X1    g04997(.A1(new_n5110_), .A2(new_n4925_), .A3(new_n4901_), .ZN(new_n5190_));
  XOR2_X1    g04998(.A1(new_n5190_), .A2(new_n4900_), .Z(new_n5191_));
  INV_X1     g04999(.I(new_n5191_), .ZN(new_n5192_));
  NOR2_X1    g05000(.A1(new_n4895_), .A2(\asqrt[36] ), .ZN(new_n5193_));
  NOR3_X1    g05001(.A1(new_n5110_), .A2(new_n5193_), .A3(new_n4924_), .ZN(new_n5194_));
  XOR2_X1    g05002(.A1(new_n5194_), .A2(new_n4886_), .Z(new_n5195_));
  INV_X1     g05003(.I(new_n5195_), .ZN(new_n5196_));
  NAND3_X1   g05004(.A1(\asqrt[33] ), .A2(new_n4887_), .A3(new_n4888_), .ZN(new_n5197_));
  NOR4_X1    g05005(.A1(new_n5107_), .A2(new_n4810_), .A3(new_n5102_), .A4(new_n5108_), .ZN(new_n5198_));
  INV_X1     g05006(.I(new_n5198_), .ZN(new_n5199_));
  AOI21_X1   g05007(.A1(new_n5197_), .A2(new_n5199_), .B(\a[68] ), .ZN(new_n5200_));
  NOR3_X1    g05008(.A1(new_n5110_), .A2(\a[66] ), .A3(\a[67] ), .ZN(new_n5201_));
  NOR3_X1    g05009(.A1(new_n5201_), .A2(new_n4584_), .A3(new_n5198_), .ZN(new_n5202_));
  NOR2_X1    g05010(.A1(new_n5202_), .A2(new_n5200_), .ZN(new_n5203_));
  NAND3_X1   g05011(.A1(new_n195_), .A2(new_n196_), .A3(new_n4887_), .ZN(new_n5204_));
  OAI21_X1   g05012(.A1(new_n5110_), .A2(new_n4887_), .B(new_n5204_), .ZN(new_n5205_));
  NAND2_X1   g05013(.A1(new_n5205_), .A2(\asqrt[34] ), .ZN(new_n5206_));
  OAI21_X1   g05014(.A1(new_n5110_), .A2(\a[66] ), .B(\a[67] ), .ZN(new_n5207_));
  NAND2_X1   g05015(.A1(new_n5207_), .A2(new_n5197_), .ZN(new_n5208_));
  NOR2_X1    g05016(.A1(new_n5205_), .A2(\asqrt[34] ), .ZN(new_n5209_));
  OAI21_X1   g05017(.A1(new_n5208_), .A2(new_n5209_), .B(new_n5206_), .ZN(new_n5210_));
  OAI21_X1   g05018(.A1(\asqrt[35] ), .A2(new_n5210_), .B(new_n5203_), .ZN(new_n5211_));
  NAND2_X1   g05019(.A1(new_n5210_), .A2(\asqrt[35] ), .ZN(new_n5212_));
  NAND3_X1   g05020(.A1(new_n5211_), .A2(new_n4224_), .A3(new_n5212_), .ZN(new_n5213_));
  NOR3_X1    g05021(.A1(new_n5110_), .A2(new_n4918_), .A3(new_n4894_), .ZN(new_n5214_));
  XOR2_X1    g05022(.A1(new_n5214_), .A2(new_n4920_), .Z(new_n5215_));
  NAND2_X1   g05023(.A1(new_n5213_), .A2(new_n5215_), .ZN(new_n5216_));
  NAND2_X1   g05024(.A1(new_n5211_), .A2(new_n5212_), .ZN(new_n5217_));
  AOI21_X1   g05025(.A1(new_n5217_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n5218_));
  AOI21_X1   g05026(.A1(new_n5218_), .A2(new_n5216_), .B(new_n5196_), .ZN(new_n5219_));
  OAI21_X1   g05027(.A1(new_n5201_), .A2(new_n5198_), .B(new_n4584_), .ZN(new_n5220_));
  NAND3_X1   g05028(.A1(new_n5197_), .A2(\a[68] ), .A3(new_n5199_), .ZN(new_n5221_));
  NAND2_X1   g05029(.A1(new_n5220_), .A2(new_n5221_), .ZN(new_n5222_));
  NAND2_X1   g05030(.A1(\asqrt[33] ), .A2(\a[66] ), .ZN(new_n5223_));
  AOI21_X1   g05031(.A1(new_n5223_), .A2(new_n5204_), .B(new_n4810_), .ZN(new_n5224_));
  AOI21_X1   g05032(.A1(\asqrt[33] ), .A2(new_n4887_), .B(new_n4888_), .ZN(new_n5225_));
  NOR2_X1    g05033(.A1(new_n5225_), .A2(new_n5201_), .ZN(new_n5226_));
  NAND3_X1   g05034(.A1(new_n5223_), .A2(new_n4810_), .A3(new_n5204_), .ZN(new_n5227_));
  AOI21_X1   g05035(.A1(new_n5226_), .A2(new_n5227_), .B(new_n5224_), .ZN(new_n5228_));
  AOI21_X1   g05036(.A1(new_n5228_), .A2(new_n4510_), .B(new_n5222_), .ZN(new_n5229_));
  NOR2_X1    g05037(.A1(new_n5228_), .A2(new_n4510_), .ZN(new_n5230_));
  OAI21_X1   g05038(.A1(new_n5229_), .A2(new_n5230_), .B(\asqrt[36] ), .ZN(new_n5231_));
  AOI21_X1   g05039(.A1(new_n5216_), .A2(new_n5231_), .B(new_n3928_), .ZN(new_n5232_));
  NOR2_X1    g05040(.A1(new_n5219_), .A2(new_n5232_), .ZN(new_n5233_));
  AOI21_X1   g05041(.A1(new_n5233_), .A2(new_n3675_), .B(new_n5192_), .ZN(new_n5234_));
  OAI21_X1   g05042(.A1(new_n5219_), .A2(new_n5232_), .B(\asqrt[38] ), .ZN(new_n5235_));
  NAND2_X1   g05043(.A1(new_n5235_), .A2(new_n3400_), .ZN(new_n5236_));
  OAI21_X1   g05044(.A1(new_n5234_), .A2(new_n5236_), .B(new_n5189_), .ZN(new_n5237_));
  INV_X1     g05045(.I(new_n5235_), .ZN(new_n5238_));
  OAI21_X1   g05046(.A1(new_n5234_), .A2(new_n5238_), .B(\asqrt[39] ), .ZN(new_n5239_));
  NAND3_X1   g05047(.A1(new_n5237_), .A2(new_n5239_), .A3(new_n3167_), .ZN(new_n5240_));
  NAND2_X1   g05048(.A1(new_n5240_), .A2(new_n5186_), .ZN(new_n5241_));
  NAND2_X1   g05049(.A1(new_n5237_), .A2(new_n5239_), .ZN(new_n5242_));
  AOI21_X1   g05050(.A1(new_n5242_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n5243_));
  AOI21_X1   g05051(.A1(new_n5243_), .A2(new_n5241_), .B(new_n5183_), .ZN(new_n5244_));
  INV_X1     g05052(.I(new_n5189_), .ZN(new_n5245_));
  NOR2_X1    g05053(.A1(new_n5229_), .A2(new_n5230_), .ZN(new_n5246_));
  INV_X1     g05054(.I(new_n5215_), .ZN(new_n5247_));
  AOI21_X1   g05055(.A1(new_n5246_), .A2(new_n4224_), .B(new_n5247_), .ZN(new_n5248_));
  NAND2_X1   g05056(.A1(new_n5231_), .A2(new_n3928_), .ZN(new_n5249_));
  OAI21_X1   g05057(.A1(new_n5248_), .A2(new_n5249_), .B(new_n5195_), .ZN(new_n5250_));
  INV_X1     g05058(.I(new_n5231_), .ZN(new_n5251_));
  OAI21_X1   g05059(.A1(new_n5248_), .A2(new_n5251_), .B(\asqrt[37] ), .ZN(new_n5252_));
  NAND3_X1   g05060(.A1(new_n5250_), .A2(new_n5252_), .A3(new_n3675_), .ZN(new_n5253_));
  NAND2_X1   g05061(.A1(new_n5253_), .A2(new_n5191_), .ZN(new_n5254_));
  NAND2_X1   g05062(.A1(new_n5250_), .A2(new_n5252_), .ZN(new_n5255_));
  AOI21_X1   g05063(.A1(new_n5255_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n5256_));
  AOI21_X1   g05064(.A1(new_n5256_), .A2(new_n5254_), .B(new_n5245_), .ZN(new_n5257_));
  AOI21_X1   g05065(.A1(new_n5254_), .A2(new_n5235_), .B(new_n3400_), .ZN(new_n5258_));
  OAI21_X1   g05066(.A1(new_n5257_), .A2(new_n5258_), .B(\asqrt[40] ), .ZN(new_n5259_));
  AOI21_X1   g05067(.A1(new_n5241_), .A2(new_n5259_), .B(new_n2912_), .ZN(new_n5260_));
  NOR2_X1    g05068(.A1(new_n5244_), .A2(new_n5260_), .ZN(new_n5261_));
  AOI21_X1   g05069(.A1(new_n5261_), .A2(new_n2699_), .B(new_n5180_), .ZN(new_n5262_));
  OAI21_X1   g05070(.A1(new_n5244_), .A2(new_n5260_), .B(\asqrt[42] ), .ZN(new_n5263_));
  NAND2_X1   g05071(.A1(new_n5263_), .A2(new_n2464_), .ZN(new_n5264_));
  OAI21_X1   g05072(.A1(new_n5262_), .A2(new_n5264_), .B(new_n5176_), .ZN(new_n5265_));
  INV_X1     g05073(.I(new_n5263_), .ZN(new_n5266_));
  OAI21_X1   g05074(.A1(new_n5262_), .A2(new_n5266_), .B(\asqrt[43] ), .ZN(new_n5267_));
  NAND3_X1   g05075(.A1(new_n5265_), .A2(new_n5267_), .A3(new_n2271_), .ZN(new_n5268_));
  NAND2_X1   g05076(.A1(new_n5268_), .A2(new_n5174_), .ZN(new_n5269_));
  NAND2_X1   g05077(.A1(new_n5265_), .A2(new_n5267_), .ZN(new_n5270_));
  AOI21_X1   g05078(.A1(new_n5270_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n5271_));
  AOI21_X1   g05079(.A1(new_n5271_), .A2(new_n5269_), .B(new_n5171_), .ZN(new_n5272_));
  INV_X1     g05080(.I(new_n5176_), .ZN(new_n5273_));
  INV_X1     g05081(.I(new_n5186_), .ZN(new_n5274_));
  NOR2_X1    g05082(.A1(new_n5257_), .A2(new_n5258_), .ZN(new_n5275_));
  AOI21_X1   g05083(.A1(new_n5275_), .A2(new_n3167_), .B(new_n5274_), .ZN(new_n5276_));
  NAND2_X1   g05084(.A1(new_n5259_), .A2(new_n2912_), .ZN(new_n5277_));
  OAI21_X1   g05085(.A1(new_n5276_), .A2(new_n5277_), .B(new_n5182_), .ZN(new_n5278_));
  INV_X1     g05086(.I(new_n5259_), .ZN(new_n5279_));
  OAI21_X1   g05087(.A1(new_n5276_), .A2(new_n5279_), .B(\asqrt[41] ), .ZN(new_n5280_));
  NAND3_X1   g05088(.A1(new_n5278_), .A2(new_n5280_), .A3(new_n2699_), .ZN(new_n5281_));
  NAND2_X1   g05089(.A1(new_n5281_), .A2(new_n5179_), .ZN(new_n5282_));
  NAND2_X1   g05090(.A1(new_n5278_), .A2(new_n5280_), .ZN(new_n5283_));
  AOI21_X1   g05091(.A1(new_n5283_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n5284_));
  AOI21_X1   g05092(.A1(new_n5284_), .A2(new_n5282_), .B(new_n5273_), .ZN(new_n5285_));
  AOI21_X1   g05093(.A1(new_n5282_), .A2(new_n5263_), .B(new_n2464_), .ZN(new_n5286_));
  OAI21_X1   g05094(.A1(new_n5285_), .A2(new_n5286_), .B(\asqrt[44] ), .ZN(new_n5287_));
  AOI21_X1   g05095(.A1(new_n5269_), .A2(new_n5287_), .B(new_n2072_), .ZN(new_n5288_));
  NOR2_X1    g05096(.A1(new_n5272_), .A2(new_n5288_), .ZN(new_n5289_));
  AOI21_X1   g05097(.A1(new_n5289_), .A2(new_n1884_), .B(new_n5168_), .ZN(new_n5290_));
  OAI21_X1   g05098(.A1(new_n5272_), .A2(new_n5288_), .B(\asqrt[46] ), .ZN(new_n5291_));
  NAND2_X1   g05099(.A1(new_n5291_), .A2(new_n1688_), .ZN(new_n5292_));
  OAI21_X1   g05100(.A1(new_n5290_), .A2(new_n5292_), .B(new_n5164_), .ZN(new_n5293_));
  INV_X1     g05101(.I(new_n5291_), .ZN(new_n5294_));
  OAI21_X1   g05102(.A1(new_n5290_), .A2(new_n5294_), .B(\asqrt[47] ), .ZN(new_n5295_));
  NAND3_X1   g05103(.A1(new_n5293_), .A2(new_n5295_), .A3(new_n1533_), .ZN(new_n5296_));
  NAND2_X1   g05104(.A1(new_n5296_), .A2(new_n5162_), .ZN(new_n5297_));
  NAND2_X1   g05105(.A1(new_n5293_), .A2(new_n5295_), .ZN(new_n5298_));
  AOI21_X1   g05106(.A1(new_n5298_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n5299_));
  AOI21_X1   g05107(.A1(new_n5299_), .A2(new_n5297_), .B(new_n5159_), .ZN(new_n5300_));
  INV_X1     g05108(.I(new_n5164_), .ZN(new_n5301_));
  INV_X1     g05109(.I(new_n5174_), .ZN(new_n5302_));
  NOR2_X1    g05110(.A1(new_n5285_), .A2(new_n5286_), .ZN(new_n5303_));
  AOI21_X1   g05111(.A1(new_n5303_), .A2(new_n2271_), .B(new_n5302_), .ZN(new_n5304_));
  NAND2_X1   g05112(.A1(new_n5287_), .A2(new_n2072_), .ZN(new_n5305_));
  OAI21_X1   g05113(.A1(new_n5304_), .A2(new_n5305_), .B(new_n5170_), .ZN(new_n5306_));
  INV_X1     g05114(.I(new_n5287_), .ZN(new_n5307_));
  OAI21_X1   g05115(.A1(new_n5304_), .A2(new_n5307_), .B(\asqrt[45] ), .ZN(new_n5308_));
  NAND3_X1   g05116(.A1(new_n5306_), .A2(new_n5308_), .A3(new_n1884_), .ZN(new_n5309_));
  NAND2_X1   g05117(.A1(new_n5309_), .A2(new_n5167_), .ZN(new_n5310_));
  NAND2_X1   g05118(.A1(new_n5306_), .A2(new_n5308_), .ZN(new_n5311_));
  AOI21_X1   g05119(.A1(new_n5311_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n5312_));
  AOI21_X1   g05120(.A1(new_n5312_), .A2(new_n5310_), .B(new_n5301_), .ZN(new_n5313_));
  AOI21_X1   g05121(.A1(new_n5310_), .A2(new_n5291_), .B(new_n1688_), .ZN(new_n5314_));
  OAI21_X1   g05122(.A1(new_n5313_), .A2(new_n5314_), .B(\asqrt[48] ), .ZN(new_n5315_));
  AOI21_X1   g05123(.A1(new_n5297_), .A2(new_n5315_), .B(new_n1368_), .ZN(new_n5316_));
  NOR2_X1    g05124(.A1(new_n5300_), .A2(new_n5316_), .ZN(new_n5317_));
  AOI21_X1   g05125(.A1(new_n5317_), .A2(new_n1228_), .B(new_n5156_), .ZN(new_n5318_));
  OAI21_X1   g05126(.A1(new_n5300_), .A2(new_n5316_), .B(\asqrt[50] ), .ZN(new_n5319_));
  NAND2_X1   g05127(.A1(new_n5319_), .A2(new_n1088_), .ZN(new_n5320_));
  OAI21_X1   g05128(.A1(new_n5318_), .A2(new_n5320_), .B(new_n5152_), .ZN(new_n5321_));
  INV_X1     g05129(.I(new_n5319_), .ZN(new_n5322_));
  OAI21_X1   g05130(.A1(new_n5318_), .A2(new_n5322_), .B(\asqrt[51] ), .ZN(new_n5323_));
  NAND3_X1   g05131(.A1(new_n5321_), .A2(new_n5323_), .A3(new_n962_), .ZN(new_n5324_));
  NAND2_X1   g05132(.A1(new_n5324_), .A2(new_n5150_), .ZN(new_n5325_));
  NAND2_X1   g05133(.A1(new_n5321_), .A2(new_n5323_), .ZN(new_n5326_));
  AOI21_X1   g05134(.A1(new_n5326_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n5327_));
  AOI21_X1   g05135(.A1(new_n5327_), .A2(new_n5325_), .B(new_n5147_), .ZN(new_n5328_));
  INV_X1     g05136(.I(new_n5152_), .ZN(new_n5329_));
  INV_X1     g05137(.I(new_n5162_), .ZN(new_n5330_));
  NOR2_X1    g05138(.A1(new_n5313_), .A2(new_n5314_), .ZN(new_n5331_));
  AOI21_X1   g05139(.A1(new_n5331_), .A2(new_n1533_), .B(new_n5330_), .ZN(new_n5332_));
  NAND2_X1   g05140(.A1(new_n5315_), .A2(new_n1368_), .ZN(new_n5333_));
  OAI21_X1   g05141(.A1(new_n5332_), .A2(new_n5333_), .B(new_n5158_), .ZN(new_n5334_));
  INV_X1     g05142(.I(new_n5315_), .ZN(new_n5335_));
  OAI21_X1   g05143(.A1(new_n5332_), .A2(new_n5335_), .B(\asqrt[49] ), .ZN(new_n5336_));
  NAND3_X1   g05144(.A1(new_n5334_), .A2(new_n5336_), .A3(new_n1228_), .ZN(new_n5337_));
  NAND2_X1   g05145(.A1(new_n5337_), .A2(new_n5155_), .ZN(new_n5338_));
  NAND2_X1   g05146(.A1(new_n5334_), .A2(new_n5336_), .ZN(new_n5339_));
  AOI21_X1   g05147(.A1(new_n5339_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n5340_));
  AOI21_X1   g05148(.A1(new_n5340_), .A2(new_n5338_), .B(new_n5329_), .ZN(new_n5341_));
  AOI21_X1   g05149(.A1(new_n5338_), .A2(new_n5319_), .B(new_n1088_), .ZN(new_n5342_));
  OAI21_X1   g05150(.A1(new_n5341_), .A2(new_n5342_), .B(\asqrt[52] ), .ZN(new_n5343_));
  AOI21_X1   g05151(.A1(new_n5325_), .A2(new_n5343_), .B(new_n842_), .ZN(new_n5344_));
  NOR2_X1    g05152(.A1(new_n5328_), .A2(new_n5344_), .ZN(new_n5345_));
  AOI21_X1   g05153(.A1(new_n5345_), .A2(new_n720_), .B(new_n5144_), .ZN(new_n5346_));
  OAI21_X1   g05154(.A1(new_n5328_), .A2(new_n5344_), .B(\asqrt[54] ), .ZN(new_n5347_));
  NAND2_X1   g05155(.A1(new_n5347_), .A2(new_n630_), .ZN(new_n5348_));
  OAI21_X1   g05156(.A1(new_n5346_), .A2(new_n5348_), .B(new_n5140_), .ZN(new_n5349_));
  INV_X1     g05157(.I(new_n5347_), .ZN(new_n5350_));
  OAI21_X1   g05158(.A1(new_n5346_), .A2(new_n5350_), .B(\asqrt[55] ), .ZN(new_n5351_));
  NAND3_X1   g05159(.A1(new_n5349_), .A2(new_n5351_), .A3(new_n545_), .ZN(new_n5352_));
  NAND2_X1   g05160(.A1(new_n5352_), .A2(new_n5138_), .ZN(new_n5353_));
  NAND2_X1   g05161(.A1(new_n5349_), .A2(new_n5351_), .ZN(new_n5354_));
  AOI21_X1   g05162(.A1(new_n5354_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n5355_));
  AOI21_X1   g05163(.A1(new_n5355_), .A2(new_n5353_), .B(new_n5135_), .ZN(new_n5356_));
  INV_X1     g05164(.I(new_n5140_), .ZN(new_n5357_));
  INV_X1     g05165(.I(new_n5150_), .ZN(new_n5358_));
  NOR2_X1    g05166(.A1(new_n5341_), .A2(new_n5342_), .ZN(new_n5359_));
  AOI21_X1   g05167(.A1(new_n5359_), .A2(new_n962_), .B(new_n5358_), .ZN(new_n5360_));
  NAND2_X1   g05168(.A1(new_n5343_), .A2(new_n842_), .ZN(new_n5361_));
  OAI21_X1   g05169(.A1(new_n5360_), .A2(new_n5361_), .B(new_n5146_), .ZN(new_n5362_));
  INV_X1     g05170(.I(new_n5343_), .ZN(new_n5363_));
  OAI21_X1   g05171(.A1(new_n5360_), .A2(new_n5363_), .B(\asqrt[53] ), .ZN(new_n5364_));
  NAND3_X1   g05172(.A1(new_n5362_), .A2(new_n5364_), .A3(new_n720_), .ZN(new_n5365_));
  NAND2_X1   g05173(.A1(new_n5365_), .A2(new_n5143_), .ZN(new_n5366_));
  NAND2_X1   g05174(.A1(new_n5362_), .A2(new_n5364_), .ZN(new_n5367_));
  AOI21_X1   g05175(.A1(new_n5367_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n5368_));
  AOI21_X1   g05176(.A1(new_n5368_), .A2(new_n5366_), .B(new_n5357_), .ZN(new_n5369_));
  AOI21_X1   g05177(.A1(new_n5366_), .A2(new_n5347_), .B(new_n630_), .ZN(new_n5370_));
  OAI21_X1   g05178(.A1(new_n5369_), .A2(new_n5370_), .B(\asqrt[56] ), .ZN(new_n5371_));
  AOI21_X1   g05179(.A1(new_n5353_), .A2(new_n5371_), .B(new_n450_), .ZN(new_n5372_));
  NOR2_X1    g05180(.A1(new_n5356_), .A2(new_n5372_), .ZN(new_n5373_));
  AOI21_X1   g05181(.A1(new_n5373_), .A2(new_n403_), .B(new_n5132_), .ZN(new_n5374_));
  OAI21_X1   g05182(.A1(new_n5356_), .A2(new_n5372_), .B(\asqrt[58] ), .ZN(new_n5375_));
  NAND2_X1   g05183(.A1(new_n5375_), .A2(new_n339_), .ZN(new_n5376_));
  OAI21_X1   g05184(.A1(new_n5374_), .A2(new_n5376_), .B(new_n5128_), .ZN(new_n5377_));
  INV_X1     g05185(.I(new_n5375_), .ZN(new_n5378_));
  OAI21_X1   g05186(.A1(new_n5374_), .A2(new_n5378_), .B(\asqrt[59] ), .ZN(new_n5379_));
  NAND3_X1   g05187(.A1(new_n5377_), .A2(new_n5379_), .A3(new_n288_), .ZN(new_n5380_));
  NAND2_X1   g05188(.A1(new_n5380_), .A2(new_n5126_), .ZN(new_n5381_));
  INV_X1     g05189(.I(new_n5128_), .ZN(new_n5382_));
  INV_X1     g05190(.I(new_n5138_), .ZN(new_n5383_));
  NOR2_X1    g05191(.A1(new_n5369_), .A2(new_n5370_), .ZN(new_n5384_));
  AOI21_X1   g05192(.A1(new_n5384_), .A2(new_n545_), .B(new_n5383_), .ZN(new_n5385_));
  NAND2_X1   g05193(.A1(new_n5371_), .A2(new_n450_), .ZN(new_n5386_));
  OAI21_X1   g05194(.A1(new_n5385_), .A2(new_n5386_), .B(new_n5134_), .ZN(new_n5387_));
  INV_X1     g05195(.I(new_n5371_), .ZN(new_n5388_));
  OAI21_X1   g05196(.A1(new_n5385_), .A2(new_n5388_), .B(\asqrt[57] ), .ZN(new_n5389_));
  NAND3_X1   g05197(.A1(new_n5387_), .A2(new_n5389_), .A3(new_n403_), .ZN(new_n5390_));
  NAND2_X1   g05198(.A1(new_n5390_), .A2(new_n5131_), .ZN(new_n5391_));
  NAND2_X1   g05199(.A1(new_n5387_), .A2(new_n5389_), .ZN(new_n5392_));
  AOI21_X1   g05200(.A1(new_n5392_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n5393_));
  AOI21_X1   g05201(.A1(new_n5393_), .A2(new_n5391_), .B(new_n5382_), .ZN(new_n5394_));
  AOI21_X1   g05202(.A1(new_n5391_), .A2(new_n5375_), .B(new_n339_), .ZN(new_n5395_));
  OAI21_X1   g05203(.A1(new_n5394_), .A2(new_n5395_), .B(\asqrt[60] ), .ZN(new_n5396_));
  AOI21_X1   g05204(.A1(new_n5381_), .A2(new_n5396_), .B(new_n242_), .ZN(new_n5397_));
  NAND3_X1   g05205(.A1(\asqrt[33] ), .A2(new_n5055_), .A3(new_n5071_), .ZN(new_n5398_));
  XOR2_X1    g05206(.A1(new_n5398_), .A2(new_n5083_), .Z(new_n5399_));
  INV_X1     g05207(.I(new_n5399_), .ZN(new_n5400_));
  NAND2_X1   g05208(.A1(new_n5377_), .A2(new_n5379_), .ZN(new_n5401_));
  AOI21_X1   g05209(.A1(new_n5401_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n5402_));
  AOI21_X1   g05210(.A1(new_n5402_), .A2(new_n5381_), .B(new_n5400_), .ZN(new_n5403_));
  OAI21_X1   g05211(.A1(new_n5403_), .A2(new_n5397_), .B(\asqrt[62] ), .ZN(new_n5404_));
  INV_X1     g05212(.I(new_n5404_), .ZN(new_n5405_));
  NOR2_X1    g05213(.A1(new_n5403_), .A2(new_n5397_), .ZN(new_n5406_));
  AOI21_X1   g05214(.A1(new_n5056_), .A2(new_n5077_), .B(new_n5072_), .ZN(new_n5407_));
  NAND2_X1   g05215(.A1(\asqrt[33] ), .A2(new_n5407_), .ZN(new_n5408_));
  XOR2_X1    g05216(.A1(new_n5408_), .A2(new_n5075_), .Z(new_n5409_));
  INV_X1     g05217(.I(new_n5409_), .ZN(new_n5410_));
  AOI21_X1   g05218(.A1(new_n5406_), .A2(new_n234_), .B(new_n5410_), .ZN(new_n5411_));
  OAI21_X1   g05219(.A1(new_n5411_), .A2(new_n5405_), .B(new_n5123_), .ZN(new_n5412_));
  OAI21_X1   g05220(.A1(new_n5412_), .A2(new_n5122_), .B(new_n193_), .ZN(new_n5413_));
  NOR2_X1    g05221(.A1(new_n5411_), .A2(new_n5405_), .ZN(new_n5414_));
  NAND2_X1   g05222(.A1(new_n5414_), .A2(new_n5122_), .ZN(new_n5415_));
  NOR2_X1    g05223(.A1(\asqrt[33] ), .A2(new_n5103_), .ZN(new_n5416_));
  INV_X1     g05224(.I(new_n5416_), .ZN(new_n5417_));
  NAND4_X1   g05225(.A1(new_n5413_), .A2(new_n5114_), .A3(new_n5415_), .A4(new_n5417_), .ZN(\asqrt[32] ));
  AOI21_X1   g05226(.A1(\asqrt[32] ), .A2(new_n195_), .B(new_n196_), .ZN(new_n5419_));
  INV_X1     g05227(.I(new_n5122_), .ZN(new_n5420_));
  INV_X1     g05228(.I(new_n5123_), .ZN(new_n5421_));
  INV_X1     g05229(.I(new_n5126_), .ZN(new_n5422_));
  NOR2_X1    g05230(.A1(new_n5394_), .A2(new_n5395_), .ZN(new_n5423_));
  AOI21_X1   g05231(.A1(new_n5423_), .A2(new_n288_), .B(new_n5422_), .ZN(new_n5424_));
  INV_X1     g05232(.I(new_n5396_), .ZN(new_n5425_));
  OAI21_X1   g05233(.A1(new_n5424_), .A2(new_n5425_), .B(\asqrt[61] ), .ZN(new_n5426_));
  NAND2_X1   g05234(.A1(new_n5396_), .A2(new_n242_), .ZN(new_n5427_));
  OAI21_X1   g05235(.A1(new_n5424_), .A2(new_n5427_), .B(new_n5399_), .ZN(new_n5428_));
  NAND3_X1   g05236(.A1(new_n5428_), .A2(new_n5426_), .A3(new_n234_), .ZN(new_n5429_));
  NAND2_X1   g05237(.A1(new_n5429_), .A2(new_n5409_), .ZN(new_n5430_));
  AOI21_X1   g05238(.A1(new_n5430_), .A2(new_n5404_), .B(new_n5421_), .ZN(new_n5431_));
  AOI21_X1   g05239(.A1(new_n5431_), .A2(new_n5420_), .B(\asqrt[63] ), .ZN(new_n5432_));
  NAND2_X1   g05240(.A1(new_n5430_), .A2(new_n5404_), .ZN(new_n5433_));
  NOR2_X1    g05241(.A1(new_n5433_), .A2(new_n5420_), .ZN(new_n5434_));
  NOR4_X1    g05242(.A1(new_n5432_), .A2(new_n5113_), .A3(new_n5434_), .A4(new_n5416_), .ZN(new_n5435_));
  NOR3_X1    g05243(.A1(new_n5435_), .A2(\a[64] ), .A3(\a[65] ), .ZN(new_n5436_));
  NOR2_X1    g05244(.A1(new_n5419_), .A2(new_n5436_), .ZN(new_n5437_));
  INV_X1     g05245(.I(\a[62] ), .ZN(new_n5438_));
  INV_X1     g05246(.I(\a[63] ), .ZN(new_n5439_));
  NAND3_X1   g05247(.A1(new_n5438_), .A2(new_n5439_), .A3(new_n195_), .ZN(new_n5440_));
  NAND2_X1   g05248(.A1(\asqrt[32] ), .A2(\a[64] ), .ZN(new_n5441_));
  AOI21_X1   g05249(.A1(new_n5441_), .A2(new_n5440_), .B(new_n5110_), .ZN(new_n5442_));
  OAI21_X1   g05250(.A1(new_n5435_), .A2(new_n195_), .B(new_n5440_), .ZN(new_n5443_));
  NOR2_X1    g05251(.A1(new_n5443_), .A2(\asqrt[33] ), .ZN(new_n5444_));
  NAND2_X1   g05252(.A1(new_n5433_), .A2(new_n5122_), .ZN(new_n5445_));
  NOR2_X1    g05253(.A1(new_n5435_), .A2(new_n5122_), .ZN(new_n5446_));
  NAND2_X1   g05254(.A1(new_n5446_), .A2(new_n5414_), .ZN(new_n5447_));
  AOI21_X1   g05255(.A1(new_n5447_), .A2(new_n5445_), .B(new_n193_), .ZN(new_n5448_));
  NAND3_X1   g05256(.A1(\asqrt[32] ), .A2(new_n5404_), .A3(new_n5429_), .ZN(new_n5449_));
  XOR2_X1    g05257(.A1(new_n5449_), .A2(new_n5409_), .Z(new_n5450_));
  INV_X1     g05258(.I(new_n5450_), .ZN(new_n5451_));
  AOI21_X1   g05259(.A1(new_n5446_), .A2(new_n5433_), .B(new_n5434_), .ZN(new_n5452_));
  INV_X1     g05260(.I(new_n5452_), .ZN(new_n5453_));
  OAI21_X1   g05261(.A1(new_n5374_), .A2(new_n5376_), .B(new_n5379_), .ZN(new_n5454_));
  NOR2_X1    g05262(.A1(new_n5435_), .A2(new_n5454_), .ZN(new_n5455_));
  XOR2_X1    g05263(.A1(new_n5455_), .A2(new_n5128_), .Z(new_n5456_));
  NAND3_X1   g05264(.A1(\asqrt[32] ), .A2(new_n5390_), .A3(new_n5375_), .ZN(new_n5457_));
  XOR2_X1    g05265(.A1(new_n5457_), .A2(new_n5132_), .Z(new_n5458_));
  OAI21_X1   g05266(.A1(new_n5385_), .A2(new_n5386_), .B(new_n5389_), .ZN(new_n5459_));
  NOR2_X1    g05267(.A1(new_n5435_), .A2(new_n5459_), .ZN(new_n5460_));
  XOR2_X1    g05268(.A1(new_n5460_), .A2(new_n5134_), .Z(new_n5461_));
  INV_X1     g05269(.I(new_n5461_), .ZN(new_n5462_));
  NAND3_X1   g05270(.A1(\asqrt[32] ), .A2(new_n5352_), .A3(new_n5371_), .ZN(new_n5463_));
  XOR2_X1    g05271(.A1(new_n5463_), .A2(new_n5383_), .Z(new_n5464_));
  INV_X1     g05272(.I(new_n5464_), .ZN(new_n5465_));
  OAI21_X1   g05273(.A1(new_n5346_), .A2(new_n5348_), .B(new_n5351_), .ZN(new_n5466_));
  NOR2_X1    g05274(.A1(new_n5435_), .A2(new_n5466_), .ZN(new_n5467_));
  XOR2_X1    g05275(.A1(new_n5467_), .A2(new_n5140_), .Z(new_n5468_));
  NAND3_X1   g05276(.A1(\asqrt[32] ), .A2(new_n5365_), .A3(new_n5347_), .ZN(new_n5469_));
  XOR2_X1    g05277(.A1(new_n5469_), .A2(new_n5144_), .Z(new_n5470_));
  OAI21_X1   g05278(.A1(new_n5360_), .A2(new_n5361_), .B(new_n5364_), .ZN(new_n5471_));
  NOR2_X1    g05279(.A1(new_n5435_), .A2(new_n5471_), .ZN(new_n5472_));
  XOR2_X1    g05280(.A1(new_n5472_), .A2(new_n5146_), .Z(new_n5473_));
  INV_X1     g05281(.I(new_n5473_), .ZN(new_n5474_));
  NAND3_X1   g05282(.A1(\asqrt[32] ), .A2(new_n5324_), .A3(new_n5343_), .ZN(new_n5475_));
  XOR2_X1    g05283(.A1(new_n5475_), .A2(new_n5358_), .Z(new_n5476_));
  INV_X1     g05284(.I(new_n5476_), .ZN(new_n5477_));
  OAI21_X1   g05285(.A1(new_n5318_), .A2(new_n5320_), .B(new_n5323_), .ZN(new_n5478_));
  NOR2_X1    g05286(.A1(new_n5435_), .A2(new_n5478_), .ZN(new_n5479_));
  XOR2_X1    g05287(.A1(new_n5479_), .A2(new_n5152_), .Z(new_n5480_));
  NAND3_X1   g05288(.A1(\asqrt[32] ), .A2(new_n5337_), .A3(new_n5319_), .ZN(new_n5481_));
  XOR2_X1    g05289(.A1(new_n5481_), .A2(new_n5156_), .Z(new_n5482_));
  OAI21_X1   g05290(.A1(new_n5332_), .A2(new_n5333_), .B(new_n5336_), .ZN(new_n5483_));
  NOR2_X1    g05291(.A1(new_n5435_), .A2(new_n5483_), .ZN(new_n5484_));
  XOR2_X1    g05292(.A1(new_n5484_), .A2(new_n5158_), .Z(new_n5485_));
  INV_X1     g05293(.I(new_n5485_), .ZN(new_n5486_));
  NAND3_X1   g05294(.A1(\asqrt[32] ), .A2(new_n5296_), .A3(new_n5315_), .ZN(new_n5487_));
  XOR2_X1    g05295(.A1(new_n5487_), .A2(new_n5330_), .Z(new_n5488_));
  INV_X1     g05296(.I(new_n5488_), .ZN(new_n5489_));
  OAI21_X1   g05297(.A1(new_n5290_), .A2(new_n5292_), .B(new_n5295_), .ZN(new_n5490_));
  NOR2_X1    g05298(.A1(new_n5435_), .A2(new_n5490_), .ZN(new_n5491_));
  XOR2_X1    g05299(.A1(new_n5491_), .A2(new_n5164_), .Z(new_n5492_));
  NAND3_X1   g05300(.A1(\asqrt[32] ), .A2(new_n5309_), .A3(new_n5291_), .ZN(new_n5493_));
  XOR2_X1    g05301(.A1(new_n5493_), .A2(new_n5168_), .Z(new_n5494_));
  OAI21_X1   g05302(.A1(new_n5304_), .A2(new_n5305_), .B(new_n5308_), .ZN(new_n5495_));
  NOR2_X1    g05303(.A1(new_n5435_), .A2(new_n5495_), .ZN(new_n5496_));
  XOR2_X1    g05304(.A1(new_n5496_), .A2(new_n5170_), .Z(new_n5497_));
  INV_X1     g05305(.I(new_n5497_), .ZN(new_n5498_));
  NAND3_X1   g05306(.A1(\asqrt[32] ), .A2(new_n5268_), .A3(new_n5287_), .ZN(new_n5499_));
  XOR2_X1    g05307(.A1(new_n5499_), .A2(new_n5302_), .Z(new_n5500_));
  INV_X1     g05308(.I(new_n5500_), .ZN(new_n5501_));
  OAI21_X1   g05309(.A1(new_n5262_), .A2(new_n5264_), .B(new_n5267_), .ZN(new_n5502_));
  NOR2_X1    g05310(.A1(new_n5435_), .A2(new_n5502_), .ZN(new_n5503_));
  XOR2_X1    g05311(.A1(new_n5503_), .A2(new_n5176_), .Z(new_n5504_));
  NAND3_X1   g05312(.A1(\asqrt[32] ), .A2(new_n5281_), .A3(new_n5263_), .ZN(new_n5505_));
  XOR2_X1    g05313(.A1(new_n5505_), .A2(new_n5180_), .Z(new_n5506_));
  OAI21_X1   g05314(.A1(new_n5276_), .A2(new_n5277_), .B(new_n5280_), .ZN(new_n5507_));
  NOR2_X1    g05315(.A1(new_n5435_), .A2(new_n5507_), .ZN(new_n5508_));
  XOR2_X1    g05316(.A1(new_n5508_), .A2(new_n5182_), .Z(new_n5509_));
  INV_X1     g05317(.I(new_n5509_), .ZN(new_n5510_));
  NAND3_X1   g05318(.A1(\asqrt[32] ), .A2(new_n5240_), .A3(new_n5259_), .ZN(new_n5511_));
  XOR2_X1    g05319(.A1(new_n5511_), .A2(new_n5274_), .Z(new_n5512_));
  INV_X1     g05320(.I(new_n5512_), .ZN(new_n5513_));
  OAI21_X1   g05321(.A1(new_n5234_), .A2(new_n5236_), .B(new_n5239_), .ZN(new_n5514_));
  NOR2_X1    g05322(.A1(new_n5435_), .A2(new_n5514_), .ZN(new_n5515_));
  XOR2_X1    g05323(.A1(new_n5515_), .A2(new_n5189_), .Z(new_n5516_));
  NAND3_X1   g05324(.A1(\asqrt[32] ), .A2(new_n5253_), .A3(new_n5235_), .ZN(new_n5517_));
  XOR2_X1    g05325(.A1(new_n5517_), .A2(new_n5192_), .Z(new_n5518_));
  OAI21_X1   g05326(.A1(new_n5248_), .A2(new_n5249_), .B(new_n5252_), .ZN(new_n5519_));
  NOR2_X1    g05327(.A1(new_n5435_), .A2(new_n5519_), .ZN(new_n5520_));
  XOR2_X1    g05328(.A1(new_n5520_), .A2(new_n5195_), .Z(new_n5521_));
  INV_X1     g05329(.I(new_n5521_), .ZN(new_n5522_));
  NAND3_X1   g05330(.A1(\asqrt[32] ), .A2(new_n5213_), .A3(new_n5231_), .ZN(new_n5523_));
  XOR2_X1    g05331(.A1(new_n5523_), .A2(new_n5247_), .Z(new_n5524_));
  INV_X1     g05332(.I(new_n5524_), .ZN(new_n5525_));
  NOR2_X1    g05333(.A1(new_n5210_), .A2(\asqrt[35] ), .ZN(new_n5526_));
  NOR3_X1    g05334(.A1(new_n5435_), .A2(new_n5526_), .A3(new_n5230_), .ZN(new_n5527_));
  XOR2_X1    g05335(.A1(new_n5527_), .A2(new_n5203_), .Z(new_n5528_));
  NOR4_X1    g05336(.A1(new_n5432_), .A2(new_n5110_), .A3(new_n5113_), .A4(new_n5434_), .ZN(new_n5529_));
  OAI21_X1   g05337(.A1(new_n5436_), .A2(new_n5529_), .B(new_n4887_), .ZN(new_n5530_));
  NAND3_X1   g05338(.A1(\asqrt[32] ), .A2(new_n195_), .A3(new_n196_), .ZN(new_n5531_));
  INV_X1     g05339(.I(new_n5529_), .ZN(new_n5532_));
  NAND3_X1   g05340(.A1(new_n5531_), .A2(\a[66] ), .A3(new_n5532_), .ZN(new_n5533_));
  NAND2_X1   g05341(.A1(new_n5530_), .A2(new_n5533_), .ZN(new_n5534_));
  NAND3_X1   g05342(.A1(new_n5441_), .A2(new_n5110_), .A3(new_n5440_), .ZN(new_n5535_));
  AOI21_X1   g05343(.A1(new_n5437_), .A2(new_n5535_), .B(new_n5442_), .ZN(new_n5536_));
  AOI21_X1   g05344(.A1(new_n5536_), .A2(new_n4810_), .B(new_n5534_), .ZN(new_n5537_));
  NOR2_X1    g05345(.A1(new_n5536_), .A2(new_n4810_), .ZN(new_n5538_));
  NOR3_X1    g05346(.A1(new_n5537_), .A2(\asqrt[35] ), .A3(new_n5538_), .ZN(new_n5539_));
  NOR3_X1    g05347(.A1(new_n5435_), .A2(new_n5224_), .A3(new_n5209_), .ZN(new_n5540_));
  XOR2_X1    g05348(.A1(new_n5540_), .A2(new_n5226_), .Z(new_n5541_));
  INV_X1     g05349(.I(new_n5541_), .ZN(new_n5542_));
  OAI21_X1   g05350(.A1(new_n5537_), .A2(new_n5538_), .B(\asqrt[35] ), .ZN(new_n5543_));
  OAI21_X1   g05351(.A1(new_n5539_), .A2(new_n5542_), .B(new_n5543_), .ZN(new_n5544_));
  OAI21_X1   g05352(.A1(new_n5544_), .A2(\asqrt[36] ), .B(new_n5528_), .ZN(new_n5545_));
  AOI21_X1   g05353(.A1(new_n5544_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n5546_));
  AOI21_X1   g05354(.A1(new_n5546_), .A2(new_n5545_), .B(new_n5525_), .ZN(new_n5547_));
  NAND2_X1   g05355(.A1(new_n5544_), .A2(\asqrt[36] ), .ZN(new_n5548_));
  AOI21_X1   g05356(.A1(new_n5545_), .A2(new_n5548_), .B(new_n3928_), .ZN(new_n5549_));
  NOR2_X1    g05357(.A1(new_n5547_), .A2(new_n5549_), .ZN(new_n5550_));
  AOI21_X1   g05358(.A1(new_n5550_), .A2(new_n3675_), .B(new_n5522_), .ZN(new_n5551_));
  OAI21_X1   g05359(.A1(new_n5547_), .A2(new_n5549_), .B(\asqrt[38] ), .ZN(new_n5552_));
  NAND2_X1   g05360(.A1(new_n5552_), .A2(new_n3400_), .ZN(new_n5553_));
  OAI21_X1   g05361(.A1(new_n5551_), .A2(new_n5553_), .B(new_n5518_), .ZN(new_n5554_));
  INV_X1     g05362(.I(new_n5552_), .ZN(new_n5555_));
  OAI21_X1   g05363(.A1(new_n5551_), .A2(new_n5555_), .B(\asqrt[39] ), .ZN(new_n5556_));
  NAND3_X1   g05364(.A1(new_n5554_), .A2(new_n5556_), .A3(new_n3167_), .ZN(new_n5557_));
  NAND2_X1   g05365(.A1(new_n5557_), .A2(new_n5516_), .ZN(new_n5558_));
  NAND2_X1   g05366(.A1(new_n5554_), .A2(new_n5556_), .ZN(new_n5559_));
  AOI21_X1   g05367(.A1(new_n5559_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n5560_));
  AOI21_X1   g05368(.A1(new_n5560_), .A2(new_n5558_), .B(new_n5513_), .ZN(new_n5561_));
  INV_X1     g05369(.I(new_n5518_), .ZN(new_n5562_));
  INV_X1     g05370(.I(new_n5528_), .ZN(new_n5563_));
  AOI21_X1   g05371(.A1(new_n5531_), .A2(new_n5532_), .B(\a[66] ), .ZN(new_n5564_));
  NOR3_X1    g05372(.A1(new_n5436_), .A2(new_n4887_), .A3(new_n5529_), .ZN(new_n5565_));
  NOR2_X1    g05373(.A1(new_n5565_), .A2(new_n5564_), .ZN(new_n5566_));
  OAI21_X1   g05374(.A1(new_n5435_), .A2(\a[64] ), .B(\a[65] ), .ZN(new_n5567_));
  NAND2_X1   g05375(.A1(new_n5567_), .A2(new_n5531_), .ZN(new_n5568_));
  NAND2_X1   g05376(.A1(new_n5443_), .A2(\asqrt[33] ), .ZN(new_n5569_));
  OAI21_X1   g05377(.A1(new_n5568_), .A2(new_n5444_), .B(new_n5569_), .ZN(new_n5570_));
  OAI21_X1   g05378(.A1(\asqrt[34] ), .A2(new_n5570_), .B(new_n5566_), .ZN(new_n5571_));
  NAND2_X1   g05379(.A1(new_n5570_), .A2(\asqrt[34] ), .ZN(new_n5572_));
  NAND3_X1   g05380(.A1(new_n5571_), .A2(new_n4510_), .A3(new_n5572_), .ZN(new_n5573_));
  AOI21_X1   g05381(.A1(new_n5571_), .A2(new_n5572_), .B(new_n4510_), .ZN(new_n5574_));
  AOI21_X1   g05382(.A1(new_n5573_), .A2(new_n5541_), .B(new_n5574_), .ZN(new_n5575_));
  AOI21_X1   g05383(.A1(new_n5575_), .A2(new_n4224_), .B(new_n5563_), .ZN(new_n5576_));
  OAI21_X1   g05384(.A1(new_n5575_), .A2(new_n4224_), .B(new_n3928_), .ZN(new_n5577_));
  OAI21_X1   g05385(.A1(new_n5576_), .A2(new_n5577_), .B(new_n5524_), .ZN(new_n5578_));
  NOR2_X1    g05386(.A1(new_n5575_), .A2(new_n4224_), .ZN(new_n5579_));
  OAI21_X1   g05387(.A1(new_n5576_), .A2(new_n5579_), .B(\asqrt[37] ), .ZN(new_n5580_));
  NAND3_X1   g05388(.A1(new_n5578_), .A2(new_n5580_), .A3(new_n3675_), .ZN(new_n5581_));
  NAND2_X1   g05389(.A1(new_n5581_), .A2(new_n5521_), .ZN(new_n5582_));
  NAND2_X1   g05390(.A1(new_n5578_), .A2(new_n5580_), .ZN(new_n5583_));
  AOI21_X1   g05391(.A1(new_n5583_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n5584_));
  AOI21_X1   g05392(.A1(new_n5584_), .A2(new_n5582_), .B(new_n5562_), .ZN(new_n5585_));
  AOI21_X1   g05393(.A1(new_n5582_), .A2(new_n5552_), .B(new_n3400_), .ZN(new_n5586_));
  OAI21_X1   g05394(.A1(new_n5585_), .A2(new_n5586_), .B(\asqrt[40] ), .ZN(new_n5587_));
  AOI21_X1   g05395(.A1(new_n5558_), .A2(new_n5587_), .B(new_n2912_), .ZN(new_n5588_));
  NOR2_X1    g05396(.A1(new_n5561_), .A2(new_n5588_), .ZN(new_n5589_));
  AOI21_X1   g05397(.A1(new_n5589_), .A2(new_n2699_), .B(new_n5510_), .ZN(new_n5590_));
  OAI21_X1   g05398(.A1(new_n5561_), .A2(new_n5588_), .B(\asqrt[42] ), .ZN(new_n5591_));
  NAND2_X1   g05399(.A1(new_n5591_), .A2(new_n2464_), .ZN(new_n5592_));
  OAI21_X1   g05400(.A1(new_n5590_), .A2(new_n5592_), .B(new_n5506_), .ZN(new_n5593_));
  INV_X1     g05401(.I(new_n5591_), .ZN(new_n5594_));
  OAI21_X1   g05402(.A1(new_n5590_), .A2(new_n5594_), .B(\asqrt[43] ), .ZN(new_n5595_));
  NAND3_X1   g05403(.A1(new_n5593_), .A2(new_n5595_), .A3(new_n2271_), .ZN(new_n5596_));
  NAND2_X1   g05404(.A1(new_n5596_), .A2(new_n5504_), .ZN(new_n5597_));
  NAND2_X1   g05405(.A1(new_n5593_), .A2(new_n5595_), .ZN(new_n5598_));
  AOI21_X1   g05406(.A1(new_n5598_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n5599_));
  AOI21_X1   g05407(.A1(new_n5599_), .A2(new_n5597_), .B(new_n5501_), .ZN(new_n5600_));
  INV_X1     g05408(.I(new_n5506_), .ZN(new_n5601_));
  INV_X1     g05409(.I(new_n5516_), .ZN(new_n5602_));
  NOR2_X1    g05410(.A1(new_n5585_), .A2(new_n5586_), .ZN(new_n5603_));
  AOI21_X1   g05411(.A1(new_n5603_), .A2(new_n3167_), .B(new_n5602_), .ZN(new_n5604_));
  NAND2_X1   g05412(.A1(new_n5587_), .A2(new_n2912_), .ZN(new_n5605_));
  OAI21_X1   g05413(.A1(new_n5604_), .A2(new_n5605_), .B(new_n5512_), .ZN(new_n5606_));
  INV_X1     g05414(.I(new_n5587_), .ZN(new_n5607_));
  OAI21_X1   g05415(.A1(new_n5604_), .A2(new_n5607_), .B(\asqrt[41] ), .ZN(new_n5608_));
  NAND3_X1   g05416(.A1(new_n5606_), .A2(new_n5608_), .A3(new_n2699_), .ZN(new_n5609_));
  NAND2_X1   g05417(.A1(new_n5609_), .A2(new_n5509_), .ZN(new_n5610_));
  NAND2_X1   g05418(.A1(new_n5606_), .A2(new_n5608_), .ZN(new_n5611_));
  AOI21_X1   g05419(.A1(new_n5611_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n5612_));
  AOI21_X1   g05420(.A1(new_n5612_), .A2(new_n5610_), .B(new_n5601_), .ZN(new_n5613_));
  AOI21_X1   g05421(.A1(new_n5610_), .A2(new_n5591_), .B(new_n2464_), .ZN(new_n5614_));
  OAI21_X1   g05422(.A1(new_n5613_), .A2(new_n5614_), .B(\asqrt[44] ), .ZN(new_n5615_));
  AOI21_X1   g05423(.A1(new_n5597_), .A2(new_n5615_), .B(new_n2072_), .ZN(new_n5616_));
  NOR2_X1    g05424(.A1(new_n5600_), .A2(new_n5616_), .ZN(new_n5617_));
  AOI21_X1   g05425(.A1(new_n5617_), .A2(new_n1884_), .B(new_n5498_), .ZN(new_n5618_));
  OAI21_X1   g05426(.A1(new_n5600_), .A2(new_n5616_), .B(\asqrt[46] ), .ZN(new_n5619_));
  NAND2_X1   g05427(.A1(new_n5619_), .A2(new_n1688_), .ZN(new_n5620_));
  OAI21_X1   g05428(.A1(new_n5618_), .A2(new_n5620_), .B(new_n5494_), .ZN(new_n5621_));
  INV_X1     g05429(.I(new_n5619_), .ZN(new_n5622_));
  OAI21_X1   g05430(.A1(new_n5618_), .A2(new_n5622_), .B(\asqrt[47] ), .ZN(new_n5623_));
  NAND3_X1   g05431(.A1(new_n5621_), .A2(new_n5623_), .A3(new_n1533_), .ZN(new_n5624_));
  NAND2_X1   g05432(.A1(new_n5624_), .A2(new_n5492_), .ZN(new_n5625_));
  NAND2_X1   g05433(.A1(new_n5621_), .A2(new_n5623_), .ZN(new_n5626_));
  AOI21_X1   g05434(.A1(new_n5626_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n5627_));
  AOI21_X1   g05435(.A1(new_n5627_), .A2(new_n5625_), .B(new_n5489_), .ZN(new_n5628_));
  INV_X1     g05436(.I(new_n5494_), .ZN(new_n5629_));
  INV_X1     g05437(.I(new_n5504_), .ZN(new_n5630_));
  NOR2_X1    g05438(.A1(new_n5613_), .A2(new_n5614_), .ZN(new_n5631_));
  AOI21_X1   g05439(.A1(new_n5631_), .A2(new_n2271_), .B(new_n5630_), .ZN(new_n5632_));
  NAND2_X1   g05440(.A1(new_n5615_), .A2(new_n2072_), .ZN(new_n5633_));
  OAI21_X1   g05441(.A1(new_n5632_), .A2(new_n5633_), .B(new_n5500_), .ZN(new_n5634_));
  INV_X1     g05442(.I(new_n5615_), .ZN(new_n5635_));
  OAI21_X1   g05443(.A1(new_n5632_), .A2(new_n5635_), .B(\asqrt[45] ), .ZN(new_n5636_));
  NAND3_X1   g05444(.A1(new_n5634_), .A2(new_n5636_), .A3(new_n1884_), .ZN(new_n5637_));
  NAND2_X1   g05445(.A1(new_n5637_), .A2(new_n5497_), .ZN(new_n5638_));
  NAND2_X1   g05446(.A1(new_n5634_), .A2(new_n5636_), .ZN(new_n5639_));
  AOI21_X1   g05447(.A1(new_n5639_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n5640_));
  AOI21_X1   g05448(.A1(new_n5640_), .A2(new_n5638_), .B(new_n5629_), .ZN(new_n5641_));
  AOI21_X1   g05449(.A1(new_n5638_), .A2(new_n5619_), .B(new_n1688_), .ZN(new_n5642_));
  OAI21_X1   g05450(.A1(new_n5641_), .A2(new_n5642_), .B(\asqrt[48] ), .ZN(new_n5643_));
  AOI21_X1   g05451(.A1(new_n5625_), .A2(new_n5643_), .B(new_n1368_), .ZN(new_n5644_));
  NOR2_X1    g05452(.A1(new_n5628_), .A2(new_n5644_), .ZN(new_n5645_));
  AOI21_X1   g05453(.A1(new_n5645_), .A2(new_n1228_), .B(new_n5486_), .ZN(new_n5646_));
  OAI21_X1   g05454(.A1(new_n5628_), .A2(new_n5644_), .B(\asqrt[50] ), .ZN(new_n5647_));
  NAND2_X1   g05455(.A1(new_n5647_), .A2(new_n1088_), .ZN(new_n5648_));
  OAI21_X1   g05456(.A1(new_n5646_), .A2(new_n5648_), .B(new_n5482_), .ZN(new_n5649_));
  INV_X1     g05457(.I(new_n5647_), .ZN(new_n5650_));
  OAI21_X1   g05458(.A1(new_n5646_), .A2(new_n5650_), .B(\asqrt[51] ), .ZN(new_n5651_));
  NAND3_X1   g05459(.A1(new_n5649_), .A2(new_n5651_), .A3(new_n962_), .ZN(new_n5652_));
  NAND2_X1   g05460(.A1(new_n5652_), .A2(new_n5480_), .ZN(new_n5653_));
  NAND2_X1   g05461(.A1(new_n5649_), .A2(new_n5651_), .ZN(new_n5654_));
  AOI21_X1   g05462(.A1(new_n5654_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n5655_));
  AOI21_X1   g05463(.A1(new_n5655_), .A2(new_n5653_), .B(new_n5477_), .ZN(new_n5656_));
  INV_X1     g05464(.I(new_n5482_), .ZN(new_n5657_));
  INV_X1     g05465(.I(new_n5492_), .ZN(new_n5658_));
  NOR2_X1    g05466(.A1(new_n5641_), .A2(new_n5642_), .ZN(new_n5659_));
  AOI21_X1   g05467(.A1(new_n5659_), .A2(new_n1533_), .B(new_n5658_), .ZN(new_n5660_));
  NAND2_X1   g05468(.A1(new_n5643_), .A2(new_n1368_), .ZN(new_n5661_));
  OAI21_X1   g05469(.A1(new_n5660_), .A2(new_n5661_), .B(new_n5488_), .ZN(new_n5662_));
  INV_X1     g05470(.I(new_n5643_), .ZN(new_n5663_));
  OAI21_X1   g05471(.A1(new_n5660_), .A2(new_n5663_), .B(\asqrt[49] ), .ZN(new_n5664_));
  NAND3_X1   g05472(.A1(new_n5662_), .A2(new_n5664_), .A3(new_n1228_), .ZN(new_n5665_));
  NAND2_X1   g05473(.A1(new_n5665_), .A2(new_n5485_), .ZN(new_n5666_));
  NAND2_X1   g05474(.A1(new_n5662_), .A2(new_n5664_), .ZN(new_n5667_));
  AOI21_X1   g05475(.A1(new_n5667_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n5668_));
  AOI21_X1   g05476(.A1(new_n5668_), .A2(new_n5666_), .B(new_n5657_), .ZN(new_n5669_));
  AOI21_X1   g05477(.A1(new_n5666_), .A2(new_n5647_), .B(new_n1088_), .ZN(new_n5670_));
  OAI21_X1   g05478(.A1(new_n5669_), .A2(new_n5670_), .B(\asqrt[52] ), .ZN(new_n5671_));
  AOI21_X1   g05479(.A1(new_n5653_), .A2(new_n5671_), .B(new_n842_), .ZN(new_n5672_));
  NOR2_X1    g05480(.A1(new_n5656_), .A2(new_n5672_), .ZN(new_n5673_));
  AOI21_X1   g05481(.A1(new_n5673_), .A2(new_n720_), .B(new_n5474_), .ZN(new_n5674_));
  OAI21_X1   g05482(.A1(new_n5656_), .A2(new_n5672_), .B(\asqrt[54] ), .ZN(new_n5675_));
  NAND2_X1   g05483(.A1(new_n5675_), .A2(new_n630_), .ZN(new_n5676_));
  OAI21_X1   g05484(.A1(new_n5674_), .A2(new_n5676_), .B(new_n5470_), .ZN(new_n5677_));
  INV_X1     g05485(.I(new_n5675_), .ZN(new_n5678_));
  OAI21_X1   g05486(.A1(new_n5674_), .A2(new_n5678_), .B(\asqrt[55] ), .ZN(new_n5679_));
  NAND3_X1   g05487(.A1(new_n5677_), .A2(new_n5679_), .A3(new_n545_), .ZN(new_n5680_));
  NAND2_X1   g05488(.A1(new_n5680_), .A2(new_n5468_), .ZN(new_n5681_));
  NAND2_X1   g05489(.A1(new_n5677_), .A2(new_n5679_), .ZN(new_n5682_));
  AOI21_X1   g05490(.A1(new_n5682_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n5683_));
  AOI21_X1   g05491(.A1(new_n5683_), .A2(new_n5681_), .B(new_n5465_), .ZN(new_n5684_));
  INV_X1     g05492(.I(new_n5470_), .ZN(new_n5685_));
  INV_X1     g05493(.I(new_n5480_), .ZN(new_n5686_));
  NOR2_X1    g05494(.A1(new_n5669_), .A2(new_n5670_), .ZN(new_n5687_));
  AOI21_X1   g05495(.A1(new_n5687_), .A2(new_n962_), .B(new_n5686_), .ZN(new_n5688_));
  NAND2_X1   g05496(.A1(new_n5671_), .A2(new_n842_), .ZN(new_n5689_));
  OAI21_X1   g05497(.A1(new_n5688_), .A2(new_n5689_), .B(new_n5476_), .ZN(new_n5690_));
  INV_X1     g05498(.I(new_n5671_), .ZN(new_n5691_));
  OAI21_X1   g05499(.A1(new_n5688_), .A2(new_n5691_), .B(\asqrt[53] ), .ZN(new_n5692_));
  NAND3_X1   g05500(.A1(new_n5690_), .A2(new_n5692_), .A3(new_n720_), .ZN(new_n5693_));
  NAND2_X1   g05501(.A1(new_n5693_), .A2(new_n5473_), .ZN(new_n5694_));
  NAND2_X1   g05502(.A1(new_n5690_), .A2(new_n5692_), .ZN(new_n5695_));
  AOI21_X1   g05503(.A1(new_n5695_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n5696_));
  AOI21_X1   g05504(.A1(new_n5696_), .A2(new_n5694_), .B(new_n5685_), .ZN(new_n5697_));
  AOI21_X1   g05505(.A1(new_n5694_), .A2(new_n5675_), .B(new_n630_), .ZN(new_n5698_));
  OAI21_X1   g05506(.A1(new_n5697_), .A2(new_n5698_), .B(\asqrt[56] ), .ZN(new_n5699_));
  AOI21_X1   g05507(.A1(new_n5681_), .A2(new_n5699_), .B(new_n450_), .ZN(new_n5700_));
  NOR2_X1    g05508(.A1(new_n5684_), .A2(new_n5700_), .ZN(new_n5701_));
  AOI21_X1   g05509(.A1(new_n5701_), .A2(new_n403_), .B(new_n5462_), .ZN(new_n5702_));
  OAI21_X1   g05510(.A1(new_n5684_), .A2(new_n5700_), .B(\asqrt[58] ), .ZN(new_n5703_));
  NAND2_X1   g05511(.A1(new_n5703_), .A2(new_n339_), .ZN(new_n5704_));
  OAI21_X1   g05512(.A1(new_n5702_), .A2(new_n5704_), .B(new_n5458_), .ZN(new_n5705_));
  INV_X1     g05513(.I(new_n5703_), .ZN(new_n5706_));
  OAI21_X1   g05514(.A1(new_n5702_), .A2(new_n5706_), .B(\asqrt[59] ), .ZN(new_n5707_));
  NAND3_X1   g05515(.A1(new_n5705_), .A2(new_n5707_), .A3(new_n288_), .ZN(new_n5708_));
  NAND2_X1   g05516(.A1(new_n5708_), .A2(new_n5456_), .ZN(new_n5709_));
  INV_X1     g05517(.I(new_n5458_), .ZN(new_n5710_));
  INV_X1     g05518(.I(new_n5468_), .ZN(new_n5711_));
  NOR2_X1    g05519(.A1(new_n5697_), .A2(new_n5698_), .ZN(new_n5712_));
  AOI21_X1   g05520(.A1(new_n5712_), .A2(new_n545_), .B(new_n5711_), .ZN(new_n5713_));
  NAND2_X1   g05521(.A1(new_n5699_), .A2(new_n450_), .ZN(new_n5714_));
  OAI21_X1   g05522(.A1(new_n5713_), .A2(new_n5714_), .B(new_n5464_), .ZN(new_n5715_));
  INV_X1     g05523(.I(new_n5699_), .ZN(new_n5716_));
  OAI21_X1   g05524(.A1(new_n5713_), .A2(new_n5716_), .B(\asqrt[57] ), .ZN(new_n5717_));
  NAND3_X1   g05525(.A1(new_n5715_), .A2(new_n5717_), .A3(new_n403_), .ZN(new_n5718_));
  NAND2_X1   g05526(.A1(new_n5718_), .A2(new_n5461_), .ZN(new_n5719_));
  NAND2_X1   g05527(.A1(new_n5715_), .A2(new_n5717_), .ZN(new_n5720_));
  AOI21_X1   g05528(.A1(new_n5720_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n5721_));
  AOI21_X1   g05529(.A1(new_n5721_), .A2(new_n5719_), .B(new_n5710_), .ZN(new_n5722_));
  AOI21_X1   g05530(.A1(new_n5719_), .A2(new_n5703_), .B(new_n339_), .ZN(new_n5723_));
  OAI21_X1   g05531(.A1(new_n5722_), .A2(new_n5723_), .B(\asqrt[60] ), .ZN(new_n5724_));
  AOI21_X1   g05532(.A1(new_n5709_), .A2(new_n5724_), .B(new_n242_), .ZN(new_n5725_));
  NAND3_X1   g05533(.A1(\asqrt[32] ), .A2(new_n5380_), .A3(new_n5396_), .ZN(new_n5726_));
  XOR2_X1    g05534(.A1(new_n5726_), .A2(new_n5422_), .Z(new_n5727_));
  INV_X1     g05535(.I(new_n5727_), .ZN(new_n5728_));
  NAND2_X1   g05536(.A1(new_n5705_), .A2(new_n5707_), .ZN(new_n5729_));
  AOI21_X1   g05537(.A1(new_n5729_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n5730_));
  AOI21_X1   g05538(.A1(new_n5730_), .A2(new_n5709_), .B(new_n5728_), .ZN(new_n5731_));
  OAI21_X1   g05539(.A1(new_n5731_), .A2(new_n5725_), .B(\asqrt[62] ), .ZN(new_n5732_));
  AOI21_X1   g05540(.A1(new_n5381_), .A2(new_n5402_), .B(new_n5397_), .ZN(new_n5733_));
  NAND2_X1   g05541(.A1(\asqrt[32] ), .A2(new_n5733_), .ZN(new_n5734_));
  XOR2_X1    g05542(.A1(new_n5734_), .A2(new_n5400_), .Z(new_n5735_));
  INV_X1     g05543(.I(new_n5456_), .ZN(new_n5736_));
  NOR2_X1    g05544(.A1(new_n5722_), .A2(new_n5723_), .ZN(new_n5737_));
  AOI21_X1   g05545(.A1(new_n5737_), .A2(new_n288_), .B(new_n5736_), .ZN(new_n5738_));
  INV_X1     g05546(.I(new_n5724_), .ZN(new_n5739_));
  OAI21_X1   g05547(.A1(new_n5738_), .A2(new_n5739_), .B(\asqrt[61] ), .ZN(new_n5740_));
  NAND2_X1   g05548(.A1(new_n5724_), .A2(new_n242_), .ZN(new_n5741_));
  OAI21_X1   g05549(.A1(new_n5738_), .A2(new_n5741_), .B(new_n5727_), .ZN(new_n5742_));
  NAND3_X1   g05550(.A1(new_n5742_), .A2(new_n5740_), .A3(new_n234_), .ZN(new_n5743_));
  NAND2_X1   g05551(.A1(new_n5743_), .A2(new_n5735_), .ZN(new_n5744_));
  AOI21_X1   g05552(.A1(new_n5744_), .A2(new_n5732_), .B(new_n5453_), .ZN(new_n5745_));
  AOI21_X1   g05553(.A1(new_n5745_), .A2(new_n5451_), .B(\asqrt[63] ), .ZN(new_n5746_));
  NAND2_X1   g05554(.A1(new_n5744_), .A2(new_n5732_), .ZN(new_n5747_));
  NOR2_X1    g05555(.A1(new_n5747_), .A2(new_n5451_), .ZN(new_n5748_));
  NOR2_X1    g05556(.A1(\asqrt[32] ), .A2(new_n5420_), .ZN(new_n5749_));
  NOR4_X1    g05557(.A1(new_n5746_), .A2(new_n5448_), .A3(new_n5748_), .A4(new_n5749_), .ZN(new_n5750_));
  NOR3_X1    g05558(.A1(new_n5750_), .A2(new_n5442_), .A3(new_n5444_), .ZN(new_n5751_));
  XOR2_X1    g05559(.A1(new_n5751_), .A2(new_n5437_), .Z(new_n5752_));
  INV_X1     g05560(.I(new_n5752_), .ZN(new_n5753_));
  INV_X1     g05561(.I(new_n5448_), .ZN(new_n5754_));
  INV_X1     g05562(.I(new_n5732_), .ZN(new_n5755_));
  NOR2_X1    g05563(.A1(new_n5731_), .A2(new_n5725_), .ZN(new_n5756_));
  INV_X1     g05564(.I(new_n5735_), .ZN(new_n5757_));
  AOI21_X1   g05565(.A1(new_n5756_), .A2(new_n234_), .B(new_n5757_), .ZN(new_n5758_));
  OAI21_X1   g05566(.A1(new_n5758_), .A2(new_n5755_), .B(new_n5452_), .ZN(new_n5759_));
  OAI21_X1   g05567(.A1(new_n5759_), .A2(new_n5450_), .B(new_n193_), .ZN(new_n5760_));
  NOR2_X1    g05568(.A1(new_n5758_), .A2(new_n5755_), .ZN(new_n5761_));
  NAND2_X1   g05569(.A1(new_n5761_), .A2(new_n5450_), .ZN(new_n5762_));
  INV_X1     g05570(.I(new_n5749_), .ZN(new_n5763_));
  NAND4_X1   g05571(.A1(new_n5760_), .A2(new_n5754_), .A3(new_n5762_), .A4(new_n5763_), .ZN(\asqrt[31] ));
  NAND3_X1   g05572(.A1(\asqrt[31] ), .A2(new_n5438_), .A3(new_n5439_), .ZN(new_n5765_));
  NAND4_X1   g05573(.A1(new_n5760_), .A2(\asqrt[32] ), .A3(new_n5762_), .A4(new_n5754_), .ZN(new_n5766_));
  AOI21_X1   g05574(.A1(new_n5765_), .A2(new_n5766_), .B(\a[64] ), .ZN(new_n5767_));
  NOR3_X1    g05575(.A1(new_n5750_), .A2(\a[62] ), .A3(\a[63] ), .ZN(new_n5768_));
  INV_X1     g05576(.I(new_n5766_), .ZN(new_n5769_));
  NOR3_X1    g05577(.A1(new_n5768_), .A2(new_n195_), .A3(new_n5769_), .ZN(new_n5770_));
  NOR2_X1    g05578(.A1(new_n5770_), .A2(new_n5767_), .ZN(new_n5771_));
  INV_X1     g05579(.I(\a[60] ), .ZN(new_n5772_));
  INV_X1     g05580(.I(\a[61] ), .ZN(new_n5773_));
  NAND3_X1   g05581(.A1(new_n5772_), .A2(new_n5773_), .A3(new_n5438_), .ZN(new_n5774_));
  OAI21_X1   g05582(.A1(new_n5750_), .A2(new_n5438_), .B(new_n5774_), .ZN(new_n5775_));
  NAND2_X1   g05583(.A1(new_n5775_), .A2(\asqrt[32] ), .ZN(new_n5776_));
  OAI21_X1   g05584(.A1(new_n5750_), .A2(\a[62] ), .B(\a[63] ), .ZN(new_n5777_));
  NAND2_X1   g05585(.A1(new_n5777_), .A2(new_n5765_), .ZN(new_n5778_));
  NOR2_X1    g05586(.A1(new_n5775_), .A2(\asqrt[32] ), .ZN(new_n5779_));
  OAI21_X1   g05587(.A1(new_n5778_), .A2(new_n5779_), .B(new_n5776_), .ZN(new_n5780_));
  OAI21_X1   g05588(.A1(new_n5780_), .A2(\asqrt[33] ), .B(new_n5771_), .ZN(new_n5781_));
  NAND2_X1   g05589(.A1(new_n5780_), .A2(\asqrt[33] ), .ZN(new_n5782_));
  NAND3_X1   g05590(.A1(new_n5781_), .A2(new_n4810_), .A3(new_n5782_), .ZN(new_n5783_));
  OAI21_X1   g05591(.A1(new_n5768_), .A2(new_n5769_), .B(new_n195_), .ZN(new_n5784_));
  NAND3_X1   g05592(.A1(new_n5765_), .A2(\a[64] ), .A3(new_n5766_), .ZN(new_n5785_));
  NAND2_X1   g05593(.A1(new_n5784_), .A2(new_n5785_), .ZN(new_n5786_));
  NAND2_X1   g05594(.A1(\asqrt[31] ), .A2(\a[62] ), .ZN(new_n5787_));
  AOI21_X1   g05595(.A1(new_n5787_), .A2(new_n5774_), .B(new_n5435_), .ZN(new_n5788_));
  AOI21_X1   g05596(.A1(\asqrt[31] ), .A2(new_n5438_), .B(new_n5439_), .ZN(new_n5789_));
  NOR2_X1    g05597(.A1(new_n5768_), .A2(new_n5789_), .ZN(new_n5790_));
  NAND3_X1   g05598(.A1(new_n5787_), .A2(new_n5435_), .A3(new_n5774_), .ZN(new_n5791_));
  AOI21_X1   g05599(.A1(new_n5790_), .A2(new_n5791_), .B(new_n5788_), .ZN(new_n5792_));
  AOI21_X1   g05600(.A1(new_n5792_), .A2(new_n5110_), .B(new_n5786_), .ZN(new_n5793_));
  NOR2_X1    g05601(.A1(new_n5792_), .A2(new_n5110_), .ZN(new_n5794_));
  OAI21_X1   g05602(.A1(new_n5793_), .A2(new_n5794_), .B(\asqrt[34] ), .ZN(new_n5795_));
  NAND2_X1   g05603(.A1(new_n5747_), .A2(new_n5450_), .ZN(new_n5796_));
  NOR2_X1    g05604(.A1(new_n5750_), .A2(new_n5450_), .ZN(new_n5797_));
  NAND2_X1   g05605(.A1(new_n5797_), .A2(new_n5761_), .ZN(new_n5798_));
  AOI21_X1   g05606(.A1(new_n5798_), .A2(new_n5796_), .B(new_n193_), .ZN(new_n5799_));
  INV_X1     g05607(.I(new_n5799_), .ZN(new_n5800_));
  NAND3_X1   g05608(.A1(\asqrt[31] ), .A2(new_n5732_), .A3(new_n5743_), .ZN(new_n5801_));
  XOR2_X1    g05609(.A1(new_n5801_), .A2(new_n5735_), .Z(new_n5802_));
  AOI21_X1   g05610(.A1(new_n5797_), .A2(new_n5747_), .B(new_n5748_), .ZN(new_n5803_));
  OAI21_X1   g05611(.A1(new_n5702_), .A2(new_n5704_), .B(new_n5707_), .ZN(new_n5804_));
  NOR2_X1    g05612(.A1(new_n5750_), .A2(new_n5804_), .ZN(new_n5805_));
  XOR2_X1    g05613(.A1(new_n5805_), .A2(new_n5458_), .Z(new_n5806_));
  NAND3_X1   g05614(.A1(\asqrt[31] ), .A2(new_n5718_), .A3(new_n5703_), .ZN(new_n5807_));
  XOR2_X1    g05615(.A1(new_n5807_), .A2(new_n5462_), .Z(new_n5808_));
  OAI21_X1   g05616(.A1(new_n5713_), .A2(new_n5714_), .B(new_n5717_), .ZN(new_n5809_));
  NOR2_X1    g05617(.A1(new_n5750_), .A2(new_n5809_), .ZN(new_n5810_));
  XOR2_X1    g05618(.A1(new_n5810_), .A2(new_n5464_), .Z(new_n5811_));
  INV_X1     g05619(.I(new_n5811_), .ZN(new_n5812_));
  NAND3_X1   g05620(.A1(\asqrt[31] ), .A2(new_n5680_), .A3(new_n5699_), .ZN(new_n5813_));
  XOR2_X1    g05621(.A1(new_n5813_), .A2(new_n5711_), .Z(new_n5814_));
  INV_X1     g05622(.I(new_n5814_), .ZN(new_n5815_));
  OAI21_X1   g05623(.A1(new_n5674_), .A2(new_n5676_), .B(new_n5679_), .ZN(new_n5816_));
  NOR2_X1    g05624(.A1(new_n5750_), .A2(new_n5816_), .ZN(new_n5817_));
  XOR2_X1    g05625(.A1(new_n5817_), .A2(new_n5470_), .Z(new_n5818_));
  NAND3_X1   g05626(.A1(\asqrt[31] ), .A2(new_n5693_), .A3(new_n5675_), .ZN(new_n5819_));
  XOR2_X1    g05627(.A1(new_n5819_), .A2(new_n5474_), .Z(new_n5820_));
  OAI21_X1   g05628(.A1(new_n5688_), .A2(new_n5689_), .B(new_n5692_), .ZN(new_n5821_));
  NOR2_X1    g05629(.A1(new_n5750_), .A2(new_n5821_), .ZN(new_n5822_));
  XOR2_X1    g05630(.A1(new_n5822_), .A2(new_n5476_), .Z(new_n5823_));
  INV_X1     g05631(.I(new_n5823_), .ZN(new_n5824_));
  NAND3_X1   g05632(.A1(\asqrt[31] ), .A2(new_n5652_), .A3(new_n5671_), .ZN(new_n5825_));
  XOR2_X1    g05633(.A1(new_n5825_), .A2(new_n5686_), .Z(new_n5826_));
  INV_X1     g05634(.I(new_n5826_), .ZN(new_n5827_));
  OAI21_X1   g05635(.A1(new_n5646_), .A2(new_n5648_), .B(new_n5651_), .ZN(new_n5828_));
  NOR2_X1    g05636(.A1(new_n5750_), .A2(new_n5828_), .ZN(new_n5829_));
  XOR2_X1    g05637(.A1(new_n5829_), .A2(new_n5482_), .Z(new_n5830_));
  NAND3_X1   g05638(.A1(\asqrt[31] ), .A2(new_n5665_), .A3(new_n5647_), .ZN(new_n5831_));
  XOR2_X1    g05639(.A1(new_n5831_), .A2(new_n5486_), .Z(new_n5832_));
  OAI21_X1   g05640(.A1(new_n5660_), .A2(new_n5661_), .B(new_n5664_), .ZN(new_n5833_));
  NOR2_X1    g05641(.A1(new_n5750_), .A2(new_n5833_), .ZN(new_n5834_));
  XOR2_X1    g05642(.A1(new_n5834_), .A2(new_n5488_), .Z(new_n5835_));
  INV_X1     g05643(.I(new_n5835_), .ZN(new_n5836_));
  NAND3_X1   g05644(.A1(\asqrt[31] ), .A2(new_n5624_), .A3(new_n5643_), .ZN(new_n5837_));
  XOR2_X1    g05645(.A1(new_n5837_), .A2(new_n5658_), .Z(new_n5838_));
  INV_X1     g05646(.I(new_n5838_), .ZN(new_n5839_));
  OAI21_X1   g05647(.A1(new_n5618_), .A2(new_n5620_), .B(new_n5623_), .ZN(new_n5840_));
  NOR2_X1    g05648(.A1(new_n5750_), .A2(new_n5840_), .ZN(new_n5841_));
  XOR2_X1    g05649(.A1(new_n5841_), .A2(new_n5494_), .Z(new_n5842_));
  NAND3_X1   g05650(.A1(\asqrt[31] ), .A2(new_n5637_), .A3(new_n5619_), .ZN(new_n5843_));
  XOR2_X1    g05651(.A1(new_n5843_), .A2(new_n5498_), .Z(new_n5844_));
  OAI21_X1   g05652(.A1(new_n5632_), .A2(new_n5633_), .B(new_n5636_), .ZN(new_n5845_));
  NOR2_X1    g05653(.A1(new_n5750_), .A2(new_n5845_), .ZN(new_n5846_));
  XOR2_X1    g05654(.A1(new_n5846_), .A2(new_n5500_), .Z(new_n5847_));
  INV_X1     g05655(.I(new_n5847_), .ZN(new_n5848_));
  NAND3_X1   g05656(.A1(\asqrt[31] ), .A2(new_n5596_), .A3(new_n5615_), .ZN(new_n5849_));
  XOR2_X1    g05657(.A1(new_n5849_), .A2(new_n5630_), .Z(new_n5850_));
  INV_X1     g05658(.I(new_n5850_), .ZN(new_n5851_));
  OAI21_X1   g05659(.A1(new_n5590_), .A2(new_n5592_), .B(new_n5595_), .ZN(new_n5852_));
  NOR2_X1    g05660(.A1(new_n5750_), .A2(new_n5852_), .ZN(new_n5853_));
  XOR2_X1    g05661(.A1(new_n5853_), .A2(new_n5506_), .Z(new_n5854_));
  NAND3_X1   g05662(.A1(\asqrt[31] ), .A2(new_n5609_), .A3(new_n5591_), .ZN(new_n5855_));
  XOR2_X1    g05663(.A1(new_n5855_), .A2(new_n5510_), .Z(new_n5856_));
  OAI21_X1   g05664(.A1(new_n5604_), .A2(new_n5605_), .B(new_n5608_), .ZN(new_n5857_));
  NOR2_X1    g05665(.A1(new_n5750_), .A2(new_n5857_), .ZN(new_n5858_));
  XOR2_X1    g05666(.A1(new_n5858_), .A2(new_n5512_), .Z(new_n5859_));
  INV_X1     g05667(.I(new_n5859_), .ZN(new_n5860_));
  NAND3_X1   g05668(.A1(\asqrt[31] ), .A2(new_n5557_), .A3(new_n5587_), .ZN(new_n5861_));
  XOR2_X1    g05669(.A1(new_n5861_), .A2(new_n5602_), .Z(new_n5862_));
  INV_X1     g05670(.I(new_n5862_), .ZN(new_n5863_));
  OAI21_X1   g05671(.A1(new_n5551_), .A2(new_n5553_), .B(new_n5556_), .ZN(new_n5864_));
  NOR2_X1    g05672(.A1(new_n5750_), .A2(new_n5864_), .ZN(new_n5865_));
  XOR2_X1    g05673(.A1(new_n5865_), .A2(new_n5518_), .Z(new_n5866_));
  NAND3_X1   g05674(.A1(\asqrt[31] ), .A2(new_n5581_), .A3(new_n5552_), .ZN(new_n5867_));
  XOR2_X1    g05675(.A1(new_n5867_), .A2(new_n5522_), .Z(new_n5868_));
  AOI21_X1   g05676(.A1(new_n5545_), .A2(new_n5546_), .B(new_n5549_), .ZN(new_n5869_));
  NAND2_X1   g05677(.A1(\asqrt[31] ), .A2(new_n5869_), .ZN(new_n5870_));
  XOR2_X1    g05678(.A1(new_n5870_), .A2(new_n5525_), .Z(new_n5871_));
  INV_X1     g05679(.I(new_n5871_), .ZN(new_n5872_));
  NOR2_X1    g05680(.A1(new_n5544_), .A2(\asqrt[36] ), .ZN(new_n5873_));
  NOR3_X1    g05681(.A1(new_n5750_), .A2(new_n5873_), .A3(new_n5579_), .ZN(new_n5874_));
  XOR2_X1    g05682(.A1(new_n5874_), .A2(new_n5528_), .Z(new_n5875_));
  INV_X1     g05683(.I(new_n5875_), .ZN(new_n5876_));
  NOR3_X1    g05684(.A1(new_n5750_), .A2(new_n5539_), .A3(new_n5574_), .ZN(new_n5877_));
  XOR2_X1    g05685(.A1(new_n5877_), .A2(new_n5541_), .Z(new_n5878_));
  NOR2_X1    g05686(.A1(new_n5570_), .A2(\asqrt[34] ), .ZN(new_n5879_));
  NOR3_X1    g05687(.A1(new_n5750_), .A2(new_n5879_), .A3(new_n5538_), .ZN(new_n5880_));
  XOR2_X1    g05688(.A1(new_n5880_), .A2(new_n5566_), .Z(new_n5881_));
  NOR2_X1    g05689(.A1(new_n5793_), .A2(new_n5794_), .ZN(new_n5882_));
  AOI21_X1   g05690(.A1(new_n5882_), .A2(new_n4810_), .B(new_n5753_), .ZN(new_n5883_));
  NAND2_X1   g05691(.A1(new_n5795_), .A2(new_n4510_), .ZN(new_n5884_));
  OAI21_X1   g05692(.A1(new_n5883_), .A2(new_n5884_), .B(new_n5881_), .ZN(new_n5885_));
  INV_X1     g05693(.I(new_n5795_), .ZN(new_n5886_));
  OAI21_X1   g05694(.A1(new_n5883_), .A2(new_n5886_), .B(\asqrt[35] ), .ZN(new_n5887_));
  NAND3_X1   g05695(.A1(new_n5885_), .A2(new_n5887_), .A3(new_n4224_), .ZN(new_n5888_));
  NAND2_X1   g05696(.A1(new_n5888_), .A2(new_n5878_), .ZN(new_n5889_));
  NAND2_X1   g05697(.A1(new_n5885_), .A2(new_n5887_), .ZN(new_n5890_));
  AOI21_X1   g05698(.A1(new_n5890_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n5891_));
  AOI21_X1   g05699(.A1(new_n5891_), .A2(new_n5889_), .B(new_n5876_), .ZN(new_n5892_));
  INV_X1     g05700(.I(new_n5881_), .ZN(new_n5893_));
  NAND2_X1   g05701(.A1(new_n5783_), .A2(new_n5752_), .ZN(new_n5894_));
  NAND2_X1   g05702(.A1(new_n5781_), .A2(new_n5782_), .ZN(new_n5895_));
  AOI21_X1   g05703(.A1(new_n5895_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n5896_));
  AOI21_X1   g05704(.A1(new_n5896_), .A2(new_n5894_), .B(new_n5893_), .ZN(new_n5897_));
  AOI21_X1   g05705(.A1(new_n5894_), .A2(new_n5795_), .B(new_n4510_), .ZN(new_n5898_));
  OAI21_X1   g05706(.A1(new_n5897_), .A2(new_n5898_), .B(\asqrt[36] ), .ZN(new_n5899_));
  AOI21_X1   g05707(.A1(new_n5889_), .A2(new_n5899_), .B(new_n3928_), .ZN(new_n5900_));
  NOR2_X1    g05708(.A1(new_n5892_), .A2(new_n5900_), .ZN(new_n5901_));
  AOI21_X1   g05709(.A1(new_n5901_), .A2(new_n3675_), .B(new_n5872_), .ZN(new_n5902_));
  OAI21_X1   g05710(.A1(new_n5892_), .A2(new_n5900_), .B(\asqrt[38] ), .ZN(new_n5903_));
  NAND2_X1   g05711(.A1(new_n5903_), .A2(new_n3400_), .ZN(new_n5904_));
  OAI21_X1   g05712(.A1(new_n5902_), .A2(new_n5904_), .B(new_n5868_), .ZN(new_n5905_));
  INV_X1     g05713(.I(new_n5903_), .ZN(new_n5906_));
  OAI21_X1   g05714(.A1(new_n5902_), .A2(new_n5906_), .B(\asqrt[39] ), .ZN(new_n5907_));
  NAND3_X1   g05715(.A1(new_n5905_), .A2(new_n5907_), .A3(new_n3167_), .ZN(new_n5908_));
  NAND2_X1   g05716(.A1(new_n5908_), .A2(new_n5866_), .ZN(new_n5909_));
  NAND2_X1   g05717(.A1(new_n5905_), .A2(new_n5907_), .ZN(new_n5910_));
  AOI21_X1   g05718(.A1(new_n5910_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n5911_));
  AOI21_X1   g05719(.A1(new_n5911_), .A2(new_n5909_), .B(new_n5863_), .ZN(new_n5912_));
  INV_X1     g05720(.I(new_n5868_), .ZN(new_n5913_));
  INV_X1     g05721(.I(new_n5878_), .ZN(new_n5914_));
  NOR2_X1    g05722(.A1(new_n5897_), .A2(new_n5898_), .ZN(new_n5915_));
  AOI21_X1   g05723(.A1(new_n5915_), .A2(new_n4224_), .B(new_n5914_), .ZN(new_n5916_));
  NAND2_X1   g05724(.A1(new_n5899_), .A2(new_n3928_), .ZN(new_n5917_));
  OAI21_X1   g05725(.A1(new_n5916_), .A2(new_n5917_), .B(new_n5875_), .ZN(new_n5918_));
  INV_X1     g05726(.I(new_n5899_), .ZN(new_n5919_));
  OAI21_X1   g05727(.A1(new_n5916_), .A2(new_n5919_), .B(\asqrt[37] ), .ZN(new_n5920_));
  NAND3_X1   g05728(.A1(new_n5918_), .A2(new_n5920_), .A3(new_n3675_), .ZN(new_n5921_));
  NAND2_X1   g05729(.A1(new_n5921_), .A2(new_n5871_), .ZN(new_n5922_));
  NAND2_X1   g05730(.A1(new_n5918_), .A2(new_n5920_), .ZN(new_n5923_));
  AOI21_X1   g05731(.A1(new_n5923_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n5924_));
  AOI21_X1   g05732(.A1(new_n5924_), .A2(new_n5922_), .B(new_n5913_), .ZN(new_n5925_));
  AOI21_X1   g05733(.A1(new_n5922_), .A2(new_n5903_), .B(new_n3400_), .ZN(new_n5926_));
  OAI21_X1   g05734(.A1(new_n5925_), .A2(new_n5926_), .B(\asqrt[40] ), .ZN(new_n5927_));
  AOI21_X1   g05735(.A1(new_n5909_), .A2(new_n5927_), .B(new_n2912_), .ZN(new_n5928_));
  NOR2_X1    g05736(.A1(new_n5912_), .A2(new_n5928_), .ZN(new_n5929_));
  AOI21_X1   g05737(.A1(new_n5929_), .A2(new_n2699_), .B(new_n5860_), .ZN(new_n5930_));
  OAI21_X1   g05738(.A1(new_n5912_), .A2(new_n5928_), .B(\asqrt[42] ), .ZN(new_n5931_));
  NAND2_X1   g05739(.A1(new_n5931_), .A2(new_n2464_), .ZN(new_n5932_));
  OAI21_X1   g05740(.A1(new_n5930_), .A2(new_n5932_), .B(new_n5856_), .ZN(new_n5933_));
  INV_X1     g05741(.I(new_n5931_), .ZN(new_n5934_));
  OAI21_X1   g05742(.A1(new_n5930_), .A2(new_n5934_), .B(\asqrt[43] ), .ZN(new_n5935_));
  NAND3_X1   g05743(.A1(new_n5933_), .A2(new_n5935_), .A3(new_n2271_), .ZN(new_n5936_));
  NAND2_X1   g05744(.A1(new_n5936_), .A2(new_n5854_), .ZN(new_n5937_));
  NAND2_X1   g05745(.A1(new_n5933_), .A2(new_n5935_), .ZN(new_n5938_));
  AOI21_X1   g05746(.A1(new_n5938_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n5939_));
  AOI21_X1   g05747(.A1(new_n5939_), .A2(new_n5937_), .B(new_n5851_), .ZN(new_n5940_));
  INV_X1     g05748(.I(new_n5856_), .ZN(new_n5941_));
  INV_X1     g05749(.I(new_n5866_), .ZN(new_n5942_));
  NOR2_X1    g05750(.A1(new_n5925_), .A2(new_n5926_), .ZN(new_n5943_));
  AOI21_X1   g05751(.A1(new_n5943_), .A2(new_n3167_), .B(new_n5942_), .ZN(new_n5944_));
  NAND2_X1   g05752(.A1(new_n5927_), .A2(new_n2912_), .ZN(new_n5945_));
  OAI21_X1   g05753(.A1(new_n5944_), .A2(new_n5945_), .B(new_n5862_), .ZN(new_n5946_));
  INV_X1     g05754(.I(new_n5927_), .ZN(new_n5947_));
  OAI21_X1   g05755(.A1(new_n5944_), .A2(new_n5947_), .B(\asqrt[41] ), .ZN(new_n5948_));
  NAND3_X1   g05756(.A1(new_n5946_), .A2(new_n5948_), .A3(new_n2699_), .ZN(new_n5949_));
  NAND2_X1   g05757(.A1(new_n5949_), .A2(new_n5859_), .ZN(new_n5950_));
  NAND2_X1   g05758(.A1(new_n5946_), .A2(new_n5948_), .ZN(new_n5951_));
  AOI21_X1   g05759(.A1(new_n5951_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n5952_));
  AOI21_X1   g05760(.A1(new_n5952_), .A2(new_n5950_), .B(new_n5941_), .ZN(new_n5953_));
  AOI21_X1   g05761(.A1(new_n5950_), .A2(new_n5931_), .B(new_n2464_), .ZN(new_n5954_));
  OAI21_X1   g05762(.A1(new_n5953_), .A2(new_n5954_), .B(\asqrt[44] ), .ZN(new_n5955_));
  AOI21_X1   g05763(.A1(new_n5937_), .A2(new_n5955_), .B(new_n2072_), .ZN(new_n5956_));
  NOR2_X1    g05764(.A1(new_n5940_), .A2(new_n5956_), .ZN(new_n5957_));
  AOI21_X1   g05765(.A1(new_n5957_), .A2(new_n1884_), .B(new_n5848_), .ZN(new_n5958_));
  OAI21_X1   g05766(.A1(new_n5940_), .A2(new_n5956_), .B(\asqrt[46] ), .ZN(new_n5959_));
  NAND2_X1   g05767(.A1(new_n5959_), .A2(new_n1688_), .ZN(new_n5960_));
  OAI21_X1   g05768(.A1(new_n5958_), .A2(new_n5960_), .B(new_n5844_), .ZN(new_n5961_));
  INV_X1     g05769(.I(new_n5959_), .ZN(new_n5962_));
  OAI21_X1   g05770(.A1(new_n5958_), .A2(new_n5962_), .B(\asqrt[47] ), .ZN(new_n5963_));
  NAND3_X1   g05771(.A1(new_n5961_), .A2(new_n5963_), .A3(new_n1533_), .ZN(new_n5964_));
  NAND2_X1   g05772(.A1(new_n5964_), .A2(new_n5842_), .ZN(new_n5965_));
  NAND2_X1   g05773(.A1(new_n5961_), .A2(new_n5963_), .ZN(new_n5966_));
  AOI21_X1   g05774(.A1(new_n5966_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n5967_));
  AOI21_X1   g05775(.A1(new_n5967_), .A2(new_n5965_), .B(new_n5839_), .ZN(new_n5968_));
  INV_X1     g05776(.I(new_n5844_), .ZN(new_n5969_));
  INV_X1     g05777(.I(new_n5854_), .ZN(new_n5970_));
  NOR2_X1    g05778(.A1(new_n5953_), .A2(new_n5954_), .ZN(new_n5971_));
  AOI21_X1   g05779(.A1(new_n5971_), .A2(new_n2271_), .B(new_n5970_), .ZN(new_n5972_));
  NAND2_X1   g05780(.A1(new_n5955_), .A2(new_n2072_), .ZN(new_n5973_));
  OAI21_X1   g05781(.A1(new_n5972_), .A2(new_n5973_), .B(new_n5850_), .ZN(new_n5974_));
  INV_X1     g05782(.I(new_n5955_), .ZN(new_n5975_));
  OAI21_X1   g05783(.A1(new_n5972_), .A2(new_n5975_), .B(\asqrt[45] ), .ZN(new_n5976_));
  NAND3_X1   g05784(.A1(new_n5974_), .A2(new_n5976_), .A3(new_n1884_), .ZN(new_n5977_));
  NAND2_X1   g05785(.A1(new_n5977_), .A2(new_n5847_), .ZN(new_n5978_));
  NAND2_X1   g05786(.A1(new_n5974_), .A2(new_n5976_), .ZN(new_n5979_));
  AOI21_X1   g05787(.A1(new_n5979_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n5980_));
  AOI21_X1   g05788(.A1(new_n5980_), .A2(new_n5978_), .B(new_n5969_), .ZN(new_n5981_));
  AOI21_X1   g05789(.A1(new_n5978_), .A2(new_n5959_), .B(new_n1688_), .ZN(new_n5982_));
  OAI21_X1   g05790(.A1(new_n5981_), .A2(new_n5982_), .B(\asqrt[48] ), .ZN(new_n5983_));
  AOI21_X1   g05791(.A1(new_n5965_), .A2(new_n5983_), .B(new_n1368_), .ZN(new_n5984_));
  NOR2_X1    g05792(.A1(new_n5968_), .A2(new_n5984_), .ZN(new_n5985_));
  AOI21_X1   g05793(.A1(new_n5985_), .A2(new_n1228_), .B(new_n5836_), .ZN(new_n5986_));
  OAI21_X1   g05794(.A1(new_n5968_), .A2(new_n5984_), .B(\asqrt[50] ), .ZN(new_n5987_));
  NAND2_X1   g05795(.A1(new_n5987_), .A2(new_n1088_), .ZN(new_n5988_));
  OAI21_X1   g05796(.A1(new_n5986_), .A2(new_n5988_), .B(new_n5832_), .ZN(new_n5989_));
  INV_X1     g05797(.I(new_n5987_), .ZN(new_n5990_));
  OAI21_X1   g05798(.A1(new_n5986_), .A2(new_n5990_), .B(\asqrt[51] ), .ZN(new_n5991_));
  NAND3_X1   g05799(.A1(new_n5989_), .A2(new_n5991_), .A3(new_n962_), .ZN(new_n5992_));
  NAND2_X1   g05800(.A1(new_n5992_), .A2(new_n5830_), .ZN(new_n5993_));
  NAND2_X1   g05801(.A1(new_n5989_), .A2(new_n5991_), .ZN(new_n5994_));
  AOI21_X1   g05802(.A1(new_n5994_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n5995_));
  AOI21_X1   g05803(.A1(new_n5995_), .A2(new_n5993_), .B(new_n5827_), .ZN(new_n5996_));
  INV_X1     g05804(.I(new_n5832_), .ZN(new_n5997_));
  INV_X1     g05805(.I(new_n5842_), .ZN(new_n5998_));
  NOR2_X1    g05806(.A1(new_n5981_), .A2(new_n5982_), .ZN(new_n5999_));
  AOI21_X1   g05807(.A1(new_n5999_), .A2(new_n1533_), .B(new_n5998_), .ZN(new_n6000_));
  NAND2_X1   g05808(.A1(new_n5983_), .A2(new_n1368_), .ZN(new_n6001_));
  OAI21_X1   g05809(.A1(new_n6000_), .A2(new_n6001_), .B(new_n5838_), .ZN(new_n6002_));
  INV_X1     g05810(.I(new_n5983_), .ZN(new_n6003_));
  OAI21_X1   g05811(.A1(new_n6000_), .A2(new_n6003_), .B(\asqrt[49] ), .ZN(new_n6004_));
  NAND3_X1   g05812(.A1(new_n6002_), .A2(new_n6004_), .A3(new_n1228_), .ZN(new_n6005_));
  NAND2_X1   g05813(.A1(new_n6005_), .A2(new_n5835_), .ZN(new_n6006_));
  NAND2_X1   g05814(.A1(new_n6002_), .A2(new_n6004_), .ZN(new_n6007_));
  AOI21_X1   g05815(.A1(new_n6007_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n6008_));
  AOI21_X1   g05816(.A1(new_n6008_), .A2(new_n6006_), .B(new_n5997_), .ZN(new_n6009_));
  AOI21_X1   g05817(.A1(new_n6006_), .A2(new_n5987_), .B(new_n1088_), .ZN(new_n6010_));
  OAI21_X1   g05818(.A1(new_n6009_), .A2(new_n6010_), .B(\asqrt[52] ), .ZN(new_n6011_));
  AOI21_X1   g05819(.A1(new_n5993_), .A2(new_n6011_), .B(new_n842_), .ZN(new_n6012_));
  NOR2_X1    g05820(.A1(new_n5996_), .A2(new_n6012_), .ZN(new_n6013_));
  AOI21_X1   g05821(.A1(new_n6013_), .A2(new_n720_), .B(new_n5824_), .ZN(new_n6014_));
  OAI21_X1   g05822(.A1(new_n5996_), .A2(new_n6012_), .B(\asqrt[54] ), .ZN(new_n6015_));
  NAND2_X1   g05823(.A1(new_n6015_), .A2(new_n630_), .ZN(new_n6016_));
  OAI21_X1   g05824(.A1(new_n6014_), .A2(new_n6016_), .B(new_n5820_), .ZN(new_n6017_));
  INV_X1     g05825(.I(new_n6015_), .ZN(new_n6018_));
  OAI21_X1   g05826(.A1(new_n6014_), .A2(new_n6018_), .B(\asqrt[55] ), .ZN(new_n6019_));
  NAND3_X1   g05827(.A1(new_n6017_), .A2(new_n6019_), .A3(new_n545_), .ZN(new_n6020_));
  NAND2_X1   g05828(.A1(new_n6020_), .A2(new_n5818_), .ZN(new_n6021_));
  NAND2_X1   g05829(.A1(new_n6017_), .A2(new_n6019_), .ZN(new_n6022_));
  AOI21_X1   g05830(.A1(new_n6022_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n6023_));
  AOI21_X1   g05831(.A1(new_n6023_), .A2(new_n6021_), .B(new_n5815_), .ZN(new_n6024_));
  INV_X1     g05832(.I(new_n5820_), .ZN(new_n6025_));
  INV_X1     g05833(.I(new_n5830_), .ZN(new_n6026_));
  NOR2_X1    g05834(.A1(new_n6009_), .A2(new_n6010_), .ZN(new_n6027_));
  AOI21_X1   g05835(.A1(new_n6027_), .A2(new_n962_), .B(new_n6026_), .ZN(new_n6028_));
  NAND2_X1   g05836(.A1(new_n6011_), .A2(new_n842_), .ZN(new_n6029_));
  OAI21_X1   g05837(.A1(new_n6028_), .A2(new_n6029_), .B(new_n5826_), .ZN(new_n6030_));
  INV_X1     g05838(.I(new_n6011_), .ZN(new_n6031_));
  OAI21_X1   g05839(.A1(new_n6028_), .A2(new_n6031_), .B(\asqrt[53] ), .ZN(new_n6032_));
  NAND3_X1   g05840(.A1(new_n6030_), .A2(new_n6032_), .A3(new_n720_), .ZN(new_n6033_));
  NAND2_X1   g05841(.A1(new_n6033_), .A2(new_n5823_), .ZN(new_n6034_));
  NAND2_X1   g05842(.A1(new_n6030_), .A2(new_n6032_), .ZN(new_n6035_));
  AOI21_X1   g05843(.A1(new_n6035_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n6036_));
  AOI21_X1   g05844(.A1(new_n6036_), .A2(new_n6034_), .B(new_n6025_), .ZN(new_n6037_));
  AOI21_X1   g05845(.A1(new_n6034_), .A2(new_n6015_), .B(new_n630_), .ZN(new_n6038_));
  OAI21_X1   g05846(.A1(new_n6037_), .A2(new_n6038_), .B(\asqrt[56] ), .ZN(new_n6039_));
  AOI21_X1   g05847(.A1(new_n6021_), .A2(new_n6039_), .B(new_n450_), .ZN(new_n6040_));
  NOR2_X1    g05848(.A1(new_n6024_), .A2(new_n6040_), .ZN(new_n6041_));
  AOI21_X1   g05849(.A1(new_n6041_), .A2(new_n403_), .B(new_n5812_), .ZN(new_n6042_));
  OAI21_X1   g05850(.A1(new_n6024_), .A2(new_n6040_), .B(\asqrt[58] ), .ZN(new_n6043_));
  NAND2_X1   g05851(.A1(new_n6043_), .A2(new_n339_), .ZN(new_n6044_));
  OAI21_X1   g05852(.A1(new_n6042_), .A2(new_n6044_), .B(new_n5808_), .ZN(new_n6045_));
  INV_X1     g05853(.I(new_n6043_), .ZN(new_n6046_));
  OAI21_X1   g05854(.A1(new_n6042_), .A2(new_n6046_), .B(\asqrt[59] ), .ZN(new_n6047_));
  NAND3_X1   g05855(.A1(new_n6045_), .A2(new_n6047_), .A3(new_n288_), .ZN(new_n6048_));
  NAND2_X1   g05856(.A1(new_n6048_), .A2(new_n5806_), .ZN(new_n6049_));
  INV_X1     g05857(.I(new_n5808_), .ZN(new_n6050_));
  INV_X1     g05858(.I(new_n5818_), .ZN(new_n6051_));
  NOR2_X1    g05859(.A1(new_n6037_), .A2(new_n6038_), .ZN(new_n6052_));
  AOI21_X1   g05860(.A1(new_n6052_), .A2(new_n545_), .B(new_n6051_), .ZN(new_n6053_));
  NAND2_X1   g05861(.A1(new_n6039_), .A2(new_n450_), .ZN(new_n6054_));
  OAI21_X1   g05862(.A1(new_n6053_), .A2(new_n6054_), .B(new_n5814_), .ZN(new_n6055_));
  INV_X1     g05863(.I(new_n6039_), .ZN(new_n6056_));
  OAI21_X1   g05864(.A1(new_n6053_), .A2(new_n6056_), .B(\asqrt[57] ), .ZN(new_n6057_));
  NAND3_X1   g05865(.A1(new_n6055_), .A2(new_n6057_), .A3(new_n403_), .ZN(new_n6058_));
  NAND2_X1   g05866(.A1(new_n6058_), .A2(new_n5811_), .ZN(new_n6059_));
  NAND2_X1   g05867(.A1(new_n6055_), .A2(new_n6057_), .ZN(new_n6060_));
  AOI21_X1   g05868(.A1(new_n6060_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n6061_));
  AOI21_X1   g05869(.A1(new_n6061_), .A2(new_n6059_), .B(new_n6050_), .ZN(new_n6062_));
  AOI21_X1   g05870(.A1(new_n6059_), .A2(new_n6043_), .B(new_n339_), .ZN(new_n6063_));
  OAI21_X1   g05871(.A1(new_n6062_), .A2(new_n6063_), .B(\asqrt[60] ), .ZN(new_n6064_));
  AOI21_X1   g05872(.A1(new_n6049_), .A2(new_n6064_), .B(new_n242_), .ZN(new_n6065_));
  NAND3_X1   g05873(.A1(\asqrt[31] ), .A2(new_n5708_), .A3(new_n5724_), .ZN(new_n6066_));
  XOR2_X1    g05874(.A1(new_n6066_), .A2(new_n5736_), .Z(new_n6067_));
  INV_X1     g05875(.I(new_n6067_), .ZN(new_n6068_));
  NAND2_X1   g05876(.A1(new_n6045_), .A2(new_n6047_), .ZN(new_n6069_));
  AOI21_X1   g05877(.A1(new_n6069_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n6070_));
  AOI21_X1   g05878(.A1(new_n6070_), .A2(new_n6049_), .B(new_n6068_), .ZN(new_n6071_));
  OAI21_X1   g05879(.A1(new_n6071_), .A2(new_n6065_), .B(\asqrt[62] ), .ZN(new_n6072_));
  INV_X1     g05880(.I(new_n6072_), .ZN(new_n6073_));
  NOR2_X1    g05881(.A1(new_n6071_), .A2(new_n6065_), .ZN(new_n6074_));
  AOI21_X1   g05882(.A1(new_n5709_), .A2(new_n5730_), .B(new_n5725_), .ZN(new_n6075_));
  NAND2_X1   g05883(.A1(\asqrt[31] ), .A2(new_n6075_), .ZN(new_n6076_));
  XOR2_X1    g05884(.A1(new_n6076_), .A2(new_n5728_), .Z(new_n6077_));
  INV_X1     g05885(.I(new_n6077_), .ZN(new_n6078_));
  AOI21_X1   g05886(.A1(new_n6074_), .A2(new_n234_), .B(new_n6078_), .ZN(new_n6079_));
  OAI21_X1   g05887(.A1(new_n6079_), .A2(new_n6073_), .B(new_n5803_), .ZN(new_n6080_));
  OAI21_X1   g05888(.A1(new_n6080_), .A2(new_n5802_), .B(new_n193_), .ZN(new_n6081_));
  NOR2_X1    g05889(.A1(new_n6079_), .A2(new_n6073_), .ZN(new_n6082_));
  NAND2_X1   g05890(.A1(new_n6082_), .A2(new_n5802_), .ZN(new_n6083_));
  NOR2_X1    g05891(.A1(\asqrt[31] ), .A2(new_n5451_), .ZN(new_n6084_));
  INV_X1     g05892(.I(new_n6084_), .ZN(new_n6085_));
  NAND4_X1   g05893(.A1(new_n6081_), .A2(new_n5800_), .A3(new_n6083_), .A4(new_n6085_), .ZN(\asqrt[30] ));
  NAND3_X1   g05894(.A1(\asqrt[30] ), .A2(new_n5783_), .A3(new_n5795_), .ZN(new_n6087_));
  XOR2_X1    g05895(.A1(new_n6087_), .A2(new_n5753_), .Z(new_n6088_));
  INV_X1     g05896(.I(new_n6088_), .ZN(new_n6089_));
  INV_X1     g05897(.I(new_n5806_), .ZN(new_n6090_));
  NOR2_X1    g05898(.A1(new_n6062_), .A2(new_n6063_), .ZN(new_n6091_));
  AOI21_X1   g05899(.A1(new_n6091_), .A2(new_n288_), .B(new_n6090_), .ZN(new_n6092_));
  INV_X1     g05900(.I(new_n6064_), .ZN(new_n6093_));
  OAI21_X1   g05901(.A1(new_n6092_), .A2(new_n6093_), .B(\asqrt[61] ), .ZN(new_n6094_));
  NAND2_X1   g05902(.A1(new_n6064_), .A2(new_n242_), .ZN(new_n6095_));
  OAI21_X1   g05903(.A1(new_n6092_), .A2(new_n6095_), .B(new_n6067_), .ZN(new_n6096_));
  NAND3_X1   g05904(.A1(new_n6096_), .A2(new_n6094_), .A3(new_n234_), .ZN(new_n6097_));
  NAND2_X1   g05905(.A1(new_n6097_), .A2(new_n6077_), .ZN(new_n6098_));
  NAND2_X1   g05906(.A1(new_n6098_), .A2(new_n6072_), .ZN(new_n6099_));
  NAND2_X1   g05907(.A1(new_n6099_), .A2(new_n5802_), .ZN(new_n6100_));
  INV_X1     g05908(.I(new_n5802_), .ZN(new_n6101_));
  INV_X1     g05909(.I(new_n5803_), .ZN(new_n6102_));
  AOI21_X1   g05910(.A1(new_n6098_), .A2(new_n6072_), .B(new_n6102_), .ZN(new_n6103_));
  AOI21_X1   g05911(.A1(new_n6103_), .A2(new_n6101_), .B(\asqrt[63] ), .ZN(new_n6104_));
  NOR2_X1    g05912(.A1(new_n6099_), .A2(new_n6101_), .ZN(new_n6105_));
  NOR4_X1    g05913(.A1(new_n6104_), .A2(new_n5799_), .A3(new_n6105_), .A4(new_n6084_), .ZN(new_n6106_));
  NOR2_X1    g05914(.A1(new_n6106_), .A2(new_n5802_), .ZN(new_n6107_));
  NAND2_X1   g05915(.A1(new_n6107_), .A2(new_n6082_), .ZN(new_n6108_));
  AOI21_X1   g05916(.A1(new_n6108_), .A2(new_n6100_), .B(new_n193_), .ZN(new_n6109_));
  INV_X1     g05917(.I(new_n6109_), .ZN(new_n6110_));
  NAND3_X1   g05918(.A1(\asqrt[30] ), .A2(new_n6072_), .A3(new_n6097_), .ZN(new_n6111_));
  XOR2_X1    g05919(.A1(new_n6111_), .A2(new_n6077_), .Z(new_n6112_));
  AOI21_X1   g05920(.A1(new_n6107_), .A2(new_n6099_), .B(new_n6105_), .ZN(new_n6113_));
  OAI21_X1   g05921(.A1(new_n6042_), .A2(new_n6044_), .B(new_n6047_), .ZN(new_n6114_));
  NOR2_X1    g05922(.A1(new_n6106_), .A2(new_n6114_), .ZN(new_n6115_));
  XOR2_X1    g05923(.A1(new_n6115_), .A2(new_n5808_), .Z(new_n6116_));
  NAND3_X1   g05924(.A1(\asqrt[30] ), .A2(new_n6058_), .A3(new_n6043_), .ZN(new_n6117_));
  XOR2_X1    g05925(.A1(new_n6117_), .A2(new_n5812_), .Z(new_n6118_));
  OAI21_X1   g05926(.A1(new_n6053_), .A2(new_n6054_), .B(new_n6057_), .ZN(new_n6119_));
  NOR2_X1    g05927(.A1(new_n6106_), .A2(new_n6119_), .ZN(new_n6120_));
  XOR2_X1    g05928(.A1(new_n6120_), .A2(new_n5814_), .Z(new_n6121_));
  INV_X1     g05929(.I(new_n6121_), .ZN(new_n6122_));
  NAND3_X1   g05930(.A1(\asqrt[30] ), .A2(new_n6020_), .A3(new_n6039_), .ZN(new_n6123_));
  XOR2_X1    g05931(.A1(new_n6123_), .A2(new_n6051_), .Z(new_n6124_));
  INV_X1     g05932(.I(new_n6124_), .ZN(new_n6125_));
  OAI21_X1   g05933(.A1(new_n6014_), .A2(new_n6016_), .B(new_n6019_), .ZN(new_n6126_));
  NOR2_X1    g05934(.A1(new_n6106_), .A2(new_n6126_), .ZN(new_n6127_));
  XOR2_X1    g05935(.A1(new_n6127_), .A2(new_n5820_), .Z(new_n6128_));
  NAND3_X1   g05936(.A1(\asqrt[30] ), .A2(new_n6033_), .A3(new_n6015_), .ZN(new_n6129_));
  XOR2_X1    g05937(.A1(new_n6129_), .A2(new_n5824_), .Z(new_n6130_));
  OAI21_X1   g05938(.A1(new_n6028_), .A2(new_n6029_), .B(new_n6032_), .ZN(new_n6131_));
  NOR2_X1    g05939(.A1(new_n6106_), .A2(new_n6131_), .ZN(new_n6132_));
  XOR2_X1    g05940(.A1(new_n6132_), .A2(new_n5826_), .Z(new_n6133_));
  INV_X1     g05941(.I(new_n6133_), .ZN(new_n6134_));
  NAND3_X1   g05942(.A1(\asqrt[30] ), .A2(new_n5992_), .A3(new_n6011_), .ZN(new_n6135_));
  XOR2_X1    g05943(.A1(new_n6135_), .A2(new_n6026_), .Z(new_n6136_));
  INV_X1     g05944(.I(new_n6136_), .ZN(new_n6137_));
  OAI21_X1   g05945(.A1(new_n5986_), .A2(new_n5988_), .B(new_n5991_), .ZN(new_n6138_));
  NOR2_X1    g05946(.A1(new_n6106_), .A2(new_n6138_), .ZN(new_n6139_));
  XOR2_X1    g05947(.A1(new_n6139_), .A2(new_n5832_), .Z(new_n6140_));
  NAND3_X1   g05948(.A1(\asqrt[30] ), .A2(new_n6005_), .A3(new_n5987_), .ZN(new_n6141_));
  XOR2_X1    g05949(.A1(new_n6141_), .A2(new_n5836_), .Z(new_n6142_));
  OAI21_X1   g05950(.A1(new_n6000_), .A2(new_n6001_), .B(new_n6004_), .ZN(new_n6143_));
  NOR2_X1    g05951(.A1(new_n6106_), .A2(new_n6143_), .ZN(new_n6144_));
  XOR2_X1    g05952(.A1(new_n6144_), .A2(new_n5838_), .Z(new_n6145_));
  INV_X1     g05953(.I(new_n6145_), .ZN(new_n6146_));
  NAND3_X1   g05954(.A1(\asqrt[30] ), .A2(new_n5964_), .A3(new_n5983_), .ZN(new_n6147_));
  XOR2_X1    g05955(.A1(new_n6147_), .A2(new_n5998_), .Z(new_n6148_));
  INV_X1     g05956(.I(new_n6148_), .ZN(new_n6149_));
  OAI21_X1   g05957(.A1(new_n5958_), .A2(new_n5960_), .B(new_n5963_), .ZN(new_n6150_));
  NOR2_X1    g05958(.A1(new_n6106_), .A2(new_n6150_), .ZN(new_n6151_));
  XOR2_X1    g05959(.A1(new_n6151_), .A2(new_n5844_), .Z(new_n6152_));
  NAND3_X1   g05960(.A1(\asqrt[30] ), .A2(new_n5977_), .A3(new_n5959_), .ZN(new_n6153_));
  XOR2_X1    g05961(.A1(new_n6153_), .A2(new_n5848_), .Z(new_n6154_));
  OAI21_X1   g05962(.A1(new_n5972_), .A2(new_n5973_), .B(new_n5976_), .ZN(new_n6155_));
  NOR2_X1    g05963(.A1(new_n6106_), .A2(new_n6155_), .ZN(new_n6156_));
  XOR2_X1    g05964(.A1(new_n6156_), .A2(new_n5850_), .Z(new_n6157_));
  INV_X1     g05965(.I(new_n6157_), .ZN(new_n6158_));
  NAND3_X1   g05966(.A1(\asqrt[30] ), .A2(new_n5936_), .A3(new_n5955_), .ZN(new_n6159_));
  XOR2_X1    g05967(.A1(new_n6159_), .A2(new_n5970_), .Z(new_n6160_));
  INV_X1     g05968(.I(new_n6160_), .ZN(new_n6161_));
  OAI21_X1   g05969(.A1(new_n5930_), .A2(new_n5932_), .B(new_n5935_), .ZN(new_n6162_));
  NOR2_X1    g05970(.A1(new_n6106_), .A2(new_n6162_), .ZN(new_n6163_));
  XOR2_X1    g05971(.A1(new_n6163_), .A2(new_n5856_), .Z(new_n6164_));
  NAND3_X1   g05972(.A1(\asqrt[30] ), .A2(new_n5949_), .A3(new_n5931_), .ZN(new_n6165_));
  XOR2_X1    g05973(.A1(new_n6165_), .A2(new_n5860_), .Z(new_n6166_));
  OAI21_X1   g05974(.A1(new_n5944_), .A2(new_n5945_), .B(new_n5948_), .ZN(new_n6167_));
  NOR2_X1    g05975(.A1(new_n6106_), .A2(new_n6167_), .ZN(new_n6168_));
  XOR2_X1    g05976(.A1(new_n6168_), .A2(new_n5862_), .Z(new_n6169_));
  INV_X1     g05977(.I(new_n6169_), .ZN(new_n6170_));
  NAND3_X1   g05978(.A1(\asqrt[30] ), .A2(new_n5908_), .A3(new_n5927_), .ZN(new_n6171_));
  XOR2_X1    g05979(.A1(new_n6171_), .A2(new_n5942_), .Z(new_n6172_));
  INV_X1     g05980(.I(new_n6172_), .ZN(new_n6173_));
  OAI21_X1   g05981(.A1(new_n5902_), .A2(new_n5904_), .B(new_n5907_), .ZN(new_n6174_));
  NOR2_X1    g05982(.A1(new_n6106_), .A2(new_n6174_), .ZN(new_n6175_));
  XOR2_X1    g05983(.A1(new_n6175_), .A2(new_n5868_), .Z(new_n6176_));
  NAND3_X1   g05984(.A1(\asqrt[30] ), .A2(new_n5921_), .A3(new_n5903_), .ZN(new_n6177_));
  XOR2_X1    g05985(.A1(new_n6177_), .A2(new_n5872_), .Z(new_n6178_));
  OAI21_X1   g05986(.A1(new_n5916_), .A2(new_n5917_), .B(new_n5920_), .ZN(new_n6179_));
  NOR2_X1    g05987(.A1(new_n6106_), .A2(new_n6179_), .ZN(new_n6180_));
  XOR2_X1    g05988(.A1(new_n6180_), .A2(new_n5875_), .Z(new_n6181_));
  INV_X1     g05989(.I(new_n6181_), .ZN(new_n6182_));
  NAND3_X1   g05990(.A1(\asqrt[30] ), .A2(new_n5888_), .A3(new_n5899_), .ZN(new_n6183_));
  XOR2_X1    g05991(.A1(new_n6183_), .A2(new_n5914_), .Z(new_n6184_));
  INV_X1     g05992(.I(new_n6184_), .ZN(new_n6185_));
  OAI21_X1   g05993(.A1(new_n5883_), .A2(new_n5884_), .B(new_n5887_), .ZN(new_n6186_));
  NOR2_X1    g05994(.A1(new_n6106_), .A2(new_n6186_), .ZN(new_n6187_));
  XOR2_X1    g05995(.A1(new_n6187_), .A2(new_n5881_), .Z(new_n6188_));
  NOR2_X1    g05996(.A1(new_n5780_), .A2(\asqrt[33] ), .ZN(new_n6189_));
  NOR3_X1    g05997(.A1(new_n6106_), .A2(new_n6189_), .A3(new_n5794_), .ZN(new_n6190_));
  XOR2_X1    g05998(.A1(new_n6190_), .A2(new_n5771_), .Z(new_n6191_));
  INV_X1     g05999(.I(new_n6191_), .ZN(new_n6192_));
  NAND3_X1   g06000(.A1(\asqrt[30] ), .A2(new_n5772_), .A3(new_n5773_), .ZN(new_n6193_));
  NOR4_X1    g06001(.A1(new_n6104_), .A2(new_n5750_), .A3(new_n5799_), .A4(new_n6105_), .ZN(new_n6194_));
  INV_X1     g06002(.I(new_n6194_), .ZN(new_n6195_));
  AOI21_X1   g06003(.A1(new_n6193_), .A2(new_n6195_), .B(\a[62] ), .ZN(new_n6196_));
  NOR3_X1    g06004(.A1(new_n6106_), .A2(\a[60] ), .A3(\a[61] ), .ZN(new_n6197_));
  NOR3_X1    g06005(.A1(new_n6197_), .A2(new_n5438_), .A3(new_n6194_), .ZN(new_n6198_));
  NOR2_X1    g06006(.A1(new_n6198_), .A2(new_n6196_), .ZN(new_n6199_));
  INV_X1     g06007(.I(\a[58] ), .ZN(new_n6200_));
  INV_X1     g06008(.I(\a[59] ), .ZN(new_n6201_));
  NAND3_X1   g06009(.A1(new_n6200_), .A2(new_n6201_), .A3(new_n5772_), .ZN(new_n6202_));
  OAI21_X1   g06010(.A1(new_n6106_), .A2(new_n5772_), .B(new_n6202_), .ZN(new_n6203_));
  NAND2_X1   g06011(.A1(new_n6203_), .A2(\asqrt[31] ), .ZN(new_n6204_));
  OAI21_X1   g06012(.A1(new_n6106_), .A2(\a[60] ), .B(\a[61] ), .ZN(new_n6205_));
  NAND2_X1   g06013(.A1(new_n6205_), .A2(new_n6193_), .ZN(new_n6206_));
  NOR2_X1    g06014(.A1(new_n6203_), .A2(\asqrt[31] ), .ZN(new_n6207_));
  OAI21_X1   g06015(.A1(new_n6206_), .A2(new_n6207_), .B(new_n6204_), .ZN(new_n6208_));
  OAI21_X1   g06016(.A1(new_n6208_), .A2(\asqrt[32] ), .B(new_n6199_), .ZN(new_n6209_));
  NAND2_X1   g06017(.A1(new_n6208_), .A2(\asqrt[32] ), .ZN(new_n6210_));
  NAND3_X1   g06018(.A1(new_n6209_), .A2(new_n5110_), .A3(new_n6210_), .ZN(new_n6211_));
  NOR3_X1    g06019(.A1(new_n6106_), .A2(new_n5788_), .A3(new_n5779_), .ZN(new_n6212_));
  XOR2_X1    g06020(.A1(new_n6212_), .A2(new_n5790_), .Z(new_n6213_));
  AOI21_X1   g06021(.A1(new_n6209_), .A2(new_n6210_), .B(new_n5110_), .ZN(new_n6214_));
  AOI21_X1   g06022(.A1(new_n6211_), .A2(new_n6213_), .B(new_n6214_), .ZN(new_n6215_));
  AOI21_X1   g06023(.A1(new_n6215_), .A2(new_n4810_), .B(new_n6192_), .ZN(new_n6216_));
  OAI21_X1   g06024(.A1(new_n6215_), .A2(new_n4810_), .B(new_n4510_), .ZN(new_n6217_));
  OAI21_X1   g06025(.A1(new_n6216_), .A2(new_n6217_), .B(new_n6088_), .ZN(new_n6218_));
  NOR2_X1    g06026(.A1(new_n6215_), .A2(new_n4810_), .ZN(new_n6219_));
  OAI21_X1   g06027(.A1(new_n6216_), .A2(new_n6219_), .B(\asqrt[35] ), .ZN(new_n6220_));
  NAND3_X1   g06028(.A1(new_n6218_), .A2(new_n6220_), .A3(new_n4224_), .ZN(new_n6221_));
  NAND2_X1   g06029(.A1(new_n6221_), .A2(new_n6188_), .ZN(new_n6222_));
  NAND2_X1   g06030(.A1(new_n6218_), .A2(new_n6220_), .ZN(new_n6223_));
  AOI21_X1   g06031(.A1(new_n6223_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n6224_));
  AOI21_X1   g06032(.A1(new_n6224_), .A2(new_n6222_), .B(new_n6185_), .ZN(new_n6225_));
  OAI21_X1   g06033(.A1(new_n6197_), .A2(new_n6194_), .B(new_n5438_), .ZN(new_n6226_));
  NAND3_X1   g06034(.A1(new_n6193_), .A2(new_n6195_), .A3(\a[62] ), .ZN(new_n6227_));
  NAND2_X1   g06035(.A1(new_n6226_), .A2(new_n6227_), .ZN(new_n6228_));
  NAND2_X1   g06036(.A1(\asqrt[30] ), .A2(\a[60] ), .ZN(new_n6229_));
  AOI21_X1   g06037(.A1(new_n6229_), .A2(new_n6202_), .B(new_n5750_), .ZN(new_n6230_));
  AOI21_X1   g06038(.A1(\asqrt[30] ), .A2(new_n5772_), .B(new_n5773_), .ZN(new_n6231_));
  NOR2_X1    g06039(.A1(new_n6197_), .A2(new_n6231_), .ZN(new_n6232_));
  NAND3_X1   g06040(.A1(new_n6229_), .A2(new_n5750_), .A3(new_n6202_), .ZN(new_n6233_));
  AOI21_X1   g06041(.A1(new_n6232_), .A2(new_n6233_), .B(new_n6230_), .ZN(new_n6234_));
  AOI21_X1   g06042(.A1(new_n6234_), .A2(new_n5435_), .B(new_n6228_), .ZN(new_n6235_));
  NOR2_X1    g06043(.A1(new_n6234_), .A2(new_n5435_), .ZN(new_n6236_));
  NOR3_X1    g06044(.A1(new_n6235_), .A2(\asqrt[33] ), .A3(new_n6236_), .ZN(new_n6237_));
  INV_X1     g06045(.I(new_n6213_), .ZN(new_n6238_));
  OAI21_X1   g06046(.A1(new_n6235_), .A2(new_n6236_), .B(\asqrt[33] ), .ZN(new_n6239_));
  OAI21_X1   g06047(.A1(new_n6237_), .A2(new_n6238_), .B(new_n6239_), .ZN(new_n6240_));
  OAI21_X1   g06048(.A1(new_n6240_), .A2(\asqrt[34] ), .B(new_n6191_), .ZN(new_n6241_));
  AOI21_X1   g06049(.A1(new_n6240_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n6242_));
  AOI21_X1   g06050(.A1(new_n6242_), .A2(new_n6241_), .B(new_n6089_), .ZN(new_n6243_));
  NAND2_X1   g06051(.A1(new_n6240_), .A2(\asqrt[34] ), .ZN(new_n6244_));
  AOI21_X1   g06052(.A1(new_n6241_), .A2(new_n6244_), .B(new_n4510_), .ZN(new_n6245_));
  OAI21_X1   g06053(.A1(new_n6243_), .A2(new_n6245_), .B(\asqrt[36] ), .ZN(new_n6246_));
  AOI21_X1   g06054(.A1(new_n6222_), .A2(new_n6246_), .B(new_n3928_), .ZN(new_n6247_));
  NOR2_X1    g06055(.A1(new_n6225_), .A2(new_n6247_), .ZN(new_n6248_));
  AOI21_X1   g06056(.A1(new_n6248_), .A2(new_n3675_), .B(new_n6182_), .ZN(new_n6249_));
  OAI21_X1   g06057(.A1(new_n6225_), .A2(new_n6247_), .B(\asqrt[38] ), .ZN(new_n6250_));
  NAND2_X1   g06058(.A1(new_n6250_), .A2(new_n3400_), .ZN(new_n6251_));
  OAI21_X1   g06059(.A1(new_n6249_), .A2(new_n6251_), .B(new_n6178_), .ZN(new_n6252_));
  INV_X1     g06060(.I(new_n6250_), .ZN(new_n6253_));
  OAI21_X1   g06061(.A1(new_n6249_), .A2(new_n6253_), .B(\asqrt[39] ), .ZN(new_n6254_));
  NAND3_X1   g06062(.A1(new_n6252_), .A2(new_n6254_), .A3(new_n3167_), .ZN(new_n6255_));
  NAND2_X1   g06063(.A1(new_n6255_), .A2(new_n6176_), .ZN(new_n6256_));
  NAND2_X1   g06064(.A1(new_n6252_), .A2(new_n6254_), .ZN(new_n6257_));
  AOI21_X1   g06065(.A1(new_n6257_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n6258_));
  AOI21_X1   g06066(.A1(new_n6258_), .A2(new_n6256_), .B(new_n6173_), .ZN(new_n6259_));
  INV_X1     g06067(.I(new_n6178_), .ZN(new_n6260_));
  INV_X1     g06068(.I(new_n6188_), .ZN(new_n6261_));
  NOR2_X1    g06069(.A1(new_n6243_), .A2(new_n6245_), .ZN(new_n6262_));
  AOI21_X1   g06070(.A1(new_n6262_), .A2(new_n4224_), .B(new_n6261_), .ZN(new_n6263_));
  NAND2_X1   g06071(.A1(new_n6246_), .A2(new_n3928_), .ZN(new_n6264_));
  OAI21_X1   g06072(.A1(new_n6263_), .A2(new_n6264_), .B(new_n6184_), .ZN(new_n6265_));
  INV_X1     g06073(.I(new_n6246_), .ZN(new_n6266_));
  OAI21_X1   g06074(.A1(new_n6263_), .A2(new_n6266_), .B(\asqrt[37] ), .ZN(new_n6267_));
  NAND3_X1   g06075(.A1(new_n6265_), .A2(new_n6267_), .A3(new_n3675_), .ZN(new_n6268_));
  NAND2_X1   g06076(.A1(new_n6268_), .A2(new_n6181_), .ZN(new_n6269_));
  NAND2_X1   g06077(.A1(new_n6265_), .A2(new_n6267_), .ZN(new_n6270_));
  AOI21_X1   g06078(.A1(new_n6270_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n6271_));
  AOI21_X1   g06079(.A1(new_n6271_), .A2(new_n6269_), .B(new_n6260_), .ZN(new_n6272_));
  AOI21_X1   g06080(.A1(new_n6269_), .A2(new_n6250_), .B(new_n3400_), .ZN(new_n6273_));
  OAI21_X1   g06081(.A1(new_n6272_), .A2(new_n6273_), .B(\asqrt[40] ), .ZN(new_n6274_));
  AOI21_X1   g06082(.A1(new_n6256_), .A2(new_n6274_), .B(new_n2912_), .ZN(new_n6275_));
  NOR2_X1    g06083(.A1(new_n6259_), .A2(new_n6275_), .ZN(new_n6276_));
  AOI21_X1   g06084(.A1(new_n6276_), .A2(new_n2699_), .B(new_n6170_), .ZN(new_n6277_));
  OAI21_X1   g06085(.A1(new_n6259_), .A2(new_n6275_), .B(\asqrt[42] ), .ZN(new_n6278_));
  NAND2_X1   g06086(.A1(new_n6278_), .A2(new_n2464_), .ZN(new_n6279_));
  OAI21_X1   g06087(.A1(new_n6277_), .A2(new_n6279_), .B(new_n6166_), .ZN(new_n6280_));
  INV_X1     g06088(.I(new_n6278_), .ZN(new_n6281_));
  OAI21_X1   g06089(.A1(new_n6277_), .A2(new_n6281_), .B(\asqrt[43] ), .ZN(new_n6282_));
  NAND3_X1   g06090(.A1(new_n6280_), .A2(new_n6282_), .A3(new_n2271_), .ZN(new_n6283_));
  NAND2_X1   g06091(.A1(new_n6283_), .A2(new_n6164_), .ZN(new_n6284_));
  NAND2_X1   g06092(.A1(new_n6280_), .A2(new_n6282_), .ZN(new_n6285_));
  AOI21_X1   g06093(.A1(new_n6285_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n6286_));
  AOI21_X1   g06094(.A1(new_n6286_), .A2(new_n6284_), .B(new_n6161_), .ZN(new_n6287_));
  INV_X1     g06095(.I(new_n6166_), .ZN(new_n6288_));
  INV_X1     g06096(.I(new_n6176_), .ZN(new_n6289_));
  NOR2_X1    g06097(.A1(new_n6272_), .A2(new_n6273_), .ZN(new_n6290_));
  AOI21_X1   g06098(.A1(new_n6290_), .A2(new_n3167_), .B(new_n6289_), .ZN(new_n6291_));
  NAND2_X1   g06099(.A1(new_n6274_), .A2(new_n2912_), .ZN(new_n6292_));
  OAI21_X1   g06100(.A1(new_n6291_), .A2(new_n6292_), .B(new_n6172_), .ZN(new_n6293_));
  INV_X1     g06101(.I(new_n6274_), .ZN(new_n6294_));
  OAI21_X1   g06102(.A1(new_n6291_), .A2(new_n6294_), .B(\asqrt[41] ), .ZN(new_n6295_));
  NAND3_X1   g06103(.A1(new_n6293_), .A2(new_n6295_), .A3(new_n2699_), .ZN(new_n6296_));
  NAND2_X1   g06104(.A1(new_n6296_), .A2(new_n6169_), .ZN(new_n6297_));
  NAND2_X1   g06105(.A1(new_n6293_), .A2(new_n6295_), .ZN(new_n6298_));
  AOI21_X1   g06106(.A1(new_n6298_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n6299_));
  AOI21_X1   g06107(.A1(new_n6299_), .A2(new_n6297_), .B(new_n6288_), .ZN(new_n6300_));
  AOI21_X1   g06108(.A1(new_n6297_), .A2(new_n6278_), .B(new_n2464_), .ZN(new_n6301_));
  OAI21_X1   g06109(.A1(new_n6300_), .A2(new_n6301_), .B(\asqrt[44] ), .ZN(new_n6302_));
  AOI21_X1   g06110(.A1(new_n6284_), .A2(new_n6302_), .B(new_n2072_), .ZN(new_n6303_));
  NOR2_X1    g06111(.A1(new_n6287_), .A2(new_n6303_), .ZN(new_n6304_));
  AOI21_X1   g06112(.A1(new_n6304_), .A2(new_n1884_), .B(new_n6158_), .ZN(new_n6305_));
  OAI21_X1   g06113(.A1(new_n6287_), .A2(new_n6303_), .B(\asqrt[46] ), .ZN(new_n6306_));
  NAND2_X1   g06114(.A1(new_n6306_), .A2(new_n1688_), .ZN(new_n6307_));
  OAI21_X1   g06115(.A1(new_n6305_), .A2(new_n6307_), .B(new_n6154_), .ZN(new_n6308_));
  INV_X1     g06116(.I(new_n6306_), .ZN(new_n6309_));
  OAI21_X1   g06117(.A1(new_n6305_), .A2(new_n6309_), .B(\asqrt[47] ), .ZN(new_n6310_));
  NAND3_X1   g06118(.A1(new_n6308_), .A2(new_n6310_), .A3(new_n1533_), .ZN(new_n6311_));
  NAND2_X1   g06119(.A1(new_n6311_), .A2(new_n6152_), .ZN(new_n6312_));
  NAND2_X1   g06120(.A1(new_n6308_), .A2(new_n6310_), .ZN(new_n6313_));
  AOI21_X1   g06121(.A1(new_n6313_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n6314_));
  AOI21_X1   g06122(.A1(new_n6314_), .A2(new_n6312_), .B(new_n6149_), .ZN(new_n6315_));
  INV_X1     g06123(.I(new_n6154_), .ZN(new_n6316_));
  INV_X1     g06124(.I(new_n6164_), .ZN(new_n6317_));
  NOR2_X1    g06125(.A1(new_n6300_), .A2(new_n6301_), .ZN(new_n6318_));
  AOI21_X1   g06126(.A1(new_n6318_), .A2(new_n2271_), .B(new_n6317_), .ZN(new_n6319_));
  NAND2_X1   g06127(.A1(new_n6302_), .A2(new_n2072_), .ZN(new_n6320_));
  OAI21_X1   g06128(.A1(new_n6319_), .A2(new_n6320_), .B(new_n6160_), .ZN(new_n6321_));
  INV_X1     g06129(.I(new_n6302_), .ZN(new_n6322_));
  OAI21_X1   g06130(.A1(new_n6319_), .A2(new_n6322_), .B(\asqrt[45] ), .ZN(new_n6323_));
  NAND3_X1   g06131(.A1(new_n6321_), .A2(new_n6323_), .A3(new_n1884_), .ZN(new_n6324_));
  NAND2_X1   g06132(.A1(new_n6324_), .A2(new_n6157_), .ZN(new_n6325_));
  NAND2_X1   g06133(.A1(new_n6321_), .A2(new_n6323_), .ZN(new_n6326_));
  AOI21_X1   g06134(.A1(new_n6326_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n6327_));
  AOI21_X1   g06135(.A1(new_n6327_), .A2(new_n6325_), .B(new_n6316_), .ZN(new_n6328_));
  AOI21_X1   g06136(.A1(new_n6325_), .A2(new_n6306_), .B(new_n1688_), .ZN(new_n6329_));
  OAI21_X1   g06137(.A1(new_n6328_), .A2(new_n6329_), .B(\asqrt[48] ), .ZN(new_n6330_));
  AOI21_X1   g06138(.A1(new_n6312_), .A2(new_n6330_), .B(new_n1368_), .ZN(new_n6331_));
  NOR2_X1    g06139(.A1(new_n6315_), .A2(new_n6331_), .ZN(new_n6332_));
  AOI21_X1   g06140(.A1(new_n6332_), .A2(new_n1228_), .B(new_n6146_), .ZN(new_n6333_));
  OAI21_X1   g06141(.A1(new_n6315_), .A2(new_n6331_), .B(\asqrt[50] ), .ZN(new_n6334_));
  NAND2_X1   g06142(.A1(new_n6334_), .A2(new_n1088_), .ZN(new_n6335_));
  OAI21_X1   g06143(.A1(new_n6333_), .A2(new_n6335_), .B(new_n6142_), .ZN(new_n6336_));
  INV_X1     g06144(.I(new_n6334_), .ZN(new_n6337_));
  OAI21_X1   g06145(.A1(new_n6333_), .A2(new_n6337_), .B(\asqrt[51] ), .ZN(new_n6338_));
  NAND3_X1   g06146(.A1(new_n6336_), .A2(new_n6338_), .A3(new_n962_), .ZN(new_n6339_));
  NAND2_X1   g06147(.A1(new_n6339_), .A2(new_n6140_), .ZN(new_n6340_));
  NAND2_X1   g06148(.A1(new_n6336_), .A2(new_n6338_), .ZN(new_n6341_));
  AOI21_X1   g06149(.A1(new_n6341_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n6342_));
  AOI21_X1   g06150(.A1(new_n6342_), .A2(new_n6340_), .B(new_n6137_), .ZN(new_n6343_));
  INV_X1     g06151(.I(new_n6142_), .ZN(new_n6344_));
  INV_X1     g06152(.I(new_n6152_), .ZN(new_n6345_));
  NOR2_X1    g06153(.A1(new_n6328_), .A2(new_n6329_), .ZN(new_n6346_));
  AOI21_X1   g06154(.A1(new_n6346_), .A2(new_n1533_), .B(new_n6345_), .ZN(new_n6347_));
  NAND2_X1   g06155(.A1(new_n6330_), .A2(new_n1368_), .ZN(new_n6348_));
  OAI21_X1   g06156(.A1(new_n6347_), .A2(new_n6348_), .B(new_n6148_), .ZN(new_n6349_));
  INV_X1     g06157(.I(new_n6330_), .ZN(new_n6350_));
  OAI21_X1   g06158(.A1(new_n6347_), .A2(new_n6350_), .B(\asqrt[49] ), .ZN(new_n6351_));
  NAND3_X1   g06159(.A1(new_n6349_), .A2(new_n6351_), .A3(new_n1228_), .ZN(new_n6352_));
  NAND2_X1   g06160(.A1(new_n6352_), .A2(new_n6145_), .ZN(new_n6353_));
  NAND2_X1   g06161(.A1(new_n6349_), .A2(new_n6351_), .ZN(new_n6354_));
  AOI21_X1   g06162(.A1(new_n6354_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n6355_));
  AOI21_X1   g06163(.A1(new_n6355_), .A2(new_n6353_), .B(new_n6344_), .ZN(new_n6356_));
  AOI21_X1   g06164(.A1(new_n6353_), .A2(new_n6334_), .B(new_n1088_), .ZN(new_n6357_));
  OAI21_X1   g06165(.A1(new_n6356_), .A2(new_n6357_), .B(\asqrt[52] ), .ZN(new_n6358_));
  AOI21_X1   g06166(.A1(new_n6340_), .A2(new_n6358_), .B(new_n842_), .ZN(new_n6359_));
  NOR2_X1    g06167(.A1(new_n6343_), .A2(new_n6359_), .ZN(new_n6360_));
  AOI21_X1   g06168(.A1(new_n6360_), .A2(new_n720_), .B(new_n6134_), .ZN(new_n6361_));
  OAI21_X1   g06169(.A1(new_n6343_), .A2(new_n6359_), .B(\asqrt[54] ), .ZN(new_n6362_));
  NAND2_X1   g06170(.A1(new_n6362_), .A2(new_n630_), .ZN(new_n6363_));
  OAI21_X1   g06171(.A1(new_n6361_), .A2(new_n6363_), .B(new_n6130_), .ZN(new_n6364_));
  INV_X1     g06172(.I(new_n6362_), .ZN(new_n6365_));
  OAI21_X1   g06173(.A1(new_n6361_), .A2(new_n6365_), .B(\asqrt[55] ), .ZN(new_n6366_));
  NAND3_X1   g06174(.A1(new_n6364_), .A2(new_n6366_), .A3(new_n545_), .ZN(new_n6367_));
  NAND2_X1   g06175(.A1(new_n6367_), .A2(new_n6128_), .ZN(new_n6368_));
  NAND2_X1   g06176(.A1(new_n6364_), .A2(new_n6366_), .ZN(new_n6369_));
  AOI21_X1   g06177(.A1(new_n6369_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n6370_));
  AOI21_X1   g06178(.A1(new_n6370_), .A2(new_n6368_), .B(new_n6125_), .ZN(new_n6371_));
  INV_X1     g06179(.I(new_n6130_), .ZN(new_n6372_));
  INV_X1     g06180(.I(new_n6140_), .ZN(new_n6373_));
  NOR2_X1    g06181(.A1(new_n6356_), .A2(new_n6357_), .ZN(new_n6374_));
  AOI21_X1   g06182(.A1(new_n6374_), .A2(new_n962_), .B(new_n6373_), .ZN(new_n6375_));
  NAND2_X1   g06183(.A1(new_n6358_), .A2(new_n842_), .ZN(new_n6376_));
  OAI21_X1   g06184(.A1(new_n6375_), .A2(new_n6376_), .B(new_n6136_), .ZN(new_n6377_));
  INV_X1     g06185(.I(new_n6358_), .ZN(new_n6378_));
  OAI21_X1   g06186(.A1(new_n6375_), .A2(new_n6378_), .B(\asqrt[53] ), .ZN(new_n6379_));
  NAND3_X1   g06187(.A1(new_n6377_), .A2(new_n6379_), .A3(new_n720_), .ZN(new_n6380_));
  NAND2_X1   g06188(.A1(new_n6380_), .A2(new_n6133_), .ZN(new_n6381_));
  NAND2_X1   g06189(.A1(new_n6377_), .A2(new_n6379_), .ZN(new_n6382_));
  AOI21_X1   g06190(.A1(new_n6382_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n6383_));
  AOI21_X1   g06191(.A1(new_n6383_), .A2(new_n6381_), .B(new_n6372_), .ZN(new_n6384_));
  AOI21_X1   g06192(.A1(new_n6381_), .A2(new_n6362_), .B(new_n630_), .ZN(new_n6385_));
  OAI21_X1   g06193(.A1(new_n6384_), .A2(new_n6385_), .B(\asqrt[56] ), .ZN(new_n6386_));
  AOI21_X1   g06194(.A1(new_n6368_), .A2(new_n6386_), .B(new_n450_), .ZN(new_n6387_));
  NOR2_X1    g06195(.A1(new_n6371_), .A2(new_n6387_), .ZN(new_n6388_));
  AOI21_X1   g06196(.A1(new_n6388_), .A2(new_n403_), .B(new_n6122_), .ZN(new_n6389_));
  OAI21_X1   g06197(.A1(new_n6371_), .A2(new_n6387_), .B(\asqrt[58] ), .ZN(new_n6390_));
  NAND2_X1   g06198(.A1(new_n6390_), .A2(new_n339_), .ZN(new_n6391_));
  OAI21_X1   g06199(.A1(new_n6389_), .A2(new_n6391_), .B(new_n6118_), .ZN(new_n6392_));
  INV_X1     g06200(.I(new_n6390_), .ZN(new_n6393_));
  OAI21_X1   g06201(.A1(new_n6389_), .A2(new_n6393_), .B(\asqrt[59] ), .ZN(new_n6394_));
  NAND3_X1   g06202(.A1(new_n6392_), .A2(new_n6394_), .A3(new_n288_), .ZN(new_n6395_));
  NAND2_X1   g06203(.A1(new_n6395_), .A2(new_n6116_), .ZN(new_n6396_));
  INV_X1     g06204(.I(new_n6118_), .ZN(new_n6397_));
  INV_X1     g06205(.I(new_n6128_), .ZN(new_n6398_));
  NOR2_X1    g06206(.A1(new_n6384_), .A2(new_n6385_), .ZN(new_n6399_));
  AOI21_X1   g06207(.A1(new_n6399_), .A2(new_n545_), .B(new_n6398_), .ZN(new_n6400_));
  NAND2_X1   g06208(.A1(new_n6386_), .A2(new_n450_), .ZN(new_n6401_));
  OAI21_X1   g06209(.A1(new_n6400_), .A2(new_n6401_), .B(new_n6124_), .ZN(new_n6402_));
  INV_X1     g06210(.I(new_n6386_), .ZN(new_n6403_));
  OAI21_X1   g06211(.A1(new_n6400_), .A2(new_n6403_), .B(\asqrt[57] ), .ZN(new_n6404_));
  NAND3_X1   g06212(.A1(new_n6402_), .A2(new_n6404_), .A3(new_n403_), .ZN(new_n6405_));
  NAND2_X1   g06213(.A1(new_n6405_), .A2(new_n6121_), .ZN(new_n6406_));
  NAND2_X1   g06214(.A1(new_n6402_), .A2(new_n6404_), .ZN(new_n6407_));
  AOI21_X1   g06215(.A1(new_n6407_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n6408_));
  AOI21_X1   g06216(.A1(new_n6408_), .A2(new_n6406_), .B(new_n6397_), .ZN(new_n6409_));
  AOI21_X1   g06217(.A1(new_n6406_), .A2(new_n6390_), .B(new_n339_), .ZN(new_n6410_));
  OAI21_X1   g06218(.A1(new_n6409_), .A2(new_n6410_), .B(\asqrt[60] ), .ZN(new_n6411_));
  AOI21_X1   g06219(.A1(new_n6396_), .A2(new_n6411_), .B(new_n242_), .ZN(new_n6412_));
  NAND3_X1   g06220(.A1(\asqrt[30] ), .A2(new_n6048_), .A3(new_n6064_), .ZN(new_n6413_));
  XOR2_X1    g06221(.A1(new_n6413_), .A2(new_n6090_), .Z(new_n6414_));
  INV_X1     g06222(.I(new_n6414_), .ZN(new_n6415_));
  NAND2_X1   g06223(.A1(new_n6392_), .A2(new_n6394_), .ZN(new_n6416_));
  AOI21_X1   g06224(.A1(new_n6416_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n6417_));
  AOI21_X1   g06225(.A1(new_n6417_), .A2(new_n6396_), .B(new_n6415_), .ZN(new_n6418_));
  OAI21_X1   g06226(.A1(new_n6418_), .A2(new_n6412_), .B(\asqrt[62] ), .ZN(new_n6419_));
  INV_X1     g06227(.I(new_n6419_), .ZN(new_n6420_));
  NOR2_X1    g06228(.A1(new_n6418_), .A2(new_n6412_), .ZN(new_n6421_));
  AOI21_X1   g06229(.A1(new_n6049_), .A2(new_n6070_), .B(new_n6065_), .ZN(new_n6422_));
  NAND2_X1   g06230(.A1(\asqrt[30] ), .A2(new_n6422_), .ZN(new_n6423_));
  XOR2_X1    g06231(.A1(new_n6423_), .A2(new_n6068_), .Z(new_n6424_));
  INV_X1     g06232(.I(new_n6424_), .ZN(new_n6425_));
  AOI21_X1   g06233(.A1(new_n6421_), .A2(new_n234_), .B(new_n6425_), .ZN(new_n6426_));
  OAI21_X1   g06234(.A1(new_n6426_), .A2(new_n6420_), .B(new_n6113_), .ZN(new_n6427_));
  OAI21_X1   g06235(.A1(new_n6427_), .A2(new_n6112_), .B(new_n193_), .ZN(new_n6428_));
  NOR2_X1    g06236(.A1(new_n6426_), .A2(new_n6420_), .ZN(new_n6429_));
  NAND2_X1   g06237(.A1(new_n6429_), .A2(new_n6112_), .ZN(new_n6430_));
  NOR2_X1    g06238(.A1(\asqrt[30] ), .A2(new_n6101_), .ZN(new_n6431_));
  INV_X1     g06239(.I(new_n6431_), .ZN(new_n6432_));
  NAND4_X1   g06240(.A1(new_n6428_), .A2(new_n6110_), .A3(new_n6430_), .A4(new_n6432_), .ZN(\asqrt[29] ));
  AOI21_X1   g06241(.A1(new_n6241_), .A2(new_n6242_), .B(new_n6245_), .ZN(new_n6434_));
  NAND2_X1   g06242(.A1(\asqrt[29] ), .A2(new_n6434_), .ZN(new_n6435_));
  XOR2_X1    g06243(.A1(new_n6435_), .A2(new_n6089_), .Z(new_n6436_));
  INV_X1     g06244(.I(new_n6436_), .ZN(new_n6437_));
  NOR2_X1    g06245(.A1(new_n6240_), .A2(\asqrt[34] ), .ZN(new_n6438_));
  INV_X1     g06246(.I(new_n6112_), .ZN(new_n6439_));
  INV_X1     g06247(.I(new_n6113_), .ZN(new_n6440_));
  INV_X1     g06248(.I(new_n6116_), .ZN(new_n6441_));
  NOR2_X1    g06249(.A1(new_n6409_), .A2(new_n6410_), .ZN(new_n6442_));
  AOI21_X1   g06250(.A1(new_n6442_), .A2(new_n288_), .B(new_n6441_), .ZN(new_n6443_));
  INV_X1     g06251(.I(new_n6411_), .ZN(new_n6444_));
  OAI21_X1   g06252(.A1(new_n6443_), .A2(new_n6444_), .B(\asqrt[61] ), .ZN(new_n6445_));
  NAND2_X1   g06253(.A1(new_n6411_), .A2(new_n242_), .ZN(new_n6446_));
  OAI21_X1   g06254(.A1(new_n6443_), .A2(new_n6446_), .B(new_n6414_), .ZN(new_n6447_));
  NAND3_X1   g06255(.A1(new_n6447_), .A2(new_n6445_), .A3(new_n234_), .ZN(new_n6448_));
  NAND2_X1   g06256(.A1(new_n6448_), .A2(new_n6424_), .ZN(new_n6449_));
  AOI21_X1   g06257(.A1(new_n6449_), .A2(new_n6419_), .B(new_n6440_), .ZN(new_n6450_));
  AOI21_X1   g06258(.A1(new_n6450_), .A2(new_n6439_), .B(\asqrt[63] ), .ZN(new_n6451_));
  NAND2_X1   g06259(.A1(new_n6449_), .A2(new_n6419_), .ZN(new_n6452_));
  NOR2_X1    g06260(.A1(new_n6452_), .A2(new_n6439_), .ZN(new_n6453_));
  NOR4_X1    g06261(.A1(new_n6451_), .A2(new_n6109_), .A3(new_n6453_), .A4(new_n6431_), .ZN(new_n6454_));
  NOR3_X1    g06262(.A1(new_n6454_), .A2(new_n6438_), .A3(new_n6219_), .ZN(new_n6455_));
  XOR2_X1    g06263(.A1(new_n6455_), .A2(new_n6191_), .Z(new_n6456_));
  NOR3_X1    g06264(.A1(new_n6454_), .A2(new_n6237_), .A3(new_n6214_), .ZN(new_n6457_));
  XOR2_X1    g06265(.A1(new_n6457_), .A2(new_n6213_), .Z(new_n6458_));
  INV_X1     g06266(.I(new_n6458_), .ZN(new_n6459_));
  NOR2_X1    g06267(.A1(new_n6208_), .A2(\asqrt[32] ), .ZN(new_n6460_));
  NOR3_X1    g06268(.A1(new_n6454_), .A2(new_n6460_), .A3(new_n6236_), .ZN(new_n6461_));
  XOR2_X1    g06269(.A1(new_n6461_), .A2(new_n6199_), .Z(new_n6462_));
  INV_X1     g06270(.I(new_n6462_), .ZN(new_n6463_));
  NAND3_X1   g06271(.A1(\asqrt[29] ), .A2(new_n6200_), .A3(new_n6201_), .ZN(new_n6464_));
  NOR4_X1    g06272(.A1(new_n6451_), .A2(new_n6106_), .A3(new_n6109_), .A4(new_n6453_), .ZN(new_n6465_));
  INV_X1     g06273(.I(new_n6465_), .ZN(new_n6466_));
  AOI21_X1   g06274(.A1(new_n6464_), .A2(new_n6466_), .B(\a[60] ), .ZN(new_n6467_));
  NOR3_X1    g06275(.A1(new_n6454_), .A2(\a[58] ), .A3(\a[59] ), .ZN(new_n6468_));
  NOR3_X1    g06276(.A1(new_n6468_), .A2(new_n5772_), .A3(new_n6465_), .ZN(new_n6469_));
  NOR2_X1    g06277(.A1(new_n6469_), .A2(new_n6467_), .ZN(new_n6470_));
  INV_X1     g06278(.I(\a[56] ), .ZN(new_n6471_));
  INV_X1     g06279(.I(\a[57] ), .ZN(new_n6472_));
  NAND3_X1   g06280(.A1(new_n6471_), .A2(new_n6472_), .A3(new_n6200_), .ZN(new_n6473_));
  OAI21_X1   g06281(.A1(new_n6454_), .A2(new_n6200_), .B(new_n6473_), .ZN(new_n6474_));
  NAND2_X1   g06282(.A1(new_n6474_), .A2(\asqrt[30] ), .ZN(new_n6475_));
  OAI21_X1   g06283(.A1(new_n6454_), .A2(\a[58] ), .B(\a[59] ), .ZN(new_n6476_));
  NAND2_X1   g06284(.A1(new_n6476_), .A2(new_n6464_), .ZN(new_n6477_));
  NOR2_X1    g06285(.A1(new_n6474_), .A2(\asqrt[30] ), .ZN(new_n6478_));
  OAI21_X1   g06286(.A1(new_n6477_), .A2(new_n6478_), .B(new_n6475_), .ZN(new_n6479_));
  OAI21_X1   g06287(.A1(\asqrt[31] ), .A2(new_n6479_), .B(new_n6470_), .ZN(new_n6480_));
  NAND2_X1   g06288(.A1(new_n6479_), .A2(\asqrt[31] ), .ZN(new_n6481_));
  NAND3_X1   g06289(.A1(new_n6480_), .A2(new_n5435_), .A3(new_n6481_), .ZN(new_n6482_));
  NOR3_X1    g06290(.A1(new_n6454_), .A2(new_n6230_), .A3(new_n6207_), .ZN(new_n6483_));
  XOR2_X1    g06291(.A1(new_n6483_), .A2(new_n6232_), .Z(new_n6484_));
  NAND2_X1   g06292(.A1(new_n6482_), .A2(new_n6484_), .ZN(new_n6485_));
  NAND2_X1   g06293(.A1(new_n6480_), .A2(new_n6481_), .ZN(new_n6486_));
  AOI21_X1   g06294(.A1(new_n6486_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n6487_));
  AOI21_X1   g06295(.A1(new_n6487_), .A2(new_n6485_), .B(new_n6463_), .ZN(new_n6488_));
  OAI21_X1   g06296(.A1(new_n6468_), .A2(new_n6465_), .B(new_n5772_), .ZN(new_n6489_));
  NAND3_X1   g06297(.A1(new_n6464_), .A2(\a[60] ), .A3(new_n6466_), .ZN(new_n6490_));
  NAND2_X1   g06298(.A1(new_n6489_), .A2(new_n6490_), .ZN(new_n6491_));
  NAND2_X1   g06299(.A1(\asqrt[29] ), .A2(\a[58] ), .ZN(new_n6492_));
  AOI21_X1   g06300(.A1(new_n6492_), .A2(new_n6473_), .B(new_n6106_), .ZN(new_n6493_));
  AOI21_X1   g06301(.A1(\asqrt[29] ), .A2(new_n6200_), .B(new_n6201_), .ZN(new_n6494_));
  NOR2_X1    g06302(.A1(new_n6494_), .A2(new_n6468_), .ZN(new_n6495_));
  NAND3_X1   g06303(.A1(new_n6492_), .A2(new_n6106_), .A3(new_n6473_), .ZN(new_n6496_));
  AOI21_X1   g06304(.A1(new_n6495_), .A2(new_n6496_), .B(new_n6493_), .ZN(new_n6497_));
  AOI21_X1   g06305(.A1(new_n6497_), .A2(new_n5750_), .B(new_n6491_), .ZN(new_n6498_));
  NOR2_X1    g06306(.A1(new_n6497_), .A2(new_n5750_), .ZN(new_n6499_));
  OAI21_X1   g06307(.A1(new_n6498_), .A2(new_n6499_), .B(\asqrt[32] ), .ZN(new_n6500_));
  AOI21_X1   g06308(.A1(new_n6485_), .A2(new_n6500_), .B(new_n5110_), .ZN(new_n6501_));
  NOR2_X1    g06309(.A1(new_n6488_), .A2(new_n6501_), .ZN(new_n6502_));
  AOI21_X1   g06310(.A1(new_n6502_), .A2(new_n4810_), .B(new_n6459_), .ZN(new_n6503_));
  OAI21_X1   g06311(.A1(new_n6488_), .A2(new_n6501_), .B(\asqrt[34] ), .ZN(new_n6504_));
  NAND2_X1   g06312(.A1(new_n6504_), .A2(new_n4510_), .ZN(new_n6505_));
  OAI21_X1   g06313(.A1(new_n6503_), .A2(new_n6505_), .B(new_n6456_), .ZN(new_n6506_));
  INV_X1     g06314(.I(new_n6504_), .ZN(new_n6507_));
  OAI21_X1   g06315(.A1(new_n6503_), .A2(new_n6507_), .B(\asqrt[35] ), .ZN(new_n6508_));
  NAND3_X1   g06316(.A1(new_n6506_), .A2(new_n6508_), .A3(new_n4224_), .ZN(new_n6509_));
  INV_X1     g06317(.I(new_n6456_), .ZN(new_n6510_));
  NOR2_X1    g06318(.A1(new_n6498_), .A2(new_n6499_), .ZN(new_n6511_));
  INV_X1     g06319(.I(new_n6484_), .ZN(new_n6512_));
  AOI21_X1   g06320(.A1(new_n6511_), .A2(new_n5435_), .B(new_n6512_), .ZN(new_n6513_));
  NAND2_X1   g06321(.A1(new_n6500_), .A2(new_n5110_), .ZN(new_n6514_));
  OAI21_X1   g06322(.A1(new_n6513_), .A2(new_n6514_), .B(new_n6462_), .ZN(new_n6515_));
  INV_X1     g06323(.I(new_n6500_), .ZN(new_n6516_));
  OAI21_X1   g06324(.A1(new_n6513_), .A2(new_n6516_), .B(\asqrt[33] ), .ZN(new_n6517_));
  NAND3_X1   g06325(.A1(new_n6515_), .A2(new_n6517_), .A3(new_n4810_), .ZN(new_n6518_));
  NAND2_X1   g06326(.A1(new_n6518_), .A2(new_n6458_), .ZN(new_n6519_));
  NAND2_X1   g06327(.A1(new_n6515_), .A2(new_n6517_), .ZN(new_n6520_));
  AOI21_X1   g06328(.A1(new_n6520_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n6521_));
  AOI21_X1   g06329(.A1(new_n6521_), .A2(new_n6519_), .B(new_n6510_), .ZN(new_n6522_));
  AOI21_X1   g06330(.A1(new_n6519_), .A2(new_n6504_), .B(new_n4510_), .ZN(new_n6523_));
  OAI21_X1   g06331(.A1(new_n6522_), .A2(new_n6523_), .B(\asqrt[36] ), .ZN(new_n6524_));
  NAND2_X1   g06332(.A1(new_n6452_), .A2(new_n6112_), .ZN(new_n6525_));
  NOR2_X1    g06333(.A1(new_n6454_), .A2(new_n6112_), .ZN(new_n6526_));
  NAND2_X1   g06334(.A1(new_n6526_), .A2(new_n6429_), .ZN(new_n6527_));
  AOI21_X1   g06335(.A1(new_n6527_), .A2(new_n6525_), .B(new_n193_), .ZN(new_n6528_));
  INV_X1     g06336(.I(new_n6528_), .ZN(new_n6529_));
  NAND3_X1   g06337(.A1(\asqrt[29] ), .A2(new_n6419_), .A3(new_n6448_), .ZN(new_n6530_));
  XOR2_X1    g06338(.A1(new_n6530_), .A2(new_n6424_), .Z(new_n6531_));
  AOI21_X1   g06339(.A1(new_n6526_), .A2(new_n6452_), .B(new_n6453_), .ZN(new_n6532_));
  OAI21_X1   g06340(.A1(new_n6389_), .A2(new_n6391_), .B(new_n6394_), .ZN(new_n6533_));
  NOR2_X1    g06341(.A1(new_n6454_), .A2(new_n6533_), .ZN(new_n6534_));
  XOR2_X1    g06342(.A1(new_n6534_), .A2(new_n6118_), .Z(new_n6535_));
  NAND3_X1   g06343(.A1(\asqrt[29] ), .A2(new_n6405_), .A3(new_n6390_), .ZN(new_n6536_));
  XOR2_X1    g06344(.A1(new_n6536_), .A2(new_n6122_), .Z(new_n6537_));
  OAI21_X1   g06345(.A1(new_n6400_), .A2(new_n6401_), .B(new_n6404_), .ZN(new_n6538_));
  NOR2_X1    g06346(.A1(new_n6454_), .A2(new_n6538_), .ZN(new_n6539_));
  XOR2_X1    g06347(.A1(new_n6539_), .A2(new_n6124_), .Z(new_n6540_));
  INV_X1     g06348(.I(new_n6540_), .ZN(new_n6541_));
  NAND3_X1   g06349(.A1(\asqrt[29] ), .A2(new_n6367_), .A3(new_n6386_), .ZN(new_n6542_));
  XOR2_X1    g06350(.A1(new_n6542_), .A2(new_n6398_), .Z(new_n6543_));
  INV_X1     g06351(.I(new_n6543_), .ZN(new_n6544_));
  OAI21_X1   g06352(.A1(new_n6361_), .A2(new_n6363_), .B(new_n6366_), .ZN(new_n6545_));
  NOR2_X1    g06353(.A1(new_n6454_), .A2(new_n6545_), .ZN(new_n6546_));
  XOR2_X1    g06354(.A1(new_n6546_), .A2(new_n6130_), .Z(new_n6547_));
  NAND3_X1   g06355(.A1(\asqrt[29] ), .A2(new_n6380_), .A3(new_n6362_), .ZN(new_n6548_));
  XOR2_X1    g06356(.A1(new_n6548_), .A2(new_n6134_), .Z(new_n6549_));
  OAI21_X1   g06357(.A1(new_n6375_), .A2(new_n6376_), .B(new_n6379_), .ZN(new_n6550_));
  NOR2_X1    g06358(.A1(new_n6454_), .A2(new_n6550_), .ZN(new_n6551_));
  XOR2_X1    g06359(.A1(new_n6551_), .A2(new_n6136_), .Z(new_n6552_));
  INV_X1     g06360(.I(new_n6552_), .ZN(new_n6553_));
  NAND3_X1   g06361(.A1(\asqrt[29] ), .A2(new_n6339_), .A3(new_n6358_), .ZN(new_n6554_));
  XOR2_X1    g06362(.A1(new_n6554_), .A2(new_n6373_), .Z(new_n6555_));
  INV_X1     g06363(.I(new_n6555_), .ZN(new_n6556_));
  OAI21_X1   g06364(.A1(new_n6333_), .A2(new_n6335_), .B(new_n6338_), .ZN(new_n6557_));
  NOR2_X1    g06365(.A1(new_n6454_), .A2(new_n6557_), .ZN(new_n6558_));
  XOR2_X1    g06366(.A1(new_n6558_), .A2(new_n6142_), .Z(new_n6559_));
  NAND3_X1   g06367(.A1(\asqrt[29] ), .A2(new_n6352_), .A3(new_n6334_), .ZN(new_n6560_));
  XOR2_X1    g06368(.A1(new_n6560_), .A2(new_n6146_), .Z(new_n6561_));
  OAI21_X1   g06369(.A1(new_n6347_), .A2(new_n6348_), .B(new_n6351_), .ZN(new_n6562_));
  NOR2_X1    g06370(.A1(new_n6454_), .A2(new_n6562_), .ZN(new_n6563_));
  XOR2_X1    g06371(.A1(new_n6563_), .A2(new_n6148_), .Z(new_n6564_));
  INV_X1     g06372(.I(new_n6564_), .ZN(new_n6565_));
  NAND3_X1   g06373(.A1(\asqrt[29] ), .A2(new_n6311_), .A3(new_n6330_), .ZN(new_n6566_));
  XOR2_X1    g06374(.A1(new_n6566_), .A2(new_n6345_), .Z(new_n6567_));
  INV_X1     g06375(.I(new_n6567_), .ZN(new_n6568_));
  OAI21_X1   g06376(.A1(new_n6305_), .A2(new_n6307_), .B(new_n6310_), .ZN(new_n6569_));
  NOR2_X1    g06377(.A1(new_n6454_), .A2(new_n6569_), .ZN(new_n6570_));
  XOR2_X1    g06378(.A1(new_n6570_), .A2(new_n6154_), .Z(new_n6571_));
  NAND3_X1   g06379(.A1(\asqrt[29] ), .A2(new_n6324_), .A3(new_n6306_), .ZN(new_n6572_));
  XOR2_X1    g06380(.A1(new_n6572_), .A2(new_n6158_), .Z(new_n6573_));
  OAI21_X1   g06381(.A1(new_n6319_), .A2(new_n6320_), .B(new_n6323_), .ZN(new_n6574_));
  NOR2_X1    g06382(.A1(new_n6454_), .A2(new_n6574_), .ZN(new_n6575_));
  XOR2_X1    g06383(.A1(new_n6575_), .A2(new_n6160_), .Z(new_n6576_));
  INV_X1     g06384(.I(new_n6576_), .ZN(new_n6577_));
  NAND3_X1   g06385(.A1(\asqrt[29] ), .A2(new_n6283_), .A3(new_n6302_), .ZN(new_n6578_));
  XOR2_X1    g06386(.A1(new_n6578_), .A2(new_n6317_), .Z(new_n6579_));
  INV_X1     g06387(.I(new_n6579_), .ZN(new_n6580_));
  OAI21_X1   g06388(.A1(new_n6277_), .A2(new_n6279_), .B(new_n6282_), .ZN(new_n6581_));
  NOR2_X1    g06389(.A1(new_n6454_), .A2(new_n6581_), .ZN(new_n6582_));
  XOR2_X1    g06390(.A1(new_n6582_), .A2(new_n6166_), .Z(new_n6583_));
  NAND3_X1   g06391(.A1(\asqrt[29] ), .A2(new_n6296_), .A3(new_n6278_), .ZN(new_n6584_));
  XOR2_X1    g06392(.A1(new_n6584_), .A2(new_n6170_), .Z(new_n6585_));
  OAI21_X1   g06393(.A1(new_n6291_), .A2(new_n6292_), .B(new_n6295_), .ZN(new_n6586_));
  NOR2_X1    g06394(.A1(new_n6454_), .A2(new_n6586_), .ZN(new_n6587_));
  XOR2_X1    g06395(.A1(new_n6587_), .A2(new_n6172_), .Z(new_n6588_));
  INV_X1     g06396(.I(new_n6588_), .ZN(new_n6589_));
  NAND3_X1   g06397(.A1(\asqrt[29] ), .A2(new_n6255_), .A3(new_n6274_), .ZN(new_n6590_));
  XOR2_X1    g06398(.A1(new_n6590_), .A2(new_n6289_), .Z(new_n6591_));
  INV_X1     g06399(.I(new_n6591_), .ZN(new_n6592_));
  OAI21_X1   g06400(.A1(new_n6249_), .A2(new_n6251_), .B(new_n6254_), .ZN(new_n6593_));
  NOR2_X1    g06401(.A1(new_n6454_), .A2(new_n6593_), .ZN(new_n6594_));
  XOR2_X1    g06402(.A1(new_n6594_), .A2(new_n6178_), .Z(new_n6595_));
  NAND3_X1   g06403(.A1(\asqrt[29] ), .A2(new_n6268_), .A3(new_n6250_), .ZN(new_n6596_));
  XOR2_X1    g06404(.A1(new_n6596_), .A2(new_n6182_), .Z(new_n6597_));
  OAI21_X1   g06405(.A1(new_n6263_), .A2(new_n6264_), .B(new_n6267_), .ZN(new_n6598_));
  NOR2_X1    g06406(.A1(new_n6454_), .A2(new_n6598_), .ZN(new_n6599_));
  XOR2_X1    g06407(.A1(new_n6599_), .A2(new_n6184_), .Z(new_n6600_));
  INV_X1     g06408(.I(new_n6600_), .ZN(new_n6601_));
  NAND3_X1   g06409(.A1(\asqrt[29] ), .A2(new_n6221_), .A3(new_n6246_), .ZN(new_n6602_));
  XOR2_X1    g06410(.A1(new_n6602_), .A2(new_n6261_), .Z(new_n6603_));
  INV_X1     g06411(.I(new_n6603_), .ZN(new_n6604_));
  NAND2_X1   g06412(.A1(new_n6509_), .A2(new_n6436_), .ZN(new_n6605_));
  NAND2_X1   g06413(.A1(new_n6506_), .A2(new_n6508_), .ZN(new_n6606_));
  AOI21_X1   g06414(.A1(new_n6606_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n6607_));
  AOI21_X1   g06415(.A1(new_n6607_), .A2(new_n6605_), .B(new_n6604_), .ZN(new_n6608_));
  AOI21_X1   g06416(.A1(new_n6605_), .A2(new_n6524_), .B(new_n3928_), .ZN(new_n6609_));
  NOR2_X1    g06417(.A1(new_n6608_), .A2(new_n6609_), .ZN(new_n6610_));
  AOI21_X1   g06418(.A1(new_n6610_), .A2(new_n3675_), .B(new_n6601_), .ZN(new_n6611_));
  OAI21_X1   g06419(.A1(new_n6608_), .A2(new_n6609_), .B(\asqrt[38] ), .ZN(new_n6612_));
  NAND2_X1   g06420(.A1(new_n6612_), .A2(new_n3400_), .ZN(new_n6613_));
  OAI21_X1   g06421(.A1(new_n6611_), .A2(new_n6613_), .B(new_n6597_), .ZN(new_n6614_));
  INV_X1     g06422(.I(new_n6612_), .ZN(new_n6615_));
  OAI21_X1   g06423(.A1(new_n6611_), .A2(new_n6615_), .B(\asqrt[39] ), .ZN(new_n6616_));
  NAND3_X1   g06424(.A1(new_n6614_), .A2(new_n6616_), .A3(new_n3167_), .ZN(new_n6617_));
  NAND2_X1   g06425(.A1(new_n6617_), .A2(new_n6595_), .ZN(new_n6618_));
  NAND2_X1   g06426(.A1(new_n6614_), .A2(new_n6616_), .ZN(new_n6619_));
  AOI21_X1   g06427(.A1(new_n6619_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n6620_));
  AOI21_X1   g06428(.A1(new_n6620_), .A2(new_n6618_), .B(new_n6592_), .ZN(new_n6621_));
  INV_X1     g06429(.I(new_n6597_), .ZN(new_n6622_));
  NOR2_X1    g06430(.A1(new_n6522_), .A2(new_n6523_), .ZN(new_n6623_));
  AOI21_X1   g06431(.A1(new_n6623_), .A2(new_n4224_), .B(new_n6437_), .ZN(new_n6624_));
  NAND2_X1   g06432(.A1(new_n6524_), .A2(new_n3928_), .ZN(new_n6625_));
  OAI21_X1   g06433(.A1(new_n6624_), .A2(new_n6625_), .B(new_n6603_), .ZN(new_n6626_));
  INV_X1     g06434(.I(new_n6524_), .ZN(new_n6627_));
  OAI21_X1   g06435(.A1(new_n6624_), .A2(new_n6627_), .B(\asqrt[37] ), .ZN(new_n6628_));
  NAND3_X1   g06436(.A1(new_n6626_), .A2(new_n6628_), .A3(new_n3675_), .ZN(new_n6629_));
  NAND2_X1   g06437(.A1(new_n6629_), .A2(new_n6600_), .ZN(new_n6630_));
  NAND2_X1   g06438(.A1(new_n6626_), .A2(new_n6628_), .ZN(new_n6631_));
  AOI21_X1   g06439(.A1(new_n6631_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n6632_));
  AOI21_X1   g06440(.A1(new_n6632_), .A2(new_n6630_), .B(new_n6622_), .ZN(new_n6633_));
  AOI21_X1   g06441(.A1(new_n6630_), .A2(new_n6612_), .B(new_n3400_), .ZN(new_n6634_));
  OAI21_X1   g06442(.A1(new_n6633_), .A2(new_n6634_), .B(\asqrt[40] ), .ZN(new_n6635_));
  AOI21_X1   g06443(.A1(new_n6618_), .A2(new_n6635_), .B(new_n2912_), .ZN(new_n6636_));
  NOR2_X1    g06444(.A1(new_n6621_), .A2(new_n6636_), .ZN(new_n6637_));
  AOI21_X1   g06445(.A1(new_n6637_), .A2(new_n2699_), .B(new_n6589_), .ZN(new_n6638_));
  OAI21_X1   g06446(.A1(new_n6621_), .A2(new_n6636_), .B(\asqrt[42] ), .ZN(new_n6639_));
  NAND2_X1   g06447(.A1(new_n6639_), .A2(new_n2464_), .ZN(new_n6640_));
  OAI21_X1   g06448(.A1(new_n6638_), .A2(new_n6640_), .B(new_n6585_), .ZN(new_n6641_));
  INV_X1     g06449(.I(new_n6639_), .ZN(new_n6642_));
  OAI21_X1   g06450(.A1(new_n6638_), .A2(new_n6642_), .B(\asqrt[43] ), .ZN(new_n6643_));
  NAND3_X1   g06451(.A1(new_n6641_), .A2(new_n6643_), .A3(new_n2271_), .ZN(new_n6644_));
  NAND2_X1   g06452(.A1(new_n6644_), .A2(new_n6583_), .ZN(new_n6645_));
  NAND2_X1   g06453(.A1(new_n6641_), .A2(new_n6643_), .ZN(new_n6646_));
  AOI21_X1   g06454(.A1(new_n6646_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n6647_));
  AOI21_X1   g06455(.A1(new_n6647_), .A2(new_n6645_), .B(new_n6580_), .ZN(new_n6648_));
  INV_X1     g06456(.I(new_n6585_), .ZN(new_n6649_));
  INV_X1     g06457(.I(new_n6595_), .ZN(new_n6650_));
  NOR2_X1    g06458(.A1(new_n6633_), .A2(new_n6634_), .ZN(new_n6651_));
  AOI21_X1   g06459(.A1(new_n6651_), .A2(new_n3167_), .B(new_n6650_), .ZN(new_n6652_));
  NAND2_X1   g06460(.A1(new_n6635_), .A2(new_n2912_), .ZN(new_n6653_));
  OAI21_X1   g06461(.A1(new_n6652_), .A2(new_n6653_), .B(new_n6591_), .ZN(new_n6654_));
  INV_X1     g06462(.I(new_n6635_), .ZN(new_n6655_));
  OAI21_X1   g06463(.A1(new_n6652_), .A2(new_n6655_), .B(\asqrt[41] ), .ZN(new_n6656_));
  NAND3_X1   g06464(.A1(new_n6654_), .A2(new_n6656_), .A3(new_n2699_), .ZN(new_n6657_));
  NAND2_X1   g06465(.A1(new_n6657_), .A2(new_n6588_), .ZN(new_n6658_));
  NAND2_X1   g06466(.A1(new_n6654_), .A2(new_n6656_), .ZN(new_n6659_));
  AOI21_X1   g06467(.A1(new_n6659_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n6660_));
  AOI21_X1   g06468(.A1(new_n6660_), .A2(new_n6658_), .B(new_n6649_), .ZN(new_n6661_));
  AOI21_X1   g06469(.A1(new_n6658_), .A2(new_n6639_), .B(new_n2464_), .ZN(new_n6662_));
  OAI21_X1   g06470(.A1(new_n6661_), .A2(new_n6662_), .B(\asqrt[44] ), .ZN(new_n6663_));
  AOI21_X1   g06471(.A1(new_n6645_), .A2(new_n6663_), .B(new_n2072_), .ZN(new_n6664_));
  NOR2_X1    g06472(.A1(new_n6648_), .A2(new_n6664_), .ZN(new_n6665_));
  AOI21_X1   g06473(.A1(new_n6665_), .A2(new_n1884_), .B(new_n6577_), .ZN(new_n6666_));
  OAI21_X1   g06474(.A1(new_n6648_), .A2(new_n6664_), .B(\asqrt[46] ), .ZN(new_n6667_));
  NAND2_X1   g06475(.A1(new_n6667_), .A2(new_n1688_), .ZN(new_n6668_));
  OAI21_X1   g06476(.A1(new_n6666_), .A2(new_n6668_), .B(new_n6573_), .ZN(new_n6669_));
  INV_X1     g06477(.I(new_n6667_), .ZN(new_n6670_));
  OAI21_X1   g06478(.A1(new_n6666_), .A2(new_n6670_), .B(\asqrt[47] ), .ZN(new_n6671_));
  NAND3_X1   g06479(.A1(new_n6669_), .A2(new_n6671_), .A3(new_n1533_), .ZN(new_n6672_));
  NAND2_X1   g06480(.A1(new_n6672_), .A2(new_n6571_), .ZN(new_n6673_));
  NAND2_X1   g06481(.A1(new_n6669_), .A2(new_n6671_), .ZN(new_n6674_));
  AOI21_X1   g06482(.A1(new_n6674_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n6675_));
  AOI21_X1   g06483(.A1(new_n6675_), .A2(new_n6673_), .B(new_n6568_), .ZN(new_n6676_));
  INV_X1     g06484(.I(new_n6573_), .ZN(new_n6677_));
  INV_X1     g06485(.I(new_n6583_), .ZN(new_n6678_));
  NOR2_X1    g06486(.A1(new_n6661_), .A2(new_n6662_), .ZN(new_n6679_));
  AOI21_X1   g06487(.A1(new_n6679_), .A2(new_n2271_), .B(new_n6678_), .ZN(new_n6680_));
  NAND2_X1   g06488(.A1(new_n6663_), .A2(new_n2072_), .ZN(new_n6681_));
  OAI21_X1   g06489(.A1(new_n6680_), .A2(new_n6681_), .B(new_n6579_), .ZN(new_n6682_));
  INV_X1     g06490(.I(new_n6663_), .ZN(new_n6683_));
  OAI21_X1   g06491(.A1(new_n6680_), .A2(new_n6683_), .B(\asqrt[45] ), .ZN(new_n6684_));
  NAND3_X1   g06492(.A1(new_n6682_), .A2(new_n6684_), .A3(new_n1884_), .ZN(new_n6685_));
  NAND2_X1   g06493(.A1(new_n6685_), .A2(new_n6576_), .ZN(new_n6686_));
  NAND2_X1   g06494(.A1(new_n6682_), .A2(new_n6684_), .ZN(new_n6687_));
  AOI21_X1   g06495(.A1(new_n6687_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n6688_));
  AOI21_X1   g06496(.A1(new_n6688_), .A2(new_n6686_), .B(new_n6677_), .ZN(new_n6689_));
  AOI21_X1   g06497(.A1(new_n6686_), .A2(new_n6667_), .B(new_n1688_), .ZN(new_n6690_));
  OAI21_X1   g06498(.A1(new_n6689_), .A2(new_n6690_), .B(\asqrt[48] ), .ZN(new_n6691_));
  AOI21_X1   g06499(.A1(new_n6673_), .A2(new_n6691_), .B(new_n1368_), .ZN(new_n6692_));
  NOR2_X1    g06500(.A1(new_n6676_), .A2(new_n6692_), .ZN(new_n6693_));
  AOI21_X1   g06501(.A1(new_n6693_), .A2(new_n1228_), .B(new_n6565_), .ZN(new_n6694_));
  OAI21_X1   g06502(.A1(new_n6676_), .A2(new_n6692_), .B(\asqrt[50] ), .ZN(new_n6695_));
  NAND2_X1   g06503(.A1(new_n6695_), .A2(new_n1088_), .ZN(new_n6696_));
  OAI21_X1   g06504(.A1(new_n6694_), .A2(new_n6696_), .B(new_n6561_), .ZN(new_n6697_));
  INV_X1     g06505(.I(new_n6695_), .ZN(new_n6698_));
  OAI21_X1   g06506(.A1(new_n6694_), .A2(new_n6698_), .B(\asqrt[51] ), .ZN(new_n6699_));
  NAND3_X1   g06507(.A1(new_n6697_), .A2(new_n6699_), .A3(new_n962_), .ZN(new_n6700_));
  NAND2_X1   g06508(.A1(new_n6700_), .A2(new_n6559_), .ZN(new_n6701_));
  NAND2_X1   g06509(.A1(new_n6697_), .A2(new_n6699_), .ZN(new_n6702_));
  AOI21_X1   g06510(.A1(new_n6702_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n6703_));
  AOI21_X1   g06511(.A1(new_n6703_), .A2(new_n6701_), .B(new_n6556_), .ZN(new_n6704_));
  INV_X1     g06512(.I(new_n6561_), .ZN(new_n6705_));
  INV_X1     g06513(.I(new_n6571_), .ZN(new_n6706_));
  NOR2_X1    g06514(.A1(new_n6689_), .A2(new_n6690_), .ZN(new_n6707_));
  AOI21_X1   g06515(.A1(new_n6707_), .A2(new_n1533_), .B(new_n6706_), .ZN(new_n6708_));
  NAND2_X1   g06516(.A1(new_n6691_), .A2(new_n1368_), .ZN(new_n6709_));
  OAI21_X1   g06517(.A1(new_n6708_), .A2(new_n6709_), .B(new_n6567_), .ZN(new_n6710_));
  INV_X1     g06518(.I(new_n6691_), .ZN(new_n6711_));
  OAI21_X1   g06519(.A1(new_n6708_), .A2(new_n6711_), .B(\asqrt[49] ), .ZN(new_n6712_));
  NAND3_X1   g06520(.A1(new_n6710_), .A2(new_n6712_), .A3(new_n1228_), .ZN(new_n6713_));
  NAND2_X1   g06521(.A1(new_n6713_), .A2(new_n6564_), .ZN(new_n6714_));
  NAND2_X1   g06522(.A1(new_n6710_), .A2(new_n6712_), .ZN(new_n6715_));
  AOI21_X1   g06523(.A1(new_n6715_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n6716_));
  AOI21_X1   g06524(.A1(new_n6716_), .A2(new_n6714_), .B(new_n6705_), .ZN(new_n6717_));
  AOI21_X1   g06525(.A1(new_n6714_), .A2(new_n6695_), .B(new_n1088_), .ZN(new_n6718_));
  OAI21_X1   g06526(.A1(new_n6717_), .A2(new_n6718_), .B(\asqrt[52] ), .ZN(new_n6719_));
  AOI21_X1   g06527(.A1(new_n6701_), .A2(new_n6719_), .B(new_n842_), .ZN(new_n6720_));
  NOR2_X1    g06528(.A1(new_n6704_), .A2(new_n6720_), .ZN(new_n6721_));
  AOI21_X1   g06529(.A1(new_n6721_), .A2(new_n720_), .B(new_n6553_), .ZN(new_n6722_));
  OAI21_X1   g06530(.A1(new_n6704_), .A2(new_n6720_), .B(\asqrt[54] ), .ZN(new_n6723_));
  NAND2_X1   g06531(.A1(new_n6723_), .A2(new_n630_), .ZN(new_n6724_));
  OAI21_X1   g06532(.A1(new_n6722_), .A2(new_n6724_), .B(new_n6549_), .ZN(new_n6725_));
  INV_X1     g06533(.I(new_n6723_), .ZN(new_n6726_));
  OAI21_X1   g06534(.A1(new_n6722_), .A2(new_n6726_), .B(\asqrt[55] ), .ZN(new_n6727_));
  NAND3_X1   g06535(.A1(new_n6725_), .A2(new_n6727_), .A3(new_n545_), .ZN(new_n6728_));
  NAND2_X1   g06536(.A1(new_n6728_), .A2(new_n6547_), .ZN(new_n6729_));
  NAND2_X1   g06537(.A1(new_n6725_), .A2(new_n6727_), .ZN(new_n6730_));
  AOI21_X1   g06538(.A1(new_n6730_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n6731_));
  AOI21_X1   g06539(.A1(new_n6731_), .A2(new_n6729_), .B(new_n6544_), .ZN(new_n6732_));
  INV_X1     g06540(.I(new_n6549_), .ZN(new_n6733_));
  INV_X1     g06541(.I(new_n6559_), .ZN(new_n6734_));
  NOR2_X1    g06542(.A1(new_n6717_), .A2(new_n6718_), .ZN(new_n6735_));
  AOI21_X1   g06543(.A1(new_n6735_), .A2(new_n962_), .B(new_n6734_), .ZN(new_n6736_));
  NAND2_X1   g06544(.A1(new_n6719_), .A2(new_n842_), .ZN(new_n6737_));
  OAI21_X1   g06545(.A1(new_n6736_), .A2(new_n6737_), .B(new_n6555_), .ZN(new_n6738_));
  INV_X1     g06546(.I(new_n6719_), .ZN(new_n6739_));
  OAI21_X1   g06547(.A1(new_n6736_), .A2(new_n6739_), .B(\asqrt[53] ), .ZN(new_n6740_));
  NAND3_X1   g06548(.A1(new_n6738_), .A2(new_n6740_), .A3(new_n720_), .ZN(new_n6741_));
  NAND2_X1   g06549(.A1(new_n6741_), .A2(new_n6552_), .ZN(new_n6742_));
  NAND2_X1   g06550(.A1(new_n6738_), .A2(new_n6740_), .ZN(new_n6743_));
  AOI21_X1   g06551(.A1(new_n6743_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n6744_));
  AOI21_X1   g06552(.A1(new_n6744_), .A2(new_n6742_), .B(new_n6733_), .ZN(new_n6745_));
  AOI21_X1   g06553(.A1(new_n6742_), .A2(new_n6723_), .B(new_n630_), .ZN(new_n6746_));
  OAI21_X1   g06554(.A1(new_n6745_), .A2(new_n6746_), .B(\asqrt[56] ), .ZN(new_n6747_));
  AOI21_X1   g06555(.A1(new_n6729_), .A2(new_n6747_), .B(new_n450_), .ZN(new_n6748_));
  NOR2_X1    g06556(.A1(new_n6732_), .A2(new_n6748_), .ZN(new_n6749_));
  AOI21_X1   g06557(.A1(new_n6749_), .A2(new_n403_), .B(new_n6541_), .ZN(new_n6750_));
  OAI21_X1   g06558(.A1(new_n6732_), .A2(new_n6748_), .B(\asqrt[58] ), .ZN(new_n6751_));
  NAND2_X1   g06559(.A1(new_n6751_), .A2(new_n339_), .ZN(new_n6752_));
  OAI21_X1   g06560(.A1(new_n6750_), .A2(new_n6752_), .B(new_n6537_), .ZN(new_n6753_));
  INV_X1     g06561(.I(new_n6751_), .ZN(new_n6754_));
  OAI21_X1   g06562(.A1(new_n6750_), .A2(new_n6754_), .B(\asqrt[59] ), .ZN(new_n6755_));
  NAND3_X1   g06563(.A1(new_n6753_), .A2(new_n6755_), .A3(new_n288_), .ZN(new_n6756_));
  NAND2_X1   g06564(.A1(new_n6756_), .A2(new_n6535_), .ZN(new_n6757_));
  INV_X1     g06565(.I(new_n6537_), .ZN(new_n6758_));
  INV_X1     g06566(.I(new_n6547_), .ZN(new_n6759_));
  NOR2_X1    g06567(.A1(new_n6745_), .A2(new_n6746_), .ZN(new_n6760_));
  AOI21_X1   g06568(.A1(new_n6760_), .A2(new_n545_), .B(new_n6759_), .ZN(new_n6761_));
  NAND2_X1   g06569(.A1(new_n6747_), .A2(new_n450_), .ZN(new_n6762_));
  OAI21_X1   g06570(.A1(new_n6761_), .A2(new_n6762_), .B(new_n6543_), .ZN(new_n6763_));
  INV_X1     g06571(.I(new_n6747_), .ZN(new_n6764_));
  OAI21_X1   g06572(.A1(new_n6761_), .A2(new_n6764_), .B(\asqrt[57] ), .ZN(new_n6765_));
  NAND3_X1   g06573(.A1(new_n6763_), .A2(new_n6765_), .A3(new_n403_), .ZN(new_n6766_));
  NAND2_X1   g06574(.A1(new_n6766_), .A2(new_n6540_), .ZN(new_n6767_));
  NAND2_X1   g06575(.A1(new_n6763_), .A2(new_n6765_), .ZN(new_n6768_));
  AOI21_X1   g06576(.A1(new_n6768_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n6769_));
  AOI21_X1   g06577(.A1(new_n6769_), .A2(new_n6767_), .B(new_n6758_), .ZN(new_n6770_));
  AOI21_X1   g06578(.A1(new_n6767_), .A2(new_n6751_), .B(new_n339_), .ZN(new_n6771_));
  OAI21_X1   g06579(.A1(new_n6770_), .A2(new_n6771_), .B(\asqrt[60] ), .ZN(new_n6772_));
  AOI21_X1   g06580(.A1(new_n6757_), .A2(new_n6772_), .B(new_n242_), .ZN(new_n6773_));
  NAND3_X1   g06581(.A1(\asqrt[29] ), .A2(new_n6395_), .A3(new_n6411_), .ZN(new_n6774_));
  XOR2_X1    g06582(.A1(new_n6774_), .A2(new_n6441_), .Z(new_n6775_));
  INV_X1     g06583(.I(new_n6775_), .ZN(new_n6776_));
  NAND2_X1   g06584(.A1(new_n6753_), .A2(new_n6755_), .ZN(new_n6777_));
  AOI21_X1   g06585(.A1(new_n6777_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n6778_));
  AOI21_X1   g06586(.A1(new_n6778_), .A2(new_n6757_), .B(new_n6776_), .ZN(new_n6779_));
  OAI21_X1   g06587(.A1(new_n6779_), .A2(new_n6773_), .B(\asqrt[62] ), .ZN(new_n6780_));
  INV_X1     g06588(.I(new_n6780_), .ZN(new_n6781_));
  NOR2_X1    g06589(.A1(new_n6779_), .A2(new_n6773_), .ZN(new_n6782_));
  AOI21_X1   g06590(.A1(new_n6396_), .A2(new_n6417_), .B(new_n6412_), .ZN(new_n6783_));
  NAND2_X1   g06591(.A1(\asqrt[29] ), .A2(new_n6783_), .ZN(new_n6784_));
  XOR2_X1    g06592(.A1(new_n6784_), .A2(new_n6415_), .Z(new_n6785_));
  INV_X1     g06593(.I(new_n6785_), .ZN(new_n6786_));
  AOI21_X1   g06594(.A1(new_n6782_), .A2(new_n234_), .B(new_n6786_), .ZN(new_n6787_));
  OAI21_X1   g06595(.A1(new_n6787_), .A2(new_n6781_), .B(new_n6532_), .ZN(new_n6788_));
  OAI21_X1   g06596(.A1(new_n6788_), .A2(new_n6531_), .B(new_n193_), .ZN(new_n6789_));
  NOR2_X1    g06597(.A1(new_n6787_), .A2(new_n6781_), .ZN(new_n6790_));
  NAND2_X1   g06598(.A1(new_n6790_), .A2(new_n6531_), .ZN(new_n6791_));
  NOR2_X1    g06599(.A1(\asqrt[29] ), .A2(new_n6439_), .ZN(new_n6792_));
  INV_X1     g06600(.I(new_n6792_), .ZN(new_n6793_));
  NAND4_X1   g06601(.A1(new_n6789_), .A2(new_n6529_), .A3(new_n6791_), .A4(new_n6793_), .ZN(\asqrt[28] ));
  NAND3_X1   g06602(.A1(\asqrt[28] ), .A2(new_n6509_), .A3(new_n6524_), .ZN(new_n6795_));
  XOR2_X1    g06603(.A1(new_n6795_), .A2(new_n6437_), .Z(new_n6796_));
  INV_X1     g06604(.I(new_n6535_), .ZN(new_n6797_));
  NOR2_X1    g06605(.A1(new_n6770_), .A2(new_n6771_), .ZN(new_n6798_));
  AOI21_X1   g06606(.A1(new_n6798_), .A2(new_n288_), .B(new_n6797_), .ZN(new_n6799_));
  INV_X1     g06607(.I(new_n6772_), .ZN(new_n6800_));
  OAI21_X1   g06608(.A1(new_n6799_), .A2(new_n6800_), .B(\asqrt[61] ), .ZN(new_n6801_));
  NAND2_X1   g06609(.A1(new_n6772_), .A2(new_n242_), .ZN(new_n6802_));
  OAI21_X1   g06610(.A1(new_n6799_), .A2(new_n6802_), .B(new_n6775_), .ZN(new_n6803_));
  NAND3_X1   g06611(.A1(new_n6803_), .A2(new_n6801_), .A3(new_n234_), .ZN(new_n6804_));
  NAND2_X1   g06612(.A1(new_n6804_), .A2(new_n6785_), .ZN(new_n6805_));
  NAND2_X1   g06613(.A1(new_n6805_), .A2(new_n6780_), .ZN(new_n6806_));
  NAND2_X1   g06614(.A1(new_n6806_), .A2(new_n6531_), .ZN(new_n6807_));
  INV_X1     g06615(.I(new_n6531_), .ZN(new_n6808_));
  INV_X1     g06616(.I(new_n6532_), .ZN(new_n6809_));
  AOI21_X1   g06617(.A1(new_n6805_), .A2(new_n6780_), .B(new_n6809_), .ZN(new_n6810_));
  AOI21_X1   g06618(.A1(new_n6810_), .A2(new_n6808_), .B(\asqrt[63] ), .ZN(new_n6811_));
  NOR2_X1    g06619(.A1(new_n6806_), .A2(new_n6808_), .ZN(new_n6812_));
  NOR4_X1    g06620(.A1(new_n6811_), .A2(new_n6528_), .A3(new_n6812_), .A4(new_n6792_), .ZN(new_n6813_));
  NOR2_X1    g06621(.A1(new_n6813_), .A2(new_n6531_), .ZN(new_n6814_));
  NAND2_X1   g06622(.A1(new_n6814_), .A2(new_n6790_), .ZN(new_n6815_));
  AOI21_X1   g06623(.A1(new_n6815_), .A2(new_n6807_), .B(new_n193_), .ZN(new_n6816_));
  NAND3_X1   g06624(.A1(\asqrt[28] ), .A2(new_n6780_), .A3(new_n6804_), .ZN(new_n6817_));
  XOR2_X1    g06625(.A1(new_n6817_), .A2(new_n6785_), .Z(new_n6818_));
  INV_X1     g06626(.I(new_n6818_), .ZN(new_n6819_));
  AOI21_X1   g06627(.A1(new_n6814_), .A2(new_n6806_), .B(new_n6812_), .ZN(new_n6820_));
  INV_X1     g06628(.I(new_n6820_), .ZN(new_n6821_));
  OAI21_X1   g06629(.A1(new_n6750_), .A2(new_n6752_), .B(new_n6755_), .ZN(new_n6822_));
  NOR2_X1    g06630(.A1(new_n6813_), .A2(new_n6822_), .ZN(new_n6823_));
  XOR2_X1    g06631(.A1(new_n6823_), .A2(new_n6537_), .Z(new_n6824_));
  NAND3_X1   g06632(.A1(\asqrt[28] ), .A2(new_n6766_), .A3(new_n6751_), .ZN(new_n6825_));
  XOR2_X1    g06633(.A1(new_n6825_), .A2(new_n6541_), .Z(new_n6826_));
  OAI21_X1   g06634(.A1(new_n6761_), .A2(new_n6762_), .B(new_n6765_), .ZN(new_n6827_));
  NOR2_X1    g06635(.A1(new_n6813_), .A2(new_n6827_), .ZN(new_n6828_));
  XOR2_X1    g06636(.A1(new_n6828_), .A2(new_n6543_), .Z(new_n6829_));
  INV_X1     g06637(.I(new_n6829_), .ZN(new_n6830_));
  NAND3_X1   g06638(.A1(\asqrt[28] ), .A2(new_n6728_), .A3(new_n6747_), .ZN(new_n6831_));
  XOR2_X1    g06639(.A1(new_n6831_), .A2(new_n6759_), .Z(new_n6832_));
  INV_X1     g06640(.I(new_n6832_), .ZN(new_n6833_));
  OAI21_X1   g06641(.A1(new_n6722_), .A2(new_n6724_), .B(new_n6727_), .ZN(new_n6834_));
  NOR2_X1    g06642(.A1(new_n6813_), .A2(new_n6834_), .ZN(new_n6835_));
  XOR2_X1    g06643(.A1(new_n6835_), .A2(new_n6549_), .Z(new_n6836_));
  NAND3_X1   g06644(.A1(\asqrt[28] ), .A2(new_n6741_), .A3(new_n6723_), .ZN(new_n6837_));
  XOR2_X1    g06645(.A1(new_n6837_), .A2(new_n6553_), .Z(new_n6838_));
  OAI21_X1   g06646(.A1(new_n6736_), .A2(new_n6737_), .B(new_n6740_), .ZN(new_n6839_));
  NOR2_X1    g06647(.A1(new_n6813_), .A2(new_n6839_), .ZN(new_n6840_));
  XOR2_X1    g06648(.A1(new_n6840_), .A2(new_n6555_), .Z(new_n6841_));
  INV_X1     g06649(.I(new_n6841_), .ZN(new_n6842_));
  NAND3_X1   g06650(.A1(\asqrt[28] ), .A2(new_n6700_), .A3(new_n6719_), .ZN(new_n6843_));
  XOR2_X1    g06651(.A1(new_n6843_), .A2(new_n6734_), .Z(new_n6844_));
  INV_X1     g06652(.I(new_n6844_), .ZN(new_n6845_));
  OAI21_X1   g06653(.A1(new_n6694_), .A2(new_n6696_), .B(new_n6699_), .ZN(new_n6846_));
  NOR2_X1    g06654(.A1(new_n6813_), .A2(new_n6846_), .ZN(new_n6847_));
  XOR2_X1    g06655(.A1(new_n6847_), .A2(new_n6561_), .Z(new_n6848_));
  NAND3_X1   g06656(.A1(\asqrt[28] ), .A2(new_n6713_), .A3(new_n6695_), .ZN(new_n6849_));
  XOR2_X1    g06657(.A1(new_n6849_), .A2(new_n6565_), .Z(new_n6850_));
  OAI21_X1   g06658(.A1(new_n6708_), .A2(new_n6709_), .B(new_n6712_), .ZN(new_n6851_));
  NOR2_X1    g06659(.A1(new_n6813_), .A2(new_n6851_), .ZN(new_n6852_));
  XOR2_X1    g06660(.A1(new_n6852_), .A2(new_n6567_), .Z(new_n6853_));
  INV_X1     g06661(.I(new_n6853_), .ZN(new_n6854_));
  NAND3_X1   g06662(.A1(\asqrt[28] ), .A2(new_n6672_), .A3(new_n6691_), .ZN(new_n6855_));
  XOR2_X1    g06663(.A1(new_n6855_), .A2(new_n6706_), .Z(new_n6856_));
  INV_X1     g06664(.I(new_n6856_), .ZN(new_n6857_));
  OAI21_X1   g06665(.A1(new_n6666_), .A2(new_n6668_), .B(new_n6671_), .ZN(new_n6858_));
  NOR2_X1    g06666(.A1(new_n6813_), .A2(new_n6858_), .ZN(new_n6859_));
  XOR2_X1    g06667(.A1(new_n6859_), .A2(new_n6573_), .Z(new_n6860_));
  NAND3_X1   g06668(.A1(\asqrt[28] ), .A2(new_n6685_), .A3(new_n6667_), .ZN(new_n6861_));
  XOR2_X1    g06669(.A1(new_n6861_), .A2(new_n6577_), .Z(new_n6862_));
  OAI21_X1   g06670(.A1(new_n6680_), .A2(new_n6681_), .B(new_n6684_), .ZN(new_n6863_));
  NOR2_X1    g06671(.A1(new_n6813_), .A2(new_n6863_), .ZN(new_n6864_));
  XOR2_X1    g06672(.A1(new_n6864_), .A2(new_n6579_), .Z(new_n6865_));
  INV_X1     g06673(.I(new_n6865_), .ZN(new_n6866_));
  NAND3_X1   g06674(.A1(\asqrt[28] ), .A2(new_n6644_), .A3(new_n6663_), .ZN(new_n6867_));
  XOR2_X1    g06675(.A1(new_n6867_), .A2(new_n6678_), .Z(new_n6868_));
  INV_X1     g06676(.I(new_n6868_), .ZN(new_n6869_));
  OAI21_X1   g06677(.A1(new_n6638_), .A2(new_n6640_), .B(new_n6643_), .ZN(new_n6870_));
  NOR2_X1    g06678(.A1(new_n6813_), .A2(new_n6870_), .ZN(new_n6871_));
  XOR2_X1    g06679(.A1(new_n6871_), .A2(new_n6585_), .Z(new_n6872_));
  NAND3_X1   g06680(.A1(\asqrt[28] ), .A2(new_n6657_), .A3(new_n6639_), .ZN(new_n6873_));
  XOR2_X1    g06681(.A1(new_n6873_), .A2(new_n6589_), .Z(new_n6874_));
  OAI21_X1   g06682(.A1(new_n6652_), .A2(new_n6653_), .B(new_n6656_), .ZN(new_n6875_));
  NOR2_X1    g06683(.A1(new_n6813_), .A2(new_n6875_), .ZN(new_n6876_));
  XOR2_X1    g06684(.A1(new_n6876_), .A2(new_n6591_), .Z(new_n6877_));
  INV_X1     g06685(.I(new_n6877_), .ZN(new_n6878_));
  NAND3_X1   g06686(.A1(\asqrt[28] ), .A2(new_n6617_), .A3(new_n6635_), .ZN(new_n6879_));
  XOR2_X1    g06687(.A1(new_n6879_), .A2(new_n6650_), .Z(new_n6880_));
  INV_X1     g06688(.I(new_n6880_), .ZN(new_n6881_));
  OAI21_X1   g06689(.A1(new_n6611_), .A2(new_n6613_), .B(new_n6616_), .ZN(new_n6882_));
  NOR2_X1    g06690(.A1(new_n6813_), .A2(new_n6882_), .ZN(new_n6883_));
  XOR2_X1    g06691(.A1(new_n6883_), .A2(new_n6597_), .Z(new_n6884_));
  NAND3_X1   g06692(.A1(\asqrt[28] ), .A2(new_n6629_), .A3(new_n6612_), .ZN(new_n6885_));
  XOR2_X1    g06693(.A1(new_n6885_), .A2(new_n6601_), .Z(new_n6886_));
  OAI21_X1   g06694(.A1(new_n6624_), .A2(new_n6625_), .B(new_n6628_), .ZN(new_n6887_));
  NOR2_X1    g06695(.A1(new_n6813_), .A2(new_n6887_), .ZN(new_n6888_));
  XOR2_X1    g06696(.A1(new_n6888_), .A2(new_n6603_), .Z(new_n6889_));
  INV_X1     g06697(.I(new_n6889_), .ZN(new_n6890_));
  INV_X1     g06698(.I(new_n6796_), .ZN(new_n6891_));
  OAI21_X1   g06699(.A1(new_n6503_), .A2(new_n6505_), .B(new_n6508_), .ZN(new_n6892_));
  NOR2_X1    g06700(.A1(new_n6813_), .A2(new_n6892_), .ZN(new_n6893_));
  XOR2_X1    g06701(.A1(new_n6893_), .A2(new_n6456_), .Z(new_n6894_));
  NAND3_X1   g06702(.A1(\asqrt[28] ), .A2(new_n6518_), .A3(new_n6504_), .ZN(new_n6895_));
  XOR2_X1    g06703(.A1(new_n6895_), .A2(new_n6459_), .Z(new_n6896_));
  OAI21_X1   g06704(.A1(new_n6513_), .A2(new_n6514_), .B(new_n6517_), .ZN(new_n6897_));
  NOR2_X1    g06705(.A1(new_n6813_), .A2(new_n6897_), .ZN(new_n6898_));
  XOR2_X1    g06706(.A1(new_n6898_), .A2(new_n6462_), .Z(new_n6899_));
  INV_X1     g06707(.I(new_n6899_), .ZN(new_n6900_));
  NAND3_X1   g06708(.A1(\asqrt[28] ), .A2(new_n6482_), .A3(new_n6500_), .ZN(new_n6901_));
  XOR2_X1    g06709(.A1(new_n6901_), .A2(new_n6512_), .Z(new_n6902_));
  INV_X1     g06710(.I(new_n6902_), .ZN(new_n6903_));
  NOR2_X1    g06711(.A1(new_n6479_), .A2(\asqrt[31] ), .ZN(new_n6904_));
  NOR3_X1    g06712(.A1(new_n6813_), .A2(new_n6904_), .A3(new_n6499_), .ZN(new_n6905_));
  XOR2_X1    g06713(.A1(new_n6905_), .A2(new_n6470_), .Z(new_n6906_));
  NOR3_X1    g06714(.A1(new_n6813_), .A2(\a[56] ), .A3(\a[57] ), .ZN(new_n6907_));
  NOR4_X1    g06715(.A1(new_n6811_), .A2(new_n6454_), .A3(new_n6528_), .A4(new_n6812_), .ZN(new_n6908_));
  OAI21_X1   g06716(.A1(new_n6907_), .A2(new_n6908_), .B(new_n6200_), .ZN(new_n6909_));
  NAND3_X1   g06717(.A1(\asqrt[28] ), .A2(new_n6471_), .A3(new_n6472_), .ZN(new_n6910_));
  INV_X1     g06718(.I(new_n6908_), .ZN(new_n6911_));
  NAND3_X1   g06719(.A1(new_n6910_), .A2(\a[58] ), .A3(new_n6911_), .ZN(new_n6912_));
  NAND2_X1   g06720(.A1(new_n6909_), .A2(new_n6912_), .ZN(new_n6913_));
  INV_X1     g06721(.I(\a[54] ), .ZN(new_n6914_));
  INV_X1     g06722(.I(\a[55] ), .ZN(new_n6915_));
  NAND3_X1   g06723(.A1(new_n6914_), .A2(new_n6915_), .A3(new_n6471_), .ZN(new_n6916_));
  NAND2_X1   g06724(.A1(\asqrt[28] ), .A2(\a[56] ), .ZN(new_n6917_));
  AOI21_X1   g06725(.A1(new_n6917_), .A2(new_n6916_), .B(new_n6454_), .ZN(new_n6918_));
  AOI21_X1   g06726(.A1(\asqrt[28] ), .A2(new_n6471_), .B(new_n6472_), .ZN(new_n6919_));
  NOR2_X1    g06727(.A1(new_n6907_), .A2(new_n6919_), .ZN(new_n6920_));
  NAND3_X1   g06728(.A1(new_n6917_), .A2(new_n6454_), .A3(new_n6916_), .ZN(new_n6921_));
  AOI21_X1   g06729(.A1(new_n6920_), .A2(new_n6921_), .B(new_n6918_), .ZN(new_n6922_));
  AOI21_X1   g06730(.A1(new_n6922_), .A2(new_n6106_), .B(new_n6913_), .ZN(new_n6923_));
  NOR2_X1    g06731(.A1(new_n6922_), .A2(new_n6106_), .ZN(new_n6924_));
  NOR3_X1    g06732(.A1(new_n6923_), .A2(\asqrt[31] ), .A3(new_n6924_), .ZN(new_n6925_));
  NOR3_X1    g06733(.A1(new_n6813_), .A2(new_n6493_), .A3(new_n6478_), .ZN(new_n6926_));
  XOR2_X1    g06734(.A1(new_n6926_), .A2(new_n6495_), .Z(new_n6927_));
  INV_X1     g06735(.I(new_n6927_), .ZN(new_n6928_));
  OAI21_X1   g06736(.A1(new_n6923_), .A2(new_n6924_), .B(\asqrt[31] ), .ZN(new_n6929_));
  OAI21_X1   g06737(.A1(new_n6925_), .A2(new_n6928_), .B(new_n6929_), .ZN(new_n6930_));
  OAI21_X1   g06738(.A1(new_n6930_), .A2(\asqrt[32] ), .B(new_n6906_), .ZN(new_n6931_));
  AOI21_X1   g06739(.A1(new_n6930_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n6932_));
  AOI21_X1   g06740(.A1(new_n6932_), .A2(new_n6931_), .B(new_n6903_), .ZN(new_n6933_));
  NAND2_X1   g06741(.A1(new_n6930_), .A2(\asqrt[32] ), .ZN(new_n6934_));
  AOI21_X1   g06742(.A1(new_n6931_), .A2(new_n6934_), .B(new_n5110_), .ZN(new_n6935_));
  NOR2_X1    g06743(.A1(new_n6933_), .A2(new_n6935_), .ZN(new_n6936_));
  AOI21_X1   g06744(.A1(new_n6936_), .A2(new_n4810_), .B(new_n6900_), .ZN(new_n6937_));
  OAI21_X1   g06745(.A1(new_n6933_), .A2(new_n6935_), .B(\asqrt[34] ), .ZN(new_n6938_));
  NAND2_X1   g06746(.A1(new_n6938_), .A2(new_n4510_), .ZN(new_n6939_));
  OAI21_X1   g06747(.A1(new_n6937_), .A2(new_n6939_), .B(new_n6896_), .ZN(new_n6940_));
  INV_X1     g06748(.I(new_n6938_), .ZN(new_n6941_));
  OAI21_X1   g06749(.A1(new_n6937_), .A2(new_n6941_), .B(\asqrt[35] ), .ZN(new_n6942_));
  NAND3_X1   g06750(.A1(new_n6940_), .A2(new_n6942_), .A3(new_n4224_), .ZN(new_n6943_));
  NAND2_X1   g06751(.A1(new_n6943_), .A2(new_n6894_), .ZN(new_n6944_));
  NAND2_X1   g06752(.A1(new_n6940_), .A2(new_n6942_), .ZN(new_n6945_));
  AOI21_X1   g06753(.A1(new_n6945_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n6946_));
  AOI21_X1   g06754(.A1(new_n6946_), .A2(new_n6944_), .B(new_n6891_), .ZN(new_n6947_));
  INV_X1     g06755(.I(new_n6896_), .ZN(new_n6948_));
  INV_X1     g06756(.I(new_n6906_), .ZN(new_n6949_));
  AOI21_X1   g06757(.A1(new_n6910_), .A2(new_n6911_), .B(\a[58] ), .ZN(new_n6950_));
  NOR3_X1    g06758(.A1(new_n6907_), .A2(new_n6200_), .A3(new_n6908_), .ZN(new_n6951_));
  NOR2_X1    g06759(.A1(new_n6951_), .A2(new_n6950_), .ZN(new_n6952_));
  OAI21_X1   g06760(.A1(new_n6813_), .A2(new_n6471_), .B(new_n6916_), .ZN(new_n6953_));
  NAND2_X1   g06761(.A1(new_n6953_), .A2(\asqrt[29] ), .ZN(new_n6954_));
  OAI21_X1   g06762(.A1(new_n6813_), .A2(\a[56] ), .B(\a[57] ), .ZN(new_n6955_));
  NAND2_X1   g06763(.A1(new_n6955_), .A2(new_n6910_), .ZN(new_n6956_));
  NOR2_X1    g06764(.A1(new_n6953_), .A2(\asqrt[29] ), .ZN(new_n6957_));
  OAI21_X1   g06765(.A1(new_n6956_), .A2(new_n6957_), .B(new_n6954_), .ZN(new_n6958_));
  OAI21_X1   g06766(.A1(\asqrt[30] ), .A2(new_n6958_), .B(new_n6952_), .ZN(new_n6959_));
  NAND2_X1   g06767(.A1(new_n6958_), .A2(\asqrt[30] ), .ZN(new_n6960_));
  NAND3_X1   g06768(.A1(new_n6959_), .A2(new_n5750_), .A3(new_n6960_), .ZN(new_n6961_));
  AOI21_X1   g06769(.A1(new_n6959_), .A2(new_n6960_), .B(new_n5750_), .ZN(new_n6962_));
  AOI21_X1   g06770(.A1(new_n6961_), .A2(new_n6927_), .B(new_n6962_), .ZN(new_n6963_));
  AOI21_X1   g06771(.A1(new_n6963_), .A2(new_n5435_), .B(new_n6949_), .ZN(new_n6964_));
  OAI21_X1   g06772(.A1(new_n6963_), .A2(new_n5435_), .B(new_n5110_), .ZN(new_n6965_));
  OAI21_X1   g06773(.A1(new_n6964_), .A2(new_n6965_), .B(new_n6902_), .ZN(new_n6966_));
  NOR2_X1    g06774(.A1(new_n6963_), .A2(new_n5435_), .ZN(new_n6967_));
  OAI21_X1   g06775(.A1(new_n6964_), .A2(new_n6967_), .B(\asqrt[33] ), .ZN(new_n6968_));
  NAND3_X1   g06776(.A1(new_n6966_), .A2(new_n6968_), .A3(new_n4810_), .ZN(new_n6969_));
  NAND2_X1   g06777(.A1(new_n6969_), .A2(new_n6899_), .ZN(new_n6970_));
  NAND2_X1   g06778(.A1(new_n6966_), .A2(new_n6968_), .ZN(new_n6971_));
  AOI21_X1   g06779(.A1(new_n6971_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n6972_));
  AOI21_X1   g06780(.A1(new_n6972_), .A2(new_n6970_), .B(new_n6948_), .ZN(new_n6973_));
  AOI21_X1   g06781(.A1(new_n6970_), .A2(new_n6938_), .B(new_n4510_), .ZN(new_n6974_));
  OAI21_X1   g06782(.A1(new_n6973_), .A2(new_n6974_), .B(\asqrt[36] ), .ZN(new_n6975_));
  AOI21_X1   g06783(.A1(new_n6944_), .A2(new_n6975_), .B(new_n3928_), .ZN(new_n6976_));
  NOR2_X1    g06784(.A1(new_n6947_), .A2(new_n6976_), .ZN(new_n6977_));
  AOI21_X1   g06785(.A1(new_n6977_), .A2(new_n3675_), .B(new_n6890_), .ZN(new_n6978_));
  OAI21_X1   g06786(.A1(new_n6947_), .A2(new_n6976_), .B(\asqrt[38] ), .ZN(new_n6979_));
  NAND2_X1   g06787(.A1(new_n6979_), .A2(new_n3400_), .ZN(new_n6980_));
  OAI21_X1   g06788(.A1(new_n6978_), .A2(new_n6980_), .B(new_n6886_), .ZN(new_n6981_));
  INV_X1     g06789(.I(new_n6979_), .ZN(new_n6982_));
  OAI21_X1   g06790(.A1(new_n6978_), .A2(new_n6982_), .B(\asqrt[39] ), .ZN(new_n6983_));
  NAND3_X1   g06791(.A1(new_n6981_), .A2(new_n6983_), .A3(new_n3167_), .ZN(new_n6984_));
  NAND2_X1   g06792(.A1(new_n6984_), .A2(new_n6884_), .ZN(new_n6985_));
  NAND2_X1   g06793(.A1(new_n6981_), .A2(new_n6983_), .ZN(new_n6986_));
  AOI21_X1   g06794(.A1(new_n6986_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n6987_));
  AOI21_X1   g06795(.A1(new_n6987_), .A2(new_n6985_), .B(new_n6881_), .ZN(new_n6988_));
  INV_X1     g06796(.I(new_n6886_), .ZN(new_n6989_));
  INV_X1     g06797(.I(new_n6894_), .ZN(new_n6990_));
  NOR2_X1    g06798(.A1(new_n6973_), .A2(new_n6974_), .ZN(new_n6991_));
  AOI21_X1   g06799(.A1(new_n6991_), .A2(new_n4224_), .B(new_n6990_), .ZN(new_n6992_));
  NAND2_X1   g06800(.A1(new_n6975_), .A2(new_n3928_), .ZN(new_n6993_));
  OAI21_X1   g06801(.A1(new_n6992_), .A2(new_n6993_), .B(new_n6796_), .ZN(new_n6994_));
  INV_X1     g06802(.I(new_n6975_), .ZN(new_n6995_));
  OAI21_X1   g06803(.A1(new_n6992_), .A2(new_n6995_), .B(\asqrt[37] ), .ZN(new_n6996_));
  NAND3_X1   g06804(.A1(new_n6994_), .A2(new_n6996_), .A3(new_n3675_), .ZN(new_n6997_));
  NAND2_X1   g06805(.A1(new_n6997_), .A2(new_n6889_), .ZN(new_n6998_));
  NAND2_X1   g06806(.A1(new_n6994_), .A2(new_n6996_), .ZN(new_n6999_));
  AOI21_X1   g06807(.A1(new_n6999_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n7000_));
  AOI21_X1   g06808(.A1(new_n7000_), .A2(new_n6998_), .B(new_n6989_), .ZN(new_n7001_));
  AOI21_X1   g06809(.A1(new_n6998_), .A2(new_n6979_), .B(new_n3400_), .ZN(new_n7002_));
  OAI21_X1   g06810(.A1(new_n7001_), .A2(new_n7002_), .B(\asqrt[40] ), .ZN(new_n7003_));
  AOI21_X1   g06811(.A1(new_n6985_), .A2(new_n7003_), .B(new_n2912_), .ZN(new_n7004_));
  NOR2_X1    g06812(.A1(new_n6988_), .A2(new_n7004_), .ZN(new_n7005_));
  AOI21_X1   g06813(.A1(new_n7005_), .A2(new_n2699_), .B(new_n6878_), .ZN(new_n7006_));
  OAI21_X1   g06814(.A1(new_n6988_), .A2(new_n7004_), .B(\asqrt[42] ), .ZN(new_n7007_));
  NAND2_X1   g06815(.A1(new_n7007_), .A2(new_n2464_), .ZN(new_n7008_));
  OAI21_X1   g06816(.A1(new_n7006_), .A2(new_n7008_), .B(new_n6874_), .ZN(new_n7009_));
  INV_X1     g06817(.I(new_n7007_), .ZN(new_n7010_));
  OAI21_X1   g06818(.A1(new_n7006_), .A2(new_n7010_), .B(\asqrt[43] ), .ZN(new_n7011_));
  NAND3_X1   g06819(.A1(new_n7009_), .A2(new_n7011_), .A3(new_n2271_), .ZN(new_n7012_));
  NAND2_X1   g06820(.A1(new_n7012_), .A2(new_n6872_), .ZN(new_n7013_));
  NAND2_X1   g06821(.A1(new_n7009_), .A2(new_n7011_), .ZN(new_n7014_));
  AOI21_X1   g06822(.A1(new_n7014_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n7015_));
  AOI21_X1   g06823(.A1(new_n7015_), .A2(new_n7013_), .B(new_n6869_), .ZN(new_n7016_));
  INV_X1     g06824(.I(new_n6874_), .ZN(new_n7017_));
  INV_X1     g06825(.I(new_n6884_), .ZN(new_n7018_));
  NOR2_X1    g06826(.A1(new_n7001_), .A2(new_n7002_), .ZN(new_n7019_));
  AOI21_X1   g06827(.A1(new_n7019_), .A2(new_n3167_), .B(new_n7018_), .ZN(new_n7020_));
  NAND2_X1   g06828(.A1(new_n7003_), .A2(new_n2912_), .ZN(new_n7021_));
  OAI21_X1   g06829(.A1(new_n7020_), .A2(new_n7021_), .B(new_n6880_), .ZN(new_n7022_));
  INV_X1     g06830(.I(new_n7003_), .ZN(new_n7023_));
  OAI21_X1   g06831(.A1(new_n7020_), .A2(new_n7023_), .B(\asqrt[41] ), .ZN(new_n7024_));
  NAND3_X1   g06832(.A1(new_n7022_), .A2(new_n7024_), .A3(new_n2699_), .ZN(new_n7025_));
  NAND2_X1   g06833(.A1(new_n7025_), .A2(new_n6877_), .ZN(new_n7026_));
  NAND2_X1   g06834(.A1(new_n7022_), .A2(new_n7024_), .ZN(new_n7027_));
  AOI21_X1   g06835(.A1(new_n7027_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n7028_));
  AOI21_X1   g06836(.A1(new_n7028_), .A2(new_n7026_), .B(new_n7017_), .ZN(new_n7029_));
  AOI21_X1   g06837(.A1(new_n7026_), .A2(new_n7007_), .B(new_n2464_), .ZN(new_n7030_));
  OAI21_X1   g06838(.A1(new_n7029_), .A2(new_n7030_), .B(\asqrt[44] ), .ZN(new_n7031_));
  AOI21_X1   g06839(.A1(new_n7013_), .A2(new_n7031_), .B(new_n2072_), .ZN(new_n7032_));
  NOR2_X1    g06840(.A1(new_n7016_), .A2(new_n7032_), .ZN(new_n7033_));
  AOI21_X1   g06841(.A1(new_n7033_), .A2(new_n1884_), .B(new_n6866_), .ZN(new_n7034_));
  OAI21_X1   g06842(.A1(new_n7016_), .A2(new_n7032_), .B(\asqrt[46] ), .ZN(new_n7035_));
  NAND2_X1   g06843(.A1(new_n7035_), .A2(new_n1688_), .ZN(new_n7036_));
  OAI21_X1   g06844(.A1(new_n7034_), .A2(new_n7036_), .B(new_n6862_), .ZN(new_n7037_));
  INV_X1     g06845(.I(new_n7035_), .ZN(new_n7038_));
  OAI21_X1   g06846(.A1(new_n7034_), .A2(new_n7038_), .B(\asqrt[47] ), .ZN(new_n7039_));
  NAND3_X1   g06847(.A1(new_n7037_), .A2(new_n7039_), .A3(new_n1533_), .ZN(new_n7040_));
  NAND2_X1   g06848(.A1(new_n7040_), .A2(new_n6860_), .ZN(new_n7041_));
  NAND2_X1   g06849(.A1(new_n7037_), .A2(new_n7039_), .ZN(new_n7042_));
  AOI21_X1   g06850(.A1(new_n7042_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n7043_));
  AOI21_X1   g06851(.A1(new_n7043_), .A2(new_n7041_), .B(new_n6857_), .ZN(new_n7044_));
  INV_X1     g06852(.I(new_n6862_), .ZN(new_n7045_));
  INV_X1     g06853(.I(new_n6872_), .ZN(new_n7046_));
  NOR2_X1    g06854(.A1(new_n7029_), .A2(new_n7030_), .ZN(new_n7047_));
  AOI21_X1   g06855(.A1(new_n7047_), .A2(new_n2271_), .B(new_n7046_), .ZN(new_n7048_));
  NAND2_X1   g06856(.A1(new_n7031_), .A2(new_n2072_), .ZN(new_n7049_));
  OAI21_X1   g06857(.A1(new_n7048_), .A2(new_n7049_), .B(new_n6868_), .ZN(new_n7050_));
  INV_X1     g06858(.I(new_n7031_), .ZN(new_n7051_));
  OAI21_X1   g06859(.A1(new_n7048_), .A2(new_n7051_), .B(\asqrt[45] ), .ZN(new_n7052_));
  NAND3_X1   g06860(.A1(new_n7050_), .A2(new_n7052_), .A3(new_n1884_), .ZN(new_n7053_));
  NAND2_X1   g06861(.A1(new_n7053_), .A2(new_n6865_), .ZN(new_n7054_));
  NAND2_X1   g06862(.A1(new_n7050_), .A2(new_n7052_), .ZN(new_n7055_));
  AOI21_X1   g06863(.A1(new_n7055_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n7056_));
  AOI21_X1   g06864(.A1(new_n7056_), .A2(new_n7054_), .B(new_n7045_), .ZN(new_n7057_));
  AOI21_X1   g06865(.A1(new_n7054_), .A2(new_n7035_), .B(new_n1688_), .ZN(new_n7058_));
  OAI21_X1   g06866(.A1(new_n7057_), .A2(new_n7058_), .B(\asqrt[48] ), .ZN(new_n7059_));
  AOI21_X1   g06867(.A1(new_n7041_), .A2(new_n7059_), .B(new_n1368_), .ZN(new_n7060_));
  NOR2_X1    g06868(.A1(new_n7044_), .A2(new_n7060_), .ZN(new_n7061_));
  AOI21_X1   g06869(.A1(new_n7061_), .A2(new_n1228_), .B(new_n6854_), .ZN(new_n7062_));
  OAI21_X1   g06870(.A1(new_n7044_), .A2(new_n7060_), .B(\asqrt[50] ), .ZN(new_n7063_));
  NAND2_X1   g06871(.A1(new_n7063_), .A2(new_n1088_), .ZN(new_n7064_));
  OAI21_X1   g06872(.A1(new_n7062_), .A2(new_n7064_), .B(new_n6850_), .ZN(new_n7065_));
  INV_X1     g06873(.I(new_n7063_), .ZN(new_n7066_));
  OAI21_X1   g06874(.A1(new_n7062_), .A2(new_n7066_), .B(\asqrt[51] ), .ZN(new_n7067_));
  NAND3_X1   g06875(.A1(new_n7065_), .A2(new_n7067_), .A3(new_n962_), .ZN(new_n7068_));
  NAND2_X1   g06876(.A1(new_n7068_), .A2(new_n6848_), .ZN(new_n7069_));
  NAND2_X1   g06877(.A1(new_n7065_), .A2(new_n7067_), .ZN(new_n7070_));
  AOI21_X1   g06878(.A1(new_n7070_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n7071_));
  AOI21_X1   g06879(.A1(new_n7071_), .A2(new_n7069_), .B(new_n6845_), .ZN(new_n7072_));
  INV_X1     g06880(.I(new_n6850_), .ZN(new_n7073_));
  INV_X1     g06881(.I(new_n6860_), .ZN(new_n7074_));
  NOR2_X1    g06882(.A1(new_n7057_), .A2(new_n7058_), .ZN(new_n7075_));
  AOI21_X1   g06883(.A1(new_n7075_), .A2(new_n1533_), .B(new_n7074_), .ZN(new_n7076_));
  NAND2_X1   g06884(.A1(new_n7059_), .A2(new_n1368_), .ZN(new_n7077_));
  OAI21_X1   g06885(.A1(new_n7076_), .A2(new_n7077_), .B(new_n6856_), .ZN(new_n7078_));
  INV_X1     g06886(.I(new_n7059_), .ZN(new_n7079_));
  OAI21_X1   g06887(.A1(new_n7076_), .A2(new_n7079_), .B(\asqrt[49] ), .ZN(new_n7080_));
  NAND3_X1   g06888(.A1(new_n7078_), .A2(new_n7080_), .A3(new_n1228_), .ZN(new_n7081_));
  NAND2_X1   g06889(.A1(new_n7081_), .A2(new_n6853_), .ZN(new_n7082_));
  NAND2_X1   g06890(.A1(new_n7078_), .A2(new_n7080_), .ZN(new_n7083_));
  AOI21_X1   g06891(.A1(new_n7083_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n7084_));
  AOI21_X1   g06892(.A1(new_n7084_), .A2(new_n7082_), .B(new_n7073_), .ZN(new_n7085_));
  AOI21_X1   g06893(.A1(new_n7082_), .A2(new_n7063_), .B(new_n1088_), .ZN(new_n7086_));
  OAI21_X1   g06894(.A1(new_n7085_), .A2(new_n7086_), .B(\asqrt[52] ), .ZN(new_n7087_));
  AOI21_X1   g06895(.A1(new_n7069_), .A2(new_n7087_), .B(new_n842_), .ZN(new_n7088_));
  NOR2_X1    g06896(.A1(new_n7072_), .A2(new_n7088_), .ZN(new_n7089_));
  AOI21_X1   g06897(.A1(new_n7089_), .A2(new_n720_), .B(new_n6842_), .ZN(new_n7090_));
  OAI21_X1   g06898(.A1(new_n7072_), .A2(new_n7088_), .B(\asqrt[54] ), .ZN(new_n7091_));
  NAND2_X1   g06899(.A1(new_n7091_), .A2(new_n630_), .ZN(new_n7092_));
  OAI21_X1   g06900(.A1(new_n7090_), .A2(new_n7092_), .B(new_n6838_), .ZN(new_n7093_));
  INV_X1     g06901(.I(new_n7091_), .ZN(new_n7094_));
  OAI21_X1   g06902(.A1(new_n7090_), .A2(new_n7094_), .B(\asqrt[55] ), .ZN(new_n7095_));
  NAND3_X1   g06903(.A1(new_n7093_), .A2(new_n7095_), .A3(new_n545_), .ZN(new_n7096_));
  NAND2_X1   g06904(.A1(new_n7096_), .A2(new_n6836_), .ZN(new_n7097_));
  NAND2_X1   g06905(.A1(new_n7093_), .A2(new_n7095_), .ZN(new_n7098_));
  AOI21_X1   g06906(.A1(new_n7098_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n7099_));
  AOI21_X1   g06907(.A1(new_n7099_), .A2(new_n7097_), .B(new_n6833_), .ZN(new_n7100_));
  INV_X1     g06908(.I(new_n6838_), .ZN(new_n7101_));
  INV_X1     g06909(.I(new_n6848_), .ZN(new_n7102_));
  NOR2_X1    g06910(.A1(new_n7085_), .A2(new_n7086_), .ZN(new_n7103_));
  AOI21_X1   g06911(.A1(new_n7103_), .A2(new_n962_), .B(new_n7102_), .ZN(new_n7104_));
  NAND2_X1   g06912(.A1(new_n7087_), .A2(new_n842_), .ZN(new_n7105_));
  OAI21_X1   g06913(.A1(new_n7104_), .A2(new_n7105_), .B(new_n6844_), .ZN(new_n7106_));
  INV_X1     g06914(.I(new_n7087_), .ZN(new_n7107_));
  OAI21_X1   g06915(.A1(new_n7104_), .A2(new_n7107_), .B(\asqrt[53] ), .ZN(new_n7108_));
  NAND3_X1   g06916(.A1(new_n7106_), .A2(new_n7108_), .A3(new_n720_), .ZN(new_n7109_));
  NAND2_X1   g06917(.A1(new_n7109_), .A2(new_n6841_), .ZN(new_n7110_));
  NAND2_X1   g06918(.A1(new_n7106_), .A2(new_n7108_), .ZN(new_n7111_));
  AOI21_X1   g06919(.A1(new_n7111_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n7112_));
  AOI21_X1   g06920(.A1(new_n7112_), .A2(new_n7110_), .B(new_n7101_), .ZN(new_n7113_));
  AOI21_X1   g06921(.A1(new_n7110_), .A2(new_n7091_), .B(new_n630_), .ZN(new_n7114_));
  OAI21_X1   g06922(.A1(new_n7113_), .A2(new_n7114_), .B(\asqrt[56] ), .ZN(new_n7115_));
  AOI21_X1   g06923(.A1(new_n7097_), .A2(new_n7115_), .B(new_n450_), .ZN(new_n7116_));
  NOR2_X1    g06924(.A1(new_n7100_), .A2(new_n7116_), .ZN(new_n7117_));
  AOI21_X1   g06925(.A1(new_n7117_), .A2(new_n403_), .B(new_n6830_), .ZN(new_n7118_));
  OAI21_X1   g06926(.A1(new_n7100_), .A2(new_n7116_), .B(\asqrt[58] ), .ZN(new_n7119_));
  NAND2_X1   g06927(.A1(new_n7119_), .A2(new_n339_), .ZN(new_n7120_));
  OAI21_X1   g06928(.A1(new_n7118_), .A2(new_n7120_), .B(new_n6826_), .ZN(new_n7121_));
  INV_X1     g06929(.I(new_n7119_), .ZN(new_n7122_));
  OAI21_X1   g06930(.A1(new_n7118_), .A2(new_n7122_), .B(\asqrt[59] ), .ZN(new_n7123_));
  NAND3_X1   g06931(.A1(new_n7121_), .A2(new_n7123_), .A3(new_n288_), .ZN(new_n7124_));
  NAND2_X1   g06932(.A1(new_n7124_), .A2(new_n6824_), .ZN(new_n7125_));
  INV_X1     g06933(.I(new_n6826_), .ZN(new_n7126_));
  INV_X1     g06934(.I(new_n6836_), .ZN(new_n7127_));
  NOR2_X1    g06935(.A1(new_n7113_), .A2(new_n7114_), .ZN(new_n7128_));
  AOI21_X1   g06936(.A1(new_n7128_), .A2(new_n545_), .B(new_n7127_), .ZN(new_n7129_));
  NAND2_X1   g06937(.A1(new_n7115_), .A2(new_n450_), .ZN(new_n7130_));
  OAI21_X1   g06938(.A1(new_n7129_), .A2(new_n7130_), .B(new_n6832_), .ZN(new_n7131_));
  INV_X1     g06939(.I(new_n7115_), .ZN(new_n7132_));
  OAI21_X1   g06940(.A1(new_n7129_), .A2(new_n7132_), .B(\asqrt[57] ), .ZN(new_n7133_));
  NAND3_X1   g06941(.A1(new_n7131_), .A2(new_n7133_), .A3(new_n403_), .ZN(new_n7134_));
  NAND2_X1   g06942(.A1(new_n7134_), .A2(new_n6829_), .ZN(new_n7135_));
  NAND2_X1   g06943(.A1(new_n7131_), .A2(new_n7133_), .ZN(new_n7136_));
  AOI21_X1   g06944(.A1(new_n7136_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n7137_));
  AOI21_X1   g06945(.A1(new_n7137_), .A2(new_n7135_), .B(new_n7126_), .ZN(new_n7138_));
  AOI21_X1   g06946(.A1(new_n7135_), .A2(new_n7119_), .B(new_n339_), .ZN(new_n7139_));
  OAI21_X1   g06947(.A1(new_n7138_), .A2(new_n7139_), .B(\asqrt[60] ), .ZN(new_n7140_));
  AOI21_X1   g06948(.A1(new_n7125_), .A2(new_n7140_), .B(new_n242_), .ZN(new_n7141_));
  NAND3_X1   g06949(.A1(\asqrt[28] ), .A2(new_n6756_), .A3(new_n6772_), .ZN(new_n7142_));
  XOR2_X1    g06950(.A1(new_n7142_), .A2(new_n6797_), .Z(new_n7143_));
  INV_X1     g06951(.I(new_n7143_), .ZN(new_n7144_));
  NAND2_X1   g06952(.A1(new_n7121_), .A2(new_n7123_), .ZN(new_n7145_));
  AOI21_X1   g06953(.A1(new_n7145_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n7146_));
  AOI21_X1   g06954(.A1(new_n7146_), .A2(new_n7125_), .B(new_n7144_), .ZN(new_n7147_));
  OAI21_X1   g06955(.A1(new_n7147_), .A2(new_n7141_), .B(\asqrt[62] ), .ZN(new_n7148_));
  AOI21_X1   g06956(.A1(new_n6757_), .A2(new_n6778_), .B(new_n6773_), .ZN(new_n7149_));
  NAND2_X1   g06957(.A1(\asqrt[28] ), .A2(new_n7149_), .ZN(new_n7150_));
  XOR2_X1    g06958(.A1(new_n7150_), .A2(new_n6776_), .Z(new_n7151_));
  INV_X1     g06959(.I(new_n6824_), .ZN(new_n7152_));
  NOR2_X1    g06960(.A1(new_n7138_), .A2(new_n7139_), .ZN(new_n7153_));
  AOI21_X1   g06961(.A1(new_n7153_), .A2(new_n288_), .B(new_n7152_), .ZN(new_n7154_));
  INV_X1     g06962(.I(new_n7140_), .ZN(new_n7155_));
  OAI21_X1   g06963(.A1(new_n7154_), .A2(new_n7155_), .B(\asqrt[61] ), .ZN(new_n7156_));
  NAND2_X1   g06964(.A1(new_n7140_), .A2(new_n242_), .ZN(new_n7157_));
  OAI21_X1   g06965(.A1(new_n7154_), .A2(new_n7157_), .B(new_n7143_), .ZN(new_n7158_));
  NAND3_X1   g06966(.A1(new_n7158_), .A2(new_n7156_), .A3(new_n234_), .ZN(new_n7159_));
  NAND2_X1   g06967(.A1(new_n7159_), .A2(new_n7151_), .ZN(new_n7160_));
  AOI21_X1   g06968(.A1(new_n7160_), .A2(new_n7148_), .B(new_n6821_), .ZN(new_n7161_));
  AOI21_X1   g06969(.A1(new_n7161_), .A2(new_n6819_), .B(\asqrt[63] ), .ZN(new_n7162_));
  NAND2_X1   g06970(.A1(new_n7160_), .A2(new_n7148_), .ZN(new_n7163_));
  NOR2_X1    g06971(.A1(new_n7163_), .A2(new_n6819_), .ZN(new_n7164_));
  NOR2_X1    g06972(.A1(\asqrt[28] ), .A2(new_n6808_), .ZN(new_n7165_));
  NOR4_X1    g06973(.A1(new_n7162_), .A2(new_n6816_), .A3(new_n7164_), .A4(new_n7165_), .ZN(new_n7166_));
  OAI21_X1   g06974(.A1(new_n6992_), .A2(new_n6993_), .B(new_n6996_), .ZN(new_n7167_));
  NOR2_X1    g06975(.A1(new_n7166_), .A2(new_n7167_), .ZN(new_n7168_));
  XOR2_X1    g06976(.A1(new_n7168_), .A2(new_n6796_), .Z(new_n7169_));
  INV_X1     g06977(.I(new_n7169_), .ZN(new_n7170_));
  INV_X1     g06978(.I(new_n6816_), .ZN(new_n7171_));
  INV_X1     g06979(.I(new_n7148_), .ZN(new_n7172_));
  NOR2_X1    g06980(.A1(new_n7147_), .A2(new_n7141_), .ZN(new_n7173_));
  INV_X1     g06981(.I(new_n7151_), .ZN(new_n7174_));
  AOI21_X1   g06982(.A1(new_n7173_), .A2(new_n234_), .B(new_n7174_), .ZN(new_n7175_));
  OAI21_X1   g06983(.A1(new_n7175_), .A2(new_n7172_), .B(new_n6820_), .ZN(new_n7176_));
  OAI21_X1   g06984(.A1(new_n7176_), .A2(new_n6818_), .B(new_n193_), .ZN(new_n7177_));
  NOR2_X1    g06985(.A1(new_n7175_), .A2(new_n7172_), .ZN(new_n7178_));
  NAND2_X1   g06986(.A1(new_n7178_), .A2(new_n6818_), .ZN(new_n7179_));
  INV_X1     g06987(.I(new_n7165_), .ZN(new_n7180_));
  NAND4_X1   g06988(.A1(new_n7177_), .A2(new_n7171_), .A3(new_n7179_), .A4(new_n7180_), .ZN(\asqrt[27] ));
  NAND3_X1   g06989(.A1(\asqrt[27] ), .A2(new_n6943_), .A3(new_n6975_), .ZN(new_n7182_));
  XOR2_X1    g06990(.A1(new_n7182_), .A2(new_n6990_), .Z(new_n7183_));
  OAI21_X1   g06991(.A1(new_n6937_), .A2(new_n6939_), .B(new_n6942_), .ZN(new_n7184_));
  NOR2_X1    g06992(.A1(new_n7166_), .A2(new_n7184_), .ZN(new_n7185_));
  XOR2_X1    g06993(.A1(new_n7185_), .A2(new_n6896_), .Z(new_n7186_));
  INV_X1     g06994(.I(new_n7186_), .ZN(new_n7187_));
  NAND3_X1   g06995(.A1(\asqrt[27] ), .A2(new_n6969_), .A3(new_n6938_), .ZN(new_n7188_));
  XOR2_X1    g06996(.A1(new_n7188_), .A2(new_n6900_), .Z(new_n7189_));
  INV_X1     g06997(.I(new_n7189_), .ZN(new_n7190_));
  AOI21_X1   g06998(.A1(new_n6931_), .A2(new_n6932_), .B(new_n6935_), .ZN(new_n7191_));
  NAND2_X1   g06999(.A1(\asqrt[27] ), .A2(new_n7191_), .ZN(new_n7192_));
  XOR2_X1    g07000(.A1(new_n7192_), .A2(new_n6903_), .Z(new_n7193_));
  NOR2_X1    g07001(.A1(new_n6930_), .A2(\asqrt[32] ), .ZN(new_n7194_));
  NOR3_X1    g07002(.A1(new_n7166_), .A2(new_n7194_), .A3(new_n6967_), .ZN(new_n7195_));
  XOR2_X1    g07003(.A1(new_n7195_), .A2(new_n6906_), .Z(new_n7196_));
  NOR3_X1    g07004(.A1(new_n7166_), .A2(new_n6925_), .A3(new_n6962_), .ZN(new_n7197_));
  XOR2_X1    g07005(.A1(new_n7197_), .A2(new_n6927_), .Z(new_n7198_));
  INV_X1     g07006(.I(new_n7198_), .ZN(new_n7199_));
  NOR2_X1    g07007(.A1(new_n6958_), .A2(\asqrt[30] ), .ZN(new_n7200_));
  NOR3_X1    g07008(.A1(new_n7166_), .A2(new_n7200_), .A3(new_n6924_), .ZN(new_n7201_));
  XOR2_X1    g07009(.A1(new_n7201_), .A2(new_n6952_), .Z(new_n7202_));
  INV_X1     g07010(.I(new_n7202_), .ZN(new_n7203_));
  NAND3_X1   g07011(.A1(\asqrt[27] ), .A2(new_n6914_), .A3(new_n6915_), .ZN(new_n7204_));
  NAND4_X1   g07012(.A1(new_n7177_), .A2(\asqrt[28] ), .A3(new_n7179_), .A4(new_n7171_), .ZN(new_n7205_));
  AOI21_X1   g07013(.A1(new_n7204_), .A2(new_n7205_), .B(\a[56] ), .ZN(new_n7206_));
  NOR3_X1    g07014(.A1(new_n7166_), .A2(\a[54] ), .A3(\a[55] ), .ZN(new_n7207_));
  INV_X1     g07015(.I(new_n7205_), .ZN(new_n7208_));
  NOR3_X1    g07016(.A1(new_n7207_), .A2(new_n6471_), .A3(new_n7208_), .ZN(new_n7209_));
  NOR2_X1    g07017(.A1(new_n7209_), .A2(new_n7206_), .ZN(new_n7210_));
  INV_X1     g07018(.I(\a[52] ), .ZN(new_n7211_));
  INV_X1     g07019(.I(\a[53] ), .ZN(new_n7212_));
  NAND3_X1   g07020(.A1(new_n7211_), .A2(new_n7212_), .A3(new_n6914_), .ZN(new_n7213_));
  OAI21_X1   g07021(.A1(new_n7166_), .A2(new_n6914_), .B(new_n7213_), .ZN(new_n7214_));
  NAND2_X1   g07022(.A1(new_n7214_), .A2(\asqrt[28] ), .ZN(new_n7215_));
  OAI21_X1   g07023(.A1(new_n7166_), .A2(\a[54] ), .B(\a[55] ), .ZN(new_n7216_));
  NAND2_X1   g07024(.A1(new_n7216_), .A2(new_n7204_), .ZN(new_n7217_));
  NOR2_X1    g07025(.A1(new_n7214_), .A2(\asqrt[28] ), .ZN(new_n7218_));
  OAI21_X1   g07026(.A1(new_n7217_), .A2(new_n7218_), .B(new_n7215_), .ZN(new_n7219_));
  OAI21_X1   g07027(.A1(new_n7219_), .A2(\asqrt[29] ), .B(new_n7210_), .ZN(new_n7220_));
  NAND2_X1   g07028(.A1(new_n7219_), .A2(\asqrt[29] ), .ZN(new_n7221_));
  NAND3_X1   g07029(.A1(new_n7220_), .A2(new_n6106_), .A3(new_n7221_), .ZN(new_n7222_));
  NOR3_X1    g07030(.A1(new_n7166_), .A2(new_n6918_), .A3(new_n6957_), .ZN(new_n7223_));
  XOR2_X1    g07031(.A1(new_n7223_), .A2(new_n6920_), .Z(new_n7224_));
  NAND2_X1   g07032(.A1(new_n7222_), .A2(new_n7224_), .ZN(new_n7225_));
  NAND2_X1   g07033(.A1(new_n7220_), .A2(new_n7221_), .ZN(new_n7226_));
  AOI21_X1   g07034(.A1(new_n7226_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n7227_));
  AOI21_X1   g07035(.A1(new_n7227_), .A2(new_n7225_), .B(new_n7203_), .ZN(new_n7228_));
  OAI21_X1   g07036(.A1(new_n7207_), .A2(new_n7208_), .B(new_n6471_), .ZN(new_n7229_));
  NAND3_X1   g07037(.A1(new_n7204_), .A2(\a[56] ), .A3(new_n7205_), .ZN(new_n7230_));
  NAND2_X1   g07038(.A1(new_n7229_), .A2(new_n7230_), .ZN(new_n7231_));
  NAND2_X1   g07039(.A1(\asqrt[27] ), .A2(\a[54] ), .ZN(new_n7232_));
  AOI21_X1   g07040(.A1(new_n7232_), .A2(new_n7213_), .B(new_n6813_), .ZN(new_n7233_));
  AOI21_X1   g07041(.A1(\asqrt[27] ), .A2(new_n6914_), .B(new_n6915_), .ZN(new_n7234_));
  NOR2_X1    g07042(.A1(new_n7207_), .A2(new_n7234_), .ZN(new_n7235_));
  NAND3_X1   g07043(.A1(new_n7232_), .A2(new_n6813_), .A3(new_n7213_), .ZN(new_n7236_));
  AOI21_X1   g07044(.A1(new_n7235_), .A2(new_n7236_), .B(new_n7233_), .ZN(new_n7237_));
  AOI21_X1   g07045(.A1(new_n7237_), .A2(new_n6454_), .B(new_n7231_), .ZN(new_n7238_));
  NOR2_X1    g07046(.A1(new_n7237_), .A2(new_n6454_), .ZN(new_n7239_));
  OAI21_X1   g07047(.A1(new_n7238_), .A2(new_n7239_), .B(\asqrt[30] ), .ZN(new_n7240_));
  AOI21_X1   g07048(.A1(new_n7225_), .A2(new_n7240_), .B(new_n5750_), .ZN(new_n7241_));
  NOR2_X1    g07049(.A1(new_n7228_), .A2(new_n7241_), .ZN(new_n7242_));
  AOI21_X1   g07050(.A1(new_n7242_), .A2(new_n5435_), .B(new_n7199_), .ZN(new_n7243_));
  OAI21_X1   g07051(.A1(new_n7228_), .A2(new_n7241_), .B(\asqrt[32] ), .ZN(new_n7244_));
  NAND2_X1   g07052(.A1(new_n7244_), .A2(new_n5110_), .ZN(new_n7245_));
  OAI21_X1   g07053(.A1(new_n7243_), .A2(new_n7245_), .B(new_n7196_), .ZN(new_n7246_));
  INV_X1     g07054(.I(new_n7244_), .ZN(new_n7247_));
  OAI21_X1   g07055(.A1(new_n7243_), .A2(new_n7247_), .B(\asqrt[33] ), .ZN(new_n7248_));
  NAND3_X1   g07056(.A1(new_n7246_), .A2(new_n7248_), .A3(new_n4810_), .ZN(new_n7249_));
  NAND2_X1   g07057(.A1(new_n7249_), .A2(new_n7193_), .ZN(new_n7250_));
  NAND2_X1   g07058(.A1(new_n7246_), .A2(new_n7248_), .ZN(new_n7251_));
  AOI21_X1   g07059(.A1(new_n7251_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n7252_));
  AOI21_X1   g07060(.A1(new_n7252_), .A2(new_n7250_), .B(new_n7190_), .ZN(new_n7253_));
  INV_X1     g07061(.I(new_n7196_), .ZN(new_n7254_));
  NOR2_X1    g07062(.A1(new_n7238_), .A2(new_n7239_), .ZN(new_n7255_));
  INV_X1     g07063(.I(new_n7224_), .ZN(new_n7256_));
  AOI21_X1   g07064(.A1(new_n7255_), .A2(new_n6106_), .B(new_n7256_), .ZN(new_n7257_));
  NAND2_X1   g07065(.A1(new_n7240_), .A2(new_n5750_), .ZN(new_n7258_));
  OAI21_X1   g07066(.A1(new_n7257_), .A2(new_n7258_), .B(new_n7202_), .ZN(new_n7259_));
  INV_X1     g07067(.I(new_n7240_), .ZN(new_n7260_));
  OAI21_X1   g07068(.A1(new_n7257_), .A2(new_n7260_), .B(\asqrt[31] ), .ZN(new_n7261_));
  NAND3_X1   g07069(.A1(new_n7259_), .A2(new_n7261_), .A3(new_n5435_), .ZN(new_n7262_));
  NAND2_X1   g07070(.A1(new_n7262_), .A2(new_n7198_), .ZN(new_n7263_));
  NAND2_X1   g07071(.A1(new_n7259_), .A2(new_n7261_), .ZN(new_n7264_));
  AOI21_X1   g07072(.A1(new_n7264_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n7265_));
  AOI21_X1   g07073(.A1(new_n7265_), .A2(new_n7263_), .B(new_n7254_), .ZN(new_n7266_));
  AOI21_X1   g07074(.A1(new_n7263_), .A2(new_n7244_), .B(new_n5110_), .ZN(new_n7267_));
  OAI21_X1   g07075(.A1(new_n7266_), .A2(new_n7267_), .B(\asqrt[34] ), .ZN(new_n7268_));
  AOI21_X1   g07076(.A1(new_n7250_), .A2(new_n7268_), .B(new_n4510_), .ZN(new_n7269_));
  NOR2_X1    g07077(.A1(new_n7253_), .A2(new_n7269_), .ZN(new_n7270_));
  AOI21_X1   g07078(.A1(new_n7270_), .A2(new_n4224_), .B(new_n7187_), .ZN(new_n7271_));
  OAI21_X1   g07079(.A1(new_n7253_), .A2(new_n7269_), .B(\asqrt[36] ), .ZN(new_n7272_));
  NAND2_X1   g07080(.A1(new_n7272_), .A2(new_n3928_), .ZN(new_n7273_));
  OAI21_X1   g07081(.A1(new_n7271_), .A2(new_n7273_), .B(new_n7183_), .ZN(new_n7274_));
  INV_X1     g07082(.I(new_n7272_), .ZN(new_n7275_));
  OAI21_X1   g07083(.A1(new_n7271_), .A2(new_n7275_), .B(\asqrt[37] ), .ZN(new_n7276_));
  NAND3_X1   g07084(.A1(new_n7274_), .A2(new_n7276_), .A3(new_n3675_), .ZN(new_n7277_));
  INV_X1     g07085(.I(new_n7183_), .ZN(new_n7278_));
  INV_X1     g07086(.I(new_n7193_), .ZN(new_n7279_));
  NOR2_X1    g07087(.A1(new_n7266_), .A2(new_n7267_), .ZN(new_n7280_));
  AOI21_X1   g07088(.A1(new_n7280_), .A2(new_n4810_), .B(new_n7279_), .ZN(new_n7281_));
  NAND2_X1   g07089(.A1(new_n7268_), .A2(new_n4510_), .ZN(new_n7282_));
  OAI21_X1   g07090(.A1(new_n7281_), .A2(new_n7282_), .B(new_n7189_), .ZN(new_n7283_));
  INV_X1     g07091(.I(new_n7268_), .ZN(new_n7284_));
  OAI21_X1   g07092(.A1(new_n7281_), .A2(new_n7284_), .B(\asqrt[35] ), .ZN(new_n7285_));
  NAND3_X1   g07093(.A1(new_n7283_), .A2(new_n7285_), .A3(new_n4224_), .ZN(new_n7286_));
  NAND2_X1   g07094(.A1(new_n7286_), .A2(new_n7186_), .ZN(new_n7287_));
  NAND2_X1   g07095(.A1(new_n7283_), .A2(new_n7285_), .ZN(new_n7288_));
  AOI21_X1   g07096(.A1(new_n7288_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n7289_));
  AOI21_X1   g07097(.A1(new_n7289_), .A2(new_n7287_), .B(new_n7278_), .ZN(new_n7290_));
  AOI21_X1   g07098(.A1(new_n7287_), .A2(new_n7272_), .B(new_n3928_), .ZN(new_n7291_));
  OAI21_X1   g07099(.A1(new_n7290_), .A2(new_n7291_), .B(\asqrt[38] ), .ZN(new_n7292_));
  NAND2_X1   g07100(.A1(new_n7163_), .A2(new_n6818_), .ZN(new_n7293_));
  NOR2_X1    g07101(.A1(new_n7166_), .A2(new_n6818_), .ZN(new_n7294_));
  NAND2_X1   g07102(.A1(new_n7294_), .A2(new_n7178_), .ZN(new_n7295_));
  AOI21_X1   g07103(.A1(new_n7295_), .A2(new_n7293_), .B(new_n193_), .ZN(new_n7296_));
  INV_X1     g07104(.I(new_n7296_), .ZN(new_n7297_));
  NAND3_X1   g07105(.A1(\asqrt[27] ), .A2(new_n7148_), .A3(new_n7159_), .ZN(new_n7298_));
  XOR2_X1    g07106(.A1(new_n7298_), .A2(new_n7151_), .Z(new_n7299_));
  AOI21_X1   g07107(.A1(new_n7294_), .A2(new_n7163_), .B(new_n7164_), .ZN(new_n7300_));
  OAI21_X1   g07108(.A1(new_n7118_), .A2(new_n7120_), .B(new_n7123_), .ZN(new_n7301_));
  NOR2_X1    g07109(.A1(new_n7166_), .A2(new_n7301_), .ZN(new_n7302_));
  XOR2_X1    g07110(.A1(new_n7302_), .A2(new_n6826_), .Z(new_n7303_));
  NAND3_X1   g07111(.A1(\asqrt[27] ), .A2(new_n7134_), .A3(new_n7119_), .ZN(new_n7304_));
  XOR2_X1    g07112(.A1(new_n7304_), .A2(new_n6830_), .Z(new_n7305_));
  OAI21_X1   g07113(.A1(new_n7129_), .A2(new_n7130_), .B(new_n7133_), .ZN(new_n7306_));
  NOR2_X1    g07114(.A1(new_n7166_), .A2(new_n7306_), .ZN(new_n7307_));
  XOR2_X1    g07115(.A1(new_n7307_), .A2(new_n6832_), .Z(new_n7308_));
  INV_X1     g07116(.I(new_n7308_), .ZN(new_n7309_));
  NAND3_X1   g07117(.A1(\asqrt[27] ), .A2(new_n7096_), .A3(new_n7115_), .ZN(new_n7310_));
  XOR2_X1    g07118(.A1(new_n7310_), .A2(new_n7127_), .Z(new_n7311_));
  INV_X1     g07119(.I(new_n7311_), .ZN(new_n7312_));
  OAI21_X1   g07120(.A1(new_n7090_), .A2(new_n7092_), .B(new_n7095_), .ZN(new_n7313_));
  NOR2_X1    g07121(.A1(new_n7166_), .A2(new_n7313_), .ZN(new_n7314_));
  XOR2_X1    g07122(.A1(new_n7314_), .A2(new_n6838_), .Z(new_n7315_));
  NAND3_X1   g07123(.A1(\asqrt[27] ), .A2(new_n7109_), .A3(new_n7091_), .ZN(new_n7316_));
  XOR2_X1    g07124(.A1(new_n7316_), .A2(new_n6842_), .Z(new_n7317_));
  OAI21_X1   g07125(.A1(new_n7104_), .A2(new_n7105_), .B(new_n7108_), .ZN(new_n7318_));
  NOR2_X1    g07126(.A1(new_n7166_), .A2(new_n7318_), .ZN(new_n7319_));
  XOR2_X1    g07127(.A1(new_n7319_), .A2(new_n6844_), .Z(new_n7320_));
  INV_X1     g07128(.I(new_n7320_), .ZN(new_n7321_));
  NAND3_X1   g07129(.A1(\asqrt[27] ), .A2(new_n7068_), .A3(new_n7087_), .ZN(new_n7322_));
  XOR2_X1    g07130(.A1(new_n7322_), .A2(new_n7102_), .Z(new_n7323_));
  INV_X1     g07131(.I(new_n7323_), .ZN(new_n7324_));
  OAI21_X1   g07132(.A1(new_n7062_), .A2(new_n7064_), .B(new_n7067_), .ZN(new_n7325_));
  NOR2_X1    g07133(.A1(new_n7166_), .A2(new_n7325_), .ZN(new_n7326_));
  XOR2_X1    g07134(.A1(new_n7326_), .A2(new_n6850_), .Z(new_n7327_));
  NAND3_X1   g07135(.A1(\asqrt[27] ), .A2(new_n7081_), .A3(new_n7063_), .ZN(new_n7328_));
  XOR2_X1    g07136(.A1(new_n7328_), .A2(new_n6854_), .Z(new_n7329_));
  OAI21_X1   g07137(.A1(new_n7076_), .A2(new_n7077_), .B(new_n7080_), .ZN(new_n7330_));
  NOR2_X1    g07138(.A1(new_n7166_), .A2(new_n7330_), .ZN(new_n7331_));
  XOR2_X1    g07139(.A1(new_n7331_), .A2(new_n6856_), .Z(new_n7332_));
  INV_X1     g07140(.I(new_n7332_), .ZN(new_n7333_));
  NAND3_X1   g07141(.A1(\asqrt[27] ), .A2(new_n7040_), .A3(new_n7059_), .ZN(new_n7334_));
  XOR2_X1    g07142(.A1(new_n7334_), .A2(new_n7074_), .Z(new_n7335_));
  INV_X1     g07143(.I(new_n7335_), .ZN(new_n7336_));
  OAI21_X1   g07144(.A1(new_n7034_), .A2(new_n7036_), .B(new_n7039_), .ZN(new_n7337_));
  NOR2_X1    g07145(.A1(new_n7166_), .A2(new_n7337_), .ZN(new_n7338_));
  XOR2_X1    g07146(.A1(new_n7338_), .A2(new_n6862_), .Z(new_n7339_));
  NAND3_X1   g07147(.A1(\asqrt[27] ), .A2(new_n7053_), .A3(new_n7035_), .ZN(new_n7340_));
  XOR2_X1    g07148(.A1(new_n7340_), .A2(new_n6866_), .Z(new_n7341_));
  OAI21_X1   g07149(.A1(new_n7048_), .A2(new_n7049_), .B(new_n7052_), .ZN(new_n7342_));
  NOR2_X1    g07150(.A1(new_n7166_), .A2(new_n7342_), .ZN(new_n7343_));
  XOR2_X1    g07151(.A1(new_n7343_), .A2(new_n6868_), .Z(new_n7344_));
  INV_X1     g07152(.I(new_n7344_), .ZN(new_n7345_));
  NAND3_X1   g07153(.A1(\asqrt[27] ), .A2(new_n7012_), .A3(new_n7031_), .ZN(new_n7346_));
  XOR2_X1    g07154(.A1(new_n7346_), .A2(new_n7046_), .Z(new_n7347_));
  INV_X1     g07155(.I(new_n7347_), .ZN(new_n7348_));
  OAI21_X1   g07156(.A1(new_n7006_), .A2(new_n7008_), .B(new_n7011_), .ZN(new_n7349_));
  NOR2_X1    g07157(.A1(new_n7166_), .A2(new_n7349_), .ZN(new_n7350_));
  XOR2_X1    g07158(.A1(new_n7350_), .A2(new_n6874_), .Z(new_n7351_));
  NAND3_X1   g07159(.A1(\asqrt[27] ), .A2(new_n7025_), .A3(new_n7007_), .ZN(new_n7352_));
  XOR2_X1    g07160(.A1(new_n7352_), .A2(new_n6878_), .Z(new_n7353_));
  OAI21_X1   g07161(.A1(new_n7020_), .A2(new_n7021_), .B(new_n7024_), .ZN(new_n7354_));
  NOR2_X1    g07162(.A1(new_n7166_), .A2(new_n7354_), .ZN(new_n7355_));
  XOR2_X1    g07163(.A1(new_n7355_), .A2(new_n6880_), .Z(new_n7356_));
  INV_X1     g07164(.I(new_n7356_), .ZN(new_n7357_));
  NAND3_X1   g07165(.A1(\asqrt[27] ), .A2(new_n6984_), .A3(new_n7003_), .ZN(new_n7358_));
  XOR2_X1    g07166(.A1(new_n7358_), .A2(new_n7018_), .Z(new_n7359_));
  INV_X1     g07167(.I(new_n7359_), .ZN(new_n7360_));
  OAI21_X1   g07168(.A1(new_n6978_), .A2(new_n6980_), .B(new_n6983_), .ZN(new_n7361_));
  NOR2_X1    g07169(.A1(new_n7166_), .A2(new_n7361_), .ZN(new_n7362_));
  XOR2_X1    g07170(.A1(new_n7362_), .A2(new_n6886_), .Z(new_n7363_));
  NAND3_X1   g07171(.A1(\asqrt[27] ), .A2(new_n6997_), .A3(new_n6979_), .ZN(new_n7364_));
  XOR2_X1    g07172(.A1(new_n7364_), .A2(new_n6890_), .Z(new_n7365_));
  NOR2_X1    g07173(.A1(new_n7290_), .A2(new_n7291_), .ZN(new_n7366_));
  AOI21_X1   g07174(.A1(new_n7366_), .A2(new_n3675_), .B(new_n7170_), .ZN(new_n7367_));
  NAND2_X1   g07175(.A1(new_n7292_), .A2(new_n3400_), .ZN(new_n7368_));
  OAI21_X1   g07176(.A1(new_n7367_), .A2(new_n7368_), .B(new_n7365_), .ZN(new_n7369_));
  INV_X1     g07177(.I(new_n7292_), .ZN(new_n7370_));
  OAI21_X1   g07178(.A1(new_n7367_), .A2(new_n7370_), .B(\asqrt[39] ), .ZN(new_n7371_));
  NAND3_X1   g07179(.A1(new_n7369_), .A2(new_n7371_), .A3(new_n3167_), .ZN(new_n7372_));
  NAND2_X1   g07180(.A1(new_n7372_), .A2(new_n7363_), .ZN(new_n7373_));
  NAND2_X1   g07181(.A1(new_n7369_), .A2(new_n7371_), .ZN(new_n7374_));
  AOI21_X1   g07182(.A1(new_n7374_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n7375_));
  AOI21_X1   g07183(.A1(new_n7375_), .A2(new_n7373_), .B(new_n7360_), .ZN(new_n7376_));
  INV_X1     g07184(.I(new_n7365_), .ZN(new_n7377_));
  NAND2_X1   g07185(.A1(new_n7277_), .A2(new_n7169_), .ZN(new_n7378_));
  NAND2_X1   g07186(.A1(new_n7274_), .A2(new_n7276_), .ZN(new_n7379_));
  AOI21_X1   g07187(.A1(new_n7379_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n7380_));
  AOI21_X1   g07188(.A1(new_n7380_), .A2(new_n7378_), .B(new_n7377_), .ZN(new_n7381_));
  AOI21_X1   g07189(.A1(new_n7378_), .A2(new_n7292_), .B(new_n3400_), .ZN(new_n7382_));
  OAI21_X1   g07190(.A1(new_n7381_), .A2(new_n7382_), .B(\asqrt[40] ), .ZN(new_n7383_));
  AOI21_X1   g07191(.A1(new_n7373_), .A2(new_n7383_), .B(new_n2912_), .ZN(new_n7384_));
  NOR2_X1    g07192(.A1(new_n7376_), .A2(new_n7384_), .ZN(new_n7385_));
  AOI21_X1   g07193(.A1(new_n7385_), .A2(new_n2699_), .B(new_n7357_), .ZN(new_n7386_));
  OAI21_X1   g07194(.A1(new_n7376_), .A2(new_n7384_), .B(\asqrt[42] ), .ZN(new_n7387_));
  NAND2_X1   g07195(.A1(new_n7387_), .A2(new_n2464_), .ZN(new_n7388_));
  OAI21_X1   g07196(.A1(new_n7386_), .A2(new_n7388_), .B(new_n7353_), .ZN(new_n7389_));
  INV_X1     g07197(.I(new_n7387_), .ZN(new_n7390_));
  OAI21_X1   g07198(.A1(new_n7386_), .A2(new_n7390_), .B(\asqrt[43] ), .ZN(new_n7391_));
  NAND3_X1   g07199(.A1(new_n7389_), .A2(new_n7391_), .A3(new_n2271_), .ZN(new_n7392_));
  NAND2_X1   g07200(.A1(new_n7392_), .A2(new_n7351_), .ZN(new_n7393_));
  NAND2_X1   g07201(.A1(new_n7389_), .A2(new_n7391_), .ZN(new_n7394_));
  AOI21_X1   g07202(.A1(new_n7394_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n7395_));
  AOI21_X1   g07203(.A1(new_n7395_), .A2(new_n7393_), .B(new_n7348_), .ZN(new_n7396_));
  INV_X1     g07204(.I(new_n7353_), .ZN(new_n7397_));
  INV_X1     g07205(.I(new_n7363_), .ZN(new_n7398_));
  NOR2_X1    g07206(.A1(new_n7381_), .A2(new_n7382_), .ZN(new_n7399_));
  AOI21_X1   g07207(.A1(new_n7399_), .A2(new_n3167_), .B(new_n7398_), .ZN(new_n7400_));
  NAND2_X1   g07208(.A1(new_n7383_), .A2(new_n2912_), .ZN(new_n7401_));
  OAI21_X1   g07209(.A1(new_n7400_), .A2(new_n7401_), .B(new_n7359_), .ZN(new_n7402_));
  INV_X1     g07210(.I(new_n7383_), .ZN(new_n7403_));
  OAI21_X1   g07211(.A1(new_n7400_), .A2(new_n7403_), .B(\asqrt[41] ), .ZN(new_n7404_));
  NAND3_X1   g07212(.A1(new_n7402_), .A2(new_n7404_), .A3(new_n2699_), .ZN(new_n7405_));
  NAND2_X1   g07213(.A1(new_n7405_), .A2(new_n7356_), .ZN(new_n7406_));
  NAND2_X1   g07214(.A1(new_n7402_), .A2(new_n7404_), .ZN(new_n7407_));
  AOI21_X1   g07215(.A1(new_n7407_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n7408_));
  AOI21_X1   g07216(.A1(new_n7408_), .A2(new_n7406_), .B(new_n7397_), .ZN(new_n7409_));
  AOI21_X1   g07217(.A1(new_n7406_), .A2(new_n7387_), .B(new_n2464_), .ZN(new_n7410_));
  OAI21_X1   g07218(.A1(new_n7409_), .A2(new_n7410_), .B(\asqrt[44] ), .ZN(new_n7411_));
  AOI21_X1   g07219(.A1(new_n7393_), .A2(new_n7411_), .B(new_n2072_), .ZN(new_n7412_));
  NOR2_X1    g07220(.A1(new_n7396_), .A2(new_n7412_), .ZN(new_n7413_));
  AOI21_X1   g07221(.A1(new_n7413_), .A2(new_n1884_), .B(new_n7345_), .ZN(new_n7414_));
  OAI21_X1   g07222(.A1(new_n7396_), .A2(new_n7412_), .B(\asqrt[46] ), .ZN(new_n7415_));
  NAND2_X1   g07223(.A1(new_n7415_), .A2(new_n1688_), .ZN(new_n7416_));
  OAI21_X1   g07224(.A1(new_n7414_), .A2(new_n7416_), .B(new_n7341_), .ZN(new_n7417_));
  INV_X1     g07225(.I(new_n7415_), .ZN(new_n7418_));
  OAI21_X1   g07226(.A1(new_n7414_), .A2(new_n7418_), .B(\asqrt[47] ), .ZN(new_n7419_));
  NAND3_X1   g07227(.A1(new_n7417_), .A2(new_n7419_), .A3(new_n1533_), .ZN(new_n7420_));
  NAND2_X1   g07228(.A1(new_n7420_), .A2(new_n7339_), .ZN(new_n7421_));
  NAND2_X1   g07229(.A1(new_n7417_), .A2(new_n7419_), .ZN(new_n7422_));
  AOI21_X1   g07230(.A1(new_n7422_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n7423_));
  AOI21_X1   g07231(.A1(new_n7423_), .A2(new_n7421_), .B(new_n7336_), .ZN(new_n7424_));
  INV_X1     g07232(.I(new_n7341_), .ZN(new_n7425_));
  INV_X1     g07233(.I(new_n7351_), .ZN(new_n7426_));
  NOR2_X1    g07234(.A1(new_n7409_), .A2(new_n7410_), .ZN(new_n7427_));
  AOI21_X1   g07235(.A1(new_n7427_), .A2(new_n2271_), .B(new_n7426_), .ZN(new_n7428_));
  NAND2_X1   g07236(.A1(new_n7411_), .A2(new_n2072_), .ZN(new_n7429_));
  OAI21_X1   g07237(.A1(new_n7428_), .A2(new_n7429_), .B(new_n7347_), .ZN(new_n7430_));
  INV_X1     g07238(.I(new_n7411_), .ZN(new_n7431_));
  OAI21_X1   g07239(.A1(new_n7428_), .A2(new_n7431_), .B(\asqrt[45] ), .ZN(new_n7432_));
  NAND3_X1   g07240(.A1(new_n7430_), .A2(new_n7432_), .A3(new_n1884_), .ZN(new_n7433_));
  NAND2_X1   g07241(.A1(new_n7433_), .A2(new_n7344_), .ZN(new_n7434_));
  NAND2_X1   g07242(.A1(new_n7430_), .A2(new_n7432_), .ZN(new_n7435_));
  AOI21_X1   g07243(.A1(new_n7435_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n7436_));
  AOI21_X1   g07244(.A1(new_n7436_), .A2(new_n7434_), .B(new_n7425_), .ZN(new_n7437_));
  AOI21_X1   g07245(.A1(new_n7434_), .A2(new_n7415_), .B(new_n1688_), .ZN(new_n7438_));
  OAI21_X1   g07246(.A1(new_n7437_), .A2(new_n7438_), .B(\asqrt[48] ), .ZN(new_n7439_));
  AOI21_X1   g07247(.A1(new_n7421_), .A2(new_n7439_), .B(new_n1368_), .ZN(new_n7440_));
  NOR2_X1    g07248(.A1(new_n7424_), .A2(new_n7440_), .ZN(new_n7441_));
  AOI21_X1   g07249(.A1(new_n7441_), .A2(new_n1228_), .B(new_n7333_), .ZN(new_n7442_));
  OAI21_X1   g07250(.A1(new_n7424_), .A2(new_n7440_), .B(\asqrt[50] ), .ZN(new_n7443_));
  NAND2_X1   g07251(.A1(new_n7443_), .A2(new_n1088_), .ZN(new_n7444_));
  OAI21_X1   g07252(.A1(new_n7442_), .A2(new_n7444_), .B(new_n7329_), .ZN(new_n7445_));
  INV_X1     g07253(.I(new_n7443_), .ZN(new_n7446_));
  OAI21_X1   g07254(.A1(new_n7442_), .A2(new_n7446_), .B(\asqrt[51] ), .ZN(new_n7447_));
  NAND3_X1   g07255(.A1(new_n7445_), .A2(new_n7447_), .A3(new_n962_), .ZN(new_n7448_));
  NAND2_X1   g07256(.A1(new_n7448_), .A2(new_n7327_), .ZN(new_n7449_));
  NAND2_X1   g07257(.A1(new_n7445_), .A2(new_n7447_), .ZN(new_n7450_));
  AOI21_X1   g07258(.A1(new_n7450_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n7451_));
  AOI21_X1   g07259(.A1(new_n7451_), .A2(new_n7449_), .B(new_n7324_), .ZN(new_n7452_));
  INV_X1     g07260(.I(new_n7329_), .ZN(new_n7453_));
  INV_X1     g07261(.I(new_n7339_), .ZN(new_n7454_));
  NOR2_X1    g07262(.A1(new_n7437_), .A2(new_n7438_), .ZN(new_n7455_));
  AOI21_X1   g07263(.A1(new_n7455_), .A2(new_n1533_), .B(new_n7454_), .ZN(new_n7456_));
  NAND2_X1   g07264(.A1(new_n7439_), .A2(new_n1368_), .ZN(new_n7457_));
  OAI21_X1   g07265(.A1(new_n7456_), .A2(new_n7457_), .B(new_n7335_), .ZN(new_n7458_));
  INV_X1     g07266(.I(new_n7439_), .ZN(new_n7459_));
  OAI21_X1   g07267(.A1(new_n7456_), .A2(new_n7459_), .B(\asqrt[49] ), .ZN(new_n7460_));
  NAND3_X1   g07268(.A1(new_n7458_), .A2(new_n7460_), .A3(new_n1228_), .ZN(new_n7461_));
  NAND2_X1   g07269(.A1(new_n7461_), .A2(new_n7332_), .ZN(new_n7462_));
  NAND2_X1   g07270(.A1(new_n7458_), .A2(new_n7460_), .ZN(new_n7463_));
  AOI21_X1   g07271(.A1(new_n7463_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n7464_));
  AOI21_X1   g07272(.A1(new_n7464_), .A2(new_n7462_), .B(new_n7453_), .ZN(new_n7465_));
  AOI21_X1   g07273(.A1(new_n7462_), .A2(new_n7443_), .B(new_n1088_), .ZN(new_n7466_));
  OAI21_X1   g07274(.A1(new_n7465_), .A2(new_n7466_), .B(\asqrt[52] ), .ZN(new_n7467_));
  AOI21_X1   g07275(.A1(new_n7449_), .A2(new_n7467_), .B(new_n842_), .ZN(new_n7468_));
  NOR2_X1    g07276(.A1(new_n7452_), .A2(new_n7468_), .ZN(new_n7469_));
  AOI21_X1   g07277(.A1(new_n7469_), .A2(new_n720_), .B(new_n7321_), .ZN(new_n7470_));
  OAI21_X1   g07278(.A1(new_n7452_), .A2(new_n7468_), .B(\asqrt[54] ), .ZN(new_n7471_));
  NAND2_X1   g07279(.A1(new_n7471_), .A2(new_n630_), .ZN(new_n7472_));
  OAI21_X1   g07280(.A1(new_n7470_), .A2(new_n7472_), .B(new_n7317_), .ZN(new_n7473_));
  INV_X1     g07281(.I(new_n7471_), .ZN(new_n7474_));
  OAI21_X1   g07282(.A1(new_n7470_), .A2(new_n7474_), .B(\asqrt[55] ), .ZN(new_n7475_));
  NAND3_X1   g07283(.A1(new_n7473_), .A2(new_n7475_), .A3(new_n545_), .ZN(new_n7476_));
  NAND2_X1   g07284(.A1(new_n7476_), .A2(new_n7315_), .ZN(new_n7477_));
  NAND2_X1   g07285(.A1(new_n7473_), .A2(new_n7475_), .ZN(new_n7478_));
  AOI21_X1   g07286(.A1(new_n7478_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n7479_));
  AOI21_X1   g07287(.A1(new_n7479_), .A2(new_n7477_), .B(new_n7312_), .ZN(new_n7480_));
  INV_X1     g07288(.I(new_n7317_), .ZN(new_n7481_));
  INV_X1     g07289(.I(new_n7327_), .ZN(new_n7482_));
  NOR2_X1    g07290(.A1(new_n7465_), .A2(new_n7466_), .ZN(new_n7483_));
  AOI21_X1   g07291(.A1(new_n7483_), .A2(new_n962_), .B(new_n7482_), .ZN(new_n7484_));
  NAND2_X1   g07292(.A1(new_n7467_), .A2(new_n842_), .ZN(new_n7485_));
  OAI21_X1   g07293(.A1(new_n7484_), .A2(new_n7485_), .B(new_n7323_), .ZN(new_n7486_));
  INV_X1     g07294(.I(new_n7467_), .ZN(new_n7487_));
  OAI21_X1   g07295(.A1(new_n7484_), .A2(new_n7487_), .B(\asqrt[53] ), .ZN(new_n7488_));
  NAND3_X1   g07296(.A1(new_n7486_), .A2(new_n7488_), .A3(new_n720_), .ZN(new_n7489_));
  NAND2_X1   g07297(.A1(new_n7489_), .A2(new_n7320_), .ZN(new_n7490_));
  NAND2_X1   g07298(.A1(new_n7486_), .A2(new_n7488_), .ZN(new_n7491_));
  AOI21_X1   g07299(.A1(new_n7491_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n7492_));
  AOI21_X1   g07300(.A1(new_n7492_), .A2(new_n7490_), .B(new_n7481_), .ZN(new_n7493_));
  AOI21_X1   g07301(.A1(new_n7490_), .A2(new_n7471_), .B(new_n630_), .ZN(new_n7494_));
  OAI21_X1   g07302(.A1(new_n7493_), .A2(new_n7494_), .B(\asqrt[56] ), .ZN(new_n7495_));
  AOI21_X1   g07303(.A1(new_n7477_), .A2(new_n7495_), .B(new_n450_), .ZN(new_n7496_));
  NOR2_X1    g07304(.A1(new_n7480_), .A2(new_n7496_), .ZN(new_n7497_));
  AOI21_X1   g07305(.A1(new_n7497_), .A2(new_n403_), .B(new_n7309_), .ZN(new_n7498_));
  OAI21_X1   g07306(.A1(new_n7480_), .A2(new_n7496_), .B(\asqrt[58] ), .ZN(new_n7499_));
  NAND2_X1   g07307(.A1(new_n7499_), .A2(new_n339_), .ZN(new_n7500_));
  OAI21_X1   g07308(.A1(new_n7498_), .A2(new_n7500_), .B(new_n7305_), .ZN(new_n7501_));
  INV_X1     g07309(.I(new_n7499_), .ZN(new_n7502_));
  OAI21_X1   g07310(.A1(new_n7498_), .A2(new_n7502_), .B(\asqrt[59] ), .ZN(new_n7503_));
  NAND3_X1   g07311(.A1(new_n7501_), .A2(new_n7503_), .A3(new_n288_), .ZN(new_n7504_));
  NAND2_X1   g07312(.A1(new_n7504_), .A2(new_n7303_), .ZN(new_n7505_));
  INV_X1     g07313(.I(new_n7305_), .ZN(new_n7506_));
  INV_X1     g07314(.I(new_n7315_), .ZN(new_n7507_));
  NOR2_X1    g07315(.A1(new_n7493_), .A2(new_n7494_), .ZN(new_n7508_));
  AOI21_X1   g07316(.A1(new_n7508_), .A2(new_n545_), .B(new_n7507_), .ZN(new_n7509_));
  NAND2_X1   g07317(.A1(new_n7495_), .A2(new_n450_), .ZN(new_n7510_));
  OAI21_X1   g07318(.A1(new_n7509_), .A2(new_n7510_), .B(new_n7311_), .ZN(new_n7511_));
  INV_X1     g07319(.I(new_n7495_), .ZN(new_n7512_));
  OAI21_X1   g07320(.A1(new_n7509_), .A2(new_n7512_), .B(\asqrt[57] ), .ZN(new_n7513_));
  NAND3_X1   g07321(.A1(new_n7511_), .A2(new_n7513_), .A3(new_n403_), .ZN(new_n7514_));
  NAND2_X1   g07322(.A1(new_n7514_), .A2(new_n7308_), .ZN(new_n7515_));
  NAND2_X1   g07323(.A1(new_n7511_), .A2(new_n7513_), .ZN(new_n7516_));
  AOI21_X1   g07324(.A1(new_n7516_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n7517_));
  AOI21_X1   g07325(.A1(new_n7517_), .A2(new_n7515_), .B(new_n7506_), .ZN(new_n7518_));
  AOI21_X1   g07326(.A1(new_n7515_), .A2(new_n7499_), .B(new_n339_), .ZN(new_n7519_));
  OAI21_X1   g07327(.A1(new_n7518_), .A2(new_n7519_), .B(\asqrt[60] ), .ZN(new_n7520_));
  AOI21_X1   g07328(.A1(new_n7505_), .A2(new_n7520_), .B(new_n242_), .ZN(new_n7521_));
  NAND3_X1   g07329(.A1(\asqrt[27] ), .A2(new_n7124_), .A3(new_n7140_), .ZN(new_n7522_));
  XOR2_X1    g07330(.A1(new_n7522_), .A2(new_n7152_), .Z(new_n7523_));
  INV_X1     g07331(.I(new_n7523_), .ZN(new_n7524_));
  NAND2_X1   g07332(.A1(new_n7501_), .A2(new_n7503_), .ZN(new_n7525_));
  AOI21_X1   g07333(.A1(new_n7525_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n7526_));
  AOI21_X1   g07334(.A1(new_n7526_), .A2(new_n7505_), .B(new_n7524_), .ZN(new_n7527_));
  OAI21_X1   g07335(.A1(new_n7527_), .A2(new_n7521_), .B(\asqrt[62] ), .ZN(new_n7528_));
  INV_X1     g07336(.I(new_n7528_), .ZN(new_n7529_));
  NOR2_X1    g07337(.A1(new_n7527_), .A2(new_n7521_), .ZN(new_n7530_));
  AOI21_X1   g07338(.A1(new_n7125_), .A2(new_n7146_), .B(new_n7141_), .ZN(new_n7531_));
  NAND2_X1   g07339(.A1(\asqrt[27] ), .A2(new_n7531_), .ZN(new_n7532_));
  XOR2_X1    g07340(.A1(new_n7532_), .A2(new_n7144_), .Z(new_n7533_));
  INV_X1     g07341(.I(new_n7533_), .ZN(new_n7534_));
  AOI21_X1   g07342(.A1(new_n7530_), .A2(new_n234_), .B(new_n7534_), .ZN(new_n7535_));
  OAI21_X1   g07343(.A1(new_n7535_), .A2(new_n7529_), .B(new_n7300_), .ZN(new_n7536_));
  OAI21_X1   g07344(.A1(new_n7536_), .A2(new_n7299_), .B(new_n193_), .ZN(new_n7537_));
  NOR2_X1    g07345(.A1(new_n7535_), .A2(new_n7529_), .ZN(new_n7538_));
  NAND2_X1   g07346(.A1(new_n7538_), .A2(new_n7299_), .ZN(new_n7539_));
  NOR2_X1    g07347(.A1(\asqrt[27] ), .A2(new_n6819_), .ZN(new_n7540_));
  INV_X1     g07348(.I(new_n7540_), .ZN(new_n7541_));
  NAND4_X1   g07349(.A1(new_n7537_), .A2(new_n7297_), .A3(new_n7539_), .A4(new_n7541_), .ZN(\asqrt[26] ));
  NAND3_X1   g07350(.A1(\asqrt[26] ), .A2(new_n7277_), .A3(new_n7292_), .ZN(new_n7543_));
  XOR2_X1    g07351(.A1(new_n7543_), .A2(new_n7170_), .Z(new_n7544_));
  INV_X1     g07352(.I(new_n7303_), .ZN(new_n7545_));
  NOR2_X1    g07353(.A1(new_n7518_), .A2(new_n7519_), .ZN(new_n7546_));
  AOI21_X1   g07354(.A1(new_n7546_), .A2(new_n288_), .B(new_n7545_), .ZN(new_n7547_));
  INV_X1     g07355(.I(new_n7520_), .ZN(new_n7548_));
  OAI21_X1   g07356(.A1(new_n7547_), .A2(new_n7548_), .B(\asqrt[61] ), .ZN(new_n7549_));
  NAND2_X1   g07357(.A1(new_n7520_), .A2(new_n242_), .ZN(new_n7550_));
  OAI21_X1   g07358(.A1(new_n7547_), .A2(new_n7550_), .B(new_n7523_), .ZN(new_n7551_));
  NAND3_X1   g07359(.A1(new_n7551_), .A2(new_n7549_), .A3(new_n234_), .ZN(new_n7552_));
  NAND2_X1   g07360(.A1(new_n7552_), .A2(new_n7533_), .ZN(new_n7553_));
  NAND2_X1   g07361(.A1(new_n7553_), .A2(new_n7528_), .ZN(new_n7554_));
  NAND2_X1   g07362(.A1(new_n7554_), .A2(new_n7299_), .ZN(new_n7555_));
  INV_X1     g07363(.I(new_n7299_), .ZN(new_n7556_));
  INV_X1     g07364(.I(new_n7300_), .ZN(new_n7557_));
  AOI21_X1   g07365(.A1(new_n7553_), .A2(new_n7528_), .B(new_n7557_), .ZN(new_n7558_));
  AOI21_X1   g07366(.A1(new_n7558_), .A2(new_n7556_), .B(\asqrt[63] ), .ZN(new_n7559_));
  NOR2_X1    g07367(.A1(new_n7554_), .A2(new_n7556_), .ZN(new_n7560_));
  NOR4_X1    g07368(.A1(new_n7559_), .A2(new_n7296_), .A3(new_n7560_), .A4(new_n7540_), .ZN(new_n7561_));
  NOR2_X1    g07369(.A1(new_n7561_), .A2(new_n7299_), .ZN(new_n7562_));
  NAND2_X1   g07370(.A1(new_n7562_), .A2(new_n7538_), .ZN(new_n7563_));
  AOI21_X1   g07371(.A1(new_n7563_), .A2(new_n7555_), .B(new_n193_), .ZN(new_n7564_));
  NAND3_X1   g07372(.A1(\asqrt[26] ), .A2(new_n7528_), .A3(new_n7552_), .ZN(new_n7565_));
  XOR2_X1    g07373(.A1(new_n7565_), .A2(new_n7533_), .Z(new_n7566_));
  INV_X1     g07374(.I(new_n7566_), .ZN(new_n7567_));
  AOI21_X1   g07375(.A1(new_n7562_), .A2(new_n7554_), .B(new_n7560_), .ZN(new_n7568_));
  INV_X1     g07376(.I(new_n7568_), .ZN(new_n7569_));
  OAI21_X1   g07377(.A1(new_n7498_), .A2(new_n7500_), .B(new_n7503_), .ZN(new_n7570_));
  NOR2_X1    g07378(.A1(new_n7561_), .A2(new_n7570_), .ZN(new_n7571_));
  XOR2_X1    g07379(.A1(new_n7571_), .A2(new_n7305_), .Z(new_n7572_));
  NAND3_X1   g07380(.A1(\asqrt[26] ), .A2(new_n7514_), .A3(new_n7499_), .ZN(new_n7573_));
  XOR2_X1    g07381(.A1(new_n7573_), .A2(new_n7309_), .Z(new_n7574_));
  OAI21_X1   g07382(.A1(new_n7509_), .A2(new_n7510_), .B(new_n7513_), .ZN(new_n7575_));
  NOR2_X1    g07383(.A1(new_n7561_), .A2(new_n7575_), .ZN(new_n7576_));
  XOR2_X1    g07384(.A1(new_n7576_), .A2(new_n7311_), .Z(new_n7577_));
  INV_X1     g07385(.I(new_n7577_), .ZN(new_n7578_));
  NAND3_X1   g07386(.A1(\asqrt[26] ), .A2(new_n7476_), .A3(new_n7495_), .ZN(new_n7579_));
  XOR2_X1    g07387(.A1(new_n7579_), .A2(new_n7507_), .Z(new_n7580_));
  INV_X1     g07388(.I(new_n7580_), .ZN(new_n7581_));
  OAI21_X1   g07389(.A1(new_n7470_), .A2(new_n7472_), .B(new_n7475_), .ZN(new_n7582_));
  NOR2_X1    g07390(.A1(new_n7561_), .A2(new_n7582_), .ZN(new_n7583_));
  XOR2_X1    g07391(.A1(new_n7583_), .A2(new_n7317_), .Z(new_n7584_));
  NAND3_X1   g07392(.A1(\asqrt[26] ), .A2(new_n7489_), .A3(new_n7471_), .ZN(new_n7585_));
  XOR2_X1    g07393(.A1(new_n7585_), .A2(new_n7321_), .Z(new_n7586_));
  OAI21_X1   g07394(.A1(new_n7484_), .A2(new_n7485_), .B(new_n7488_), .ZN(new_n7587_));
  NOR2_X1    g07395(.A1(new_n7561_), .A2(new_n7587_), .ZN(new_n7588_));
  XOR2_X1    g07396(.A1(new_n7588_), .A2(new_n7323_), .Z(new_n7589_));
  INV_X1     g07397(.I(new_n7589_), .ZN(new_n7590_));
  NAND3_X1   g07398(.A1(\asqrt[26] ), .A2(new_n7448_), .A3(new_n7467_), .ZN(new_n7591_));
  XOR2_X1    g07399(.A1(new_n7591_), .A2(new_n7482_), .Z(new_n7592_));
  INV_X1     g07400(.I(new_n7592_), .ZN(new_n7593_));
  OAI21_X1   g07401(.A1(new_n7442_), .A2(new_n7444_), .B(new_n7447_), .ZN(new_n7594_));
  NOR2_X1    g07402(.A1(new_n7561_), .A2(new_n7594_), .ZN(new_n7595_));
  XOR2_X1    g07403(.A1(new_n7595_), .A2(new_n7329_), .Z(new_n7596_));
  NAND3_X1   g07404(.A1(\asqrt[26] ), .A2(new_n7461_), .A3(new_n7443_), .ZN(new_n7597_));
  XOR2_X1    g07405(.A1(new_n7597_), .A2(new_n7333_), .Z(new_n7598_));
  OAI21_X1   g07406(.A1(new_n7456_), .A2(new_n7457_), .B(new_n7460_), .ZN(new_n7599_));
  NOR2_X1    g07407(.A1(new_n7561_), .A2(new_n7599_), .ZN(new_n7600_));
  XOR2_X1    g07408(.A1(new_n7600_), .A2(new_n7335_), .Z(new_n7601_));
  INV_X1     g07409(.I(new_n7601_), .ZN(new_n7602_));
  NAND3_X1   g07410(.A1(\asqrt[26] ), .A2(new_n7420_), .A3(new_n7439_), .ZN(new_n7603_));
  XOR2_X1    g07411(.A1(new_n7603_), .A2(new_n7454_), .Z(new_n7604_));
  INV_X1     g07412(.I(new_n7604_), .ZN(new_n7605_));
  OAI21_X1   g07413(.A1(new_n7414_), .A2(new_n7416_), .B(new_n7419_), .ZN(new_n7606_));
  NOR2_X1    g07414(.A1(new_n7561_), .A2(new_n7606_), .ZN(new_n7607_));
  XOR2_X1    g07415(.A1(new_n7607_), .A2(new_n7341_), .Z(new_n7608_));
  NAND3_X1   g07416(.A1(\asqrt[26] ), .A2(new_n7433_), .A3(new_n7415_), .ZN(new_n7609_));
  XOR2_X1    g07417(.A1(new_n7609_), .A2(new_n7345_), .Z(new_n7610_));
  OAI21_X1   g07418(.A1(new_n7428_), .A2(new_n7429_), .B(new_n7432_), .ZN(new_n7611_));
  NOR2_X1    g07419(.A1(new_n7561_), .A2(new_n7611_), .ZN(new_n7612_));
  XOR2_X1    g07420(.A1(new_n7612_), .A2(new_n7347_), .Z(new_n7613_));
  INV_X1     g07421(.I(new_n7613_), .ZN(new_n7614_));
  NAND3_X1   g07422(.A1(\asqrt[26] ), .A2(new_n7392_), .A3(new_n7411_), .ZN(new_n7615_));
  XOR2_X1    g07423(.A1(new_n7615_), .A2(new_n7426_), .Z(new_n7616_));
  INV_X1     g07424(.I(new_n7616_), .ZN(new_n7617_));
  OAI21_X1   g07425(.A1(new_n7386_), .A2(new_n7388_), .B(new_n7391_), .ZN(new_n7618_));
  NOR2_X1    g07426(.A1(new_n7561_), .A2(new_n7618_), .ZN(new_n7619_));
  XOR2_X1    g07427(.A1(new_n7619_), .A2(new_n7353_), .Z(new_n7620_));
  NAND3_X1   g07428(.A1(\asqrt[26] ), .A2(new_n7405_), .A3(new_n7387_), .ZN(new_n7621_));
  XOR2_X1    g07429(.A1(new_n7621_), .A2(new_n7357_), .Z(new_n7622_));
  OAI21_X1   g07430(.A1(new_n7400_), .A2(new_n7401_), .B(new_n7404_), .ZN(new_n7623_));
  NOR2_X1    g07431(.A1(new_n7561_), .A2(new_n7623_), .ZN(new_n7624_));
  XOR2_X1    g07432(.A1(new_n7624_), .A2(new_n7359_), .Z(new_n7625_));
  INV_X1     g07433(.I(new_n7625_), .ZN(new_n7626_));
  NAND3_X1   g07434(.A1(\asqrt[26] ), .A2(new_n7372_), .A3(new_n7383_), .ZN(new_n7627_));
  XOR2_X1    g07435(.A1(new_n7627_), .A2(new_n7398_), .Z(new_n7628_));
  INV_X1     g07436(.I(new_n7628_), .ZN(new_n7629_));
  OAI21_X1   g07437(.A1(new_n7367_), .A2(new_n7368_), .B(new_n7371_), .ZN(new_n7630_));
  NOR2_X1    g07438(.A1(new_n7561_), .A2(new_n7630_), .ZN(new_n7631_));
  XOR2_X1    g07439(.A1(new_n7631_), .A2(new_n7365_), .Z(new_n7632_));
  OAI21_X1   g07440(.A1(new_n7271_), .A2(new_n7273_), .B(new_n7276_), .ZN(new_n7633_));
  NOR2_X1    g07441(.A1(new_n7561_), .A2(new_n7633_), .ZN(new_n7634_));
  XOR2_X1    g07442(.A1(new_n7634_), .A2(new_n7183_), .Z(new_n7635_));
  INV_X1     g07443(.I(new_n7635_), .ZN(new_n7636_));
  NAND3_X1   g07444(.A1(\asqrt[26] ), .A2(new_n7286_), .A3(new_n7272_), .ZN(new_n7637_));
  XOR2_X1    g07445(.A1(new_n7637_), .A2(new_n7187_), .Z(new_n7638_));
  INV_X1     g07446(.I(new_n7638_), .ZN(new_n7639_));
  OAI21_X1   g07447(.A1(new_n7281_), .A2(new_n7282_), .B(new_n7285_), .ZN(new_n7640_));
  NOR2_X1    g07448(.A1(new_n7561_), .A2(new_n7640_), .ZN(new_n7641_));
  XOR2_X1    g07449(.A1(new_n7641_), .A2(new_n7189_), .Z(new_n7642_));
  NAND3_X1   g07450(.A1(\asqrt[26] ), .A2(new_n7249_), .A3(new_n7268_), .ZN(new_n7643_));
  XOR2_X1    g07451(.A1(new_n7643_), .A2(new_n7279_), .Z(new_n7644_));
  OAI21_X1   g07452(.A1(new_n7243_), .A2(new_n7245_), .B(new_n7248_), .ZN(new_n7645_));
  NOR2_X1    g07453(.A1(new_n7561_), .A2(new_n7645_), .ZN(new_n7646_));
  XOR2_X1    g07454(.A1(new_n7646_), .A2(new_n7196_), .Z(new_n7647_));
  INV_X1     g07455(.I(new_n7647_), .ZN(new_n7648_));
  NAND3_X1   g07456(.A1(\asqrt[26] ), .A2(new_n7262_), .A3(new_n7244_), .ZN(new_n7649_));
  XOR2_X1    g07457(.A1(new_n7649_), .A2(new_n7199_), .Z(new_n7650_));
  INV_X1     g07458(.I(new_n7650_), .ZN(new_n7651_));
  OAI21_X1   g07459(.A1(new_n7257_), .A2(new_n7258_), .B(new_n7261_), .ZN(new_n7652_));
  NOR2_X1    g07460(.A1(new_n7561_), .A2(new_n7652_), .ZN(new_n7653_));
  XOR2_X1    g07461(.A1(new_n7653_), .A2(new_n7202_), .Z(new_n7654_));
  NAND3_X1   g07462(.A1(\asqrt[26] ), .A2(new_n7222_), .A3(new_n7240_), .ZN(new_n7655_));
  XOR2_X1    g07463(.A1(new_n7655_), .A2(new_n7256_), .Z(new_n7656_));
  NOR2_X1    g07464(.A1(new_n7219_), .A2(\asqrt[29] ), .ZN(new_n7657_));
  NOR3_X1    g07465(.A1(new_n7561_), .A2(new_n7657_), .A3(new_n7239_), .ZN(new_n7658_));
  XOR2_X1    g07466(.A1(new_n7658_), .A2(new_n7210_), .Z(new_n7659_));
  INV_X1     g07467(.I(new_n7659_), .ZN(new_n7660_));
  NAND3_X1   g07468(.A1(\asqrt[26] ), .A2(new_n7211_), .A3(new_n7212_), .ZN(new_n7661_));
  NOR4_X1    g07469(.A1(new_n7559_), .A2(new_n7166_), .A3(new_n7296_), .A4(new_n7560_), .ZN(new_n7662_));
  INV_X1     g07470(.I(new_n7662_), .ZN(new_n7663_));
  AOI21_X1   g07471(.A1(new_n7661_), .A2(new_n7663_), .B(\a[54] ), .ZN(new_n7664_));
  NOR3_X1    g07472(.A1(new_n7561_), .A2(\a[52] ), .A3(\a[53] ), .ZN(new_n7665_));
  NOR3_X1    g07473(.A1(new_n7665_), .A2(new_n6914_), .A3(new_n7662_), .ZN(new_n7666_));
  NOR2_X1    g07474(.A1(new_n7666_), .A2(new_n7664_), .ZN(new_n7667_));
  INV_X1     g07475(.I(\a[50] ), .ZN(new_n7668_));
  INV_X1     g07476(.I(\a[51] ), .ZN(new_n7669_));
  NAND3_X1   g07477(.A1(new_n7668_), .A2(new_n7669_), .A3(new_n7211_), .ZN(new_n7670_));
  OAI21_X1   g07478(.A1(new_n7561_), .A2(new_n7211_), .B(new_n7670_), .ZN(new_n7671_));
  NAND2_X1   g07479(.A1(new_n7671_), .A2(\asqrt[27] ), .ZN(new_n7672_));
  OAI21_X1   g07480(.A1(new_n7561_), .A2(\a[52] ), .B(\a[53] ), .ZN(new_n7673_));
  NAND2_X1   g07481(.A1(new_n7673_), .A2(new_n7661_), .ZN(new_n7674_));
  NOR2_X1    g07482(.A1(new_n7671_), .A2(\asqrt[27] ), .ZN(new_n7675_));
  OAI21_X1   g07483(.A1(new_n7674_), .A2(new_n7675_), .B(new_n7672_), .ZN(new_n7676_));
  OAI21_X1   g07484(.A1(new_n7676_), .A2(\asqrt[28] ), .B(new_n7667_), .ZN(new_n7677_));
  NAND2_X1   g07485(.A1(new_n7676_), .A2(\asqrt[28] ), .ZN(new_n7678_));
  NAND3_X1   g07486(.A1(new_n7677_), .A2(new_n6454_), .A3(new_n7678_), .ZN(new_n7679_));
  NOR3_X1    g07487(.A1(new_n7561_), .A2(new_n7233_), .A3(new_n7218_), .ZN(new_n7680_));
  XOR2_X1    g07488(.A1(new_n7680_), .A2(new_n7235_), .Z(new_n7681_));
  AOI21_X1   g07489(.A1(new_n7677_), .A2(new_n7678_), .B(new_n6454_), .ZN(new_n7682_));
  AOI21_X1   g07490(.A1(new_n7679_), .A2(new_n7681_), .B(new_n7682_), .ZN(new_n7683_));
  AOI21_X1   g07491(.A1(new_n7683_), .A2(new_n6106_), .B(new_n7660_), .ZN(new_n7684_));
  OAI21_X1   g07492(.A1(new_n7683_), .A2(new_n6106_), .B(new_n5750_), .ZN(new_n7685_));
  OAI21_X1   g07493(.A1(new_n7684_), .A2(new_n7685_), .B(new_n7656_), .ZN(new_n7686_));
  NOR2_X1    g07494(.A1(new_n7683_), .A2(new_n6106_), .ZN(new_n7687_));
  OAI21_X1   g07495(.A1(new_n7684_), .A2(new_n7687_), .B(\asqrt[31] ), .ZN(new_n7688_));
  NAND3_X1   g07496(.A1(new_n7686_), .A2(new_n7688_), .A3(new_n5435_), .ZN(new_n7689_));
  NAND2_X1   g07497(.A1(new_n7689_), .A2(new_n7654_), .ZN(new_n7690_));
  NAND2_X1   g07498(.A1(new_n7686_), .A2(new_n7688_), .ZN(new_n7691_));
  AOI21_X1   g07499(.A1(new_n7691_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n7692_));
  AOI21_X1   g07500(.A1(new_n7692_), .A2(new_n7690_), .B(new_n7651_), .ZN(new_n7693_));
  INV_X1     g07501(.I(new_n7656_), .ZN(new_n7694_));
  OAI21_X1   g07502(.A1(new_n7665_), .A2(new_n7662_), .B(new_n6914_), .ZN(new_n7695_));
  NAND3_X1   g07503(.A1(new_n7661_), .A2(new_n7663_), .A3(\a[54] ), .ZN(new_n7696_));
  NAND2_X1   g07504(.A1(new_n7695_), .A2(new_n7696_), .ZN(new_n7697_));
  NAND2_X1   g07505(.A1(\asqrt[26] ), .A2(\a[52] ), .ZN(new_n7698_));
  AOI21_X1   g07506(.A1(new_n7698_), .A2(new_n7670_), .B(new_n7166_), .ZN(new_n7699_));
  AOI21_X1   g07507(.A1(\asqrt[26] ), .A2(new_n7211_), .B(new_n7212_), .ZN(new_n7700_));
  NOR2_X1    g07508(.A1(new_n7665_), .A2(new_n7700_), .ZN(new_n7701_));
  NAND3_X1   g07509(.A1(new_n7698_), .A2(new_n7166_), .A3(new_n7670_), .ZN(new_n7702_));
  AOI21_X1   g07510(.A1(new_n7701_), .A2(new_n7702_), .B(new_n7699_), .ZN(new_n7703_));
  AOI21_X1   g07511(.A1(new_n7703_), .A2(new_n6813_), .B(new_n7697_), .ZN(new_n7704_));
  NOR2_X1    g07512(.A1(new_n7703_), .A2(new_n6813_), .ZN(new_n7705_));
  NOR3_X1    g07513(.A1(new_n7704_), .A2(\asqrt[29] ), .A3(new_n7705_), .ZN(new_n7706_));
  INV_X1     g07514(.I(new_n7681_), .ZN(new_n7707_));
  OAI21_X1   g07515(.A1(new_n7704_), .A2(new_n7705_), .B(\asqrt[29] ), .ZN(new_n7708_));
  OAI21_X1   g07516(.A1(new_n7706_), .A2(new_n7707_), .B(new_n7708_), .ZN(new_n7709_));
  OAI21_X1   g07517(.A1(new_n7709_), .A2(\asqrt[30] ), .B(new_n7659_), .ZN(new_n7710_));
  AOI21_X1   g07518(.A1(new_n7709_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n7711_));
  AOI21_X1   g07519(.A1(new_n7711_), .A2(new_n7710_), .B(new_n7694_), .ZN(new_n7712_));
  NAND2_X1   g07520(.A1(new_n7709_), .A2(\asqrt[30] ), .ZN(new_n7713_));
  AOI21_X1   g07521(.A1(new_n7710_), .A2(new_n7713_), .B(new_n5750_), .ZN(new_n7714_));
  OAI21_X1   g07522(.A1(new_n7712_), .A2(new_n7714_), .B(\asqrt[32] ), .ZN(new_n7715_));
  AOI21_X1   g07523(.A1(new_n7690_), .A2(new_n7715_), .B(new_n5110_), .ZN(new_n7716_));
  NOR2_X1    g07524(.A1(new_n7693_), .A2(new_n7716_), .ZN(new_n7717_));
  AOI21_X1   g07525(.A1(new_n7717_), .A2(new_n4810_), .B(new_n7648_), .ZN(new_n7718_));
  OAI21_X1   g07526(.A1(new_n7693_), .A2(new_n7716_), .B(\asqrt[34] ), .ZN(new_n7719_));
  NAND2_X1   g07527(.A1(new_n7719_), .A2(new_n4510_), .ZN(new_n7720_));
  OAI21_X1   g07528(.A1(new_n7718_), .A2(new_n7720_), .B(new_n7644_), .ZN(new_n7721_));
  INV_X1     g07529(.I(new_n7719_), .ZN(new_n7722_));
  OAI21_X1   g07530(.A1(new_n7718_), .A2(new_n7722_), .B(\asqrt[35] ), .ZN(new_n7723_));
  NAND3_X1   g07531(.A1(new_n7721_), .A2(new_n7723_), .A3(new_n4224_), .ZN(new_n7724_));
  NAND2_X1   g07532(.A1(new_n7724_), .A2(new_n7642_), .ZN(new_n7725_));
  NAND2_X1   g07533(.A1(new_n7721_), .A2(new_n7723_), .ZN(new_n7726_));
  AOI21_X1   g07534(.A1(new_n7726_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n7727_));
  AOI21_X1   g07535(.A1(new_n7727_), .A2(new_n7725_), .B(new_n7639_), .ZN(new_n7728_));
  INV_X1     g07536(.I(new_n7644_), .ZN(new_n7729_));
  INV_X1     g07537(.I(new_n7654_), .ZN(new_n7730_));
  NOR2_X1    g07538(.A1(new_n7712_), .A2(new_n7714_), .ZN(new_n7731_));
  AOI21_X1   g07539(.A1(new_n7731_), .A2(new_n5435_), .B(new_n7730_), .ZN(new_n7732_));
  NAND2_X1   g07540(.A1(new_n7715_), .A2(new_n5110_), .ZN(new_n7733_));
  OAI21_X1   g07541(.A1(new_n7732_), .A2(new_n7733_), .B(new_n7650_), .ZN(new_n7734_));
  INV_X1     g07542(.I(new_n7715_), .ZN(new_n7735_));
  OAI21_X1   g07543(.A1(new_n7732_), .A2(new_n7735_), .B(\asqrt[33] ), .ZN(new_n7736_));
  NAND3_X1   g07544(.A1(new_n7734_), .A2(new_n7736_), .A3(new_n4810_), .ZN(new_n7737_));
  NAND2_X1   g07545(.A1(new_n7737_), .A2(new_n7647_), .ZN(new_n7738_));
  NAND2_X1   g07546(.A1(new_n7734_), .A2(new_n7736_), .ZN(new_n7739_));
  AOI21_X1   g07547(.A1(new_n7739_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n7740_));
  AOI21_X1   g07548(.A1(new_n7740_), .A2(new_n7738_), .B(new_n7729_), .ZN(new_n7741_));
  AOI21_X1   g07549(.A1(new_n7738_), .A2(new_n7719_), .B(new_n4510_), .ZN(new_n7742_));
  OAI21_X1   g07550(.A1(new_n7741_), .A2(new_n7742_), .B(\asqrt[36] ), .ZN(new_n7743_));
  AOI21_X1   g07551(.A1(new_n7725_), .A2(new_n7743_), .B(new_n3928_), .ZN(new_n7744_));
  NOR2_X1    g07552(.A1(new_n7728_), .A2(new_n7744_), .ZN(new_n7745_));
  AOI21_X1   g07553(.A1(new_n7745_), .A2(new_n3675_), .B(new_n7636_), .ZN(new_n7746_));
  OAI21_X1   g07554(.A1(new_n7728_), .A2(new_n7744_), .B(\asqrt[38] ), .ZN(new_n7747_));
  NAND2_X1   g07555(.A1(new_n7747_), .A2(new_n3400_), .ZN(new_n7748_));
  OAI21_X1   g07556(.A1(new_n7746_), .A2(new_n7748_), .B(new_n7544_), .ZN(new_n7749_));
  INV_X1     g07557(.I(new_n7747_), .ZN(new_n7750_));
  OAI21_X1   g07558(.A1(new_n7746_), .A2(new_n7750_), .B(\asqrt[39] ), .ZN(new_n7751_));
  NAND3_X1   g07559(.A1(new_n7749_), .A2(new_n7751_), .A3(new_n3167_), .ZN(new_n7752_));
  NAND2_X1   g07560(.A1(new_n7752_), .A2(new_n7632_), .ZN(new_n7753_));
  NAND2_X1   g07561(.A1(new_n7749_), .A2(new_n7751_), .ZN(new_n7754_));
  AOI21_X1   g07562(.A1(new_n7754_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n7755_));
  AOI21_X1   g07563(.A1(new_n7755_), .A2(new_n7753_), .B(new_n7629_), .ZN(new_n7756_));
  INV_X1     g07564(.I(new_n7544_), .ZN(new_n7757_));
  INV_X1     g07565(.I(new_n7642_), .ZN(new_n7758_));
  NOR2_X1    g07566(.A1(new_n7741_), .A2(new_n7742_), .ZN(new_n7759_));
  AOI21_X1   g07567(.A1(new_n7759_), .A2(new_n4224_), .B(new_n7758_), .ZN(new_n7760_));
  NAND2_X1   g07568(.A1(new_n7743_), .A2(new_n3928_), .ZN(new_n7761_));
  OAI21_X1   g07569(.A1(new_n7760_), .A2(new_n7761_), .B(new_n7638_), .ZN(new_n7762_));
  INV_X1     g07570(.I(new_n7743_), .ZN(new_n7763_));
  OAI21_X1   g07571(.A1(new_n7760_), .A2(new_n7763_), .B(\asqrt[37] ), .ZN(new_n7764_));
  NAND3_X1   g07572(.A1(new_n7762_), .A2(new_n7764_), .A3(new_n3675_), .ZN(new_n7765_));
  NAND2_X1   g07573(.A1(new_n7765_), .A2(new_n7635_), .ZN(new_n7766_));
  NAND2_X1   g07574(.A1(new_n7762_), .A2(new_n7764_), .ZN(new_n7767_));
  AOI21_X1   g07575(.A1(new_n7767_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n7768_));
  AOI21_X1   g07576(.A1(new_n7768_), .A2(new_n7766_), .B(new_n7757_), .ZN(new_n7769_));
  AOI21_X1   g07577(.A1(new_n7766_), .A2(new_n7747_), .B(new_n3400_), .ZN(new_n7770_));
  OAI21_X1   g07578(.A1(new_n7769_), .A2(new_n7770_), .B(\asqrt[40] ), .ZN(new_n7771_));
  AOI21_X1   g07579(.A1(new_n7753_), .A2(new_n7771_), .B(new_n2912_), .ZN(new_n7772_));
  NOR2_X1    g07580(.A1(new_n7756_), .A2(new_n7772_), .ZN(new_n7773_));
  AOI21_X1   g07581(.A1(new_n7773_), .A2(new_n2699_), .B(new_n7626_), .ZN(new_n7774_));
  OAI21_X1   g07582(.A1(new_n7756_), .A2(new_n7772_), .B(\asqrt[42] ), .ZN(new_n7775_));
  NAND2_X1   g07583(.A1(new_n7775_), .A2(new_n2464_), .ZN(new_n7776_));
  OAI21_X1   g07584(.A1(new_n7774_), .A2(new_n7776_), .B(new_n7622_), .ZN(new_n7777_));
  INV_X1     g07585(.I(new_n7775_), .ZN(new_n7778_));
  OAI21_X1   g07586(.A1(new_n7774_), .A2(new_n7778_), .B(\asqrt[43] ), .ZN(new_n7779_));
  NAND3_X1   g07587(.A1(new_n7777_), .A2(new_n7779_), .A3(new_n2271_), .ZN(new_n7780_));
  NAND2_X1   g07588(.A1(new_n7780_), .A2(new_n7620_), .ZN(new_n7781_));
  NAND2_X1   g07589(.A1(new_n7777_), .A2(new_n7779_), .ZN(new_n7782_));
  AOI21_X1   g07590(.A1(new_n7782_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n7783_));
  AOI21_X1   g07591(.A1(new_n7783_), .A2(new_n7781_), .B(new_n7617_), .ZN(new_n7784_));
  INV_X1     g07592(.I(new_n7622_), .ZN(new_n7785_));
  INV_X1     g07593(.I(new_n7632_), .ZN(new_n7786_));
  NOR2_X1    g07594(.A1(new_n7769_), .A2(new_n7770_), .ZN(new_n7787_));
  AOI21_X1   g07595(.A1(new_n7787_), .A2(new_n3167_), .B(new_n7786_), .ZN(new_n7788_));
  NAND2_X1   g07596(.A1(new_n7771_), .A2(new_n2912_), .ZN(new_n7789_));
  OAI21_X1   g07597(.A1(new_n7788_), .A2(new_n7789_), .B(new_n7628_), .ZN(new_n7790_));
  INV_X1     g07598(.I(new_n7771_), .ZN(new_n7791_));
  OAI21_X1   g07599(.A1(new_n7788_), .A2(new_n7791_), .B(\asqrt[41] ), .ZN(new_n7792_));
  NAND3_X1   g07600(.A1(new_n7790_), .A2(new_n7792_), .A3(new_n2699_), .ZN(new_n7793_));
  NAND2_X1   g07601(.A1(new_n7793_), .A2(new_n7625_), .ZN(new_n7794_));
  NAND2_X1   g07602(.A1(new_n7790_), .A2(new_n7792_), .ZN(new_n7795_));
  AOI21_X1   g07603(.A1(new_n7795_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n7796_));
  AOI21_X1   g07604(.A1(new_n7796_), .A2(new_n7794_), .B(new_n7785_), .ZN(new_n7797_));
  AOI21_X1   g07605(.A1(new_n7794_), .A2(new_n7775_), .B(new_n2464_), .ZN(new_n7798_));
  OAI21_X1   g07606(.A1(new_n7797_), .A2(new_n7798_), .B(\asqrt[44] ), .ZN(new_n7799_));
  AOI21_X1   g07607(.A1(new_n7781_), .A2(new_n7799_), .B(new_n2072_), .ZN(new_n7800_));
  NOR2_X1    g07608(.A1(new_n7784_), .A2(new_n7800_), .ZN(new_n7801_));
  AOI21_X1   g07609(.A1(new_n7801_), .A2(new_n1884_), .B(new_n7614_), .ZN(new_n7802_));
  OAI21_X1   g07610(.A1(new_n7784_), .A2(new_n7800_), .B(\asqrt[46] ), .ZN(new_n7803_));
  NAND2_X1   g07611(.A1(new_n7803_), .A2(new_n1688_), .ZN(new_n7804_));
  OAI21_X1   g07612(.A1(new_n7802_), .A2(new_n7804_), .B(new_n7610_), .ZN(new_n7805_));
  INV_X1     g07613(.I(new_n7803_), .ZN(new_n7806_));
  OAI21_X1   g07614(.A1(new_n7802_), .A2(new_n7806_), .B(\asqrt[47] ), .ZN(new_n7807_));
  NAND3_X1   g07615(.A1(new_n7805_), .A2(new_n7807_), .A3(new_n1533_), .ZN(new_n7808_));
  NAND2_X1   g07616(.A1(new_n7808_), .A2(new_n7608_), .ZN(new_n7809_));
  NAND2_X1   g07617(.A1(new_n7805_), .A2(new_n7807_), .ZN(new_n7810_));
  AOI21_X1   g07618(.A1(new_n7810_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n7811_));
  AOI21_X1   g07619(.A1(new_n7811_), .A2(new_n7809_), .B(new_n7605_), .ZN(new_n7812_));
  INV_X1     g07620(.I(new_n7610_), .ZN(new_n7813_));
  INV_X1     g07621(.I(new_n7620_), .ZN(new_n7814_));
  NOR2_X1    g07622(.A1(new_n7797_), .A2(new_n7798_), .ZN(new_n7815_));
  AOI21_X1   g07623(.A1(new_n7815_), .A2(new_n2271_), .B(new_n7814_), .ZN(new_n7816_));
  NAND2_X1   g07624(.A1(new_n7799_), .A2(new_n2072_), .ZN(new_n7817_));
  OAI21_X1   g07625(.A1(new_n7816_), .A2(new_n7817_), .B(new_n7616_), .ZN(new_n7818_));
  INV_X1     g07626(.I(new_n7799_), .ZN(new_n7819_));
  OAI21_X1   g07627(.A1(new_n7816_), .A2(new_n7819_), .B(\asqrt[45] ), .ZN(new_n7820_));
  NAND3_X1   g07628(.A1(new_n7818_), .A2(new_n7820_), .A3(new_n1884_), .ZN(new_n7821_));
  NAND2_X1   g07629(.A1(new_n7821_), .A2(new_n7613_), .ZN(new_n7822_));
  NAND2_X1   g07630(.A1(new_n7818_), .A2(new_n7820_), .ZN(new_n7823_));
  AOI21_X1   g07631(.A1(new_n7823_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n7824_));
  AOI21_X1   g07632(.A1(new_n7824_), .A2(new_n7822_), .B(new_n7813_), .ZN(new_n7825_));
  AOI21_X1   g07633(.A1(new_n7822_), .A2(new_n7803_), .B(new_n1688_), .ZN(new_n7826_));
  OAI21_X1   g07634(.A1(new_n7825_), .A2(new_n7826_), .B(\asqrt[48] ), .ZN(new_n7827_));
  AOI21_X1   g07635(.A1(new_n7809_), .A2(new_n7827_), .B(new_n1368_), .ZN(new_n7828_));
  NOR2_X1    g07636(.A1(new_n7812_), .A2(new_n7828_), .ZN(new_n7829_));
  AOI21_X1   g07637(.A1(new_n7829_), .A2(new_n1228_), .B(new_n7602_), .ZN(new_n7830_));
  OAI21_X1   g07638(.A1(new_n7812_), .A2(new_n7828_), .B(\asqrt[50] ), .ZN(new_n7831_));
  NAND2_X1   g07639(.A1(new_n7831_), .A2(new_n1088_), .ZN(new_n7832_));
  OAI21_X1   g07640(.A1(new_n7830_), .A2(new_n7832_), .B(new_n7598_), .ZN(new_n7833_));
  INV_X1     g07641(.I(new_n7831_), .ZN(new_n7834_));
  OAI21_X1   g07642(.A1(new_n7830_), .A2(new_n7834_), .B(\asqrt[51] ), .ZN(new_n7835_));
  NAND3_X1   g07643(.A1(new_n7833_), .A2(new_n7835_), .A3(new_n962_), .ZN(new_n7836_));
  NAND2_X1   g07644(.A1(new_n7836_), .A2(new_n7596_), .ZN(new_n7837_));
  NAND2_X1   g07645(.A1(new_n7833_), .A2(new_n7835_), .ZN(new_n7838_));
  AOI21_X1   g07646(.A1(new_n7838_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n7839_));
  AOI21_X1   g07647(.A1(new_n7839_), .A2(new_n7837_), .B(new_n7593_), .ZN(new_n7840_));
  INV_X1     g07648(.I(new_n7598_), .ZN(new_n7841_));
  INV_X1     g07649(.I(new_n7608_), .ZN(new_n7842_));
  NOR2_X1    g07650(.A1(new_n7825_), .A2(new_n7826_), .ZN(new_n7843_));
  AOI21_X1   g07651(.A1(new_n7843_), .A2(new_n1533_), .B(new_n7842_), .ZN(new_n7844_));
  NAND2_X1   g07652(.A1(new_n7827_), .A2(new_n1368_), .ZN(new_n7845_));
  OAI21_X1   g07653(.A1(new_n7844_), .A2(new_n7845_), .B(new_n7604_), .ZN(new_n7846_));
  INV_X1     g07654(.I(new_n7827_), .ZN(new_n7847_));
  OAI21_X1   g07655(.A1(new_n7844_), .A2(new_n7847_), .B(\asqrt[49] ), .ZN(new_n7848_));
  NAND3_X1   g07656(.A1(new_n7846_), .A2(new_n7848_), .A3(new_n1228_), .ZN(new_n7849_));
  NAND2_X1   g07657(.A1(new_n7849_), .A2(new_n7601_), .ZN(new_n7850_));
  NAND2_X1   g07658(.A1(new_n7846_), .A2(new_n7848_), .ZN(new_n7851_));
  AOI21_X1   g07659(.A1(new_n7851_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n7852_));
  AOI21_X1   g07660(.A1(new_n7852_), .A2(new_n7850_), .B(new_n7841_), .ZN(new_n7853_));
  AOI21_X1   g07661(.A1(new_n7850_), .A2(new_n7831_), .B(new_n1088_), .ZN(new_n7854_));
  OAI21_X1   g07662(.A1(new_n7853_), .A2(new_n7854_), .B(\asqrt[52] ), .ZN(new_n7855_));
  AOI21_X1   g07663(.A1(new_n7837_), .A2(new_n7855_), .B(new_n842_), .ZN(new_n7856_));
  NOR2_X1    g07664(.A1(new_n7840_), .A2(new_n7856_), .ZN(new_n7857_));
  AOI21_X1   g07665(.A1(new_n7857_), .A2(new_n720_), .B(new_n7590_), .ZN(new_n7858_));
  OAI21_X1   g07666(.A1(new_n7840_), .A2(new_n7856_), .B(\asqrt[54] ), .ZN(new_n7859_));
  NAND2_X1   g07667(.A1(new_n7859_), .A2(new_n630_), .ZN(new_n7860_));
  OAI21_X1   g07668(.A1(new_n7858_), .A2(new_n7860_), .B(new_n7586_), .ZN(new_n7861_));
  INV_X1     g07669(.I(new_n7859_), .ZN(new_n7862_));
  OAI21_X1   g07670(.A1(new_n7858_), .A2(new_n7862_), .B(\asqrt[55] ), .ZN(new_n7863_));
  NAND3_X1   g07671(.A1(new_n7861_), .A2(new_n7863_), .A3(new_n545_), .ZN(new_n7864_));
  NAND2_X1   g07672(.A1(new_n7864_), .A2(new_n7584_), .ZN(new_n7865_));
  NAND2_X1   g07673(.A1(new_n7861_), .A2(new_n7863_), .ZN(new_n7866_));
  AOI21_X1   g07674(.A1(new_n7866_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n7867_));
  AOI21_X1   g07675(.A1(new_n7867_), .A2(new_n7865_), .B(new_n7581_), .ZN(new_n7868_));
  INV_X1     g07676(.I(new_n7586_), .ZN(new_n7869_));
  INV_X1     g07677(.I(new_n7596_), .ZN(new_n7870_));
  NOR2_X1    g07678(.A1(new_n7853_), .A2(new_n7854_), .ZN(new_n7871_));
  AOI21_X1   g07679(.A1(new_n7871_), .A2(new_n962_), .B(new_n7870_), .ZN(new_n7872_));
  NAND2_X1   g07680(.A1(new_n7855_), .A2(new_n842_), .ZN(new_n7873_));
  OAI21_X1   g07681(.A1(new_n7872_), .A2(new_n7873_), .B(new_n7592_), .ZN(new_n7874_));
  INV_X1     g07682(.I(new_n7855_), .ZN(new_n7875_));
  OAI21_X1   g07683(.A1(new_n7872_), .A2(new_n7875_), .B(\asqrt[53] ), .ZN(new_n7876_));
  NAND3_X1   g07684(.A1(new_n7874_), .A2(new_n7876_), .A3(new_n720_), .ZN(new_n7877_));
  NAND2_X1   g07685(.A1(new_n7877_), .A2(new_n7589_), .ZN(new_n7878_));
  NAND2_X1   g07686(.A1(new_n7874_), .A2(new_n7876_), .ZN(new_n7879_));
  AOI21_X1   g07687(.A1(new_n7879_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n7880_));
  AOI21_X1   g07688(.A1(new_n7880_), .A2(new_n7878_), .B(new_n7869_), .ZN(new_n7881_));
  AOI21_X1   g07689(.A1(new_n7878_), .A2(new_n7859_), .B(new_n630_), .ZN(new_n7882_));
  OAI21_X1   g07690(.A1(new_n7881_), .A2(new_n7882_), .B(\asqrt[56] ), .ZN(new_n7883_));
  AOI21_X1   g07691(.A1(new_n7865_), .A2(new_n7883_), .B(new_n450_), .ZN(new_n7884_));
  NOR2_X1    g07692(.A1(new_n7868_), .A2(new_n7884_), .ZN(new_n7885_));
  AOI21_X1   g07693(.A1(new_n7885_), .A2(new_n403_), .B(new_n7578_), .ZN(new_n7886_));
  OAI21_X1   g07694(.A1(new_n7868_), .A2(new_n7884_), .B(\asqrt[58] ), .ZN(new_n7887_));
  NAND2_X1   g07695(.A1(new_n7887_), .A2(new_n339_), .ZN(new_n7888_));
  OAI21_X1   g07696(.A1(new_n7886_), .A2(new_n7888_), .B(new_n7574_), .ZN(new_n7889_));
  INV_X1     g07697(.I(new_n7887_), .ZN(new_n7890_));
  OAI21_X1   g07698(.A1(new_n7886_), .A2(new_n7890_), .B(\asqrt[59] ), .ZN(new_n7891_));
  NAND3_X1   g07699(.A1(new_n7889_), .A2(new_n7891_), .A3(new_n288_), .ZN(new_n7892_));
  NAND2_X1   g07700(.A1(new_n7892_), .A2(new_n7572_), .ZN(new_n7893_));
  INV_X1     g07701(.I(new_n7574_), .ZN(new_n7894_));
  INV_X1     g07702(.I(new_n7584_), .ZN(new_n7895_));
  NOR2_X1    g07703(.A1(new_n7881_), .A2(new_n7882_), .ZN(new_n7896_));
  AOI21_X1   g07704(.A1(new_n7896_), .A2(new_n545_), .B(new_n7895_), .ZN(new_n7897_));
  NAND2_X1   g07705(.A1(new_n7883_), .A2(new_n450_), .ZN(new_n7898_));
  OAI21_X1   g07706(.A1(new_n7897_), .A2(new_n7898_), .B(new_n7580_), .ZN(new_n7899_));
  INV_X1     g07707(.I(new_n7883_), .ZN(new_n7900_));
  OAI21_X1   g07708(.A1(new_n7897_), .A2(new_n7900_), .B(\asqrt[57] ), .ZN(new_n7901_));
  NAND3_X1   g07709(.A1(new_n7899_), .A2(new_n7901_), .A3(new_n403_), .ZN(new_n7902_));
  NAND2_X1   g07710(.A1(new_n7902_), .A2(new_n7577_), .ZN(new_n7903_));
  NAND2_X1   g07711(.A1(new_n7899_), .A2(new_n7901_), .ZN(new_n7904_));
  AOI21_X1   g07712(.A1(new_n7904_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n7905_));
  AOI21_X1   g07713(.A1(new_n7905_), .A2(new_n7903_), .B(new_n7894_), .ZN(new_n7906_));
  AOI21_X1   g07714(.A1(new_n7903_), .A2(new_n7887_), .B(new_n339_), .ZN(new_n7907_));
  OAI21_X1   g07715(.A1(new_n7906_), .A2(new_n7907_), .B(\asqrt[60] ), .ZN(new_n7908_));
  AOI21_X1   g07716(.A1(new_n7893_), .A2(new_n7908_), .B(new_n242_), .ZN(new_n7909_));
  NAND3_X1   g07717(.A1(\asqrt[26] ), .A2(new_n7504_), .A3(new_n7520_), .ZN(new_n7910_));
  XOR2_X1    g07718(.A1(new_n7910_), .A2(new_n7545_), .Z(new_n7911_));
  INV_X1     g07719(.I(new_n7911_), .ZN(new_n7912_));
  NAND2_X1   g07720(.A1(new_n7889_), .A2(new_n7891_), .ZN(new_n7913_));
  AOI21_X1   g07721(.A1(new_n7913_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n7914_));
  AOI21_X1   g07722(.A1(new_n7914_), .A2(new_n7893_), .B(new_n7912_), .ZN(new_n7915_));
  OAI21_X1   g07723(.A1(new_n7915_), .A2(new_n7909_), .B(\asqrt[62] ), .ZN(new_n7916_));
  AOI21_X1   g07724(.A1(new_n7505_), .A2(new_n7526_), .B(new_n7521_), .ZN(new_n7917_));
  NAND2_X1   g07725(.A1(\asqrt[26] ), .A2(new_n7917_), .ZN(new_n7918_));
  XOR2_X1    g07726(.A1(new_n7918_), .A2(new_n7524_), .Z(new_n7919_));
  INV_X1     g07727(.I(new_n7572_), .ZN(new_n7920_));
  NOR2_X1    g07728(.A1(new_n7906_), .A2(new_n7907_), .ZN(new_n7921_));
  AOI21_X1   g07729(.A1(new_n7921_), .A2(new_n288_), .B(new_n7920_), .ZN(new_n7922_));
  INV_X1     g07730(.I(new_n7908_), .ZN(new_n7923_));
  OAI21_X1   g07731(.A1(new_n7922_), .A2(new_n7923_), .B(\asqrt[61] ), .ZN(new_n7924_));
  NAND2_X1   g07732(.A1(new_n7908_), .A2(new_n242_), .ZN(new_n7925_));
  OAI21_X1   g07733(.A1(new_n7922_), .A2(new_n7925_), .B(new_n7911_), .ZN(new_n7926_));
  NAND3_X1   g07734(.A1(new_n7926_), .A2(new_n7924_), .A3(new_n234_), .ZN(new_n7927_));
  NAND2_X1   g07735(.A1(new_n7927_), .A2(new_n7919_), .ZN(new_n7928_));
  AOI21_X1   g07736(.A1(new_n7928_), .A2(new_n7916_), .B(new_n7569_), .ZN(new_n7929_));
  AOI21_X1   g07737(.A1(new_n7929_), .A2(new_n7567_), .B(\asqrt[63] ), .ZN(new_n7930_));
  NAND2_X1   g07738(.A1(new_n7928_), .A2(new_n7916_), .ZN(new_n7931_));
  NOR2_X1    g07739(.A1(new_n7931_), .A2(new_n7567_), .ZN(new_n7932_));
  NOR2_X1    g07740(.A1(\asqrt[26] ), .A2(new_n7556_), .ZN(new_n7933_));
  NOR4_X1    g07741(.A1(new_n7930_), .A2(new_n7564_), .A3(new_n7932_), .A4(new_n7933_), .ZN(new_n7934_));
  OAI21_X1   g07742(.A1(new_n7746_), .A2(new_n7748_), .B(new_n7751_), .ZN(new_n7935_));
  NOR2_X1    g07743(.A1(new_n7934_), .A2(new_n7935_), .ZN(new_n7936_));
  XOR2_X1    g07744(.A1(new_n7936_), .A2(new_n7544_), .Z(new_n7937_));
  INV_X1     g07745(.I(new_n7937_), .ZN(new_n7938_));
  INV_X1     g07746(.I(new_n7564_), .ZN(new_n7939_));
  INV_X1     g07747(.I(new_n7916_), .ZN(new_n7940_));
  NOR2_X1    g07748(.A1(new_n7915_), .A2(new_n7909_), .ZN(new_n7941_));
  INV_X1     g07749(.I(new_n7919_), .ZN(new_n7942_));
  AOI21_X1   g07750(.A1(new_n7941_), .A2(new_n234_), .B(new_n7942_), .ZN(new_n7943_));
  OAI21_X1   g07751(.A1(new_n7943_), .A2(new_n7940_), .B(new_n7568_), .ZN(new_n7944_));
  OAI21_X1   g07752(.A1(new_n7944_), .A2(new_n7566_), .B(new_n193_), .ZN(new_n7945_));
  NOR2_X1    g07753(.A1(new_n7943_), .A2(new_n7940_), .ZN(new_n7946_));
  NAND2_X1   g07754(.A1(new_n7946_), .A2(new_n7566_), .ZN(new_n7947_));
  INV_X1     g07755(.I(new_n7933_), .ZN(new_n7948_));
  NAND4_X1   g07756(.A1(new_n7945_), .A2(new_n7939_), .A3(new_n7947_), .A4(new_n7948_), .ZN(\asqrt[25] ));
  NAND3_X1   g07757(.A1(\asqrt[25] ), .A2(new_n7765_), .A3(new_n7747_), .ZN(new_n7950_));
  XOR2_X1    g07758(.A1(new_n7950_), .A2(new_n7636_), .Z(new_n7951_));
  OAI21_X1   g07759(.A1(new_n7760_), .A2(new_n7761_), .B(new_n7764_), .ZN(new_n7952_));
  NOR2_X1    g07760(.A1(new_n7934_), .A2(new_n7952_), .ZN(new_n7953_));
  XOR2_X1    g07761(.A1(new_n7953_), .A2(new_n7638_), .Z(new_n7954_));
  INV_X1     g07762(.I(new_n7954_), .ZN(new_n7955_));
  NAND3_X1   g07763(.A1(\asqrt[25] ), .A2(new_n7724_), .A3(new_n7743_), .ZN(new_n7956_));
  XOR2_X1    g07764(.A1(new_n7956_), .A2(new_n7758_), .Z(new_n7957_));
  INV_X1     g07765(.I(new_n7957_), .ZN(new_n7958_));
  OAI21_X1   g07766(.A1(new_n7718_), .A2(new_n7720_), .B(new_n7723_), .ZN(new_n7959_));
  NOR2_X1    g07767(.A1(new_n7934_), .A2(new_n7959_), .ZN(new_n7960_));
  XOR2_X1    g07768(.A1(new_n7960_), .A2(new_n7644_), .Z(new_n7961_));
  NAND3_X1   g07769(.A1(\asqrt[25] ), .A2(new_n7737_), .A3(new_n7719_), .ZN(new_n7962_));
  XOR2_X1    g07770(.A1(new_n7962_), .A2(new_n7648_), .Z(new_n7963_));
  OAI21_X1   g07771(.A1(new_n7732_), .A2(new_n7733_), .B(new_n7736_), .ZN(new_n7964_));
  NOR2_X1    g07772(.A1(new_n7934_), .A2(new_n7964_), .ZN(new_n7965_));
  XOR2_X1    g07773(.A1(new_n7965_), .A2(new_n7650_), .Z(new_n7966_));
  INV_X1     g07774(.I(new_n7966_), .ZN(new_n7967_));
  NAND3_X1   g07775(.A1(\asqrt[25] ), .A2(new_n7689_), .A3(new_n7715_), .ZN(new_n7968_));
  XOR2_X1    g07776(.A1(new_n7968_), .A2(new_n7730_), .Z(new_n7969_));
  INV_X1     g07777(.I(new_n7969_), .ZN(new_n7970_));
  AOI21_X1   g07778(.A1(new_n7710_), .A2(new_n7711_), .B(new_n7714_), .ZN(new_n7971_));
  NAND2_X1   g07779(.A1(\asqrt[25] ), .A2(new_n7971_), .ZN(new_n7972_));
  XOR2_X1    g07780(.A1(new_n7972_), .A2(new_n7694_), .Z(new_n7973_));
  NOR2_X1    g07781(.A1(new_n7709_), .A2(\asqrt[30] ), .ZN(new_n7974_));
  NOR3_X1    g07782(.A1(new_n7934_), .A2(new_n7974_), .A3(new_n7687_), .ZN(new_n7975_));
  XOR2_X1    g07783(.A1(new_n7975_), .A2(new_n7659_), .Z(new_n7976_));
  NOR3_X1    g07784(.A1(new_n7934_), .A2(new_n7706_), .A3(new_n7682_), .ZN(new_n7977_));
  XOR2_X1    g07785(.A1(new_n7977_), .A2(new_n7681_), .Z(new_n7978_));
  INV_X1     g07786(.I(new_n7978_), .ZN(new_n7979_));
  NOR2_X1    g07787(.A1(new_n7676_), .A2(\asqrt[28] ), .ZN(new_n7980_));
  NOR3_X1    g07788(.A1(new_n7934_), .A2(new_n7980_), .A3(new_n7705_), .ZN(new_n7981_));
  XOR2_X1    g07789(.A1(new_n7981_), .A2(new_n7667_), .Z(new_n7982_));
  INV_X1     g07790(.I(new_n7982_), .ZN(new_n7983_));
  NAND3_X1   g07791(.A1(\asqrt[25] ), .A2(new_n7668_), .A3(new_n7669_), .ZN(new_n7984_));
  NOR4_X1    g07792(.A1(new_n7930_), .A2(new_n7561_), .A3(new_n7564_), .A4(new_n7932_), .ZN(new_n7985_));
  INV_X1     g07793(.I(new_n7985_), .ZN(new_n7986_));
  AOI21_X1   g07794(.A1(new_n7984_), .A2(new_n7986_), .B(\a[52] ), .ZN(new_n7987_));
  NOR3_X1    g07795(.A1(new_n7934_), .A2(\a[50] ), .A3(\a[51] ), .ZN(new_n7988_));
  NOR3_X1    g07796(.A1(new_n7988_), .A2(new_n7211_), .A3(new_n7985_), .ZN(new_n7989_));
  NOR2_X1    g07797(.A1(new_n7989_), .A2(new_n7987_), .ZN(new_n7990_));
  INV_X1     g07798(.I(\a[48] ), .ZN(new_n7991_));
  INV_X1     g07799(.I(\a[49] ), .ZN(new_n7992_));
  NAND3_X1   g07800(.A1(new_n7991_), .A2(new_n7992_), .A3(new_n7668_), .ZN(new_n7993_));
  OAI21_X1   g07801(.A1(new_n7934_), .A2(new_n7668_), .B(new_n7993_), .ZN(new_n7994_));
  NAND2_X1   g07802(.A1(new_n7994_), .A2(\asqrt[26] ), .ZN(new_n7995_));
  OAI21_X1   g07803(.A1(new_n7934_), .A2(\a[50] ), .B(\a[51] ), .ZN(new_n7996_));
  NAND2_X1   g07804(.A1(new_n7996_), .A2(new_n7984_), .ZN(new_n7997_));
  NOR2_X1    g07805(.A1(new_n7994_), .A2(\asqrt[26] ), .ZN(new_n7998_));
  OAI21_X1   g07806(.A1(new_n7997_), .A2(new_n7998_), .B(new_n7995_), .ZN(new_n7999_));
  OAI21_X1   g07807(.A1(\asqrt[27] ), .A2(new_n7999_), .B(new_n7990_), .ZN(new_n8000_));
  NAND2_X1   g07808(.A1(new_n7999_), .A2(\asqrt[27] ), .ZN(new_n8001_));
  NAND3_X1   g07809(.A1(new_n8000_), .A2(new_n6813_), .A3(new_n8001_), .ZN(new_n8002_));
  NOR3_X1    g07810(.A1(new_n7934_), .A2(new_n7699_), .A3(new_n7675_), .ZN(new_n8003_));
  XOR2_X1    g07811(.A1(new_n8003_), .A2(new_n7701_), .Z(new_n8004_));
  NAND2_X1   g07812(.A1(new_n8002_), .A2(new_n8004_), .ZN(new_n8005_));
  NAND2_X1   g07813(.A1(new_n8000_), .A2(new_n8001_), .ZN(new_n8006_));
  AOI21_X1   g07814(.A1(new_n8006_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n8007_));
  AOI21_X1   g07815(.A1(new_n8007_), .A2(new_n8005_), .B(new_n7983_), .ZN(new_n8008_));
  OAI21_X1   g07816(.A1(new_n7988_), .A2(new_n7985_), .B(new_n7211_), .ZN(new_n8009_));
  NAND3_X1   g07817(.A1(new_n7984_), .A2(\a[52] ), .A3(new_n7986_), .ZN(new_n8010_));
  NAND2_X1   g07818(.A1(new_n8009_), .A2(new_n8010_), .ZN(new_n8011_));
  NAND2_X1   g07819(.A1(\asqrt[25] ), .A2(\a[50] ), .ZN(new_n8012_));
  AOI21_X1   g07820(.A1(new_n8012_), .A2(new_n7993_), .B(new_n7561_), .ZN(new_n8013_));
  AOI21_X1   g07821(.A1(\asqrt[25] ), .A2(new_n7668_), .B(new_n7669_), .ZN(new_n8014_));
  NOR2_X1    g07822(.A1(new_n8014_), .A2(new_n7988_), .ZN(new_n8015_));
  NAND3_X1   g07823(.A1(new_n8012_), .A2(new_n7561_), .A3(new_n7993_), .ZN(new_n8016_));
  AOI21_X1   g07824(.A1(new_n8015_), .A2(new_n8016_), .B(new_n8013_), .ZN(new_n8017_));
  AOI21_X1   g07825(.A1(new_n8017_), .A2(new_n7166_), .B(new_n8011_), .ZN(new_n8018_));
  NOR2_X1    g07826(.A1(new_n8017_), .A2(new_n7166_), .ZN(new_n8019_));
  OAI21_X1   g07827(.A1(new_n8018_), .A2(new_n8019_), .B(\asqrt[28] ), .ZN(new_n8020_));
  AOI21_X1   g07828(.A1(new_n8005_), .A2(new_n8020_), .B(new_n6454_), .ZN(new_n8021_));
  NOR2_X1    g07829(.A1(new_n8008_), .A2(new_n8021_), .ZN(new_n8022_));
  AOI21_X1   g07830(.A1(new_n8022_), .A2(new_n6106_), .B(new_n7979_), .ZN(new_n8023_));
  OAI21_X1   g07831(.A1(new_n8008_), .A2(new_n8021_), .B(\asqrt[30] ), .ZN(new_n8024_));
  NAND2_X1   g07832(.A1(new_n8024_), .A2(new_n5750_), .ZN(new_n8025_));
  OAI21_X1   g07833(.A1(new_n8023_), .A2(new_n8025_), .B(new_n7976_), .ZN(new_n8026_));
  INV_X1     g07834(.I(new_n8024_), .ZN(new_n8027_));
  OAI21_X1   g07835(.A1(new_n8023_), .A2(new_n8027_), .B(\asqrt[31] ), .ZN(new_n8028_));
  NAND3_X1   g07836(.A1(new_n8026_), .A2(new_n8028_), .A3(new_n5435_), .ZN(new_n8029_));
  NAND2_X1   g07837(.A1(new_n8029_), .A2(new_n7973_), .ZN(new_n8030_));
  NAND2_X1   g07838(.A1(new_n8026_), .A2(new_n8028_), .ZN(new_n8031_));
  AOI21_X1   g07839(.A1(new_n8031_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n8032_));
  AOI21_X1   g07840(.A1(new_n8032_), .A2(new_n8030_), .B(new_n7970_), .ZN(new_n8033_));
  INV_X1     g07841(.I(new_n7976_), .ZN(new_n8034_));
  NOR2_X1    g07842(.A1(new_n8018_), .A2(new_n8019_), .ZN(new_n8035_));
  INV_X1     g07843(.I(new_n8004_), .ZN(new_n8036_));
  AOI21_X1   g07844(.A1(new_n8035_), .A2(new_n6813_), .B(new_n8036_), .ZN(new_n8037_));
  NAND2_X1   g07845(.A1(new_n8020_), .A2(new_n6454_), .ZN(new_n8038_));
  OAI21_X1   g07846(.A1(new_n8037_), .A2(new_n8038_), .B(new_n7982_), .ZN(new_n8039_));
  INV_X1     g07847(.I(new_n8020_), .ZN(new_n8040_));
  OAI21_X1   g07848(.A1(new_n8037_), .A2(new_n8040_), .B(\asqrt[29] ), .ZN(new_n8041_));
  NAND3_X1   g07849(.A1(new_n8039_), .A2(new_n8041_), .A3(new_n6106_), .ZN(new_n8042_));
  NAND2_X1   g07850(.A1(new_n8042_), .A2(new_n7978_), .ZN(new_n8043_));
  NAND2_X1   g07851(.A1(new_n8039_), .A2(new_n8041_), .ZN(new_n8044_));
  AOI21_X1   g07852(.A1(new_n8044_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n8045_));
  AOI21_X1   g07853(.A1(new_n8045_), .A2(new_n8043_), .B(new_n8034_), .ZN(new_n8046_));
  AOI21_X1   g07854(.A1(new_n8043_), .A2(new_n8024_), .B(new_n5750_), .ZN(new_n8047_));
  OAI21_X1   g07855(.A1(new_n8046_), .A2(new_n8047_), .B(\asqrt[32] ), .ZN(new_n8048_));
  AOI21_X1   g07856(.A1(new_n8030_), .A2(new_n8048_), .B(new_n5110_), .ZN(new_n8049_));
  NOR2_X1    g07857(.A1(new_n8033_), .A2(new_n8049_), .ZN(new_n8050_));
  AOI21_X1   g07858(.A1(new_n8050_), .A2(new_n4810_), .B(new_n7967_), .ZN(new_n8051_));
  OAI21_X1   g07859(.A1(new_n8033_), .A2(new_n8049_), .B(\asqrt[34] ), .ZN(new_n8052_));
  NAND2_X1   g07860(.A1(new_n8052_), .A2(new_n4510_), .ZN(new_n8053_));
  OAI21_X1   g07861(.A1(new_n8051_), .A2(new_n8053_), .B(new_n7963_), .ZN(new_n8054_));
  INV_X1     g07862(.I(new_n8052_), .ZN(new_n8055_));
  OAI21_X1   g07863(.A1(new_n8051_), .A2(new_n8055_), .B(\asqrt[35] ), .ZN(new_n8056_));
  NAND3_X1   g07864(.A1(new_n8054_), .A2(new_n8056_), .A3(new_n4224_), .ZN(new_n8057_));
  NAND2_X1   g07865(.A1(new_n8057_), .A2(new_n7961_), .ZN(new_n8058_));
  NAND2_X1   g07866(.A1(new_n8054_), .A2(new_n8056_), .ZN(new_n8059_));
  AOI21_X1   g07867(.A1(new_n8059_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n8060_));
  AOI21_X1   g07868(.A1(new_n8060_), .A2(new_n8058_), .B(new_n7958_), .ZN(new_n8061_));
  INV_X1     g07869(.I(new_n7963_), .ZN(new_n8062_));
  INV_X1     g07870(.I(new_n7973_), .ZN(new_n8063_));
  NOR2_X1    g07871(.A1(new_n8046_), .A2(new_n8047_), .ZN(new_n8064_));
  AOI21_X1   g07872(.A1(new_n8064_), .A2(new_n5435_), .B(new_n8063_), .ZN(new_n8065_));
  NAND2_X1   g07873(.A1(new_n8048_), .A2(new_n5110_), .ZN(new_n8066_));
  OAI21_X1   g07874(.A1(new_n8065_), .A2(new_n8066_), .B(new_n7969_), .ZN(new_n8067_));
  INV_X1     g07875(.I(new_n8048_), .ZN(new_n8068_));
  OAI21_X1   g07876(.A1(new_n8065_), .A2(new_n8068_), .B(\asqrt[33] ), .ZN(new_n8069_));
  NAND3_X1   g07877(.A1(new_n8067_), .A2(new_n8069_), .A3(new_n4810_), .ZN(new_n8070_));
  NAND2_X1   g07878(.A1(new_n8070_), .A2(new_n7966_), .ZN(new_n8071_));
  NAND2_X1   g07879(.A1(new_n8067_), .A2(new_n8069_), .ZN(new_n8072_));
  AOI21_X1   g07880(.A1(new_n8072_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n8073_));
  AOI21_X1   g07881(.A1(new_n8073_), .A2(new_n8071_), .B(new_n8062_), .ZN(new_n8074_));
  AOI21_X1   g07882(.A1(new_n8071_), .A2(new_n8052_), .B(new_n4510_), .ZN(new_n8075_));
  OAI21_X1   g07883(.A1(new_n8074_), .A2(new_n8075_), .B(\asqrt[36] ), .ZN(new_n8076_));
  AOI21_X1   g07884(.A1(new_n8058_), .A2(new_n8076_), .B(new_n3928_), .ZN(new_n8077_));
  NOR2_X1    g07885(.A1(new_n8061_), .A2(new_n8077_), .ZN(new_n8078_));
  AOI21_X1   g07886(.A1(new_n8078_), .A2(new_n3675_), .B(new_n7955_), .ZN(new_n8079_));
  OAI21_X1   g07887(.A1(new_n8061_), .A2(new_n8077_), .B(\asqrt[38] ), .ZN(new_n8080_));
  NAND2_X1   g07888(.A1(new_n8080_), .A2(new_n3400_), .ZN(new_n8081_));
  OAI21_X1   g07889(.A1(new_n8079_), .A2(new_n8081_), .B(new_n7951_), .ZN(new_n8082_));
  INV_X1     g07890(.I(new_n8080_), .ZN(new_n8083_));
  OAI21_X1   g07891(.A1(new_n8079_), .A2(new_n8083_), .B(\asqrt[39] ), .ZN(new_n8084_));
  NAND3_X1   g07892(.A1(new_n8082_), .A2(new_n8084_), .A3(new_n3167_), .ZN(new_n8085_));
  INV_X1     g07893(.I(new_n7951_), .ZN(new_n8086_));
  INV_X1     g07894(.I(new_n7961_), .ZN(new_n8087_));
  NOR2_X1    g07895(.A1(new_n8074_), .A2(new_n8075_), .ZN(new_n8088_));
  AOI21_X1   g07896(.A1(new_n8088_), .A2(new_n4224_), .B(new_n8087_), .ZN(new_n8089_));
  NAND2_X1   g07897(.A1(new_n8076_), .A2(new_n3928_), .ZN(new_n8090_));
  OAI21_X1   g07898(.A1(new_n8089_), .A2(new_n8090_), .B(new_n7957_), .ZN(new_n8091_));
  INV_X1     g07899(.I(new_n8076_), .ZN(new_n8092_));
  OAI21_X1   g07900(.A1(new_n8089_), .A2(new_n8092_), .B(\asqrt[37] ), .ZN(new_n8093_));
  NAND3_X1   g07901(.A1(new_n8091_), .A2(new_n8093_), .A3(new_n3675_), .ZN(new_n8094_));
  NAND2_X1   g07902(.A1(new_n8094_), .A2(new_n7954_), .ZN(new_n8095_));
  NAND2_X1   g07903(.A1(new_n8091_), .A2(new_n8093_), .ZN(new_n8096_));
  AOI21_X1   g07904(.A1(new_n8096_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n8097_));
  AOI21_X1   g07905(.A1(new_n8097_), .A2(new_n8095_), .B(new_n8086_), .ZN(new_n8098_));
  AOI21_X1   g07906(.A1(new_n8095_), .A2(new_n8080_), .B(new_n3400_), .ZN(new_n8099_));
  OAI21_X1   g07907(.A1(new_n8098_), .A2(new_n8099_), .B(\asqrt[40] ), .ZN(new_n8100_));
  NAND2_X1   g07908(.A1(new_n7931_), .A2(new_n7566_), .ZN(new_n8101_));
  NOR2_X1    g07909(.A1(new_n7934_), .A2(new_n7566_), .ZN(new_n8102_));
  NAND2_X1   g07910(.A1(new_n8102_), .A2(new_n7946_), .ZN(new_n8103_));
  AOI21_X1   g07911(.A1(new_n8103_), .A2(new_n8101_), .B(new_n193_), .ZN(new_n8104_));
  INV_X1     g07912(.I(new_n8104_), .ZN(new_n8105_));
  NAND3_X1   g07913(.A1(\asqrt[25] ), .A2(new_n7916_), .A3(new_n7927_), .ZN(new_n8106_));
  XOR2_X1    g07914(.A1(new_n8106_), .A2(new_n7919_), .Z(new_n8107_));
  AOI21_X1   g07915(.A1(new_n8102_), .A2(new_n7931_), .B(new_n7932_), .ZN(new_n8108_));
  OAI21_X1   g07916(.A1(new_n7886_), .A2(new_n7888_), .B(new_n7891_), .ZN(new_n8109_));
  NOR2_X1    g07917(.A1(new_n7934_), .A2(new_n8109_), .ZN(new_n8110_));
  XOR2_X1    g07918(.A1(new_n8110_), .A2(new_n7574_), .Z(new_n8111_));
  NAND3_X1   g07919(.A1(\asqrt[25] ), .A2(new_n7902_), .A3(new_n7887_), .ZN(new_n8112_));
  XOR2_X1    g07920(.A1(new_n8112_), .A2(new_n7578_), .Z(new_n8113_));
  OAI21_X1   g07921(.A1(new_n7897_), .A2(new_n7898_), .B(new_n7901_), .ZN(new_n8114_));
  NOR2_X1    g07922(.A1(new_n7934_), .A2(new_n8114_), .ZN(new_n8115_));
  XOR2_X1    g07923(.A1(new_n8115_), .A2(new_n7580_), .Z(new_n8116_));
  INV_X1     g07924(.I(new_n8116_), .ZN(new_n8117_));
  NAND3_X1   g07925(.A1(\asqrt[25] ), .A2(new_n7864_), .A3(new_n7883_), .ZN(new_n8118_));
  XOR2_X1    g07926(.A1(new_n8118_), .A2(new_n7895_), .Z(new_n8119_));
  INV_X1     g07927(.I(new_n8119_), .ZN(new_n8120_));
  OAI21_X1   g07928(.A1(new_n7858_), .A2(new_n7860_), .B(new_n7863_), .ZN(new_n8121_));
  NOR2_X1    g07929(.A1(new_n7934_), .A2(new_n8121_), .ZN(new_n8122_));
  XOR2_X1    g07930(.A1(new_n8122_), .A2(new_n7586_), .Z(new_n8123_));
  NAND3_X1   g07931(.A1(\asqrt[25] ), .A2(new_n7877_), .A3(new_n7859_), .ZN(new_n8124_));
  XOR2_X1    g07932(.A1(new_n8124_), .A2(new_n7590_), .Z(new_n8125_));
  OAI21_X1   g07933(.A1(new_n7872_), .A2(new_n7873_), .B(new_n7876_), .ZN(new_n8126_));
  NOR2_X1    g07934(.A1(new_n7934_), .A2(new_n8126_), .ZN(new_n8127_));
  XOR2_X1    g07935(.A1(new_n8127_), .A2(new_n7592_), .Z(new_n8128_));
  INV_X1     g07936(.I(new_n8128_), .ZN(new_n8129_));
  NAND3_X1   g07937(.A1(\asqrt[25] ), .A2(new_n7836_), .A3(new_n7855_), .ZN(new_n8130_));
  XOR2_X1    g07938(.A1(new_n8130_), .A2(new_n7870_), .Z(new_n8131_));
  INV_X1     g07939(.I(new_n8131_), .ZN(new_n8132_));
  OAI21_X1   g07940(.A1(new_n7830_), .A2(new_n7832_), .B(new_n7835_), .ZN(new_n8133_));
  NOR2_X1    g07941(.A1(new_n7934_), .A2(new_n8133_), .ZN(new_n8134_));
  XOR2_X1    g07942(.A1(new_n8134_), .A2(new_n7598_), .Z(new_n8135_));
  NAND3_X1   g07943(.A1(\asqrt[25] ), .A2(new_n7849_), .A3(new_n7831_), .ZN(new_n8136_));
  XOR2_X1    g07944(.A1(new_n8136_), .A2(new_n7602_), .Z(new_n8137_));
  OAI21_X1   g07945(.A1(new_n7844_), .A2(new_n7845_), .B(new_n7848_), .ZN(new_n8138_));
  NOR2_X1    g07946(.A1(new_n7934_), .A2(new_n8138_), .ZN(new_n8139_));
  XOR2_X1    g07947(.A1(new_n8139_), .A2(new_n7604_), .Z(new_n8140_));
  INV_X1     g07948(.I(new_n8140_), .ZN(new_n8141_));
  NAND3_X1   g07949(.A1(\asqrt[25] ), .A2(new_n7808_), .A3(new_n7827_), .ZN(new_n8142_));
  XOR2_X1    g07950(.A1(new_n8142_), .A2(new_n7842_), .Z(new_n8143_));
  INV_X1     g07951(.I(new_n8143_), .ZN(new_n8144_));
  OAI21_X1   g07952(.A1(new_n7802_), .A2(new_n7804_), .B(new_n7807_), .ZN(new_n8145_));
  NOR2_X1    g07953(.A1(new_n7934_), .A2(new_n8145_), .ZN(new_n8146_));
  XOR2_X1    g07954(.A1(new_n8146_), .A2(new_n7610_), .Z(new_n8147_));
  NAND3_X1   g07955(.A1(\asqrt[25] ), .A2(new_n7821_), .A3(new_n7803_), .ZN(new_n8148_));
  XOR2_X1    g07956(.A1(new_n8148_), .A2(new_n7614_), .Z(new_n8149_));
  OAI21_X1   g07957(.A1(new_n7816_), .A2(new_n7817_), .B(new_n7820_), .ZN(new_n8150_));
  NOR2_X1    g07958(.A1(new_n7934_), .A2(new_n8150_), .ZN(new_n8151_));
  XOR2_X1    g07959(.A1(new_n8151_), .A2(new_n7616_), .Z(new_n8152_));
  INV_X1     g07960(.I(new_n8152_), .ZN(new_n8153_));
  NAND3_X1   g07961(.A1(\asqrt[25] ), .A2(new_n7780_), .A3(new_n7799_), .ZN(new_n8154_));
  XOR2_X1    g07962(.A1(new_n8154_), .A2(new_n7814_), .Z(new_n8155_));
  INV_X1     g07963(.I(new_n8155_), .ZN(new_n8156_));
  OAI21_X1   g07964(.A1(new_n7774_), .A2(new_n7776_), .B(new_n7779_), .ZN(new_n8157_));
  NOR2_X1    g07965(.A1(new_n7934_), .A2(new_n8157_), .ZN(new_n8158_));
  XOR2_X1    g07966(.A1(new_n8158_), .A2(new_n7622_), .Z(new_n8159_));
  NAND3_X1   g07967(.A1(\asqrt[25] ), .A2(new_n7793_), .A3(new_n7775_), .ZN(new_n8160_));
  XOR2_X1    g07968(.A1(new_n8160_), .A2(new_n7626_), .Z(new_n8161_));
  OAI21_X1   g07969(.A1(new_n7788_), .A2(new_n7789_), .B(new_n7792_), .ZN(new_n8162_));
  NOR2_X1    g07970(.A1(new_n7934_), .A2(new_n8162_), .ZN(new_n8163_));
  XOR2_X1    g07971(.A1(new_n8163_), .A2(new_n7628_), .Z(new_n8164_));
  INV_X1     g07972(.I(new_n8164_), .ZN(new_n8165_));
  NAND3_X1   g07973(.A1(\asqrt[25] ), .A2(new_n7752_), .A3(new_n7771_), .ZN(new_n8166_));
  XOR2_X1    g07974(.A1(new_n8166_), .A2(new_n7786_), .Z(new_n8167_));
  INV_X1     g07975(.I(new_n8167_), .ZN(new_n8168_));
  NAND2_X1   g07976(.A1(new_n8085_), .A2(new_n7937_), .ZN(new_n8169_));
  NAND2_X1   g07977(.A1(new_n8082_), .A2(new_n8084_), .ZN(new_n8170_));
  AOI21_X1   g07978(.A1(new_n8170_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n8171_));
  AOI21_X1   g07979(.A1(new_n8171_), .A2(new_n8169_), .B(new_n8168_), .ZN(new_n8172_));
  AOI21_X1   g07980(.A1(new_n8169_), .A2(new_n8100_), .B(new_n2912_), .ZN(new_n8173_));
  NOR2_X1    g07981(.A1(new_n8172_), .A2(new_n8173_), .ZN(new_n8174_));
  AOI21_X1   g07982(.A1(new_n8174_), .A2(new_n2699_), .B(new_n8165_), .ZN(new_n8175_));
  OAI21_X1   g07983(.A1(new_n8172_), .A2(new_n8173_), .B(\asqrt[42] ), .ZN(new_n8176_));
  NAND2_X1   g07984(.A1(new_n8176_), .A2(new_n2464_), .ZN(new_n8177_));
  OAI21_X1   g07985(.A1(new_n8175_), .A2(new_n8177_), .B(new_n8161_), .ZN(new_n8178_));
  INV_X1     g07986(.I(new_n8176_), .ZN(new_n8179_));
  OAI21_X1   g07987(.A1(new_n8175_), .A2(new_n8179_), .B(\asqrt[43] ), .ZN(new_n8180_));
  NAND3_X1   g07988(.A1(new_n8178_), .A2(new_n8180_), .A3(new_n2271_), .ZN(new_n8181_));
  NAND2_X1   g07989(.A1(new_n8181_), .A2(new_n8159_), .ZN(new_n8182_));
  NAND2_X1   g07990(.A1(new_n8178_), .A2(new_n8180_), .ZN(new_n8183_));
  AOI21_X1   g07991(.A1(new_n8183_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n8184_));
  AOI21_X1   g07992(.A1(new_n8184_), .A2(new_n8182_), .B(new_n8156_), .ZN(new_n8185_));
  INV_X1     g07993(.I(new_n8161_), .ZN(new_n8186_));
  NOR2_X1    g07994(.A1(new_n8098_), .A2(new_n8099_), .ZN(new_n8187_));
  AOI21_X1   g07995(.A1(new_n8187_), .A2(new_n3167_), .B(new_n7938_), .ZN(new_n8188_));
  NAND2_X1   g07996(.A1(new_n8100_), .A2(new_n2912_), .ZN(new_n8189_));
  OAI21_X1   g07997(.A1(new_n8188_), .A2(new_n8189_), .B(new_n8167_), .ZN(new_n8190_));
  INV_X1     g07998(.I(new_n8100_), .ZN(new_n8191_));
  OAI21_X1   g07999(.A1(new_n8188_), .A2(new_n8191_), .B(\asqrt[41] ), .ZN(new_n8192_));
  NAND3_X1   g08000(.A1(new_n8190_), .A2(new_n8192_), .A3(new_n2699_), .ZN(new_n8193_));
  NAND2_X1   g08001(.A1(new_n8193_), .A2(new_n8164_), .ZN(new_n8194_));
  NAND2_X1   g08002(.A1(new_n8190_), .A2(new_n8192_), .ZN(new_n8195_));
  AOI21_X1   g08003(.A1(new_n8195_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n8196_));
  AOI21_X1   g08004(.A1(new_n8196_), .A2(new_n8194_), .B(new_n8186_), .ZN(new_n8197_));
  AOI21_X1   g08005(.A1(new_n8194_), .A2(new_n8176_), .B(new_n2464_), .ZN(new_n8198_));
  OAI21_X1   g08006(.A1(new_n8197_), .A2(new_n8198_), .B(\asqrt[44] ), .ZN(new_n8199_));
  AOI21_X1   g08007(.A1(new_n8182_), .A2(new_n8199_), .B(new_n2072_), .ZN(new_n8200_));
  NOR2_X1    g08008(.A1(new_n8185_), .A2(new_n8200_), .ZN(new_n8201_));
  AOI21_X1   g08009(.A1(new_n8201_), .A2(new_n1884_), .B(new_n8153_), .ZN(new_n8202_));
  OAI21_X1   g08010(.A1(new_n8185_), .A2(new_n8200_), .B(\asqrt[46] ), .ZN(new_n8203_));
  NAND2_X1   g08011(.A1(new_n8203_), .A2(new_n1688_), .ZN(new_n8204_));
  OAI21_X1   g08012(.A1(new_n8202_), .A2(new_n8204_), .B(new_n8149_), .ZN(new_n8205_));
  INV_X1     g08013(.I(new_n8203_), .ZN(new_n8206_));
  OAI21_X1   g08014(.A1(new_n8202_), .A2(new_n8206_), .B(\asqrt[47] ), .ZN(new_n8207_));
  NAND3_X1   g08015(.A1(new_n8205_), .A2(new_n8207_), .A3(new_n1533_), .ZN(new_n8208_));
  NAND2_X1   g08016(.A1(new_n8208_), .A2(new_n8147_), .ZN(new_n8209_));
  NAND2_X1   g08017(.A1(new_n8205_), .A2(new_n8207_), .ZN(new_n8210_));
  AOI21_X1   g08018(.A1(new_n8210_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n8211_));
  AOI21_X1   g08019(.A1(new_n8211_), .A2(new_n8209_), .B(new_n8144_), .ZN(new_n8212_));
  INV_X1     g08020(.I(new_n8149_), .ZN(new_n8213_));
  INV_X1     g08021(.I(new_n8159_), .ZN(new_n8214_));
  NOR2_X1    g08022(.A1(new_n8197_), .A2(new_n8198_), .ZN(new_n8215_));
  AOI21_X1   g08023(.A1(new_n8215_), .A2(new_n2271_), .B(new_n8214_), .ZN(new_n8216_));
  NAND2_X1   g08024(.A1(new_n8199_), .A2(new_n2072_), .ZN(new_n8217_));
  OAI21_X1   g08025(.A1(new_n8216_), .A2(new_n8217_), .B(new_n8155_), .ZN(new_n8218_));
  INV_X1     g08026(.I(new_n8199_), .ZN(new_n8219_));
  OAI21_X1   g08027(.A1(new_n8216_), .A2(new_n8219_), .B(\asqrt[45] ), .ZN(new_n8220_));
  NAND3_X1   g08028(.A1(new_n8218_), .A2(new_n8220_), .A3(new_n1884_), .ZN(new_n8221_));
  NAND2_X1   g08029(.A1(new_n8221_), .A2(new_n8152_), .ZN(new_n8222_));
  NAND2_X1   g08030(.A1(new_n8218_), .A2(new_n8220_), .ZN(new_n8223_));
  AOI21_X1   g08031(.A1(new_n8223_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n8224_));
  AOI21_X1   g08032(.A1(new_n8224_), .A2(new_n8222_), .B(new_n8213_), .ZN(new_n8225_));
  AOI21_X1   g08033(.A1(new_n8222_), .A2(new_n8203_), .B(new_n1688_), .ZN(new_n8226_));
  OAI21_X1   g08034(.A1(new_n8225_), .A2(new_n8226_), .B(\asqrt[48] ), .ZN(new_n8227_));
  AOI21_X1   g08035(.A1(new_n8209_), .A2(new_n8227_), .B(new_n1368_), .ZN(new_n8228_));
  NOR2_X1    g08036(.A1(new_n8212_), .A2(new_n8228_), .ZN(new_n8229_));
  AOI21_X1   g08037(.A1(new_n8229_), .A2(new_n1228_), .B(new_n8141_), .ZN(new_n8230_));
  OAI21_X1   g08038(.A1(new_n8212_), .A2(new_n8228_), .B(\asqrt[50] ), .ZN(new_n8231_));
  NAND2_X1   g08039(.A1(new_n8231_), .A2(new_n1088_), .ZN(new_n8232_));
  OAI21_X1   g08040(.A1(new_n8230_), .A2(new_n8232_), .B(new_n8137_), .ZN(new_n8233_));
  INV_X1     g08041(.I(new_n8231_), .ZN(new_n8234_));
  OAI21_X1   g08042(.A1(new_n8230_), .A2(new_n8234_), .B(\asqrt[51] ), .ZN(new_n8235_));
  NAND3_X1   g08043(.A1(new_n8233_), .A2(new_n8235_), .A3(new_n962_), .ZN(new_n8236_));
  NAND2_X1   g08044(.A1(new_n8236_), .A2(new_n8135_), .ZN(new_n8237_));
  NAND2_X1   g08045(.A1(new_n8233_), .A2(new_n8235_), .ZN(new_n8238_));
  AOI21_X1   g08046(.A1(new_n8238_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n8239_));
  AOI21_X1   g08047(.A1(new_n8239_), .A2(new_n8237_), .B(new_n8132_), .ZN(new_n8240_));
  INV_X1     g08048(.I(new_n8137_), .ZN(new_n8241_));
  INV_X1     g08049(.I(new_n8147_), .ZN(new_n8242_));
  NOR2_X1    g08050(.A1(new_n8225_), .A2(new_n8226_), .ZN(new_n8243_));
  AOI21_X1   g08051(.A1(new_n8243_), .A2(new_n1533_), .B(new_n8242_), .ZN(new_n8244_));
  NAND2_X1   g08052(.A1(new_n8227_), .A2(new_n1368_), .ZN(new_n8245_));
  OAI21_X1   g08053(.A1(new_n8244_), .A2(new_n8245_), .B(new_n8143_), .ZN(new_n8246_));
  INV_X1     g08054(.I(new_n8227_), .ZN(new_n8247_));
  OAI21_X1   g08055(.A1(new_n8244_), .A2(new_n8247_), .B(\asqrt[49] ), .ZN(new_n8248_));
  NAND3_X1   g08056(.A1(new_n8246_), .A2(new_n8248_), .A3(new_n1228_), .ZN(new_n8249_));
  NAND2_X1   g08057(.A1(new_n8249_), .A2(new_n8140_), .ZN(new_n8250_));
  NAND2_X1   g08058(.A1(new_n8246_), .A2(new_n8248_), .ZN(new_n8251_));
  AOI21_X1   g08059(.A1(new_n8251_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n8252_));
  AOI21_X1   g08060(.A1(new_n8252_), .A2(new_n8250_), .B(new_n8241_), .ZN(new_n8253_));
  AOI21_X1   g08061(.A1(new_n8250_), .A2(new_n8231_), .B(new_n1088_), .ZN(new_n8254_));
  OAI21_X1   g08062(.A1(new_n8253_), .A2(new_n8254_), .B(\asqrt[52] ), .ZN(new_n8255_));
  AOI21_X1   g08063(.A1(new_n8237_), .A2(new_n8255_), .B(new_n842_), .ZN(new_n8256_));
  NOR2_X1    g08064(.A1(new_n8240_), .A2(new_n8256_), .ZN(new_n8257_));
  AOI21_X1   g08065(.A1(new_n8257_), .A2(new_n720_), .B(new_n8129_), .ZN(new_n8258_));
  OAI21_X1   g08066(.A1(new_n8240_), .A2(new_n8256_), .B(\asqrt[54] ), .ZN(new_n8259_));
  NAND2_X1   g08067(.A1(new_n8259_), .A2(new_n630_), .ZN(new_n8260_));
  OAI21_X1   g08068(.A1(new_n8258_), .A2(new_n8260_), .B(new_n8125_), .ZN(new_n8261_));
  INV_X1     g08069(.I(new_n8259_), .ZN(new_n8262_));
  OAI21_X1   g08070(.A1(new_n8258_), .A2(new_n8262_), .B(\asqrt[55] ), .ZN(new_n8263_));
  NAND3_X1   g08071(.A1(new_n8261_), .A2(new_n8263_), .A3(new_n545_), .ZN(new_n8264_));
  NAND2_X1   g08072(.A1(new_n8264_), .A2(new_n8123_), .ZN(new_n8265_));
  NAND2_X1   g08073(.A1(new_n8261_), .A2(new_n8263_), .ZN(new_n8266_));
  AOI21_X1   g08074(.A1(new_n8266_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n8267_));
  AOI21_X1   g08075(.A1(new_n8267_), .A2(new_n8265_), .B(new_n8120_), .ZN(new_n8268_));
  INV_X1     g08076(.I(new_n8125_), .ZN(new_n8269_));
  INV_X1     g08077(.I(new_n8135_), .ZN(new_n8270_));
  NOR2_X1    g08078(.A1(new_n8253_), .A2(new_n8254_), .ZN(new_n8271_));
  AOI21_X1   g08079(.A1(new_n8271_), .A2(new_n962_), .B(new_n8270_), .ZN(new_n8272_));
  NAND2_X1   g08080(.A1(new_n8255_), .A2(new_n842_), .ZN(new_n8273_));
  OAI21_X1   g08081(.A1(new_n8272_), .A2(new_n8273_), .B(new_n8131_), .ZN(new_n8274_));
  INV_X1     g08082(.I(new_n8255_), .ZN(new_n8275_));
  OAI21_X1   g08083(.A1(new_n8272_), .A2(new_n8275_), .B(\asqrt[53] ), .ZN(new_n8276_));
  NAND3_X1   g08084(.A1(new_n8274_), .A2(new_n8276_), .A3(new_n720_), .ZN(new_n8277_));
  NAND2_X1   g08085(.A1(new_n8277_), .A2(new_n8128_), .ZN(new_n8278_));
  NAND2_X1   g08086(.A1(new_n8274_), .A2(new_n8276_), .ZN(new_n8279_));
  AOI21_X1   g08087(.A1(new_n8279_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n8280_));
  AOI21_X1   g08088(.A1(new_n8280_), .A2(new_n8278_), .B(new_n8269_), .ZN(new_n8281_));
  AOI21_X1   g08089(.A1(new_n8278_), .A2(new_n8259_), .B(new_n630_), .ZN(new_n8282_));
  OAI21_X1   g08090(.A1(new_n8281_), .A2(new_n8282_), .B(\asqrt[56] ), .ZN(new_n8283_));
  AOI21_X1   g08091(.A1(new_n8265_), .A2(new_n8283_), .B(new_n450_), .ZN(new_n8284_));
  NOR2_X1    g08092(.A1(new_n8268_), .A2(new_n8284_), .ZN(new_n8285_));
  AOI21_X1   g08093(.A1(new_n8285_), .A2(new_n403_), .B(new_n8117_), .ZN(new_n8286_));
  OAI21_X1   g08094(.A1(new_n8268_), .A2(new_n8284_), .B(\asqrt[58] ), .ZN(new_n8287_));
  NAND2_X1   g08095(.A1(new_n8287_), .A2(new_n339_), .ZN(new_n8288_));
  OAI21_X1   g08096(.A1(new_n8286_), .A2(new_n8288_), .B(new_n8113_), .ZN(new_n8289_));
  INV_X1     g08097(.I(new_n8287_), .ZN(new_n8290_));
  OAI21_X1   g08098(.A1(new_n8286_), .A2(new_n8290_), .B(\asqrt[59] ), .ZN(new_n8291_));
  NAND3_X1   g08099(.A1(new_n8289_), .A2(new_n8291_), .A3(new_n288_), .ZN(new_n8292_));
  NAND2_X1   g08100(.A1(new_n8292_), .A2(new_n8111_), .ZN(new_n8293_));
  INV_X1     g08101(.I(new_n8113_), .ZN(new_n8294_));
  INV_X1     g08102(.I(new_n8123_), .ZN(new_n8295_));
  NOR2_X1    g08103(.A1(new_n8281_), .A2(new_n8282_), .ZN(new_n8296_));
  AOI21_X1   g08104(.A1(new_n8296_), .A2(new_n545_), .B(new_n8295_), .ZN(new_n8297_));
  NAND2_X1   g08105(.A1(new_n8283_), .A2(new_n450_), .ZN(new_n8298_));
  OAI21_X1   g08106(.A1(new_n8297_), .A2(new_n8298_), .B(new_n8119_), .ZN(new_n8299_));
  INV_X1     g08107(.I(new_n8283_), .ZN(new_n8300_));
  OAI21_X1   g08108(.A1(new_n8297_), .A2(new_n8300_), .B(\asqrt[57] ), .ZN(new_n8301_));
  NAND3_X1   g08109(.A1(new_n8299_), .A2(new_n8301_), .A3(new_n403_), .ZN(new_n8302_));
  NAND2_X1   g08110(.A1(new_n8302_), .A2(new_n8116_), .ZN(new_n8303_));
  NAND2_X1   g08111(.A1(new_n8299_), .A2(new_n8301_), .ZN(new_n8304_));
  AOI21_X1   g08112(.A1(new_n8304_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n8305_));
  AOI21_X1   g08113(.A1(new_n8305_), .A2(new_n8303_), .B(new_n8294_), .ZN(new_n8306_));
  AOI21_X1   g08114(.A1(new_n8303_), .A2(new_n8287_), .B(new_n339_), .ZN(new_n8307_));
  OAI21_X1   g08115(.A1(new_n8306_), .A2(new_n8307_), .B(\asqrt[60] ), .ZN(new_n8308_));
  AOI21_X1   g08116(.A1(new_n8293_), .A2(new_n8308_), .B(new_n242_), .ZN(new_n8309_));
  NAND3_X1   g08117(.A1(\asqrt[25] ), .A2(new_n7892_), .A3(new_n7908_), .ZN(new_n8310_));
  XOR2_X1    g08118(.A1(new_n8310_), .A2(new_n7920_), .Z(new_n8311_));
  INV_X1     g08119(.I(new_n8311_), .ZN(new_n8312_));
  NAND2_X1   g08120(.A1(new_n8289_), .A2(new_n8291_), .ZN(new_n8313_));
  AOI21_X1   g08121(.A1(new_n8313_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n8314_));
  AOI21_X1   g08122(.A1(new_n8314_), .A2(new_n8293_), .B(new_n8312_), .ZN(new_n8315_));
  OAI21_X1   g08123(.A1(new_n8315_), .A2(new_n8309_), .B(\asqrt[62] ), .ZN(new_n8316_));
  INV_X1     g08124(.I(new_n8316_), .ZN(new_n8317_));
  NOR2_X1    g08125(.A1(new_n8315_), .A2(new_n8309_), .ZN(new_n8318_));
  AOI21_X1   g08126(.A1(new_n7893_), .A2(new_n7914_), .B(new_n7909_), .ZN(new_n8319_));
  NAND2_X1   g08127(.A1(\asqrt[25] ), .A2(new_n8319_), .ZN(new_n8320_));
  XOR2_X1    g08128(.A1(new_n8320_), .A2(new_n7912_), .Z(new_n8321_));
  INV_X1     g08129(.I(new_n8321_), .ZN(new_n8322_));
  AOI21_X1   g08130(.A1(new_n8318_), .A2(new_n234_), .B(new_n8322_), .ZN(new_n8323_));
  OAI21_X1   g08131(.A1(new_n8323_), .A2(new_n8317_), .B(new_n8108_), .ZN(new_n8324_));
  OAI21_X1   g08132(.A1(new_n8324_), .A2(new_n8107_), .B(new_n193_), .ZN(new_n8325_));
  NOR2_X1    g08133(.A1(new_n8323_), .A2(new_n8317_), .ZN(new_n8326_));
  NAND2_X1   g08134(.A1(new_n8326_), .A2(new_n8107_), .ZN(new_n8327_));
  NOR2_X1    g08135(.A1(\asqrt[25] ), .A2(new_n7567_), .ZN(new_n8328_));
  INV_X1     g08136(.I(new_n8328_), .ZN(new_n8329_));
  NAND4_X1   g08137(.A1(new_n8325_), .A2(new_n8105_), .A3(new_n8327_), .A4(new_n8329_), .ZN(\asqrt[24] ));
  NAND3_X1   g08138(.A1(\asqrt[24] ), .A2(new_n8085_), .A3(new_n8100_), .ZN(new_n8331_));
  XOR2_X1    g08139(.A1(new_n8331_), .A2(new_n7938_), .Z(new_n8332_));
  INV_X1     g08140(.I(new_n8111_), .ZN(new_n8333_));
  NOR2_X1    g08141(.A1(new_n8306_), .A2(new_n8307_), .ZN(new_n8334_));
  AOI21_X1   g08142(.A1(new_n8334_), .A2(new_n288_), .B(new_n8333_), .ZN(new_n8335_));
  INV_X1     g08143(.I(new_n8308_), .ZN(new_n8336_));
  OAI21_X1   g08144(.A1(new_n8335_), .A2(new_n8336_), .B(\asqrt[61] ), .ZN(new_n8337_));
  NAND2_X1   g08145(.A1(new_n8308_), .A2(new_n242_), .ZN(new_n8338_));
  OAI21_X1   g08146(.A1(new_n8335_), .A2(new_n8338_), .B(new_n8311_), .ZN(new_n8339_));
  NAND3_X1   g08147(.A1(new_n8339_), .A2(new_n8337_), .A3(new_n234_), .ZN(new_n8340_));
  NAND2_X1   g08148(.A1(new_n8340_), .A2(new_n8321_), .ZN(new_n8341_));
  NAND2_X1   g08149(.A1(new_n8341_), .A2(new_n8316_), .ZN(new_n8342_));
  NAND2_X1   g08150(.A1(new_n8342_), .A2(new_n8107_), .ZN(new_n8343_));
  INV_X1     g08151(.I(new_n8107_), .ZN(new_n8344_));
  INV_X1     g08152(.I(new_n8108_), .ZN(new_n8345_));
  AOI21_X1   g08153(.A1(new_n8341_), .A2(new_n8316_), .B(new_n8345_), .ZN(new_n8346_));
  AOI21_X1   g08154(.A1(new_n8346_), .A2(new_n8344_), .B(\asqrt[63] ), .ZN(new_n8347_));
  NOR2_X1    g08155(.A1(new_n8342_), .A2(new_n8344_), .ZN(new_n8348_));
  NOR4_X1    g08156(.A1(new_n8347_), .A2(new_n8104_), .A3(new_n8348_), .A4(new_n8328_), .ZN(new_n8349_));
  NOR2_X1    g08157(.A1(new_n8349_), .A2(new_n8107_), .ZN(new_n8350_));
  NAND2_X1   g08158(.A1(new_n8350_), .A2(new_n8326_), .ZN(new_n8351_));
  AOI21_X1   g08159(.A1(new_n8351_), .A2(new_n8343_), .B(new_n193_), .ZN(new_n8352_));
  NAND3_X1   g08160(.A1(\asqrt[24] ), .A2(new_n8316_), .A3(new_n8340_), .ZN(new_n8353_));
  XOR2_X1    g08161(.A1(new_n8353_), .A2(new_n8321_), .Z(new_n8354_));
  INV_X1     g08162(.I(new_n8354_), .ZN(new_n8355_));
  AOI21_X1   g08163(.A1(new_n8350_), .A2(new_n8342_), .B(new_n8348_), .ZN(new_n8356_));
  INV_X1     g08164(.I(new_n8356_), .ZN(new_n8357_));
  OAI21_X1   g08165(.A1(new_n8286_), .A2(new_n8288_), .B(new_n8291_), .ZN(new_n8358_));
  NOR2_X1    g08166(.A1(new_n8349_), .A2(new_n8358_), .ZN(new_n8359_));
  XOR2_X1    g08167(.A1(new_n8359_), .A2(new_n8113_), .Z(new_n8360_));
  NAND3_X1   g08168(.A1(\asqrt[24] ), .A2(new_n8302_), .A3(new_n8287_), .ZN(new_n8361_));
  XOR2_X1    g08169(.A1(new_n8361_), .A2(new_n8117_), .Z(new_n8362_));
  OAI21_X1   g08170(.A1(new_n8297_), .A2(new_n8298_), .B(new_n8301_), .ZN(new_n8363_));
  NOR2_X1    g08171(.A1(new_n8349_), .A2(new_n8363_), .ZN(new_n8364_));
  XOR2_X1    g08172(.A1(new_n8364_), .A2(new_n8119_), .Z(new_n8365_));
  INV_X1     g08173(.I(new_n8365_), .ZN(new_n8366_));
  NAND3_X1   g08174(.A1(\asqrt[24] ), .A2(new_n8264_), .A3(new_n8283_), .ZN(new_n8367_));
  XOR2_X1    g08175(.A1(new_n8367_), .A2(new_n8295_), .Z(new_n8368_));
  INV_X1     g08176(.I(new_n8368_), .ZN(new_n8369_));
  OAI21_X1   g08177(.A1(new_n8258_), .A2(new_n8260_), .B(new_n8263_), .ZN(new_n8370_));
  NOR2_X1    g08178(.A1(new_n8349_), .A2(new_n8370_), .ZN(new_n8371_));
  XOR2_X1    g08179(.A1(new_n8371_), .A2(new_n8125_), .Z(new_n8372_));
  NAND3_X1   g08180(.A1(\asqrt[24] ), .A2(new_n8277_), .A3(new_n8259_), .ZN(new_n8373_));
  XOR2_X1    g08181(.A1(new_n8373_), .A2(new_n8129_), .Z(new_n8374_));
  OAI21_X1   g08182(.A1(new_n8272_), .A2(new_n8273_), .B(new_n8276_), .ZN(new_n8375_));
  NOR2_X1    g08183(.A1(new_n8349_), .A2(new_n8375_), .ZN(new_n8376_));
  XOR2_X1    g08184(.A1(new_n8376_), .A2(new_n8131_), .Z(new_n8377_));
  INV_X1     g08185(.I(new_n8377_), .ZN(new_n8378_));
  NAND3_X1   g08186(.A1(\asqrt[24] ), .A2(new_n8236_), .A3(new_n8255_), .ZN(new_n8379_));
  XOR2_X1    g08187(.A1(new_n8379_), .A2(new_n8270_), .Z(new_n8380_));
  INV_X1     g08188(.I(new_n8380_), .ZN(new_n8381_));
  OAI21_X1   g08189(.A1(new_n8230_), .A2(new_n8232_), .B(new_n8235_), .ZN(new_n8382_));
  NOR2_X1    g08190(.A1(new_n8349_), .A2(new_n8382_), .ZN(new_n8383_));
  XOR2_X1    g08191(.A1(new_n8383_), .A2(new_n8137_), .Z(new_n8384_));
  NAND3_X1   g08192(.A1(\asqrt[24] ), .A2(new_n8249_), .A3(new_n8231_), .ZN(new_n8385_));
  XOR2_X1    g08193(.A1(new_n8385_), .A2(new_n8141_), .Z(new_n8386_));
  OAI21_X1   g08194(.A1(new_n8244_), .A2(new_n8245_), .B(new_n8248_), .ZN(new_n8387_));
  NOR2_X1    g08195(.A1(new_n8349_), .A2(new_n8387_), .ZN(new_n8388_));
  XOR2_X1    g08196(.A1(new_n8388_), .A2(new_n8143_), .Z(new_n8389_));
  INV_X1     g08197(.I(new_n8389_), .ZN(new_n8390_));
  NAND3_X1   g08198(.A1(\asqrt[24] ), .A2(new_n8208_), .A3(new_n8227_), .ZN(new_n8391_));
  XOR2_X1    g08199(.A1(new_n8391_), .A2(new_n8242_), .Z(new_n8392_));
  INV_X1     g08200(.I(new_n8392_), .ZN(new_n8393_));
  OAI21_X1   g08201(.A1(new_n8202_), .A2(new_n8204_), .B(new_n8207_), .ZN(new_n8394_));
  NOR2_X1    g08202(.A1(new_n8349_), .A2(new_n8394_), .ZN(new_n8395_));
  XOR2_X1    g08203(.A1(new_n8395_), .A2(new_n8149_), .Z(new_n8396_));
  NAND3_X1   g08204(.A1(\asqrt[24] ), .A2(new_n8221_), .A3(new_n8203_), .ZN(new_n8397_));
  XOR2_X1    g08205(.A1(new_n8397_), .A2(new_n8153_), .Z(new_n8398_));
  OAI21_X1   g08206(.A1(new_n8216_), .A2(new_n8217_), .B(new_n8220_), .ZN(new_n8399_));
  NOR2_X1    g08207(.A1(new_n8349_), .A2(new_n8399_), .ZN(new_n8400_));
  XOR2_X1    g08208(.A1(new_n8400_), .A2(new_n8155_), .Z(new_n8401_));
  INV_X1     g08209(.I(new_n8401_), .ZN(new_n8402_));
  NAND3_X1   g08210(.A1(\asqrt[24] ), .A2(new_n8181_), .A3(new_n8199_), .ZN(new_n8403_));
  XOR2_X1    g08211(.A1(new_n8403_), .A2(new_n8214_), .Z(new_n8404_));
  INV_X1     g08212(.I(new_n8404_), .ZN(new_n8405_));
  OAI21_X1   g08213(.A1(new_n8175_), .A2(new_n8177_), .B(new_n8180_), .ZN(new_n8406_));
  NOR2_X1    g08214(.A1(new_n8349_), .A2(new_n8406_), .ZN(new_n8407_));
  XOR2_X1    g08215(.A1(new_n8407_), .A2(new_n8161_), .Z(new_n8408_));
  NAND3_X1   g08216(.A1(\asqrt[24] ), .A2(new_n8193_), .A3(new_n8176_), .ZN(new_n8409_));
  XOR2_X1    g08217(.A1(new_n8409_), .A2(new_n8165_), .Z(new_n8410_));
  OAI21_X1   g08218(.A1(new_n8188_), .A2(new_n8189_), .B(new_n8192_), .ZN(new_n8411_));
  NOR2_X1    g08219(.A1(new_n8349_), .A2(new_n8411_), .ZN(new_n8412_));
  XOR2_X1    g08220(.A1(new_n8412_), .A2(new_n8167_), .Z(new_n8413_));
  INV_X1     g08221(.I(new_n8413_), .ZN(new_n8414_));
  INV_X1     g08222(.I(new_n8332_), .ZN(new_n8415_));
  OAI21_X1   g08223(.A1(new_n8079_), .A2(new_n8081_), .B(new_n8084_), .ZN(new_n8416_));
  NOR2_X1    g08224(.A1(new_n8349_), .A2(new_n8416_), .ZN(new_n8417_));
  XOR2_X1    g08225(.A1(new_n8417_), .A2(new_n7951_), .Z(new_n8418_));
  NAND3_X1   g08226(.A1(\asqrt[24] ), .A2(new_n8094_), .A3(new_n8080_), .ZN(new_n8419_));
  XOR2_X1    g08227(.A1(new_n8419_), .A2(new_n7955_), .Z(new_n8420_));
  OAI21_X1   g08228(.A1(new_n8089_), .A2(new_n8090_), .B(new_n8093_), .ZN(new_n8421_));
  NOR2_X1    g08229(.A1(new_n8349_), .A2(new_n8421_), .ZN(new_n8422_));
  XOR2_X1    g08230(.A1(new_n8422_), .A2(new_n7957_), .Z(new_n8423_));
  INV_X1     g08231(.I(new_n8423_), .ZN(new_n8424_));
  NAND3_X1   g08232(.A1(\asqrt[24] ), .A2(new_n8057_), .A3(new_n8076_), .ZN(new_n8425_));
  XOR2_X1    g08233(.A1(new_n8425_), .A2(new_n8087_), .Z(new_n8426_));
  INV_X1     g08234(.I(new_n8426_), .ZN(new_n8427_));
  OAI21_X1   g08235(.A1(new_n8051_), .A2(new_n8053_), .B(new_n8056_), .ZN(new_n8428_));
  NOR2_X1    g08236(.A1(new_n8349_), .A2(new_n8428_), .ZN(new_n8429_));
  XOR2_X1    g08237(.A1(new_n8429_), .A2(new_n7963_), .Z(new_n8430_));
  NAND3_X1   g08238(.A1(\asqrt[24] ), .A2(new_n8070_), .A3(new_n8052_), .ZN(new_n8431_));
  XOR2_X1    g08239(.A1(new_n8431_), .A2(new_n7967_), .Z(new_n8432_));
  OAI21_X1   g08240(.A1(new_n8065_), .A2(new_n8066_), .B(new_n8069_), .ZN(new_n8433_));
  NOR2_X1    g08241(.A1(new_n8349_), .A2(new_n8433_), .ZN(new_n8434_));
  XOR2_X1    g08242(.A1(new_n8434_), .A2(new_n7969_), .Z(new_n8435_));
  INV_X1     g08243(.I(new_n8435_), .ZN(new_n8436_));
  NAND3_X1   g08244(.A1(\asqrt[24] ), .A2(new_n8029_), .A3(new_n8048_), .ZN(new_n8437_));
  XOR2_X1    g08245(.A1(new_n8437_), .A2(new_n8063_), .Z(new_n8438_));
  INV_X1     g08246(.I(new_n8438_), .ZN(new_n8439_));
  OAI21_X1   g08247(.A1(new_n8023_), .A2(new_n8025_), .B(new_n8028_), .ZN(new_n8440_));
  NOR2_X1    g08248(.A1(new_n8349_), .A2(new_n8440_), .ZN(new_n8441_));
  XOR2_X1    g08249(.A1(new_n8441_), .A2(new_n7976_), .Z(new_n8442_));
  NAND3_X1   g08250(.A1(\asqrt[24] ), .A2(new_n8042_), .A3(new_n8024_), .ZN(new_n8443_));
  XOR2_X1    g08251(.A1(new_n8443_), .A2(new_n7979_), .Z(new_n8444_));
  OAI21_X1   g08252(.A1(new_n8037_), .A2(new_n8038_), .B(new_n8041_), .ZN(new_n8445_));
  NOR2_X1    g08253(.A1(new_n8349_), .A2(new_n8445_), .ZN(new_n8446_));
  XOR2_X1    g08254(.A1(new_n8446_), .A2(new_n7982_), .Z(new_n8447_));
  INV_X1     g08255(.I(new_n8447_), .ZN(new_n8448_));
  NAND3_X1   g08256(.A1(\asqrt[24] ), .A2(new_n8002_), .A3(new_n8020_), .ZN(new_n8449_));
  XOR2_X1    g08257(.A1(new_n8449_), .A2(new_n8036_), .Z(new_n8450_));
  INV_X1     g08258(.I(new_n8450_), .ZN(new_n8451_));
  NOR2_X1    g08259(.A1(new_n7999_), .A2(\asqrt[27] ), .ZN(new_n8452_));
  NOR3_X1    g08260(.A1(new_n8349_), .A2(new_n8452_), .A3(new_n8019_), .ZN(new_n8453_));
  XOR2_X1    g08261(.A1(new_n8453_), .A2(new_n7990_), .Z(new_n8454_));
  NOR3_X1    g08262(.A1(new_n8349_), .A2(\a[48] ), .A3(\a[49] ), .ZN(new_n8455_));
  NOR4_X1    g08263(.A1(new_n8347_), .A2(new_n7934_), .A3(new_n8104_), .A4(new_n8348_), .ZN(new_n8456_));
  OAI21_X1   g08264(.A1(new_n8455_), .A2(new_n8456_), .B(new_n7668_), .ZN(new_n8457_));
  NAND3_X1   g08265(.A1(\asqrt[24] ), .A2(new_n7991_), .A3(new_n7992_), .ZN(new_n8458_));
  INV_X1     g08266(.I(new_n8456_), .ZN(new_n8459_));
  NAND3_X1   g08267(.A1(new_n8458_), .A2(\a[50] ), .A3(new_n8459_), .ZN(new_n8460_));
  NAND2_X1   g08268(.A1(new_n8457_), .A2(new_n8460_), .ZN(new_n8461_));
  INV_X1     g08269(.I(\a[46] ), .ZN(new_n8462_));
  INV_X1     g08270(.I(\a[47] ), .ZN(new_n8463_));
  NAND3_X1   g08271(.A1(new_n8462_), .A2(new_n8463_), .A3(new_n7991_), .ZN(new_n8464_));
  NAND2_X1   g08272(.A1(\asqrt[24] ), .A2(\a[48] ), .ZN(new_n8465_));
  AOI21_X1   g08273(.A1(new_n8465_), .A2(new_n8464_), .B(new_n7934_), .ZN(new_n8466_));
  AOI21_X1   g08274(.A1(\asqrt[24] ), .A2(new_n7991_), .B(new_n7992_), .ZN(new_n8467_));
  NOR2_X1    g08275(.A1(new_n8455_), .A2(new_n8467_), .ZN(new_n8468_));
  NAND3_X1   g08276(.A1(new_n8465_), .A2(new_n7934_), .A3(new_n8464_), .ZN(new_n8469_));
  AOI21_X1   g08277(.A1(new_n8468_), .A2(new_n8469_), .B(new_n8466_), .ZN(new_n8470_));
  AOI21_X1   g08278(.A1(new_n8470_), .A2(new_n7561_), .B(new_n8461_), .ZN(new_n8471_));
  NOR2_X1    g08279(.A1(new_n8470_), .A2(new_n7561_), .ZN(new_n8472_));
  NOR3_X1    g08280(.A1(new_n8471_), .A2(\asqrt[27] ), .A3(new_n8472_), .ZN(new_n8473_));
  NOR3_X1    g08281(.A1(new_n8349_), .A2(new_n8013_), .A3(new_n7998_), .ZN(new_n8474_));
  XOR2_X1    g08282(.A1(new_n8474_), .A2(new_n8015_), .Z(new_n8475_));
  INV_X1     g08283(.I(new_n8475_), .ZN(new_n8476_));
  OAI21_X1   g08284(.A1(new_n8471_), .A2(new_n8472_), .B(\asqrt[27] ), .ZN(new_n8477_));
  OAI21_X1   g08285(.A1(new_n8473_), .A2(new_n8476_), .B(new_n8477_), .ZN(new_n8478_));
  OAI21_X1   g08286(.A1(new_n8478_), .A2(\asqrt[28] ), .B(new_n8454_), .ZN(new_n8479_));
  AOI21_X1   g08287(.A1(new_n8478_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n8480_));
  AOI21_X1   g08288(.A1(new_n8480_), .A2(new_n8479_), .B(new_n8451_), .ZN(new_n8481_));
  NAND2_X1   g08289(.A1(new_n8478_), .A2(\asqrt[28] ), .ZN(new_n8482_));
  AOI21_X1   g08290(.A1(new_n8479_), .A2(new_n8482_), .B(new_n6454_), .ZN(new_n8483_));
  NOR2_X1    g08291(.A1(new_n8481_), .A2(new_n8483_), .ZN(new_n8484_));
  AOI21_X1   g08292(.A1(new_n8484_), .A2(new_n6106_), .B(new_n8448_), .ZN(new_n8485_));
  OAI21_X1   g08293(.A1(new_n8481_), .A2(new_n8483_), .B(\asqrt[30] ), .ZN(new_n8486_));
  NAND2_X1   g08294(.A1(new_n8486_), .A2(new_n5750_), .ZN(new_n8487_));
  OAI21_X1   g08295(.A1(new_n8485_), .A2(new_n8487_), .B(new_n8444_), .ZN(new_n8488_));
  INV_X1     g08296(.I(new_n8486_), .ZN(new_n8489_));
  OAI21_X1   g08297(.A1(new_n8485_), .A2(new_n8489_), .B(\asqrt[31] ), .ZN(new_n8490_));
  NAND3_X1   g08298(.A1(new_n8488_), .A2(new_n8490_), .A3(new_n5435_), .ZN(new_n8491_));
  NAND2_X1   g08299(.A1(new_n8491_), .A2(new_n8442_), .ZN(new_n8492_));
  NAND2_X1   g08300(.A1(new_n8488_), .A2(new_n8490_), .ZN(new_n8493_));
  AOI21_X1   g08301(.A1(new_n8493_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n8494_));
  AOI21_X1   g08302(.A1(new_n8494_), .A2(new_n8492_), .B(new_n8439_), .ZN(new_n8495_));
  INV_X1     g08303(.I(new_n8444_), .ZN(new_n8496_));
  INV_X1     g08304(.I(new_n8454_), .ZN(new_n8497_));
  AOI21_X1   g08305(.A1(new_n8458_), .A2(new_n8459_), .B(\a[50] ), .ZN(new_n8498_));
  NOR3_X1    g08306(.A1(new_n8455_), .A2(new_n7668_), .A3(new_n8456_), .ZN(new_n8499_));
  NOR2_X1    g08307(.A1(new_n8499_), .A2(new_n8498_), .ZN(new_n8500_));
  OAI21_X1   g08308(.A1(new_n8349_), .A2(new_n7991_), .B(new_n8464_), .ZN(new_n8501_));
  NAND2_X1   g08309(.A1(new_n8501_), .A2(\asqrt[25] ), .ZN(new_n8502_));
  OAI21_X1   g08310(.A1(new_n8349_), .A2(\a[48] ), .B(\a[49] ), .ZN(new_n8503_));
  NAND2_X1   g08311(.A1(new_n8503_), .A2(new_n8458_), .ZN(new_n8504_));
  NOR2_X1    g08312(.A1(new_n8501_), .A2(\asqrt[25] ), .ZN(new_n8505_));
  OAI21_X1   g08313(.A1(new_n8504_), .A2(new_n8505_), .B(new_n8502_), .ZN(new_n8506_));
  OAI21_X1   g08314(.A1(\asqrt[26] ), .A2(new_n8506_), .B(new_n8500_), .ZN(new_n8507_));
  NAND2_X1   g08315(.A1(new_n8506_), .A2(\asqrt[26] ), .ZN(new_n8508_));
  NAND3_X1   g08316(.A1(new_n8507_), .A2(new_n7166_), .A3(new_n8508_), .ZN(new_n8509_));
  AOI21_X1   g08317(.A1(new_n8507_), .A2(new_n8508_), .B(new_n7166_), .ZN(new_n8510_));
  AOI21_X1   g08318(.A1(new_n8509_), .A2(new_n8475_), .B(new_n8510_), .ZN(new_n8511_));
  AOI21_X1   g08319(.A1(new_n8511_), .A2(new_n6813_), .B(new_n8497_), .ZN(new_n8512_));
  OAI21_X1   g08320(.A1(new_n8511_), .A2(new_n6813_), .B(new_n6454_), .ZN(new_n8513_));
  OAI21_X1   g08321(.A1(new_n8512_), .A2(new_n8513_), .B(new_n8450_), .ZN(new_n8514_));
  NOR2_X1    g08322(.A1(new_n8511_), .A2(new_n6813_), .ZN(new_n8515_));
  OAI21_X1   g08323(.A1(new_n8512_), .A2(new_n8515_), .B(\asqrt[29] ), .ZN(new_n8516_));
  NAND3_X1   g08324(.A1(new_n8514_), .A2(new_n8516_), .A3(new_n6106_), .ZN(new_n8517_));
  NAND2_X1   g08325(.A1(new_n8517_), .A2(new_n8447_), .ZN(new_n8518_));
  NAND2_X1   g08326(.A1(new_n8514_), .A2(new_n8516_), .ZN(new_n8519_));
  AOI21_X1   g08327(.A1(new_n8519_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n8520_));
  AOI21_X1   g08328(.A1(new_n8520_), .A2(new_n8518_), .B(new_n8496_), .ZN(new_n8521_));
  AOI21_X1   g08329(.A1(new_n8518_), .A2(new_n8486_), .B(new_n5750_), .ZN(new_n8522_));
  OAI21_X1   g08330(.A1(new_n8521_), .A2(new_n8522_), .B(\asqrt[32] ), .ZN(new_n8523_));
  AOI21_X1   g08331(.A1(new_n8492_), .A2(new_n8523_), .B(new_n5110_), .ZN(new_n8524_));
  NOR2_X1    g08332(.A1(new_n8495_), .A2(new_n8524_), .ZN(new_n8525_));
  AOI21_X1   g08333(.A1(new_n8525_), .A2(new_n4810_), .B(new_n8436_), .ZN(new_n8526_));
  OAI21_X1   g08334(.A1(new_n8495_), .A2(new_n8524_), .B(\asqrt[34] ), .ZN(new_n8527_));
  NAND2_X1   g08335(.A1(new_n8527_), .A2(new_n4510_), .ZN(new_n8528_));
  OAI21_X1   g08336(.A1(new_n8526_), .A2(new_n8528_), .B(new_n8432_), .ZN(new_n8529_));
  INV_X1     g08337(.I(new_n8527_), .ZN(new_n8530_));
  OAI21_X1   g08338(.A1(new_n8526_), .A2(new_n8530_), .B(\asqrt[35] ), .ZN(new_n8531_));
  NAND3_X1   g08339(.A1(new_n8529_), .A2(new_n8531_), .A3(new_n4224_), .ZN(new_n8532_));
  NAND2_X1   g08340(.A1(new_n8532_), .A2(new_n8430_), .ZN(new_n8533_));
  NAND2_X1   g08341(.A1(new_n8529_), .A2(new_n8531_), .ZN(new_n8534_));
  AOI21_X1   g08342(.A1(new_n8534_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n8535_));
  AOI21_X1   g08343(.A1(new_n8535_), .A2(new_n8533_), .B(new_n8427_), .ZN(new_n8536_));
  INV_X1     g08344(.I(new_n8432_), .ZN(new_n8537_));
  INV_X1     g08345(.I(new_n8442_), .ZN(new_n8538_));
  NOR2_X1    g08346(.A1(new_n8521_), .A2(new_n8522_), .ZN(new_n8539_));
  AOI21_X1   g08347(.A1(new_n8539_), .A2(new_n5435_), .B(new_n8538_), .ZN(new_n8540_));
  NAND2_X1   g08348(.A1(new_n8523_), .A2(new_n5110_), .ZN(new_n8541_));
  OAI21_X1   g08349(.A1(new_n8540_), .A2(new_n8541_), .B(new_n8438_), .ZN(new_n8542_));
  INV_X1     g08350(.I(new_n8523_), .ZN(new_n8543_));
  OAI21_X1   g08351(.A1(new_n8540_), .A2(new_n8543_), .B(\asqrt[33] ), .ZN(new_n8544_));
  NAND3_X1   g08352(.A1(new_n8542_), .A2(new_n8544_), .A3(new_n4810_), .ZN(new_n8545_));
  NAND2_X1   g08353(.A1(new_n8545_), .A2(new_n8435_), .ZN(new_n8546_));
  NAND2_X1   g08354(.A1(new_n8542_), .A2(new_n8544_), .ZN(new_n8547_));
  AOI21_X1   g08355(.A1(new_n8547_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n8548_));
  AOI21_X1   g08356(.A1(new_n8548_), .A2(new_n8546_), .B(new_n8537_), .ZN(new_n8549_));
  AOI21_X1   g08357(.A1(new_n8546_), .A2(new_n8527_), .B(new_n4510_), .ZN(new_n8550_));
  OAI21_X1   g08358(.A1(new_n8549_), .A2(new_n8550_), .B(\asqrt[36] ), .ZN(new_n8551_));
  AOI21_X1   g08359(.A1(new_n8533_), .A2(new_n8551_), .B(new_n3928_), .ZN(new_n8552_));
  NOR2_X1    g08360(.A1(new_n8536_), .A2(new_n8552_), .ZN(new_n8553_));
  AOI21_X1   g08361(.A1(new_n8553_), .A2(new_n3675_), .B(new_n8424_), .ZN(new_n8554_));
  OAI21_X1   g08362(.A1(new_n8536_), .A2(new_n8552_), .B(\asqrt[38] ), .ZN(new_n8555_));
  NAND2_X1   g08363(.A1(new_n8555_), .A2(new_n3400_), .ZN(new_n8556_));
  OAI21_X1   g08364(.A1(new_n8554_), .A2(new_n8556_), .B(new_n8420_), .ZN(new_n8557_));
  INV_X1     g08365(.I(new_n8555_), .ZN(new_n8558_));
  OAI21_X1   g08366(.A1(new_n8554_), .A2(new_n8558_), .B(\asqrt[39] ), .ZN(new_n8559_));
  NAND3_X1   g08367(.A1(new_n8557_), .A2(new_n8559_), .A3(new_n3167_), .ZN(new_n8560_));
  NAND2_X1   g08368(.A1(new_n8560_), .A2(new_n8418_), .ZN(new_n8561_));
  NAND2_X1   g08369(.A1(new_n8557_), .A2(new_n8559_), .ZN(new_n8562_));
  AOI21_X1   g08370(.A1(new_n8562_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n8563_));
  AOI21_X1   g08371(.A1(new_n8563_), .A2(new_n8561_), .B(new_n8415_), .ZN(new_n8564_));
  INV_X1     g08372(.I(new_n8420_), .ZN(new_n8565_));
  INV_X1     g08373(.I(new_n8430_), .ZN(new_n8566_));
  NOR2_X1    g08374(.A1(new_n8549_), .A2(new_n8550_), .ZN(new_n8567_));
  AOI21_X1   g08375(.A1(new_n8567_), .A2(new_n4224_), .B(new_n8566_), .ZN(new_n8568_));
  NAND2_X1   g08376(.A1(new_n8551_), .A2(new_n3928_), .ZN(new_n8569_));
  OAI21_X1   g08377(.A1(new_n8568_), .A2(new_n8569_), .B(new_n8426_), .ZN(new_n8570_));
  INV_X1     g08378(.I(new_n8551_), .ZN(new_n8571_));
  OAI21_X1   g08379(.A1(new_n8568_), .A2(new_n8571_), .B(\asqrt[37] ), .ZN(new_n8572_));
  NAND3_X1   g08380(.A1(new_n8570_), .A2(new_n8572_), .A3(new_n3675_), .ZN(new_n8573_));
  NAND2_X1   g08381(.A1(new_n8573_), .A2(new_n8423_), .ZN(new_n8574_));
  NAND2_X1   g08382(.A1(new_n8570_), .A2(new_n8572_), .ZN(new_n8575_));
  AOI21_X1   g08383(.A1(new_n8575_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n8576_));
  AOI21_X1   g08384(.A1(new_n8576_), .A2(new_n8574_), .B(new_n8565_), .ZN(new_n8577_));
  AOI21_X1   g08385(.A1(new_n8574_), .A2(new_n8555_), .B(new_n3400_), .ZN(new_n8578_));
  OAI21_X1   g08386(.A1(new_n8577_), .A2(new_n8578_), .B(\asqrt[40] ), .ZN(new_n8579_));
  AOI21_X1   g08387(.A1(new_n8561_), .A2(new_n8579_), .B(new_n2912_), .ZN(new_n8580_));
  NOR2_X1    g08388(.A1(new_n8564_), .A2(new_n8580_), .ZN(new_n8581_));
  AOI21_X1   g08389(.A1(new_n8581_), .A2(new_n2699_), .B(new_n8414_), .ZN(new_n8582_));
  OAI21_X1   g08390(.A1(new_n8564_), .A2(new_n8580_), .B(\asqrt[42] ), .ZN(new_n8583_));
  NAND2_X1   g08391(.A1(new_n8583_), .A2(new_n2464_), .ZN(new_n8584_));
  OAI21_X1   g08392(.A1(new_n8582_), .A2(new_n8584_), .B(new_n8410_), .ZN(new_n8585_));
  INV_X1     g08393(.I(new_n8583_), .ZN(new_n8586_));
  OAI21_X1   g08394(.A1(new_n8582_), .A2(new_n8586_), .B(\asqrt[43] ), .ZN(new_n8587_));
  NAND3_X1   g08395(.A1(new_n8585_), .A2(new_n8587_), .A3(new_n2271_), .ZN(new_n8588_));
  NAND2_X1   g08396(.A1(new_n8588_), .A2(new_n8408_), .ZN(new_n8589_));
  NAND2_X1   g08397(.A1(new_n8585_), .A2(new_n8587_), .ZN(new_n8590_));
  AOI21_X1   g08398(.A1(new_n8590_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n8591_));
  AOI21_X1   g08399(.A1(new_n8591_), .A2(new_n8589_), .B(new_n8405_), .ZN(new_n8592_));
  INV_X1     g08400(.I(new_n8410_), .ZN(new_n8593_));
  INV_X1     g08401(.I(new_n8418_), .ZN(new_n8594_));
  NOR2_X1    g08402(.A1(new_n8577_), .A2(new_n8578_), .ZN(new_n8595_));
  AOI21_X1   g08403(.A1(new_n8595_), .A2(new_n3167_), .B(new_n8594_), .ZN(new_n8596_));
  NAND2_X1   g08404(.A1(new_n8579_), .A2(new_n2912_), .ZN(new_n8597_));
  OAI21_X1   g08405(.A1(new_n8596_), .A2(new_n8597_), .B(new_n8332_), .ZN(new_n8598_));
  INV_X1     g08406(.I(new_n8579_), .ZN(new_n8599_));
  OAI21_X1   g08407(.A1(new_n8596_), .A2(new_n8599_), .B(\asqrt[41] ), .ZN(new_n8600_));
  NAND3_X1   g08408(.A1(new_n8598_), .A2(new_n8600_), .A3(new_n2699_), .ZN(new_n8601_));
  NAND2_X1   g08409(.A1(new_n8601_), .A2(new_n8413_), .ZN(new_n8602_));
  NAND2_X1   g08410(.A1(new_n8598_), .A2(new_n8600_), .ZN(new_n8603_));
  AOI21_X1   g08411(.A1(new_n8603_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n8604_));
  AOI21_X1   g08412(.A1(new_n8604_), .A2(new_n8602_), .B(new_n8593_), .ZN(new_n8605_));
  AOI21_X1   g08413(.A1(new_n8602_), .A2(new_n8583_), .B(new_n2464_), .ZN(new_n8606_));
  OAI21_X1   g08414(.A1(new_n8605_), .A2(new_n8606_), .B(\asqrt[44] ), .ZN(new_n8607_));
  AOI21_X1   g08415(.A1(new_n8589_), .A2(new_n8607_), .B(new_n2072_), .ZN(new_n8608_));
  NOR2_X1    g08416(.A1(new_n8592_), .A2(new_n8608_), .ZN(new_n8609_));
  AOI21_X1   g08417(.A1(new_n8609_), .A2(new_n1884_), .B(new_n8402_), .ZN(new_n8610_));
  OAI21_X1   g08418(.A1(new_n8592_), .A2(new_n8608_), .B(\asqrt[46] ), .ZN(new_n8611_));
  NAND2_X1   g08419(.A1(new_n8611_), .A2(new_n1688_), .ZN(new_n8612_));
  OAI21_X1   g08420(.A1(new_n8610_), .A2(new_n8612_), .B(new_n8398_), .ZN(new_n8613_));
  INV_X1     g08421(.I(new_n8611_), .ZN(new_n8614_));
  OAI21_X1   g08422(.A1(new_n8610_), .A2(new_n8614_), .B(\asqrt[47] ), .ZN(new_n8615_));
  NAND3_X1   g08423(.A1(new_n8613_), .A2(new_n8615_), .A3(new_n1533_), .ZN(new_n8616_));
  NAND2_X1   g08424(.A1(new_n8616_), .A2(new_n8396_), .ZN(new_n8617_));
  NAND2_X1   g08425(.A1(new_n8613_), .A2(new_n8615_), .ZN(new_n8618_));
  AOI21_X1   g08426(.A1(new_n8618_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n8619_));
  AOI21_X1   g08427(.A1(new_n8619_), .A2(new_n8617_), .B(new_n8393_), .ZN(new_n8620_));
  INV_X1     g08428(.I(new_n8398_), .ZN(new_n8621_));
  INV_X1     g08429(.I(new_n8408_), .ZN(new_n8622_));
  NOR2_X1    g08430(.A1(new_n8605_), .A2(new_n8606_), .ZN(new_n8623_));
  AOI21_X1   g08431(.A1(new_n8623_), .A2(new_n2271_), .B(new_n8622_), .ZN(new_n8624_));
  NAND2_X1   g08432(.A1(new_n8607_), .A2(new_n2072_), .ZN(new_n8625_));
  OAI21_X1   g08433(.A1(new_n8624_), .A2(new_n8625_), .B(new_n8404_), .ZN(new_n8626_));
  INV_X1     g08434(.I(new_n8607_), .ZN(new_n8627_));
  OAI21_X1   g08435(.A1(new_n8624_), .A2(new_n8627_), .B(\asqrt[45] ), .ZN(new_n8628_));
  NAND3_X1   g08436(.A1(new_n8626_), .A2(new_n8628_), .A3(new_n1884_), .ZN(new_n8629_));
  NAND2_X1   g08437(.A1(new_n8629_), .A2(new_n8401_), .ZN(new_n8630_));
  NAND2_X1   g08438(.A1(new_n8626_), .A2(new_n8628_), .ZN(new_n8631_));
  AOI21_X1   g08439(.A1(new_n8631_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n8632_));
  AOI21_X1   g08440(.A1(new_n8632_), .A2(new_n8630_), .B(new_n8621_), .ZN(new_n8633_));
  AOI21_X1   g08441(.A1(new_n8630_), .A2(new_n8611_), .B(new_n1688_), .ZN(new_n8634_));
  OAI21_X1   g08442(.A1(new_n8633_), .A2(new_n8634_), .B(\asqrt[48] ), .ZN(new_n8635_));
  AOI21_X1   g08443(.A1(new_n8617_), .A2(new_n8635_), .B(new_n1368_), .ZN(new_n8636_));
  NOR2_X1    g08444(.A1(new_n8620_), .A2(new_n8636_), .ZN(new_n8637_));
  AOI21_X1   g08445(.A1(new_n8637_), .A2(new_n1228_), .B(new_n8390_), .ZN(new_n8638_));
  OAI21_X1   g08446(.A1(new_n8620_), .A2(new_n8636_), .B(\asqrt[50] ), .ZN(new_n8639_));
  NAND2_X1   g08447(.A1(new_n8639_), .A2(new_n1088_), .ZN(new_n8640_));
  OAI21_X1   g08448(.A1(new_n8638_), .A2(new_n8640_), .B(new_n8386_), .ZN(new_n8641_));
  INV_X1     g08449(.I(new_n8639_), .ZN(new_n8642_));
  OAI21_X1   g08450(.A1(new_n8638_), .A2(new_n8642_), .B(\asqrt[51] ), .ZN(new_n8643_));
  NAND3_X1   g08451(.A1(new_n8641_), .A2(new_n8643_), .A3(new_n962_), .ZN(new_n8644_));
  NAND2_X1   g08452(.A1(new_n8644_), .A2(new_n8384_), .ZN(new_n8645_));
  NAND2_X1   g08453(.A1(new_n8641_), .A2(new_n8643_), .ZN(new_n8646_));
  AOI21_X1   g08454(.A1(new_n8646_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n8647_));
  AOI21_X1   g08455(.A1(new_n8647_), .A2(new_n8645_), .B(new_n8381_), .ZN(new_n8648_));
  INV_X1     g08456(.I(new_n8386_), .ZN(new_n8649_));
  INV_X1     g08457(.I(new_n8396_), .ZN(new_n8650_));
  NOR2_X1    g08458(.A1(new_n8633_), .A2(new_n8634_), .ZN(new_n8651_));
  AOI21_X1   g08459(.A1(new_n8651_), .A2(new_n1533_), .B(new_n8650_), .ZN(new_n8652_));
  NAND2_X1   g08460(.A1(new_n8635_), .A2(new_n1368_), .ZN(new_n8653_));
  OAI21_X1   g08461(.A1(new_n8652_), .A2(new_n8653_), .B(new_n8392_), .ZN(new_n8654_));
  INV_X1     g08462(.I(new_n8635_), .ZN(new_n8655_));
  OAI21_X1   g08463(.A1(new_n8652_), .A2(new_n8655_), .B(\asqrt[49] ), .ZN(new_n8656_));
  NAND3_X1   g08464(.A1(new_n8654_), .A2(new_n8656_), .A3(new_n1228_), .ZN(new_n8657_));
  NAND2_X1   g08465(.A1(new_n8657_), .A2(new_n8389_), .ZN(new_n8658_));
  NAND2_X1   g08466(.A1(new_n8654_), .A2(new_n8656_), .ZN(new_n8659_));
  AOI21_X1   g08467(.A1(new_n8659_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n8660_));
  AOI21_X1   g08468(.A1(new_n8660_), .A2(new_n8658_), .B(new_n8649_), .ZN(new_n8661_));
  AOI21_X1   g08469(.A1(new_n8658_), .A2(new_n8639_), .B(new_n1088_), .ZN(new_n8662_));
  OAI21_X1   g08470(.A1(new_n8661_), .A2(new_n8662_), .B(\asqrt[52] ), .ZN(new_n8663_));
  AOI21_X1   g08471(.A1(new_n8645_), .A2(new_n8663_), .B(new_n842_), .ZN(new_n8664_));
  NOR2_X1    g08472(.A1(new_n8648_), .A2(new_n8664_), .ZN(new_n8665_));
  AOI21_X1   g08473(.A1(new_n8665_), .A2(new_n720_), .B(new_n8378_), .ZN(new_n8666_));
  OAI21_X1   g08474(.A1(new_n8648_), .A2(new_n8664_), .B(\asqrt[54] ), .ZN(new_n8667_));
  NAND2_X1   g08475(.A1(new_n8667_), .A2(new_n630_), .ZN(new_n8668_));
  OAI21_X1   g08476(.A1(new_n8666_), .A2(new_n8668_), .B(new_n8374_), .ZN(new_n8669_));
  INV_X1     g08477(.I(new_n8667_), .ZN(new_n8670_));
  OAI21_X1   g08478(.A1(new_n8666_), .A2(new_n8670_), .B(\asqrt[55] ), .ZN(new_n8671_));
  NAND3_X1   g08479(.A1(new_n8669_), .A2(new_n8671_), .A3(new_n545_), .ZN(new_n8672_));
  NAND2_X1   g08480(.A1(new_n8672_), .A2(new_n8372_), .ZN(new_n8673_));
  NAND2_X1   g08481(.A1(new_n8669_), .A2(new_n8671_), .ZN(new_n8674_));
  AOI21_X1   g08482(.A1(new_n8674_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n8675_));
  AOI21_X1   g08483(.A1(new_n8675_), .A2(new_n8673_), .B(new_n8369_), .ZN(new_n8676_));
  INV_X1     g08484(.I(new_n8374_), .ZN(new_n8677_));
  INV_X1     g08485(.I(new_n8384_), .ZN(new_n8678_));
  NOR2_X1    g08486(.A1(new_n8661_), .A2(new_n8662_), .ZN(new_n8679_));
  AOI21_X1   g08487(.A1(new_n8679_), .A2(new_n962_), .B(new_n8678_), .ZN(new_n8680_));
  NAND2_X1   g08488(.A1(new_n8663_), .A2(new_n842_), .ZN(new_n8681_));
  OAI21_X1   g08489(.A1(new_n8680_), .A2(new_n8681_), .B(new_n8380_), .ZN(new_n8682_));
  INV_X1     g08490(.I(new_n8663_), .ZN(new_n8683_));
  OAI21_X1   g08491(.A1(new_n8680_), .A2(new_n8683_), .B(\asqrt[53] ), .ZN(new_n8684_));
  NAND3_X1   g08492(.A1(new_n8682_), .A2(new_n8684_), .A3(new_n720_), .ZN(new_n8685_));
  NAND2_X1   g08493(.A1(new_n8685_), .A2(new_n8377_), .ZN(new_n8686_));
  NAND2_X1   g08494(.A1(new_n8682_), .A2(new_n8684_), .ZN(new_n8687_));
  AOI21_X1   g08495(.A1(new_n8687_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n8688_));
  AOI21_X1   g08496(.A1(new_n8688_), .A2(new_n8686_), .B(new_n8677_), .ZN(new_n8689_));
  AOI21_X1   g08497(.A1(new_n8686_), .A2(new_n8667_), .B(new_n630_), .ZN(new_n8690_));
  OAI21_X1   g08498(.A1(new_n8689_), .A2(new_n8690_), .B(\asqrt[56] ), .ZN(new_n8691_));
  AOI21_X1   g08499(.A1(new_n8673_), .A2(new_n8691_), .B(new_n450_), .ZN(new_n8692_));
  NOR2_X1    g08500(.A1(new_n8676_), .A2(new_n8692_), .ZN(new_n8693_));
  AOI21_X1   g08501(.A1(new_n8693_), .A2(new_n403_), .B(new_n8366_), .ZN(new_n8694_));
  OAI21_X1   g08502(.A1(new_n8676_), .A2(new_n8692_), .B(\asqrt[58] ), .ZN(new_n8695_));
  NAND2_X1   g08503(.A1(new_n8695_), .A2(new_n339_), .ZN(new_n8696_));
  OAI21_X1   g08504(.A1(new_n8694_), .A2(new_n8696_), .B(new_n8362_), .ZN(new_n8697_));
  INV_X1     g08505(.I(new_n8695_), .ZN(new_n8698_));
  OAI21_X1   g08506(.A1(new_n8694_), .A2(new_n8698_), .B(\asqrt[59] ), .ZN(new_n8699_));
  NAND3_X1   g08507(.A1(new_n8697_), .A2(new_n8699_), .A3(new_n288_), .ZN(new_n8700_));
  NAND2_X1   g08508(.A1(new_n8700_), .A2(new_n8360_), .ZN(new_n8701_));
  INV_X1     g08509(.I(new_n8362_), .ZN(new_n8702_));
  INV_X1     g08510(.I(new_n8372_), .ZN(new_n8703_));
  NOR2_X1    g08511(.A1(new_n8689_), .A2(new_n8690_), .ZN(new_n8704_));
  AOI21_X1   g08512(.A1(new_n8704_), .A2(new_n545_), .B(new_n8703_), .ZN(new_n8705_));
  NAND2_X1   g08513(.A1(new_n8691_), .A2(new_n450_), .ZN(new_n8706_));
  OAI21_X1   g08514(.A1(new_n8705_), .A2(new_n8706_), .B(new_n8368_), .ZN(new_n8707_));
  INV_X1     g08515(.I(new_n8691_), .ZN(new_n8708_));
  OAI21_X1   g08516(.A1(new_n8705_), .A2(new_n8708_), .B(\asqrt[57] ), .ZN(new_n8709_));
  NAND3_X1   g08517(.A1(new_n8707_), .A2(new_n8709_), .A3(new_n403_), .ZN(new_n8710_));
  NAND2_X1   g08518(.A1(new_n8710_), .A2(new_n8365_), .ZN(new_n8711_));
  NAND2_X1   g08519(.A1(new_n8707_), .A2(new_n8709_), .ZN(new_n8712_));
  AOI21_X1   g08520(.A1(new_n8712_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n8713_));
  AOI21_X1   g08521(.A1(new_n8713_), .A2(new_n8711_), .B(new_n8702_), .ZN(new_n8714_));
  AOI21_X1   g08522(.A1(new_n8711_), .A2(new_n8695_), .B(new_n339_), .ZN(new_n8715_));
  OAI21_X1   g08523(.A1(new_n8714_), .A2(new_n8715_), .B(\asqrt[60] ), .ZN(new_n8716_));
  AOI21_X1   g08524(.A1(new_n8701_), .A2(new_n8716_), .B(new_n242_), .ZN(new_n8717_));
  NAND3_X1   g08525(.A1(\asqrt[24] ), .A2(new_n8292_), .A3(new_n8308_), .ZN(new_n8718_));
  XOR2_X1    g08526(.A1(new_n8718_), .A2(new_n8333_), .Z(new_n8719_));
  INV_X1     g08527(.I(new_n8719_), .ZN(new_n8720_));
  NAND2_X1   g08528(.A1(new_n8697_), .A2(new_n8699_), .ZN(new_n8721_));
  AOI21_X1   g08529(.A1(new_n8721_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n8722_));
  AOI21_X1   g08530(.A1(new_n8722_), .A2(new_n8701_), .B(new_n8720_), .ZN(new_n8723_));
  OAI21_X1   g08531(.A1(new_n8723_), .A2(new_n8717_), .B(\asqrt[62] ), .ZN(new_n8724_));
  AOI21_X1   g08532(.A1(new_n8293_), .A2(new_n8314_), .B(new_n8309_), .ZN(new_n8725_));
  NAND2_X1   g08533(.A1(\asqrt[24] ), .A2(new_n8725_), .ZN(new_n8726_));
  XOR2_X1    g08534(.A1(new_n8726_), .A2(new_n8312_), .Z(new_n8727_));
  INV_X1     g08535(.I(new_n8360_), .ZN(new_n8728_));
  NOR2_X1    g08536(.A1(new_n8714_), .A2(new_n8715_), .ZN(new_n8729_));
  AOI21_X1   g08537(.A1(new_n8729_), .A2(new_n288_), .B(new_n8728_), .ZN(new_n8730_));
  INV_X1     g08538(.I(new_n8716_), .ZN(new_n8731_));
  OAI21_X1   g08539(.A1(new_n8730_), .A2(new_n8731_), .B(\asqrt[61] ), .ZN(new_n8732_));
  NAND2_X1   g08540(.A1(new_n8716_), .A2(new_n242_), .ZN(new_n8733_));
  OAI21_X1   g08541(.A1(new_n8730_), .A2(new_n8733_), .B(new_n8719_), .ZN(new_n8734_));
  NAND3_X1   g08542(.A1(new_n8734_), .A2(new_n8732_), .A3(new_n234_), .ZN(new_n8735_));
  NAND2_X1   g08543(.A1(new_n8735_), .A2(new_n8727_), .ZN(new_n8736_));
  AOI21_X1   g08544(.A1(new_n8736_), .A2(new_n8724_), .B(new_n8357_), .ZN(new_n8737_));
  AOI21_X1   g08545(.A1(new_n8737_), .A2(new_n8355_), .B(\asqrt[63] ), .ZN(new_n8738_));
  NAND2_X1   g08546(.A1(new_n8736_), .A2(new_n8724_), .ZN(new_n8739_));
  NOR2_X1    g08547(.A1(new_n8739_), .A2(new_n8355_), .ZN(new_n8740_));
  NOR2_X1    g08548(.A1(\asqrt[24] ), .A2(new_n8344_), .ZN(new_n8741_));
  NOR4_X1    g08549(.A1(new_n8738_), .A2(new_n8352_), .A3(new_n8740_), .A4(new_n8741_), .ZN(new_n8742_));
  OAI21_X1   g08550(.A1(new_n8596_), .A2(new_n8597_), .B(new_n8600_), .ZN(new_n8743_));
  NOR2_X1    g08551(.A1(new_n8742_), .A2(new_n8743_), .ZN(new_n8744_));
  XOR2_X1    g08552(.A1(new_n8744_), .A2(new_n8332_), .Z(new_n8745_));
  INV_X1     g08553(.I(new_n8745_), .ZN(new_n8746_));
  INV_X1     g08554(.I(new_n8352_), .ZN(new_n8747_));
  INV_X1     g08555(.I(new_n8724_), .ZN(new_n8748_));
  NOR2_X1    g08556(.A1(new_n8723_), .A2(new_n8717_), .ZN(new_n8749_));
  INV_X1     g08557(.I(new_n8727_), .ZN(new_n8750_));
  AOI21_X1   g08558(.A1(new_n8749_), .A2(new_n234_), .B(new_n8750_), .ZN(new_n8751_));
  OAI21_X1   g08559(.A1(new_n8751_), .A2(new_n8748_), .B(new_n8356_), .ZN(new_n8752_));
  OAI21_X1   g08560(.A1(new_n8752_), .A2(new_n8354_), .B(new_n193_), .ZN(new_n8753_));
  NOR2_X1    g08561(.A1(new_n8751_), .A2(new_n8748_), .ZN(new_n8754_));
  NAND2_X1   g08562(.A1(new_n8754_), .A2(new_n8354_), .ZN(new_n8755_));
  INV_X1     g08563(.I(new_n8741_), .ZN(new_n8756_));
  NAND4_X1   g08564(.A1(new_n8753_), .A2(new_n8747_), .A3(new_n8755_), .A4(new_n8756_), .ZN(\asqrt[23] ));
  NAND3_X1   g08565(.A1(\asqrt[23] ), .A2(new_n8560_), .A3(new_n8579_), .ZN(new_n8758_));
  XOR2_X1    g08566(.A1(new_n8758_), .A2(new_n8594_), .Z(new_n8759_));
  OAI21_X1   g08567(.A1(new_n8554_), .A2(new_n8556_), .B(new_n8559_), .ZN(new_n8760_));
  NOR2_X1    g08568(.A1(new_n8742_), .A2(new_n8760_), .ZN(new_n8761_));
  XOR2_X1    g08569(.A1(new_n8761_), .A2(new_n8420_), .Z(new_n8762_));
  INV_X1     g08570(.I(new_n8762_), .ZN(new_n8763_));
  NAND3_X1   g08571(.A1(\asqrt[23] ), .A2(new_n8573_), .A3(new_n8555_), .ZN(new_n8764_));
  XOR2_X1    g08572(.A1(new_n8764_), .A2(new_n8424_), .Z(new_n8765_));
  INV_X1     g08573(.I(new_n8765_), .ZN(new_n8766_));
  OAI21_X1   g08574(.A1(new_n8568_), .A2(new_n8569_), .B(new_n8572_), .ZN(new_n8767_));
  NOR2_X1    g08575(.A1(new_n8742_), .A2(new_n8767_), .ZN(new_n8768_));
  XOR2_X1    g08576(.A1(new_n8768_), .A2(new_n8426_), .Z(new_n8769_));
  NAND3_X1   g08577(.A1(\asqrt[23] ), .A2(new_n8532_), .A3(new_n8551_), .ZN(new_n8770_));
  XOR2_X1    g08578(.A1(new_n8770_), .A2(new_n8566_), .Z(new_n8771_));
  OAI21_X1   g08579(.A1(new_n8526_), .A2(new_n8528_), .B(new_n8531_), .ZN(new_n8772_));
  NOR2_X1    g08580(.A1(new_n8742_), .A2(new_n8772_), .ZN(new_n8773_));
  XOR2_X1    g08581(.A1(new_n8773_), .A2(new_n8432_), .Z(new_n8774_));
  INV_X1     g08582(.I(new_n8774_), .ZN(new_n8775_));
  NAND3_X1   g08583(.A1(\asqrt[23] ), .A2(new_n8545_), .A3(new_n8527_), .ZN(new_n8776_));
  XOR2_X1    g08584(.A1(new_n8776_), .A2(new_n8436_), .Z(new_n8777_));
  INV_X1     g08585(.I(new_n8777_), .ZN(new_n8778_));
  OAI21_X1   g08586(.A1(new_n8540_), .A2(new_n8541_), .B(new_n8544_), .ZN(new_n8779_));
  NOR2_X1    g08587(.A1(new_n8742_), .A2(new_n8779_), .ZN(new_n8780_));
  XOR2_X1    g08588(.A1(new_n8780_), .A2(new_n8438_), .Z(new_n8781_));
  NAND3_X1   g08589(.A1(\asqrt[23] ), .A2(new_n8491_), .A3(new_n8523_), .ZN(new_n8782_));
  XOR2_X1    g08590(.A1(new_n8782_), .A2(new_n8538_), .Z(new_n8783_));
  OAI21_X1   g08591(.A1(new_n8485_), .A2(new_n8487_), .B(new_n8490_), .ZN(new_n8784_));
  NOR2_X1    g08592(.A1(new_n8742_), .A2(new_n8784_), .ZN(new_n8785_));
  XOR2_X1    g08593(.A1(new_n8785_), .A2(new_n8444_), .Z(new_n8786_));
  INV_X1     g08594(.I(new_n8786_), .ZN(new_n8787_));
  NAND3_X1   g08595(.A1(\asqrt[23] ), .A2(new_n8517_), .A3(new_n8486_), .ZN(new_n8788_));
  XOR2_X1    g08596(.A1(new_n8788_), .A2(new_n8448_), .Z(new_n8789_));
  INV_X1     g08597(.I(new_n8789_), .ZN(new_n8790_));
  AOI21_X1   g08598(.A1(new_n8479_), .A2(new_n8480_), .B(new_n8483_), .ZN(new_n8791_));
  NAND2_X1   g08599(.A1(\asqrt[23] ), .A2(new_n8791_), .ZN(new_n8792_));
  XOR2_X1    g08600(.A1(new_n8792_), .A2(new_n8451_), .Z(new_n8793_));
  NOR2_X1    g08601(.A1(new_n8478_), .A2(\asqrt[28] ), .ZN(new_n8794_));
  NOR3_X1    g08602(.A1(new_n8742_), .A2(new_n8794_), .A3(new_n8515_), .ZN(new_n8795_));
  XOR2_X1    g08603(.A1(new_n8795_), .A2(new_n8454_), .Z(new_n8796_));
  NOR3_X1    g08604(.A1(new_n8742_), .A2(new_n8473_), .A3(new_n8510_), .ZN(new_n8797_));
  XOR2_X1    g08605(.A1(new_n8797_), .A2(new_n8475_), .Z(new_n8798_));
  INV_X1     g08606(.I(new_n8798_), .ZN(new_n8799_));
  NOR2_X1    g08607(.A1(new_n8506_), .A2(\asqrt[26] ), .ZN(new_n8800_));
  NOR3_X1    g08608(.A1(new_n8742_), .A2(new_n8800_), .A3(new_n8472_), .ZN(new_n8801_));
  XOR2_X1    g08609(.A1(new_n8801_), .A2(new_n8500_), .Z(new_n8802_));
  INV_X1     g08610(.I(new_n8802_), .ZN(new_n8803_));
  NAND3_X1   g08611(.A1(\asqrt[23] ), .A2(new_n8462_), .A3(new_n8463_), .ZN(new_n8804_));
  NAND4_X1   g08612(.A1(new_n8753_), .A2(\asqrt[24] ), .A3(new_n8755_), .A4(new_n8747_), .ZN(new_n8805_));
  AOI21_X1   g08613(.A1(new_n8804_), .A2(new_n8805_), .B(\a[48] ), .ZN(new_n8806_));
  NOR3_X1    g08614(.A1(new_n8742_), .A2(\a[46] ), .A3(\a[47] ), .ZN(new_n8807_));
  INV_X1     g08615(.I(new_n8805_), .ZN(new_n8808_));
  NOR3_X1    g08616(.A1(new_n8807_), .A2(new_n7991_), .A3(new_n8808_), .ZN(new_n8809_));
  NOR2_X1    g08617(.A1(new_n8809_), .A2(new_n8806_), .ZN(new_n8810_));
  INV_X1     g08618(.I(\a[44] ), .ZN(new_n8811_));
  INV_X1     g08619(.I(\a[45] ), .ZN(new_n8812_));
  NAND3_X1   g08620(.A1(new_n8811_), .A2(new_n8812_), .A3(new_n8462_), .ZN(new_n8813_));
  OAI21_X1   g08621(.A1(new_n8742_), .A2(new_n8462_), .B(new_n8813_), .ZN(new_n8814_));
  NAND2_X1   g08622(.A1(new_n8814_), .A2(\asqrt[24] ), .ZN(new_n8815_));
  OAI21_X1   g08623(.A1(new_n8742_), .A2(\a[46] ), .B(\a[47] ), .ZN(new_n8816_));
  NAND2_X1   g08624(.A1(new_n8816_), .A2(new_n8804_), .ZN(new_n8817_));
  NOR2_X1    g08625(.A1(new_n8814_), .A2(\asqrt[24] ), .ZN(new_n8818_));
  OAI21_X1   g08626(.A1(new_n8817_), .A2(new_n8818_), .B(new_n8815_), .ZN(new_n8819_));
  OAI21_X1   g08627(.A1(new_n8819_), .A2(\asqrt[25] ), .B(new_n8810_), .ZN(new_n8820_));
  NAND2_X1   g08628(.A1(new_n8819_), .A2(\asqrt[25] ), .ZN(new_n8821_));
  NAND3_X1   g08629(.A1(new_n8820_), .A2(new_n7561_), .A3(new_n8821_), .ZN(new_n8822_));
  NOR3_X1    g08630(.A1(new_n8742_), .A2(new_n8466_), .A3(new_n8505_), .ZN(new_n8823_));
  XOR2_X1    g08631(.A1(new_n8823_), .A2(new_n8468_), .Z(new_n8824_));
  NAND2_X1   g08632(.A1(new_n8822_), .A2(new_n8824_), .ZN(new_n8825_));
  NAND2_X1   g08633(.A1(new_n8820_), .A2(new_n8821_), .ZN(new_n8826_));
  AOI21_X1   g08634(.A1(new_n8826_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n8827_));
  AOI21_X1   g08635(.A1(new_n8827_), .A2(new_n8825_), .B(new_n8803_), .ZN(new_n8828_));
  OAI21_X1   g08636(.A1(new_n8807_), .A2(new_n8808_), .B(new_n7991_), .ZN(new_n8829_));
  NAND3_X1   g08637(.A1(new_n8804_), .A2(\a[48] ), .A3(new_n8805_), .ZN(new_n8830_));
  NAND2_X1   g08638(.A1(new_n8829_), .A2(new_n8830_), .ZN(new_n8831_));
  NAND2_X1   g08639(.A1(\asqrt[23] ), .A2(\a[46] ), .ZN(new_n8832_));
  AOI21_X1   g08640(.A1(new_n8832_), .A2(new_n8813_), .B(new_n8349_), .ZN(new_n8833_));
  AOI21_X1   g08641(.A1(\asqrt[23] ), .A2(new_n8462_), .B(new_n8463_), .ZN(new_n8834_));
  NOR2_X1    g08642(.A1(new_n8807_), .A2(new_n8834_), .ZN(new_n8835_));
  NAND3_X1   g08643(.A1(new_n8832_), .A2(new_n8349_), .A3(new_n8813_), .ZN(new_n8836_));
  AOI21_X1   g08644(.A1(new_n8835_), .A2(new_n8836_), .B(new_n8833_), .ZN(new_n8837_));
  AOI21_X1   g08645(.A1(new_n8837_), .A2(new_n7934_), .B(new_n8831_), .ZN(new_n8838_));
  NOR2_X1    g08646(.A1(new_n8837_), .A2(new_n7934_), .ZN(new_n8839_));
  OAI21_X1   g08647(.A1(new_n8838_), .A2(new_n8839_), .B(\asqrt[26] ), .ZN(new_n8840_));
  AOI21_X1   g08648(.A1(new_n8825_), .A2(new_n8840_), .B(new_n7166_), .ZN(new_n8841_));
  NOR2_X1    g08649(.A1(new_n8828_), .A2(new_n8841_), .ZN(new_n8842_));
  AOI21_X1   g08650(.A1(new_n8842_), .A2(new_n6813_), .B(new_n8799_), .ZN(new_n8843_));
  OAI21_X1   g08651(.A1(new_n8828_), .A2(new_n8841_), .B(\asqrt[28] ), .ZN(new_n8844_));
  NAND2_X1   g08652(.A1(new_n8844_), .A2(new_n6454_), .ZN(new_n8845_));
  OAI21_X1   g08653(.A1(new_n8843_), .A2(new_n8845_), .B(new_n8796_), .ZN(new_n8846_));
  INV_X1     g08654(.I(new_n8844_), .ZN(new_n8847_));
  OAI21_X1   g08655(.A1(new_n8843_), .A2(new_n8847_), .B(\asqrt[29] ), .ZN(new_n8848_));
  NAND3_X1   g08656(.A1(new_n8846_), .A2(new_n8848_), .A3(new_n6106_), .ZN(new_n8849_));
  NAND2_X1   g08657(.A1(new_n8849_), .A2(new_n8793_), .ZN(new_n8850_));
  NAND2_X1   g08658(.A1(new_n8846_), .A2(new_n8848_), .ZN(new_n8851_));
  AOI21_X1   g08659(.A1(new_n8851_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n8852_));
  AOI21_X1   g08660(.A1(new_n8852_), .A2(new_n8850_), .B(new_n8790_), .ZN(new_n8853_));
  INV_X1     g08661(.I(new_n8796_), .ZN(new_n8854_));
  NOR2_X1    g08662(.A1(new_n8838_), .A2(new_n8839_), .ZN(new_n8855_));
  INV_X1     g08663(.I(new_n8824_), .ZN(new_n8856_));
  AOI21_X1   g08664(.A1(new_n8855_), .A2(new_n7561_), .B(new_n8856_), .ZN(new_n8857_));
  NAND2_X1   g08665(.A1(new_n8840_), .A2(new_n7166_), .ZN(new_n8858_));
  OAI21_X1   g08666(.A1(new_n8857_), .A2(new_n8858_), .B(new_n8802_), .ZN(new_n8859_));
  INV_X1     g08667(.I(new_n8840_), .ZN(new_n8860_));
  OAI21_X1   g08668(.A1(new_n8857_), .A2(new_n8860_), .B(\asqrt[27] ), .ZN(new_n8861_));
  NAND3_X1   g08669(.A1(new_n8859_), .A2(new_n8861_), .A3(new_n6813_), .ZN(new_n8862_));
  NAND2_X1   g08670(.A1(new_n8862_), .A2(new_n8798_), .ZN(new_n8863_));
  NAND2_X1   g08671(.A1(new_n8859_), .A2(new_n8861_), .ZN(new_n8864_));
  AOI21_X1   g08672(.A1(new_n8864_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n8865_));
  AOI21_X1   g08673(.A1(new_n8865_), .A2(new_n8863_), .B(new_n8854_), .ZN(new_n8866_));
  AOI21_X1   g08674(.A1(new_n8863_), .A2(new_n8844_), .B(new_n6454_), .ZN(new_n8867_));
  OAI21_X1   g08675(.A1(new_n8866_), .A2(new_n8867_), .B(\asqrt[30] ), .ZN(new_n8868_));
  AOI21_X1   g08676(.A1(new_n8850_), .A2(new_n8868_), .B(new_n5750_), .ZN(new_n8869_));
  NOR2_X1    g08677(.A1(new_n8853_), .A2(new_n8869_), .ZN(new_n8870_));
  AOI21_X1   g08678(.A1(new_n8870_), .A2(new_n5435_), .B(new_n8787_), .ZN(new_n8871_));
  OAI21_X1   g08679(.A1(new_n8853_), .A2(new_n8869_), .B(\asqrt[32] ), .ZN(new_n8872_));
  NAND2_X1   g08680(.A1(new_n8872_), .A2(new_n5110_), .ZN(new_n8873_));
  OAI21_X1   g08681(.A1(new_n8871_), .A2(new_n8873_), .B(new_n8783_), .ZN(new_n8874_));
  INV_X1     g08682(.I(new_n8872_), .ZN(new_n8875_));
  OAI21_X1   g08683(.A1(new_n8871_), .A2(new_n8875_), .B(\asqrt[33] ), .ZN(new_n8876_));
  NAND3_X1   g08684(.A1(new_n8874_), .A2(new_n8876_), .A3(new_n4810_), .ZN(new_n8877_));
  NAND2_X1   g08685(.A1(new_n8877_), .A2(new_n8781_), .ZN(new_n8878_));
  NAND2_X1   g08686(.A1(new_n8874_), .A2(new_n8876_), .ZN(new_n8879_));
  AOI21_X1   g08687(.A1(new_n8879_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n8880_));
  AOI21_X1   g08688(.A1(new_n8880_), .A2(new_n8878_), .B(new_n8778_), .ZN(new_n8881_));
  INV_X1     g08689(.I(new_n8783_), .ZN(new_n8882_));
  INV_X1     g08690(.I(new_n8793_), .ZN(new_n8883_));
  NOR2_X1    g08691(.A1(new_n8866_), .A2(new_n8867_), .ZN(new_n8884_));
  AOI21_X1   g08692(.A1(new_n8884_), .A2(new_n6106_), .B(new_n8883_), .ZN(new_n8885_));
  NAND2_X1   g08693(.A1(new_n8868_), .A2(new_n5750_), .ZN(new_n8886_));
  OAI21_X1   g08694(.A1(new_n8885_), .A2(new_n8886_), .B(new_n8789_), .ZN(new_n8887_));
  INV_X1     g08695(.I(new_n8868_), .ZN(new_n8888_));
  OAI21_X1   g08696(.A1(new_n8885_), .A2(new_n8888_), .B(\asqrt[31] ), .ZN(new_n8889_));
  NAND3_X1   g08697(.A1(new_n8887_), .A2(new_n8889_), .A3(new_n5435_), .ZN(new_n8890_));
  NAND2_X1   g08698(.A1(new_n8890_), .A2(new_n8786_), .ZN(new_n8891_));
  NAND2_X1   g08699(.A1(new_n8887_), .A2(new_n8889_), .ZN(new_n8892_));
  AOI21_X1   g08700(.A1(new_n8892_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n8893_));
  AOI21_X1   g08701(.A1(new_n8893_), .A2(new_n8891_), .B(new_n8882_), .ZN(new_n8894_));
  AOI21_X1   g08702(.A1(new_n8891_), .A2(new_n8872_), .B(new_n5110_), .ZN(new_n8895_));
  OAI21_X1   g08703(.A1(new_n8894_), .A2(new_n8895_), .B(\asqrt[34] ), .ZN(new_n8896_));
  AOI21_X1   g08704(.A1(new_n8878_), .A2(new_n8896_), .B(new_n4510_), .ZN(new_n8897_));
  NOR2_X1    g08705(.A1(new_n8881_), .A2(new_n8897_), .ZN(new_n8898_));
  AOI21_X1   g08706(.A1(new_n8898_), .A2(new_n4224_), .B(new_n8775_), .ZN(new_n8899_));
  OAI21_X1   g08707(.A1(new_n8881_), .A2(new_n8897_), .B(\asqrt[36] ), .ZN(new_n8900_));
  NAND2_X1   g08708(.A1(new_n8900_), .A2(new_n3928_), .ZN(new_n8901_));
  OAI21_X1   g08709(.A1(new_n8899_), .A2(new_n8901_), .B(new_n8771_), .ZN(new_n8902_));
  INV_X1     g08710(.I(new_n8900_), .ZN(new_n8903_));
  OAI21_X1   g08711(.A1(new_n8899_), .A2(new_n8903_), .B(\asqrt[37] ), .ZN(new_n8904_));
  NAND3_X1   g08712(.A1(new_n8902_), .A2(new_n8904_), .A3(new_n3675_), .ZN(new_n8905_));
  NAND2_X1   g08713(.A1(new_n8905_), .A2(new_n8769_), .ZN(new_n8906_));
  NAND2_X1   g08714(.A1(new_n8902_), .A2(new_n8904_), .ZN(new_n8907_));
  AOI21_X1   g08715(.A1(new_n8907_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n8908_));
  AOI21_X1   g08716(.A1(new_n8908_), .A2(new_n8906_), .B(new_n8766_), .ZN(new_n8909_));
  INV_X1     g08717(.I(new_n8771_), .ZN(new_n8910_));
  INV_X1     g08718(.I(new_n8781_), .ZN(new_n8911_));
  NOR2_X1    g08719(.A1(new_n8894_), .A2(new_n8895_), .ZN(new_n8912_));
  AOI21_X1   g08720(.A1(new_n8912_), .A2(new_n4810_), .B(new_n8911_), .ZN(new_n8913_));
  NAND2_X1   g08721(.A1(new_n8896_), .A2(new_n4510_), .ZN(new_n8914_));
  OAI21_X1   g08722(.A1(new_n8913_), .A2(new_n8914_), .B(new_n8777_), .ZN(new_n8915_));
  INV_X1     g08723(.I(new_n8896_), .ZN(new_n8916_));
  OAI21_X1   g08724(.A1(new_n8913_), .A2(new_n8916_), .B(\asqrt[35] ), .ZN(new_n8917_));
  NAND3_X1   g08725(.A1(new_n8915_), .A2(new_n8917_), .A3(new_n4224_), .ZN(new_n8918_));
  NAND2_X1   g08726(.A1(new_n8918_), .A2(new_n8774_), .ZN(new_n8919_));
  NAND2_X1   g08727(.A1(new_n8915_), .A2(new_n8917_), .ZN(new_n8920_));
  AOI21_X1   g08728(.A1(new_n8920_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n8921_));
  AOI21_X1   g08729(.A1(new_n8921_), .A2(new_n8919_), .B(new_n8910_), .ZN(new_n8922_));
  AOI21_X1   g08730(.A1(new_n8919_), .A2(new_n8900_), .B(new_n3928_), .ZN(new_n8923_));
  OAI21_X1   g08731(.A1(new_n8922_), .A2(new_n8923_), .B(\asqrt[38] ), .ZN(new_n8924_));
  AOI21_X1   g08732(.A1(new_n8906_), .A2(new_n8924_), .B(new_n3400_), .ZN(new_n8925_));
  NOR2_X1    g08733(.A1(new_n8909_), .A2(new_n8925_), .ZN(new_n8926_));
  AOI21_X1   g08734(.A1(new_n8926_), .A2(new_n3167_), .B(new_n8763_), .ZN(new_n8927_));
  OAI21_X1   g08735(.A1(new_n8909_), .A2(new_n8925_), .B(\asqrt[40] ), .ZN(new_n8928_));
  NAND2_X1   g08736(.A1(new_n8928_), .A2(new_n2912_), .ZN(new_n8929_));
  OAI21_X1   g08737(.A1(new_n8927_), .A2(new_n8929_), .B(new_n8759_), .ZN(new_n8930_));
  INV_X1     g08738(.I(new_n8928_), .ZN(new_n8931_));
  OAI21_X1   g08739(.A1(new_n8927_), .A2(new_n8931_), .B(\asqrt[41] ), .ZN(new_n8932_));
  NAND3_X1   g08740(.A1(new_n8930_), .A2(new_n8932_), .A3(new_n2699_), .ZN(new_n8933_));
  INV_X1     g08741(.I(new_n8759_), .ZN(new_n8934_));
  INV_X1     g08742(.I(new_n8769_), .ZN(new_n8935_));
  NOR2_X1    g08743(.A1(new_n8922_), .A2(new_n8923_), .ZN(new_n8936_));
  AOI21_X1   g08744(.A1(new_n8936_), .A2(new_n3675_), .B(new_n8935_), .ZN(new_n8937_));
  NAND2_X1   g08745(.A1(new_n8924_), .A2(new_n3400_), .ZN(new_n8938_));
  OAI21_X1   g08746(.A1(new_n8937_), .A2(new_n8938_), .B(new_n8765_), .ZN(new_n8939_));
  INV_X1     g08747(.I(new_n8924_), .ZN(new_n8940_));
  OAI21_X1   g08748(.A1(new_n8937_), .A2(new_n8940_), .B(\asqrt[39] ), .ZN(new_n8941_));
  NAND3_X1   g08749(.A1(new_n8939_), .A2(new_n8941_), .A3(new_n3167_), .ZN(new_n8942_));
  NAND2_X1   g08750(.A1(new_n8942_), .A2(new_n8762_), .ZN(new_n8943_));
  NAND2_X1   g08751(.A1(new_n8939_), .A2(new_n8941_), .ZN(new_n8944_));
  AOI21_X1   g08752(.A1(new_n8944_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n8945_));
  AOI21_X1   g08753(.A1(new_n8945_), .A2(new_n8943_), .B(new_n8934_), .ZN(new_n8946_));
  AOI21_X1   g08754(.A1(new_n8943_), .A2(new_n8928_), .B(new_n2912_), .ZN(new_n8947_));
  OAI21_X1   g08755(.A1(new_n8946_), .A2(new_n8947_), .B(\asqrt[42] ), .ZN(new_n8948_));
  NAND2_X1   g08756(.A1(new_n8739_), .A2(new_n8354_), .ZN(new_n8949_));
  NOR2_X1    g08757(.A1(new_n8742_), .A2(new_n8354_), .ZN(new_n8950_));
  NAND2_X1   g08758(.A1(new_n8950_), .A2(new_n8754_), .ZN(new_n8951_));
  AOI21_X1   g08759(.A1(new_n8951_), .A2(new_n8949_), .B(new_n193_), .ZN(new_n8952_));
  INV_X1     g08760(.I(new_n8952_), .ZN(new_n8953_));
  NAND3_X1   g08761(.A1(\asqrt[23] ), .A2(new_n8724_), .A3(new_n8735_), .ZN(new_n8954_));
  XOR2_X1    g08762(.A1(new_n8954_), .A2(new_n8727_), .Z(new_n8955_));
  AOI21_X1   g08763(.A1(new_n8950_), .A2(new_n8739_), .B(new_n8740_), .ZN(new_n8956_));
  OAI21_X1   g08764(.A1(new_n8694_), .A2(new_n8696_), .B(new_n8699_), .ZN(new_n8957_));
  NOR2_X1    g08765(.A1(new_n8742_), .A2(new_n8957_), .ZN(new_n8958_));
  XOR2_X1    g08766(.A1(new_n8958_), .A2(new_n8362_), .Z(new_n8959_));
  NAND3_X1   g08767(.A1(\asqrt[23] ), .A2(new_n8710_), .A3(new_n8695_), .ZN(new_n8960_));
  XOR2_X1    g08768(.A1(new_n8960_), .A2(new_n8366_), .Z(new_n8961_));
  OAI21_X1   g08769(.A1(new_n8705_), .A2(new_n8706_), .B(new_n8709_), .ZN(new_n8962_));
  NOR2_X1    g08770(.A1(new_n8742_), .A2(new_n8962_), .ZN(new_n8963_));
  XOR2_X1    g08771(.A1(new_n8963_), .A2(new_n8368_), .Z(new_n8964_));
  INV_X1     g08772(.I(new_n8964_), .ZN(new_n8965_));
  NAND3_X1   g08773(.A1(\asqrt[23] ), .A2(new_n8672_), .A3(new_n8691_), .ZN(new_n8966_));
  XOR2_X1    g08774(.A1(new_n8966_), .A2(new_n8703_), .Z(new_n8967_));
  INV_X1     g08775(.I(new_n8967_), .ZN(new_n8968_));
  OAI21_X1   g08776(.A1(new_n8666_), .A2(new_n8668_), .B(new_n8671_), .ZN(new_n8969_));
  NOR2_X1    g08777(.A1(new_n8742_), .A2(new_n8969_), .ZN(new_n8970_));
  XOR2_X1    g08778(.A1(new_n8970_), .A2(new_n8374_), .Z(new_n8971_));
  NAND3_X1   g08779(.A1(\asqrt[23] ), .A2(new_n8685_), .A3(new_n8667_), .ZN(new_n8972_));
  XOR2_X1    g08780(.A1(new_n8972_), .A2(new_n8378_), .Z(new_n8973_));
  OAI21_X1   g08781(.A1(new_n8680_), .A2(new_n8681_), .B(new_n8684_), .ZN(new_n8974_));
  NOR2_X1    g08782(.A1(new_n8742_), .A2(new_n8974_), .ZN(new_n8975_));
  XOR2_X1    g08783(.A1(new_n8975_), .A2(new_n8380_), .Z(new_n8976_));
  INV_X1     g08784(.I(new_n8976_), .ZN(new_n8977_));
  NAND3_X1   g08785(.A1(\asqrt[23] ), .A2(new_n8644_), .A3(new_n8663_), .ZN(new_n8978_));
  XOR2_X1    g08786(.A1(new_n8978_), .A2(new_n8678_), .Z(new_n8979_));
  INV_X1     g08787(.I(new_n8979_), .ZN(new_n8980_));
  OAI21_X1   g08788(.A1(new_n8638_), .A2(new_n8640_), .B(new_n8643_), .ZN(new_n8981_));
  NOR2_X1    g08789(.A1(new_n8742_), .A2(new_n8981_), .ZN(new_n8982_));
  XOR2_X1    g08790(.A1(new_n8982_), .A2(new_n8386_), .Z(new_n8983_));
  NAND3_X1   g08791(.A1(\asqrt[23] ), .A2(new_n8657_), .A3(new_n8639_), .ZN(new_n8984_));
  XOR2_X1    g08792(.A1(new_n8984_), .A2(new_n8390_), .Z(new_n8985_));
  OAI21_X1   g08793(.A1(new_n8652_), .A2(new_n8653_), .B(new_n8656_), .ZN(new_n8986_));
  NOR2_X1    g08794(.A1(new_n8742_), .A2(new_n8986_), .ZN(new_n8987_));
  XOR2_X1    g08795(.A1(new_n8987_), .A2(new_n8392_), .Z(new_n8988_));
  INV_X1     g08796(.I(new_n8988_), .ZN(new_n8989_));
  NAND3_X1   g08797(.A1(\asqrt[23] ), .A2(new_n8616_), .A3(new_n8635_), .ZN(new_n8990_));
  XOR2_X1    g08798(.A1(new_n8990_), .A2(new_n8650_), .Z(new_n8991_));
  INV_X1     g08799(.I(new_n8991_), .ZN(new_n8992_));
  OAI21_X1   g08800(.A1(new_n8610_), .A2(new_n8612_), .B(new_n8615_), .ZN(new_n8993_));
  NOR2_X1    g08801(.A1(new_n8742_), .A2(new_n8993_), .ZN(new_n8994_));
  XOR2_X1    g08802(.A1(new_n8994_), .A2(new_n8398_), .Z(new_n8995_));
  NAND3_X1   g08803(.A1(\asqrt[23] ), .A2(new_n8629_), .A3(new_n8611_), .ZN(new_n8996_));
  XOR2_X1    g08804(.A1(new_n8996_), .A2(new_n8402_), .Z(new_n8997_));
  OAI21_X1   g08805(.A1(new_n8624_), .A2(new_n8625_), .B(new_n8628_), .ZN(new_n8998_));
  NOR2_X1    g08806(.A1(new_n8742_), .A2(new_n8998_), .ZN(new_n8999_));
  XOR2_X1    g08807(.A1(new_n8999_), .A2(new_n8404_), .Z(new_n9000_));
  INV_X1     g08808(.I(new_n9000_), .ZN(new_n9001_));
  NAND3_X1   g08809(.A1(\asqrt[23] ), .A2(new_n8588_), .A3(new_n8607_), .ZN(new_n9002_));
  XOR2_X1    g08810(.A1(new_n9002_), .A2(new_n8622_), .Z(new_n9003_));
  INV_X1     g08811(.I(new_n9003_), .ZN(new_n9004_));
  OAI21_X1   g08812(.A1(new_n8582_), .A2(new_n8584_), .B(new_n8587_), .ZN(new_n9005_));
  NOR2_X1    g08813(.A1(new_n8742_), .A2(new_n9005_), .ZN(new_n9006_));
  XOR2_X1    g08814(.A1(new_n9006_), .A2(new_n8410_), .Z(new_n9007_));
  NAND3_X1   g08815(.A1(\asqrt[23] ), .A2(new_n8601_), .A3(new_n8583_), .ZN(new_n9008_));
  XOR2_X1    g08816(.A1(new_n9008_), .A2(new_n8414_), .Z(new_n9009_));
  NOR2_X1    g08817(.A1(new_n8946_), .A2(new_n8947_), .ZN(new_n9010_));
  AOI21_X1   g08818(.A1(new_n9010_), .A2(new_n2699_), .B(new_n8746_), .ZN(new_n9011_));
  NAND2_X1   g08819(.A1(new_n8948_), .A2(new_n2464_), .ZN(new_n9012_));
  OAI21_X1   g08820(.A1(new_n9011_), .A2(new_n9012_), .B(new_n9009_), .ZN(new_n9013_));
  INV_X1     g08821(.I(new_n8948_), .ZN(new_n9014_));
  OAI21_X1   g08822(.A1(new_n9011_), .A2(new_n9014_), .B(\asqrt[43] ), .ZN(new_n9015_));
  NAND3_X1   g08823(.A1(new_n9013_), .A2(new_n9015_), .A3(new_n2271_), .ZN(new_n9016_));
  NAND2_X1   g08824(.A1(new_n9016_), .A2(new_n9007_), .ZN(new_n9017_));
  NAND2_X1   g08825(.A1(new_n9013_), .A2(new_n9015_), .ZN(new_n9018_));
  AOI21_X1   g08826(.A1(new_n9018_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n9019_));
  AOI21_X1   g08827(.A1(new_n9019_), .A2(new_n9017_), .B(new_n9004_), .ZN(new_n9020_));
  INV_X1     g08828(.I(new_n9009_), .ZN(new_n9021_));
  NAND2_X1   g08829(.A1(new_n8933_), .A2(new_n8745_), .ZN(new_n9022_));
  NAND2_X1   g08830(.A1(new_n8930_), .A2(new_n8932_), .ZN(new_n9023_));
  AOI21_X1   g08831(.A1(new_n9023_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n9024_));
  AOI21_X1   g08832(.A1(new_n9024_), .A2(new_n9022_), .B(new_n9021_), .ZN(new_n9025_));
  AOI21_X1   g08833(.A1(new_n9022_), .A2(new_n8948_), .B(new_n2464_), .ZN(new_n9026_));
  OAI21_X1   g08834(.A1(new_n9025_), .A2(new_n9026_), .B(\asqrt[44] ), .ZN(new_n9027_));
  AOI21_X1   g08835(.A1(new_n9017_), .A2(new_n9027_), .B(new_n2072_), .ZN(new_n9028_));
  NOR2_X1    g08836(.A1(new_n9020_), .A2(new_n9028_), .ZN(new_n9029_));
  AOI21_X1   g08837(.A1(new_n9029_), .A2(new_n1884_), .B(new_n9001_), .ZN(new_n9030_));
  OAI21_X1   g08838(.A1(new_n9020_), .A2(new_n9028_), .B(\asqrt[46] ), .ZN(new_n9031_));
  NAND2_X1   g08839(.A1(new_n9031_), .A2(new_n1688_), .ZN(new_n9032_));
  OAI21_X1   g08840(.A1(new_n9030_), .A2(new_n9032_), .B(new_n8997_), .ZN(new_n9033_));
  INV_X1     g08841(.I(new_n9031_), .ZN(new_n9034_));
  OAI21_X1   g08842(.A1(new_n9030_), .A2(new_n9034_), .B(\asqrt[47] ), .ZN(new_n9035_));
  NAND3_X1   g08843(.A1(new_n9033_), .A2(new_n9035_), .A3(new_n1533_), .ZN(new_n9036_));
  NAND2_X1   g08844(.A1(new_n9036_), .A2(new_n8995_), .ZN(new_n9037_));
  NAND2_X1   g08845(.A1(new_n9033_), .A2(new_n9035_), .ZN(new_n9038_));
  AOI21_X1   g08846(.A1(new_n9038_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n9039_));
  AOI21_X1   g08847(.A1(new_n9039_), .A2(new_n9037_), .B(new_n8992_), .ZN(new_n9040_));
  INV_X1     g08848(.I(new_n8997_), .ZN(new_n9041_));
  INV_X1     g08849(.I(new_n9007_), .ZN(new_n9042_));
  NOR2_X1    g08850(.A1(new_n9025_), .A2(new_n9026_), .ZN(new_n9043_));
  AOI21_X1   g08851(.A1(new_n9043_), .A2(new_n2271_), .B(new_n9042_), .ZN(new_n9044_));
  NAND2_X1   g08852(.A1(new_n9027_), .A2(new_n2072_), .ZN(new_n9045_));
  OAI21_X1   g08853(.A1(new_n9044_), .A2(new_n9045_), .B(new_n9003_), .ZN(new_n9046_));
  INV_X1     g08854(.I(new_n9027_), .ZN(new_n9047_));
  OAI21_X1   g08855(.A1(new_n9044_), .A2(new_n9047_), .B(\asqrt[45] ), .ZN(new_n9048_));
  NAND3_X1   g08856(.A1(new_n9046_), .A2(new_n9048_), .A3(new_n1884_), .ZN(new_n9049_));
  NAND2_X1   g08857(.A1(new_n9049_), .A2(new_n9000_), .ZN(new_n9050_));
  NAND2_X1   g08858(.A1(new_n9046_), .A2(new_n9048_), .ZN(new_n9051_));
  AOI21_X1   g08859(.A1(new_n9051_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n9052_));
  AOI21_X1   g08860(.A1(new_n9052_), .A2(new_n9050_), .B(new_n9041_), .ZN(new_n9053_));
  AOI21_X1   g08861(.A1(new_n9050_), .A2(new_n9031_), .B(new_n1688_), .ZN(new_n9054_));
  OAI21_X1   g08862(.A1(new_n9053_), .A2(new_n9054_), .B(\asqrt[48] ), .ZN(new_n9055_));
  AOI21_X1   g08863(.A1(new_n9037_), .A2(new_n9055_), .B(new_n1368_), .ZN(new_n9056_));
  NOR2_X1    g08864(.A1(new_n9040_), .A2(new_n9056_), .ZN(new_n9057_));
  AOI21_X1   g08865(.A1(new_n9057_), .A2(new_n1228_), .B(new_n8989_), .ZN(new_n9058_));
  OAI21_X1   g08866(.A1(new_n9040_), .A2(new_n9056_), .B(\asqrt[50] ), .ZN(new_n9059_));
  NAND2_X1   g08867(.A1(new_n9059_), .A2(new_n1088_), .ZN(new_n9060_));
  OAI21_X1   g08868(.A1(new_n9058_), .A2(new_n9060_), .B(new_n8985_), .ZN(new_n9061_));
  INV_X1     g08869(.I(new_n9059_), .ZN(new_n9062_));
  OAI21_X1   g08870(.A1(new_n9058_), .A2(new_n9062_), .B(\asqrt[51] ), .ZN(new_n9063_));
  NAND3_X1   g08871(.A1(new_n9061_), .A2(new_n9063_), .A3(new_n962_), .ZN(new_n9064_));
  NAND2_X1   g08872(.A1(new_n9064_), .A2(new_n8983_), .ZN(new_n9065_));
  NAND2_X1   g08873(.A1(new_n9061_), .A2(new_n9063_), .ZN(new_n9066_));
  AOI21_X1   g08874(.A1(new_n9066_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n9067_));
  AOI21_X1   g08875(.A1(new_n9067_), .A2(new_n9065_), .B(new_n8980_), .ZN(new_n9068_));
  INV_X1     g08876(.I(new_n8985_), .ZN(new_n9069_));
  INV_X1     g08877(.I(new_n8995_), .ZN(new_n9070_));
  NOR2_X1    g08878(.A1(new_n9053_), .A2(new_n9054_), .ZN(new_n9071_));
  AOI21_X1   g08879(.A1(new_n9071_), .A2(new_n1533_), .B(new_n9070_), .ZN(new_n9072_));
  NAND2_X1   g08880(.A1(new_n9055_), .A2(new_n1368_), .ZN(new_n9073_));
  OAI21_X1   g08881(.A1(new_n9072_), .A2(new_n9073_), .B(new_n8991_), .ZN(new_n9074_));
  INV_X1     g08882(.I(new_n9055_), .ZN(new_n9075_));
  OAI21_X1   g08883(.A1(new_n9072_), .A2(new_n9075_), .B(\asqrt[49] ), .ZN(new_n9076_));
  NAND3_X1   g08884(.A1(new_n9074_), .A2(new_n9076_), .A3(new_n1228_), .ZN(new_n9077_));
  NAND2_X1   g08885(.A1(new_n9077_), .A2(new_n8988_), .ZN(new_n9078_));
  NAND2_X1   g08886(.A1(new_n9074_), .A2(new_n9076_), .ZN(new_n9079_));
  AOI21_X1   g08887(.A1(new_n9079_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n9080_));
  AOI21_X1   g08888(.A1(new_n9080_), .A2(new_n9078_), .B(new_n9069_), .ZN(new_n9081_));
  AOI21_X1   g08889(.A1(new_n9078_), .A2(new_n9059_), .B(new_n1088_), .ZN(new_n9082_));
  OAI21_X1   g08890(.A1(new_n9081_), .A2(new_n9082_), .B(\asqrt[52] ), .ZN(new_n9083_));
  AOI21_X1   g08891(.A1(new_n9065_), .A2(new_n9083_), .B(new_n842_), .ZN(new_n9084_));
  NOR2_X1    g08892(.A1(new_n9068_), .A2(new_n9084_), .ZN(new_n9085_));
  AOI21_X1   g08893(.A1(new_n9085_), .A2(new_n720_), .B(new_n8977_), .ZN(new_n9086_));
  OAI21_X1   g08894(.A1(new_n9068_), .A2(new_n9084_), .B(\asqrt[54] ), .ZN(new_n9087_));
  NAND2_X1   g08895(.A1(new_n9087_), .A2(new_n630_), .ZN(new_n9088_));
  OAI21_X1   g08896(.A1(new_n9086_), .A2(new_n9088_), .B(new_n8973_), .ZN(new_n9089_));
  INV_X1     g08897(.I(new_n9087_), .ZN(new_n9090_));
  OAI21_X1   g08898(.A1(new_n9086_), .A2(new_n9090_), .B(\asqrt[55] ), .ZN(new_n9091_));
  NAND3_X1   g08899(.A1(new_n9089_), .A2(new_n9091_), .A3(new_n545_), .ZN(new_n9092_));
  NAND2_X1   g08900(.A1(new_n9092_), .A2(new_n8971_), .ZN(new_n9093_));
  NAND2_X1   g08901(.A1(new_n9089_), .A2(new_n9091_), .ZN(new_n9094_));
  AOI21_X1   g08902(.A1(new_n9094_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n9095_));
  AOI21_X1   g08903(.A1(new_n9095_), .A2(new_n9093_), .B(new_n8968_), .ZN(new_n9096_));
  INV_X1     g08904(.I(new_n8973_), .ZN(new_n9097_));
  INV_X1     g08905(.I(new_n8983_), .ZN(new_n9098_));
  NOR2_X1    g08906(.A1(new_n9081_), .A2(new_n9082_), .ZN(new_n9099_));
  AOI21_X1   g08907(.A1(new_n9099_), .A2(new_n962_), .B(new_n9098_), .ZN(new_n9100_));
  NAND2_X1   g08908(.A1(new_n9083_), .A2(new_n842_), .ZN(new_n9101_));
  OAI21_X1   g08909(.A1(new_n9100_), .A2(new_n9101_), .B(new_n8979_), .ZN(new_n9102_));
  INV_X1     g08910(.I(new_n9083_), .ZN(new_n9103_));
  OAI21_X1   g08911(.A1(new_n9100_), .A2(new_n9103_), .B(\asqrt[53] ), .ZN(new_n9104_));
  NAND3_X1   g08912(.A1(new_n9102_), .A2(new_n9104_), .A3(new_n720_), .ZN(new_n9105_));
  NAND2_X1   g08913(.A1(new_n9105_), .A2(new_n8976_), .ZN(new_n9106_));
  NAND2_X1   g08914(.A1(new_n9102_), .A2(new_n9104_), .ZN(new_n9107_));
  AOI21_X1   g08915(.A1(new_n9107_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n9108_));
  AOI21_X1   g08916(.A1(new_n9108_), .A2(new_n9106_), .B(new_n9097_), .ZN(new_n9109_));
  AOI21_X1   g08917(.A1(new_n9106_), .A2(new_n9087_), .B(new_n630_), .ZN(new_n9110_));
  OAI21_X1   g08918(.A1(new_n9109_), .A2(new_n9110_), .B(\asqrt[56] ), .ZN(new_n9111_));
  AOI21_X1   g08919(.A1(new_n9093_), .A2(new_n9111_), .B(new_n450_), .ZN(new_n9112_));
  NOR2_X1    g08920(.A1(new_n9096_), .A2(new_n9112_), .ZN(new_n9113_));
  AOI21_X1   g08921(.A1(new_n9113_), .A2(new_n403_), .B(new_n8965_), .ZN(new_n9114_));
  OAI21_X1   g08922(.A1(new_n9096_), .A2(new_n9112_), .B(\asqrt[58] ), .ZN(new_n9115_));
  NAND2_X1   g08923(.A1(new_n9115_), .A2(new_n339_), .ZN(new_n9116_));
  OAI21_X1   g08924(.A1(new_n9114_), .A2(new_n9116_), .B(new_n8961_), .ZN(new_n9117_));
  INV_X1     g08925(.I(new_n9115_), .ZN(new_n9118_));
  OAI21_X1   g08926(.A1(new_n9114_), .A2(new_n9118_), .B(\asqrt[59] ), .ZN(new_n9119_));
  NAND3_X1   g08927(.A1(new_n9117_), .A2(new_n9119_), .A3(new_n288_), .ZN(new_n9120_));
  NAND2_X1   g08928(.A1(new_n9120_), .A2(new_n8959_), .ZN(new_n9121_));
  INV_X1     g08929(.I(new_n8961_), .ZN(new_n9122_));
  INV_X1     g08930(.I(new_n8971_), .ZN(new_n9123_));
  NOR2_X1    g08931(.A1(new_n9109_), .A2(new_n9110_), .ZN(new_n9124_));
  AOI21_X1   g08932(.A1(new_n9124_), .A2(new_n545_), .B(new_n9123_), .ZN(new_n9125_));
  NAND2_X1   g08933(.A1(new_n9111_), .A2(new_n450_), .ZN(new_n9126_));
  OAI21_X1   g08934(.A1(new_n9125_), .A2(new_n9126_), .B(new_n8967_), .ZN(new_n9127_));
  INV_X1     g08935(.I(new_n9111_), .ZN(new_n9128_));
  OAI21_X1   g08936(.A1(new_n9125_), .A2(new_n9128_), .B(\asqrt[57] ), .ZN(new_n9129_));
  NAND3_X1   g08937(.A1(new_n9127_), .A2(new_n9129_), .A3(new_n403_), .ZN(new_n9130_));
  NAND2_X1   g08938(.A1(new_n9130_), .A2(new_n8964_), .ZN(new_n9131_));
  NAND2_X1   g08939(.A1(new_n9127_), .A2(new_n9129_), .ZN(new_n9132_));
  AOI21_X1   g08940(.A1(new_n9132_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n9133_));
  AOI21_X1   g08941(.A1(new_n9133_), .A2(new_n9131_), .B(new_n9122_), .ZN(new_n9134_));
  AOI21_X1   g08942(.A1(new_n9131_), .A2(new_n9115_), .B(new_n339_), .ZN(new_n9135_));
  OAI21_X1   g08943(.A1(new_n9134_), .A2(new_n9135_), .B(\asqrt[60] ), .ZN(new_n9136_));
  AOI21_X1   g08944(.A1(new_n9121_), .A2(new_n9136_), .B(new_n242_), .ZN(new_n9137_));
  NAND3_X1   g08945(.A1(\asqrt[23] ), .A2(new_n8700_), .A3(new_n8716_), .ZN(new_n9138_));
  XOR2_X1    g08946(.A1(new_n9138_), .A2(new_n8728_), .Z(new_n9139_));
  INV_X1     g08947(.I(new_n9139_), .ZN(new_n9140_));
  NAND2_X1   g08948(.A1(new_n9117_), .A2(new_n9119_), .ZN(new_n9141_));
  AOI21_X1   g08949(.A1(new_n9141_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n9142_));
  AOI21_X1   g08950(.A1(new_n9142_), .A2(new_n9121_), .B(new_n9140_), .ZN(new_n9143_));
  OAI21_X1   g08951(.A1(new_n9143_), .A2(new_n9137_), .B(\asqrt[62] ), .ZN(new_n9144_));
  INV_X1     g08952(.I(new_n9144_), .ZN(new_n9145_));
  NOR2_X1    g08953(.A1(new_n9143_), .A2(new_n9137_), .ZN(new_n9146_));
  AOI21_X1   g08954(.A1(new_n8701_), .A2(new_n8722_), .B(new_n8717_), .ZN(new_n9147_));
  NAND2_X1   g08955(.A1(\asqrt[23] ), .A2(new_n9147_), .ZN(new_n9148_));
  XOR2_X1    g08956(.A1(new_n9148_), .A2(new_n8720_), .Z(new_n9149_));
  INV_X1     g08957(.I(new_n9149_), .ZN(new_n9150_));
  AOI21_X1   g08958(.A1(new_n9146_), .A2(new_n234_), .B(new_n9150_), .ZN(new_n9151_));
  OAI21_X1   g08959(.A1(new_n9151_), .A2(new_n9145_), .B(new_n8956_), .ZN(new_n9152_));
  OAI21_X1   g08960(.A1(new_n9152_), .A2(new_n8955_), .B(new_n193_), .ZN(new_n9153_));
  NOR2_X1    g08961(.A1(new_n9151_), .A2(new_n9145_), .ZN(new_n9154_));
  NAND2_X1   g08962(.A1(new_n9154_), .A2(new_n8955_), .ZN(new_n9155_));
  NOR2_X1    g08963(.A1(\asqrt[23] ), .A2(new_n8355_), .ZN(new_n9156_));
  INV_X1     g08964(.I(new_n9156_), .ZN(new_n9157_));
  NAND4_X1   g08965(.A1(new_n9153_), .A2(new_n8953_), .A3(new_n9155_), .A4(new_n9157_), .ZN(\asqrt[22] ));
  NAND3_X1   g08966(.A1(\asqrt[22] ), .A2(new_n8933_), .A3(new_n8948_), .ZN(new_n9159_));
  XOR2_X1    g08967(.A1(new_n9159_), .A2(new_n8746_), .Z(new_n9160_));
  INV_X1     g08968(.I(new_n8959_), .ZN(new_n9161_));
  NOR2_X1    g08969(.A1(new_n9134_), .A2(new_n9135_), .ZN(new_n9162_));
  AOI21_X1   g08970(.A1(new_n9162_), .A2(new_n288_), .B(new_n9161_), .ZN(new_n9163_));
  INV_X1     g08971(.I(new_n9136_), .ZN(new_n9164_));
  OAI21_X1   g08972(.A1(new_n9163_), .A2(new_n9164_), .B(\asqrt[61] ), .ZN(new_n9165_));
  NAND2_X1   g08973(.A1(new_n9136_), .A2(new_n242_), .ZN(new_n9166_));
  OAI21_X1   g08974(.A1(new_n9163_), .A2(new_n9166_), .B(new_n9139_), .ZN(new_n9167_));
  NAND3_X1   g08975(.A1(new_n9167_), .A2(new_n9165_), .A3(new_n234_), .ZN(new_n9168_));
  NAND2_X1   g08976(.A1(new_n9168_), .A2(new_n9149_), .ZN(new_n9169_));
  NAND2_X1   g08977(.A1(new_n9169_), .A2(new_n9144_), .ZN(new_n9170_));
  NAND2_X1   g08978(.A1(new_n9170_), .A2(new_n8955_), .ZN(new_n9171_));
  INV_X1     g08979(.I(new_n8955_), .ZN(new_n9172_));
  INV_X1     g08980(.I(new_n8956_), .ZN(new_n9173_));
  AOI21_X1   g08981(.A1(new_n9169_), .A2(new_n9144_), .B(new_n9173_), .ZN(new_n9174_));
  AOI21_X1   g08982(.A1(new_n9174_), .A2(new_n9172_), .B(\asqrt[63] ), .ZN(new_n9175_));
  NOR2_X1    g08983(.A1(new_n9170_), .A2(new_n9172_), .ZN(new_n9176_));
  NOR4_X1    g08984(.A1(new_n9175_), .A2(new_n8952_), .A3(new_n9176_), .A4(new_n9156_), .ZN(new_n9177_));
  NOR2_X1    g08985(.A1(new_n9177_), .A2(new_n8955_), .ZN(new_n9178_));
  NAND2_X1   g08986(.A1(new_n9178_), .A2(new_n9154_), .ZN(new_n9179_));
  AOI21_X1   g08987(.A1(new_n9179_), .A2(new_n9171_), .B(new_n193_), .ZN(new_n9180_));
  NAND3_X1   g08988(.A1(\asqrt[22] ), .A2(new_n9144_), .A3(new_n9168_), .ZN(new_n9181_));
  XOR2_X1    g08989(.A1(new_n9181_), .A2(new_n9149_), .Z(new_n9182_));
  INV_X1     g08990(.I(new_n9182_), .ZN(new_n9183_));
  AOI21_X1   g08991(.A1(new_n9178_), .A2(new_n9170_), .B(new_n9176_), .ZN(new_n9184_));
  INV_X1     g08992(.I(new_n9184_), .ZN(new_n9185_));
  OAI21_X1   g08993(.A1(new_n9114_), .A2(new_n9116_), .B(new_n9119_), .ZN(new_n9186_));
  NOR2_X1    g08994(.A1(new_n9177_), .A2(new_n9186_), .ZN(new_n9187_));
  XOR2_X1    g08995(.A1(new_n9187_), .A2(new_n8961_), .Z(new_n9188_));
  NAND3_X1   g08996(.A1(\asqrt[22] ), .A2(new_n9130_), .A3(new_n9115_), .ZN(new_n9189_));
  XOR2_X1    g08997(.A1(new_n9189_), .A2(new_n8965_), .Z(new_n9190_));
  OAI21_X1   g08998(.A1(new_n9125_), .A2(new_n9126_), .B(new_n9129_), .ZN(new_n9191_));
  NOR2_X1    g08999(.A1(new_n9177_), .A2(new_n9191_), .ZN(new_n9192_));
  XOR2_X1    g09000(.A1(new_n9192_), .A2(new_n8967_), .Z(new_n9193_));
  INV_X1     g09001(.I(new_n9193_), .ZN(new_n9194_));
  NAND3_X1   g09002(.A1(\asqrt[22] ), .A2(new_n9092_), .A3(new_n9111_), .ZN(new_n9195_));
  XOR2_X1    g09003(.A1(new_n9195_), .A2(new_n9123_), .Z(new_n9196_));
  INV_X1     g09004(.I(new_n9196_), .ZN(new_n9197_));
  OAI21_X1   g09005(.A1(new_n9086_), .A2(new_n9088_), .B(new_n9091_), .ZN(new_n9198_));
  NOR2_X1    g09006(.A1(new_n9177_), .A2(new_n9198_), .ZN(new_n9199_));
  XOR2_X1    g09007(.A1(new_n9199_), .A2(new_n8973_), .Z(new_n9200_));
  NAND3_X1   g09008(.A1(\asqrt[22] ), .A2(new_n9105_), .A3(new_n9087_), .ZN(new_n9201_));
  XOR2_X1    g09009(.A1(new_n9201_), .A2(new_n8977_), .Z(new_n9202_));
  OAI21_X1   g09010(.A1(new_n9100_), .A2(new_n9101_), .B(new_n9104_), .ZN(new_n9203_));
  NOR2_X1    g09011(.A1(new_n9177_), .A2(new_n9203_), .ZN(new_n9204_));
  XOR2_X1    g09012(.A1(new_n9204_), .A2(new_n8979_), .Z(new_n9205_));
  INV_X1     g09013(.I(new_n9205_), .ZN(new_n9206_));
  NAND3_X1   g09014(.A1(\asqrt[22] ), .A2(new_n9064_), .A3(new_n9083_), .ZN(new_n9207_));
  XOR2_X1    g09015(.A1(new_n9207_), .A2(new_n9098_), .Z(new_n9208_));
  INV_X1     g09016(.I(new_n9208_), .ZN(new_n9209_));
  OAI21_X1   g09017(.A1(new_n9058_), .A2(new_n9060_), .B(new_n9063_), .ZN(new_n9210_));
  NOR2_X1    g09018(.A1(new_n9177_), .A2(new_n9210_), .ZN(new_n9211_));
  XOR2_X1    g09019(.A1(new_n9211_), .A2(new_n8985_), .Z(new_n9212_));
  NAND3_X1   g09020(.A1(\asqrt[22] ), .A2(new_n9077_), .A3(new_n9059_), .ZN(new_n9213_));
  XOR2_X1    g09021(.A1(new_n9213_), .A2(new_n8989_), .Z(new_n9214_));
  OAI21_X1   g09022(.A1(new_n9072_), .A2(new_n9073_), .B(new_n9076_), .ZN(new_n9215_));
  NOR2_X1    g09023(.A1(new_n9177_), .A2(new_n9215_), .ZN(new_n9216_));
  XOR2_X1    g09024(.A1(new_n9216_), .A2(new_n8991_), .Z(new_n9217_));
  INV_X1     g09025(.I(new_n9217_), .ZN(new_n9218_));
  NAND3_X1   g09026(.A1(\asqrt[22] ), .A2(new_n9036_), .A3(new_n9055_), .ZN(new_n9219_));
  XOR2_X1    g09027(.A1(new_n9219_), .A2(new_n9070_), .Z(new_n9220_));
  INV_X1     g09028(.I(new_n9220_), .ZN(new_n9221_));
  OAI21_X1   g09029(.A1(new_n9030_), .A2(new_n9032_), .B(new_n9035_), .ZN(new_n9222_));
  NOR2_X1    g09030(.A1(new_n9177_), .A2(new_n9222_), .ZN(new_n9223_));
  XOR2_X1    g09031(.A1(new_n9223_), .A2(new_n8997_), .Z(new_n9224_));
  NAND3_X1   g09032(.A1(\asqrt[22] ), .A2(new_n9049_), .A3(new_n9031_), .ZN(new_n9225_));
  XOR2_X1    g09033(.A1(new_n9225_), .A2(new_n9001_), .Z(new_n9226_));
  OAI21_X1   g09034(.A1(new_n9044_), .A2(new_n9045_), .B(new_n9048_), .ZN(new_n9227_));
  NOR2_X1    g09035(.A1(new_n9177_), .A2(new_n9227_), .ZN(new_n9228_));
  XOR2_X1    g09036(.A1(new_n9228_), .A2(new_n9003_), .Z(new_n9229_));
  INV_X1     g09037(.I(new_n9229_), .ZN(new_n9230_));
  NAND3_X1   g09038(.A1(\asqrt[22] ), .A2(new_n9016_), .A3(new_n9027_), .ZN(new_n9231_));
  XOR2_X1    g09039(.A1(new_n9231_), .A2(new_n9042_), .Z(new_n9232_));
  INV_X1     g09040(.I(new_n9232_), .ZN(new_n9233_));
  OAI21_X1   g09041(.A1(new_n9011_), .A2(new_n9012_), .B(new_n9015_), .ZN(new_n9234_));
  NOR2_X1    g09042(.A1(new_n9177_), .A2(new_n9234_), .ZN(new_n9235_));
  XOR2_X1    g09043(.A1(new_n9235_), .A2(new_n9009_), .Z(new_n9236_));
  OAI21_X1   g09044(.A1(new_n8927_), .A2(new_n8929_), .B(new_n8932_), .ZN(new_n9237_));
  NOR2_X1    g09045(.A1(new_n9177_), .A2(new_n9237_), .ZN(new_n9238_));
  XOR2_X1    g09046(.A1(new_n9238_), .A2(new_n8759_), .Z(new_n9239_));
  INV_X1     g09047(.I(new_n9239_), .ZN(new_n9240_));
  NAND3_X1   g09048(.A1(\asqrt[22] ), .A2(new_n8942_), .A3(new_n8928_), .ZN(new_n9241_));
  XOR2_X1    g09049(.A1(new_n9241_), .A2(new_n8763_), .Z(new_n9242_));
  INV_X1     g09050(.I(new_n9242_), .ZN(new_n9243_));
  OAI21_X1   g09051(.A1(new_n8937_), .A2(new_n8938_), .B(new_n8941_), .ZN(new_n9244_));
  NOR2_X1    g09052(.A1(new_n9177_), .A2(new_n9244_), .ZN(new_n9245_));
  XOR2_X1    g09053(.A1(new_n9245_), .A2(new_n8765_), .Z(new_n9246_));
  NAND3_X1   g09054(.A1(\asqrt[22] ), .A2(new_n8905_), .A3(new_n8924_), .ZN(new_n9247_));
  XOR2_X1    g09055(.A1(new_n9247_), .A2(new_n8935_), .Z(new_n9248_));
  OAI21_X1   g09056(.A1(new_n8899_), .A2(new_n8901_), .B(new_n8904_), .ZN(new_n9249_));
  NOR2_X1    g09057(.A1(new_n9177_), .A2(new_n9249_), .ZN(new_n9250_));
  XOR2_X1    g09058(.A1(new_n9250_), .A2(new_n8771_), .Z(new_n9251_));
  INV_X1     g09059(.I(new_n9251_), .ZN(new_n9252_));
  NAND3_X1   g09060(.A1(\asqrt[22] ), .A2(new_n8918_), .A3(new_n8900_), .ZN(new_n9253_));
  XOR2_X1    g09061(.A1(new_n9253_), .A2(new_n8775_), .Z(new_n9254_));
  INV_X1     g09062(.I(new_n9254_), .ZN(new_n9255_));
  OAI21_X1   g09063(.A1(new_n8913_), .A2(new_n8914_), .B(new_n8917_), .ZN(new_n9256_));
  NOR2_X1    g09064(.A1(new_n9177_), .A2(new_n9256_), .ZN(new_n9257_));
  XOR2_X1    g09065(.A1(new_n9257_), .A2(new_n8777_), .Z(new_n9258_));
  NAND3_X1   g09066(.A1(\asqrt[22] ), .A2(new_n8877_), .A3(new_n8896_), .ZN(new_n9259_));
  XOR2_X1    g09067(.A1(new_n9259_), .A2(new_n8911_), .Z(new_n9260_));
  OAI21_X1   g09068(.A1(new_n8871_), .A2(new_n8873_), .B(new_n8876_), .ZN(new_n9261_));
  NOR2_X1    g09069(.A1(new_n9177_), .A2(new_n9261_), .ZN(new_n9262_));
  XOR2_X1    g09070(.A1(new_n9262_), .A2(new_n8783_), .Z(new_n9263_));
  INV_X1     g09071(.I(new_n9263_), .ZN(new_n9264_));
  NAND3_X1   g09072(.A1(\asqrt[22] ), .A2(new_n8890_), .A3(new_n8872_), .ZN(new_n9265_));
  XOR2_X1    g09073(.A1(new_n9265_), .A2(new_n8787_), .Z(new_n9266_));
  INV_X1     g09074(.I(new_n9266_), .ZN(new_n9267_));
  OAI21_X1   g09075(.A1(new_n8885_), .A2(new_n8886_), .B(new_n8889_), .ZN(new_n9268_));
  NOR2_X1    g09076(.A1(new_n9177_), .A2(new_n9268_), .ZN(new_n9269_));
  XOR2_X1    g09077(.A1(new_n9269_), .A2(new_n8789_), .Z(new_n9270_));
  NAND3_X1   g09078(.A1(\asqrt[22] ), .A2(new_n8849_), .A3(new_n8868_), .ZN(new_n9271_));
  XOR2_X1    g09079(.A1(new_n9271_), .A2(new_n8883_), .Z(new_n9272_));
  OAI21_X1   g09080(.A1(new_n8843_), .A2(new_n8845_), .B(new_n8848_), .ZN(new_n9273_));
  NOR2_X1    g09081(.A1(new_n9177_), .A2(new_n9273_), .ZN(new_n9274_));
  XOR2_X1    g09082(.A1(new_n9274_), .A2(new_n8796_), .Z(new_n9275_));
  INV_X1     g09083(.I(new_n9275_), .ZN(new_n9276_));
  NAND3_X1   g09084(.A1(\asqrt[22] ), .A2(new_n8862_), .A3(new_n8844_), .ZN(new_n9277_));
  XOR2_X1    g09085(.A1(new_n9277_), .A2(new_n8799_), .Z(new_n9278_));
  INV_X1     g09086(.I(new_n9278_), .ZN(new_n9279_));
  OAI21_X1   g09087(.A1(new_n8857_), .A2(new_n8858_), .B(new_n8861_), .ZN(new_n9280_));
  NOR2_X1    g09088(.A1(new_n9177_), .A2(new_n9280_), .ZN(new_n9281_));
  XOR2_X1    g09089(.A1(new_n9281_), .A2(new_n8802_), .Z(new_n9282_));
  NAND3_X1   g09090(.A1(\asqrt[22] ), .A2(new_n8822_), .A3(new_n8840_), .ZN(new_n9283_));
  XOR2_X1    g09091(.A1(new_n9283_), .A2(new_n8856_), .Z(new_n9284_));
  NOR2_X1    g09092(.A1(new_n8819_), .A2(\asqrt[25] ), .ZN(new_n9285_));
  NOR3_X1    g09093(.A1(new_n9177_), .A2(new_n9285_), .A3(new_n8839_), .ZN(new_n9286_));
  XOR2_X1    g09094(.A1(new_n9286_), .A2(new_n8810_), .Z(new_n9287_));
  INV_X1     g09095(.I(new_n9287_), .ZN(new_n9288_));
  NAND3_X1   g09096(.A1(\asqrt[22] ), .A2(new_n8811_), .A3(new_n8812_), .ZN(new_n9289_));
  NOR4_X1    g09097(.A1(new_n9175_), .A2(new_n8742_), .A3(new_n8952_), .A4(new_n9176_), .ZN(new_n9290_));
  INV_X1     g09098(.I(new_n9290_), .ZN(new_n9291_));
  AOI21_X1   g09099(.A1(new_n9289_), .A2(new_n9291_), .B(\a[46] ), .ZN(new_n9292_));
  NOR3_X1    g09100(.A1(new_n9177_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n9293_));
  NOR3_X1    g09101(.A1(new_n9293_), .A2(new_n8462_), .A3(new_n9290_), .ZN(new_n9294_));
  NOR2_X1    g09102(.A1(new_n9294_), .A2(new_n9292_), .ZN(new_n9295_));
  INV_X1     g09103(.I(\a[42] ), .ZN(new_n9296_));
  INV_X1     g09104(.I(\a[43] ), .ZN(new_n9297_));
  NAND3_X1   g09105(.A1(new_n9296_), .A2(new_n9297_), .A3(new_n8811_), .ZN(new_n9298_));
  OAI21_X1   g09106(.A1(new_n9177_), .A2(new_n8811_), .B(new_n9298_), .ZN(new_n9299_));
  NAND2_X1   g09107(.A1(new_n9299_), .A2(\asqrt[23] ), .ZN(new_n9300_));
  OAI21_X1   g09108(.A1(new_n9177_), .A2(\a[44] ), .B(\a[45] ), .ZN(new_n9301_));
  NAND2_X1   g09109(.A1(new_n9301_), .A2(new_n9289_), .ZN(new_n9302_));
  NOR2_X1    g09110(.A1(new_n9299_), .A2(\asqrt[23] ), .ZN(new_n9303_));
  OAI21_X1   g09111(.A1(new_n9302_), .A2(new_n9303_), .B(new_n9300_), .ZN(new_n9304_));
  OAI21_X1   g09112(.A1(new_n9304_), .A2(\asqrt[24] ), .B(new_n9295_), .ZN(new_n9305_));
  NAND2_X1   g09113(.A1(new_n9304_), .A2(\asqrt[24] ), .ZN(new_n9306_));
  NAND3_X1   g09114(.A1(new_n9305_), .A2(new_n7934_), .A3(new_n9306_), .ZN(new_n9307_));
  NOR3_X1    g09115(.A1(new_n9177_), .A2(new_n8833_), .A3(new_n8818_), .ZN(new_n9308_));
  XOR2_X1    g09116(.A1(new_n9308_), .A2(new_n8835_), .Z(new_n9309_));
  AOI21_X1   g09117(.A1(new_n9305_), .A2(new_n9306_), .B(new_n7934_), .ZN(new_n9310_));
  AOI21_X1   g09118(.A1(new_n9307_), .A2(new_n9309_), .B(new_n9310_), .ZN(new_n9311_));
  AOI21_X1   g09119(.A1(new_n9311_), .A2(new_n7561_), .B(new_n9288_), .ZN(new_n9312_));
  OAI21_X1   g09120(.A1(new_n9311_), .A2(new_n7561_), .B(new_n7166_), .ZN(new_n9313_));
  OAI21_X1   g09121(.A1(new_n9312_), .A2(new_n9313_), .B(new_n9284_), .ZN(new_n9314_));
  NOR2_X1    g09122(.A1(new_n9311_), .A2(new_n7561_), .ZN(new_n9315_));
  OAI21_X1   g09123(.A1(new_n9312_), .A2(new_n9315_), .B(\asqrt[27] ), .ZN(new_n9316_));
  NAND3_X1   g09124(.A1(new_n9314_), .A2(new_n9316_), .A3(new_n6813_), .ZN(new_n9317_));
  NAND2_X1   g09125(.A1(new_n9317_), .A2(new_n9282_), .ZN(new_n9318_));
  NAND2_X1   g09126(.A1(new_n9314_), .A2(new_n9316_), .ZN(new_n9319_));
  AOI21_X1   g09127(.A1(new_n9319_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n9320_));
  AOI21_X1   g09128(.A1(new_n9320_), .A2(new_n9318_), .B(new_n9279_), .ZN(new_n9321_));
  INV_X1     g09129(.I(new_n9284_), .ZN(new_n9322_));
  OAI21_X1   g09130(.A1(new_n9293_), .A2(new_n9290_), .B(new_n8462_), .ZN(new_n9323_));
  NAND3_X1   g09131(.A1(new_n9289_), .A2(new_n9291_), .A3(\a[46] ), .ZN(new_n9324_));
  NAND2_X1   g09132(.A1(new_n9323_), .A2(new_n9324_), .ZN(new_n9325_));
  NAND2_X1   g09133(.A1(\asqrt[22] ), .A2(\a[44] ), .ZN(new_n9326_));
  AOI21_X1   g09134(.A1(new_n9326_), .A2(new_n9298_), .B(new_n8742_), .ZN(new_n9327_));
  AOI21_X1   g09135(.A1(\asqrt[22] ), .A2(new_n8811_), .B(new_n8812_), .ZN(new_n9328_));
  NOR2_X1    g09136(.A1(new_n9293_), .A2(new_n9328_), .ZN(new_n9329_));
  NAND3_X1   g09137(.A1(new_n9326_), .A2(new_n8742_), .A3(new_n9298_), .ZN(new_n9330_));
  AOI21_X1   g09138(.A1(new_n9329_), .A2(new_n9330_), .B(new_n9327_), .ZN(new_n9331_));
  AOI21_X1   g09139(.A1(new_n9331_), .A2(new_n8349_), .B(new_n9325_), .ZN(new_n9332_));
  NOR2_X1    g09140(.A1(new_n9331_), .A2(new_n8349_), .ZN(new_n9333_));
  NOR3_X1    g09141(.A1(new_n9332_), .A2(\asqrt[25] ), .A3(new_n9333_), .ZN(new_n9334_));
  INV_X1     g09142(.I(new_n9309_), .ZN(new_n9335_));
  OAI21_X1   g09143(.A1(new_n9332_), .A2(new_n9333_), .B(\asqrt[25] ), .ZN(new_n9336_));
  OAI21_X1   g09144(.A1(new_n9334_), .A2(new_n9335_), .B(new_n9336_), .ZN(new_n9337_));
  OAI21_X1   g09145(.A1(new_n9337_), .A2(\asqrt[26] ), .B(new_n9287_), .ZN(new_n9338_));
  AOI21_X1   g09146(.A1(new_n9337_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n9339_));
  AOI21_X1   g09147(.A1(new_n9339_), .A2(new_n9338_), .B(new_n9322_), .ZN(new_n9340_));
  NAND2_X1   g09148(.A1(new_n9337_), .A2(\asqrt[26] ), .ZN(new_n9341_));
  AOI21_X1   g09149(.A1(new_n9338_), .A2(new_n9341_), .B(new_n7166_), .ZN(new_n9342_));
  OAI21_X1   g09150(.A1(new_n9340_), .A2(new_n9342_), .B(\asqrt[28] ), .ZN(new_n9343_));
  AOI21_X1   g09151(.A1(new_n9318_), .A2(new_n9343_), .B(new_n6454_), .ZN(new_n9344_));
  NOR2_X1    g09152(.A1(new_n9321_), .A2(new_n9344_), .ZN(new_n9345_));
  AOI21_X1   g09153(.A1(new_n9345_), .A2(new_n6106_), .B(new_n9276_), .ZN(new_n9346_));
  OAI21_X1   g09154(.A1(new_n9321_), .A2(new_n9344_), .B(\asqrt[30] ), .ZN(new_n9347_));
  NAND2_X1   g09155(.A1(new_n9347_), .A2(new_n5750_), .ZN(new_n9348_));
  OAI21_X1   g09156(.A1(new_n9346_), .A2(new_n9348_), .B(new_n9272_), .ZN(new_n9349_));
  INV_X1     g09157(.I(new_n9347_), .ZN(new_n9350_));
  OAI21_X1   g09158(.A1(new_n9346_), .A2(new_n9350_), .B(\asqrt[31] ), .ZN(new_n9351_));
  NAND3_X1   g09159(.A1(new_n9349_), .A2(new_n9351_), .A3(new_n5435_), .ZN(new_n9352_));
  NAND2_X1   g09160(.A1(new_n9352_), .A2(new_n9270_), .ZN(new_n9353_));
  NAND2_X1   g09161(.A1(new_n9349_), .A2(new_n9351_), .ZN(new_n9354_));
  AOI21_X1   g09162(.A1(new_n9354_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n9355_));
  AOI21_X1   g09163(.A1(new_n9355_), .A2(new_n9353_), .B(new_n9267_), .ZN(new_n9356_));
  INV_X1     g09164(.I(new_n9272_), .ZN(new_n9357_));
  INV_X1     g09165(.I(new_n9282_), .ZN(new_n9358_));
  NOR2_X1    g09166(.A1(new_n9340_), .A2(new_n9342_), .ZN(new_n9359_));
  AOI21_X1   g09167(.A1(new_n9359_), .A2(new_n6813_), .B(new_n9358_), .ZN(new_n9360_));
  NAND2_X1   g09168(.A1(new_n9343_), .A2(new_n6454_), .ZN(new_n9361_));
  OAI21_X1   g09169(.A1(new_n9360_), .A2(new_n9361_), .B(new_n9278_), .ZN(new_n9362_));
  INV_X1     g09170(.I(new_n9343_), .ZN(new_n9363_));
  OAI21_X1   g09171(.A1(new_n9360_), .A2(new_n9363_), .B(\asqrt[29] ), .ZN(new_n9364_));
  NAND3_X1   g09172(.A1(new_n9362_), .A2(new_n9364_), .A3(new_n6106_), .ZN(new_n9365_));
  NAND2_X1   g09173(.A1(new_n9365_), .A2(new_n9275_), .ZN(new_n9366_));
  NAND2_X1   g09174(.A1(new_n9362_), .A2(new_n9364_), .ZN(new_n9367_));
  AOI21_X1   g09175(.A1(new_n9367_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n9368_));
  AOI21_X1   g09176(.A1(new_n9368_), .A2(new_n9366_), .B(new_n9357_), .ZN(new_n9369_));
  AOI21_X1   g09177(.A1(new_n9366_), .A2(new_n9347_), .B(new_n5750_), .ZN(new_n9370_));
  OAI21_X1   g09178(.A1(new_n9369_), .A2(new_n9370_), .B(\asqrt[32] ), .ZN(new_n9371_));
  AOI21_X1   g09179(.A1(new_n9353_), .A2(new_n9371_), .B(new_n5110_), .ZN(new_n9372_));
  NOR2_X1    g09180(.A1(new_n9356_), .A2(new_n9372_), .ZN(new_n9373_));
  AOI21_X1   g09181(.A1(new_n9373_), .A2(new_n4810_), .B(new_n9264_), .ZN(new_n9374_));
  OAI21_X1   g09182(.A1(new_n9356_), .A2(new_n9372_), .B(\asqrt[34] ), .ZN(new_n9375_));
  NAND2_X1   g09183(.A1(new_n9375_), .A2(new_n4510_), .ZN(new_n9376_));
  OAI21_X1   g09184(.A1(new_n9374_), .A2(new_n9376_), .B(new_n9260_), .ZN(new_n9377_));
  INV_X1     g09185(.I(new_n9375_), .ZN(new_n9378_));
  OAI21_X1   g09186(.A1(new_n9374_), .A2(new_n9378_), .B(\asqrt[35] ), .ZN(new_n9379_));
  NAND3_X1   g09187(.A1(new_n9377_), .A2(new_n9379_), .A3(new_n4224_), .ZN(new_n9380_));
  NAND2_X1   g09188(.A1(new_n9380_), .A2(new_n9258_), .ZN(new_n9381_));
  NAND2_X1   g09189(.A1(new_n9377_), .A2(new_n9379_), .ZN(new_n9382_));
  AOI21_X1   g09190(.A1(new_n9382_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n9383_));
  AOI21_X1   g09191(.A1(new_n9383_), .A2(new_n9381_), .B(new_n9255_), .ZN(new_n9384_));
  INV_X1     g09192(.I(new_n9260_), .ZN(new_n9385_));
  INV_X1     g09193(.I(new_n9270_), .ZN(new_n9386_));
  NOR2_X1    g09194(.A1(new_n9369_), .A2(new_n9370_), .ZN(new_n9387_));
  AOI21_X1   g09195(.A1(new_n9387_), .A2(new_n5435_), .B(new_n9386_), .ZN(new_n9388_));
  NAND2_X1   g09196(.A1(new_n9371_), .A2(new_n5110_), .ZN(new_n9389_));
  OAI21_X1   g09197(.A1(new_n9388_), .A2(new_n9389_), .B(new_n9266_), .ZN(new_n9390_));
  INV_X1     g09198(.I(new_n9371_), .ZN(new_n9391_));
  OAI21_X1   g09199(.A1(new_n9388_), .A2(new_n9391_), .B(\asqrt[33] ), .ZN(new_n9392_));
  NAND3_X1   g09200(.A1(new_n9390_), .A2(new_n9392_), .A3(new_n4810_), .ZN(new_n9393_));
  NAND2_X1   g09201(.A1(new_n9393_), .A2(new_n9263_), .ZN(new_n9394_));
  NAND2_X1   g09202(.A1(new_n9390_), .A2(new_n9392_), .ZN(new_n9395_));
  AOI21_X1   g09203(.A1(new_n9395_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n9396_));
  AOI21_X1   g09204(.A1(new_n9396_), .A2(new_n9394_), .B(new_n9385_), .ZN(new_n9397_));
  AOI21_X1   g09205(.A1(new_n9394_), .A2(new_n9375_), .B(new_n4510_), .ZN(new_n9398_));
  OAI21_X1   g09206(.A1(new_n9397_), .A2(new_n9398_), .B(\asqrt[36] ), .ZN(new_n9399_));
  AOI21_X1   g09207(.A1(new_n9381_), .A2(new_n9399_), .B(new_n3928_), .ZN(new_n9400_));
  NOR2_X1    g09208(.A1(new_n9384_), .A2(new_n9400_), .ZN(new_n9401_));
  AOI21_X1   g09209(.A1(new_n9401_), .A2(new_n3675_), .B(new_n9252_), .ZN(new_n9402_));
  OAI21_X1   g09210(.A1(new_n9384_), .A2(new_n9400_), .B(\asqrt[38] ), .ZN(new_n9403_));
  NAND2_X1   g09211(.A1(new_n9403_), .A2(new_n3400_), .ZN(new_n9404_));
  OAI21_X1   g09212(.A1(new_n9402_), .A2(new_n9404_), .B(new_n9248_), .ZN(new_n9405_));
  INV_X1     g09213(.I(new_n9403_), .ZN(new_n9406_));
  OAI21_X1   g09214(.A1(new_n9402_), .A2(new_n9406_), .B(\asqrt[39] ), .ZN(new_n9407_));
  NAND3_X1   g09215(.A1(new_n9405_), .A2(new_n9407_), .A3(new_n3167_), .ZN(new_n9408_));
  NAND2_X1   g09216(.A1(new_n9408_), .A2(new_n9246_), .ZN(new_n9409_));
  NAND2_X1   g09217(.A1(new_n9405_), .A2(new_n9407_), .ZN(new_n9410_));
  AOI21_X1   g09218(.A1(new_n9410_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n9411_));
  AOI21_X1   g09219(.A1(new_n9411_), .A2(new_n9409_), .B(new_n9243_), .ZN(new_n9412_));
  INV_X1     g09220(.I(new_n9248_), .ZN(new_n9413_));
  INV_X1     g09221(.I(new_n9258_), .ZN(new_n9414_));
  NOR2_X1    g09222(.A1(new_n9397_), .A2(new_n9398_), .ZN(new_n9415_));
  AOI21_X1   g09223(.A1(new_n9415_), .A2(new_n4224_), .B(new_n9414_), .ZN(new_n9416_));
  NAND2_X1   g09224(.A1(new_n9399_), .A2(new_n3928_), .ZN(new_n9417_));
  OAI21_X1   g09225(.A1(new_n9416_), .A2(new_n9417_), .B(new_n9254_), .ZN(new_n9418_));
  INV_X1     g09226(.I(new_n9399_), .ZN(new_n9419_));
  OAI21_X1   g09227(.A1(new_n9416_), .A2(new_n9419_), .B(\asqrt[37] ), .ZN(new_n9420_));
  NAND3_X1   g09228(.A1(new_n9418_), .A2(new_n9420_), .A3(new_n3675_), .ZN(new_n9421_));
  NAND2_X1   g09229(.A1(new_n9421_), .A2(new_n9251_), .ZN(new_n9422_));
  NAND2_X1   g09230(.A1(new_n9418_), .A2(new_n9420_), .ZN(new_n9423_));
  AOI21_X1   g09231(.A1(new_n9423_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n9424_));
  AOI21_X1   g09232(.A1(new_n9424_), .A2(new_n9422_), .B(new_n9413_), .ZN(new_n9425_));
  AOI21_X1   g09233(.A1(new_n9422_), .A2(new_n9403_), .B(new_n3400_), .ZN(new_n9426_));
  OAI21_X1   g09234(.A1(new_n9425_), .A2(new_n9426_), .B(\asqrt[40] ), .ZN(new_n9427_));
  AOI21_X1   g09235(.A1(new_n9409_), .A2(new_n9427_), .B(new_n2912_), .ZN(new_n9428_));
  NOR2_X1    g09236(.A1(new_n9412_), .A2(new_n9428_), .ZN(new_n9429_));
  AOI21_X1   g09237(.A1(new_n9429_), .A2(new_n2699_), .B(new_n9240_), .ZN(new_n9430_));
  OAI21_X1   g09238(.A1(new_n9412_), .A2(new_n9428_), .B(\asqrt[42] ), .ZN(new_n9431_));
  NAND2_X1   g09239(.A1(new_n9431_), .A2(new_n2464_), .ZN(new_n9432_));
  OAI21_X1   g09240(.A1(new_n9430_), .A2(new_n9432_), .B(new_n9160_), .ZN(new_n9433_));
  INV_X1     g09241(.I(new_n9431_), .ZN(new_n9434_));
  OAI21_X1   g09242(.A1(new_n9430_), .A2(new_n9434_), .B(\asqrt[43] ), .ZN(new_n9435_));
  NAND3_X1   g09243(.A1(new_n9433_), .A2(new_n9435_), .A3(new_n2271_), .ZN(new_n9436_));
  NAND2_X1   g09244(.A1(new_n9436_), .A2(new_n9236_), .ZN(new_n9437_));
  NAND2_X1   g09245(.A1(new_n9433_), .A2(new_n9435_), .ZN(new_n9438_));
  AOI21_X1   g09246(.A1(new_n9438_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n9439_));
  AOI21_X1   g09247(.A1(new_n9439_), .A2(new_n9437_), .B(new_n9233_), .ZN(new_n9440_));
  INV_X1     g09248(.I(new_n9160_), .ZN(new_n9441_));
  INV_X1     g09249(.I(new_n9246_), .ZN(new_n9442_));
  NOR2_X1    g09250(.A1(new_n9425_), .A2(new_n9426_), .ZN(new_n9443_));
  AOI21_X1   g09251(.A1(new_n9443_), .A2(new_n3167_), .B(new_n9442_), .ZN(new_n9444_));
  NAND2_X1   g09252(.A1(new_n9427_), .A2(new_n2912_), .ZN(new_n9445_));
  OAI21_X1   g09253(.A1(new_n9444_), .A2(new_n9445_), .B(new_n9242_), .ZN(new_n9446_));
  INV_X1     g09254(.I(new_n9427_), .ZN(new_n9447_));
  OAI21_X1   g09255(.A1(new_n9444_), .A2(new_n9447_), .B(\asqrt[41] ), .ZN(new_n9448_));
  NAND3_X1   g09256(.A1(new_n9446_), .A2(new_n9448_), .A3(new_n2699_), .ZN(new_n9449_));
  NAND2_X1   g09257(.A1(new_n9449_), .A2(new_n9239_), .ZN(new_n9450_));
  NAND2_X1   g09258(.A1(new_n9446_), .A2(new_n9448_), .ZN(new_n9451_));
  AOI21_X1   g09259(.A1(new_n9451_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n9452_));
  AOI21_X1   g09260(.A1(new_n9452_), .A2(new_n9450_), .B(new_n9441_), .ZN(new_n9453_));
  AOI21_X1   g09261(.A1(new_n9450_), .A2(new_n9431_), .B(new_n2464_), .ZN(new_n9454_));
  OAI21_X1   g09262(.A1(new_n9453_), .A2(new_n9454_), .B(\asqrt[44] ), .ZN(new_n9455_));
  AOI21_X1   g09263(.A1(new_n9437_), .A2(new_n9455_), .B(new_n2072_), .ZN(new_n9456_));
  NOR2_X1    g09264(.A1(new_n9440_), .A2(new_n9456_), .ZN(new_n9457_));
  AOI21_X1   g09265(.A1(new_n9457_), .A2(new_n1884_), .B(new_n9230_), .ZN(new_n9458_));
  OAI21_X1   g09266(.A1(new_n9440_), .A2(new_n9456_), .B(\asqrt[46] ), .ZN(new_n9459_));
  NAND2_X1   g09267(.A1(new_n9459_), .A2(new_n1688_), .ZN(new_n9460_));
  OAI21_X1   g09268(.A1(new_n9458_), .A2(new_n9460_), .B(new_n9226_), .ZN(new_n9461_));
  INV_X1     g09269(.I(new_n9459_), .ZN(new_n9462_));
  OAI21_X1   g09270(.A1(new_n9458_), .A2(new_n9462_), .B(\asqrt[47] ), .ZN(new_n9463_));
  NAND3_X1   g09271(.A1(new_n9461_), .A2(new_n9463_), .A3(new_n1533_), .ZN(new_n9464_));
  NAND2_X1   g09272(.A1(new_n9464_), .A2(new_n9224_), .ZN(new_n9465_));
  NAND2_X1   g09273(.A1(new_n9461_), .A2(new_n9463_), .ZN(new_n9466_));
  AOI21_X1   g09274(.A1(new_n9466_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n9467_));
  AOI21_X1   g09275(.A1(new_n9467_), .A2(new_n9465_), .B(new_n9221_), .ZN(new_n9468_));
  INV_X1     g09276(.I(new_n9226_), .ZN(new_n9469_));
  INV_X1     g09277(.I(new_n9236_), .ZN(new_n9470_));
  NOR2_X1    g09278(.A1(new_n9453_), .A2(new_n9454_), .ZN(new_n9471_));
  AOI21_X1   g09279(.A1(new_n9471_), .A2(new_n2271_), .B(new_n9470_), .ZN(new_n9472_));
  NAND2_X1   g09280(.A1(new_n9455_), .A2(new_n2072_), .ZN(new_n9473_));
  OAI21_X1   g09281(.A1(new_n9472_), .A2(new_n9473_), .B(new_n9232_), .ZN(new_n9474_));
  INV_X1     g09282(.I(new_n9455_), .ZN(new_n9475_));
  OAI21_X1   g09283(.A1(new_n9472_), .A2(new_n9475_), .B(\asqrt[45] ), .ZN(new_n9476_));
  NAND3_X1   g09284(.A1(new_n9474_), .A2(new_n9476_), .A3(new_n1884_), .ZN(new_n9477_));
  NAND2_X1   g09285(.A1(new_n9477_), .A2(new_n9229_), .ZN(new_n9478_));
  NAND2_X1   g09286(.A1(new_n9474_), .A2(new_n9476_), .ZN(new_n9479_));
  AOI21_X1   g09287(.A1(new_n9479_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n9480_));
  AOI21_X1   g09288(.A1(new_n9480_), .A2(new_n9478_), .B(new_n9469_), .ZN(new_n9481_));
  AOI21_X1   g09289(.A1(new_n9478_), .A2(new_n9459_), .B(new_n1688_), .ZN(new_n9482_));
  OAI21_X1   g09290(.A1(new_n9481_), .A2(new_n9482_), .B(\asqrt[48] ), .ZN(new_n9483_));
  AOI21_X1   g09291(.A1(new_n9465_), .A2(new_n9483_), .B(new_n1368_), .ZN(new_n9484_));
  NOR2_X1    g09292(.A1(new_n9468_), .A2(new_n9484_), .ZN(new_n9485_));
  AOI21_X1   g09293(.A1(new_n9485_), .A2(new_n1228_), .B(new_n9218_), .ZN(new_n9486_));
  OAI21_X1   g09294(.A1(new_n9468_), .A2(new_n9484_), .B(\asqrt[50] ), .ZN(new_n9487_));
  NAND2_X1   g09295(.A1(new_n9487_), .A2(new_n1088_), .ZN(new_n9488_));
  OAI21_X1   g09296(.A1(new_n9486_), .A2(new_n9488_), .B(new_n9214_), .ZN(new_n9489_));
  INV_X1     g09297(.I(new_n9487_), .ZN(new_n9490_));
  OAI21_X1   g09298(.A1(new_n9486_), .A2(new_n9490_), .B(\asqrt[51] ), .ZN(new_n9491_));
  NAND3_X1   g09299(.A1(new_n9489_), .A2(new_n9491_), .A3(new_n962_), .ZN(new_n9492_));
  NAND2_X1   g09300(.A1(new_n9492_), .A2(new_n9212_), .ZN(new_n9493_));
  NAND2_X1   g09301(.A1(new_n9489_), .A2(new_n9491_), .ZN(new_n9494_));
  AOI21_X1   g09302(.A1(new_n9494_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n9495_));
  AOI21_X1   g09303(.A1(new_n9495_), .A2(new_n9493_), .B(new_n9209_), .ZN(new_n9496_));
  INV_X1     g09304(.I(new_n9214_), .ZN(new_n9497_));
  INV_X1     g09305(.I(new_n9224_), .ZN(new_n9498_));
  NOR2_X1    g09306(.A1(new_n9481_), .A2(new_n9482_), .ZN(new_n9499_));
  AOI21_X1   g09307(.A1(new_n9499_), .A2(new_n1533_), .B(new_n9498_), .ZN(new_n9500_));
  NAND2_X1   g09308(.A1(new_n9483_), .A2(new_n1368_), .ZN(new_n9501_));
  OAI21_X1   g09309(.A1(new_n9500_), .A2(new_n9501_), .B(new_n9220_), .ZN(new_n9502_));
  INV_X1     g09310(.I(new_n9483_), .ZN(new_n9503_));
  OAI21_X1   g09311(.A1(new_n9500_), .A2(new_n9503_), .B(\asqrt[49] ), .ZN(new_n9504_));
  NAND3_X1   g09312(.A1(new_n9502_), .A2(new_n9504_), .A3(new_n1228_), .ZN(new_n9505_));
  NAND2_X1   g09313(.A1(new_n9505_), .A2(new_n9217_), .ZN(new_n9506_));
  NAND2_X1   g09314(.A1(new_n9502_), .A2(new_n9504_), .ZN(new_n9507_));
  AOI21_X1   g09315(.A1(new_n9507_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n9508_));
  AOI21_X1   g09316(.A1(new_n9508_), .A2(new_n9506_), .B(new_n9497_), .ZN(new_n9509_));
  AOI21_X1   g09317(.A1(new_n9506_), .A2(new_n9487_), .B(new_n1088_), .ZN(new_n9510_));
  OAI21_X1   g09318(.A1(new_n9509_), .A2(new_n9510_), .B(\asqrt[52] ), .ZN(new_n9511_));
  AOI21_X1   g09319(.A1(new_n9493_), .A2(new_n9511_), .B(new_n842_), .ZN(new_n9512_));
  NOR2_X1    g09320(.A1(new_n9496_), .A2(new_n9512_), .ZN(new_n9513_));
  AOI21_X1   g09321(.A1(new_n9513_), .A2(new_n720_), .B(new_n9206_), .ZN(new_n9514_));
  OAI21_X1   g09322(.A1(new_n9496_), .A2(new_n9512_), .B(\asqrt[54] ), .ZN(new_n9515_));
  NAND2_X1   g09323(.A1(new_n9515_), .A2(new_n630_), .ZN(new_n9516_));
  OAI21_X1   g09324(.A1(new_n9514_), .A2(new_n9516_), .B(new_n9202_), .ZN(new_n9517_));
  INV_X1     g09325(.I(new_n9515_), .ZN(new_n9518_));
  OAI21_X1   g09326(.A1(new_n9514_), .A2(new_n9518_), .B(\asqrt[55] ), .ZN(new_n9519_));
  NAND3_X1   g09327(.A1(new_n9517_), .A2(new_n9519_), .A3(new_n545_), .ZN(new_n9520_));
  NAND2_X1   g09328(.A1(new_n9520_), .A2(new_n9200_), .ZN(new_n9521_));
  NAND2_X1   g09329(.A1(new_n9517_), .A2(new_n9519_), .ZN(new_n9522_));
  AOI21_X1   g09330(.A1(new_n9522_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n9523_));
  AOI21_X1   g09331(.A1(new_n9523_), .A2(new_n9521_), .B(new_n9197_), .ZN(new_n9524_));
  INV_X1     g09332(.I(new_n9202_), .ZN(new_n9525_));
  INV_X1     g09333(.I(new_n9212_), .ZN(new_n9526_));
  NOR2_X1    g09334(.A1(new_n9509_), .A2(new_n9510_), .ZN(new_n9527_));
  AOI21_X1   g09335(.A1(new_n9527_), .A2(new_n962_), .B(new_n9526_), .ZN(new_n9528_));
  NAND2_X1   g09336(.A1(new_n9511_), .A2(new_n842_), .ZN(new_n9529_));
  OAI21_X1   g09337(.A1(new_n9528_), .A2(new_n9529_), .B(new_n9208_), .ZN(new_n9530_));
  INV_X1     g09338(.I(new_n9511_), .ZN(new_n9531_));
  OAI21_X1   g09339(.A1(new_n9528_), .A2(new_n9531_), .B(\asqrt[53] ), .ZN(new_n9532_));
  NAND3_X1   g09340(.A1(new_n9530_), .A2(new_n9532_), .A3(new_n720_), .ZN(new_n9533_));
  NAND2_X1   g09341(.A1(new_n9533_), .A2(new_n9205_), .ZN(new_n9534_));
  NAND2_X1   g09342(.A1(new_n9530_), .A2(new_n9532_), .ZN(new_n9535_));
  AOI21_X1   g09343(.A1(new_n9535_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n9536_));
  AOI21_X1   g09344(.A1(new_n9536_), .A2(new_n9534_), .B(new_n9525_), .ZN(new_n9537_));
  AOI21_X1   g09345(.A1(new_n9534_), .A2(new_n9515_), .B(new_n630_), .ZN(new_n9538_));
  OAI21_X1   g09346(.A1(new_n9537_), .A2(new_n9538_), .B(\asqrt[56] ), .ZN(new_n9539_));
  AOI21_X1   g09347(.A1(new_n9521_), .A2(new_n9539_), .B(new_n450_), .ZN(new_n9540_));
  NOR2_X1    g09348(.A1(new_n9524_), .A2(new_n9540_), .ZN(new_n9541_));
  AOI21_X1   g09349(.A1(new_n9541_), .A2(new_n403_), .B(new_n9194_), .ZN(new_n9542_));
  OAI21_X1   g09350(.A1(new_n9524_), .A2(new_n9540_), .B(\asqrt[58] ), .ZN(new_n9543_));
  NAND2_X1   g09351(.A1(new_n9543_), .A2(new_n339_), .ZN(new_n9544_));
  OAI21_X1   g09352(.A1(new_n9542_), .A2(new_n9544_), .B(new_n9190_), .ZN(new_n9545_));
  INV_X1     g09353(.I(new_n9543_), .ZN(new_n9546_));
  OAI21_X1   g09354(.A1(new_n9542_), .A2(new_n9546_), .B(\asqrt[59] ), .ZN(new_n9547_));
  NAND3_X1   g09355(.A1(new_n9545_), .A2(new_n9547_), .A3(new_n288_), .ZN(new_n9548_));
  NAND2_X1   g09356(.A1(new_n9548_), .A2(new_n9188_), .ZN(new_n9549_));
  INV_X1     g09357(.I(new_n9190_), .ZN(new_n9550_));
  INV_X1     g09358(.I(new_n9200_), .ZN(new_n9551_));
  NOR2_X1    g09359(.A1(new_n9537_), .A2(new_n9538_), .ZN(new_n9552_));
  AOI21_X1   g09360(.A1(new_n9552_), .A2(new_n545_), .B(new_n9551_), .ZN(new_n9553_));
  NAND2_X1   g09361(.A1(new_n9539_), .A2(new_n450_), .ZN(new_n9554_));
  OAI21_X1   g09362(.A1(new_n9553_), .A2(new_n9554_), .B(new_n9196_), .ZN(new_n9555_));
  INV_X1     g09363(.I(new_n9539_), .ZN(new_n9556_));
  OAI21_X1   g09364(.A1(new_n9553_), .A2(new_n9556_), .B(\asqrt[57] ), .ZN(new_n9557_));
  NAND3_X1   g09365(.A1(new_n9555_), .A2(new_n9557_), .A3(new_n403_), .ZN(new_n9558_));
  NAND2_X1   g09366(.A1(new_n9558_), .A2(new_n9193_), .ZN(new_n9559_));
  NAND2_X1   g09367(.A1(new_n9555_), .A2(new_n9557_), .ZN(new_n9560_));
  AOI21_X1   g09368(.A1(new_n9560_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n9561_));
  AOI21_X1   g09369(.A1(new_n9561_), .A2(new_n9559_), .B(new_n9550_), .ZN(new_n9562_));
  AOI21_X1   g09370(.A1(new_n9559_), .A2(new_n9543_), .B(new_n339_), .ZN(new_n9563_));
  OAI21_X1   g09371(.A1(new_n9562_), .A2(new_n9563_), .B(\asqrt[60] ), .ZN(new_n9564_));
  AOI21_X1   g09372(.A1(new_n9549_), .A2(new_n9564_), .B(new_n242_), .ZN(new_n9565_));
  NAND3_X1   g09373(.A1(\asqrt[22] ), .A2(new_n9120_), .A3(new_n9136_), .ZN(new_n9566_));
  XOR2_X1    g09374(.A1(new_n9566_), .A2(new_n9161_), .Z(new_n9567_));
  INV_X1     g09375(.I(new_n9567_), .ZN(new_n9568_));
  NAND2_X1   g09376(.A1(new_n9545_), .A2(new_n9547_), .ZN(new_n9569_));
  AOI21_X1   g09377(.A1(new_n9569_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n9570_));
  AOI21_X1   g09378(.A1(new_n9570_), .A2(new_n9549_), .B(new_n9568_), .ZN(new_n9571_));
  OAI21_X1   g09379(.A1(new_n9571_), .A2(new_n9565_), .B(\asqrt[62] ), .ZN(new_n9572_));
  AOI21_X1   g09380(.A1(new_n9121_), .A2(new_n9142_), .B(new_n9137_), .ZN(new_n9573_));
  NAND2_X1   g09381(.A1(\asqrt[22] ), .A2(new_n9573_), .ZN(new_n9574_));
  XOR2_X1    g09382(.A1(new_n9574_), .A2(new_n9140_), .Z(new_n9575_));
  INV_X1     g09383(.I(new_n9188_), .ZN(new_n9576_));
  NOR2_X1    g09384(.A1(new_n9562_), .A2(new_n9563_), .ZN(new_n9577_));
  AOI21_X1   g09385(.A1(new_n9577_), .A2(new_n288_), .B(new_n9576_), .ZN(new_n9578_));
  INV_X1     g09386(.I(new_n9564_), .ZN(new_n9579_));
  OAI21_X1   g09387(.A1(new_n9578_), .A2(new_n9579_), .B(\asqrt[61] ), .ZN(new_n9580_));
  NAND2_X1   g09388(.A1(new_n9564_), .A2(new_n242_), .ZN(new_n9581_));
  OAI21_X1   g09389(.A1(new_n9578_), .A2(new_n9581_), .B(new_n9567_), .ZN(new_n9582_));
  NAND3_X1   g09390(.A1(new_n9582_), .A2(new_n9580_), .A3(new_n234_), .ZN(new_n9583_));
  NAND2_X1   g09391(.A1(new_n9583_), .A2(new_n9575_), .ZN(new_n9584_));
  AOI21_X1   g09392(.A1(new_n9584_), .A2(new_n9572_), .B(new_n9185_), .ZN(new_n9585_));
  AOI21_X1   g09393(.A1(new_n9585_), .A2(new_n9183_), .B(\asqrt[63] ), .ZN(new_n9586_));
  NAND2_X1   g09394(.A1(new_n9584_), .A2(new_n9572_), .ZN(new_n9587_));
  NOR2_X1    g09395(.A1(new_n9587_), .A2(new_n9183_), .ZN(new_n9588_));
  NOR2_X1    g09396(.A1(\asqrt[22] ), .A2(new_n9172_), .ZN(new_n9589_));
  NOR4_X1    g09397(.A1(new_n9586_), .A2(new_n9180_), .A3(new_n9588_), .A4(new_n9589_), .ZN(new_n9590_));
  OAI21_X1   g09398(.A1(new_n9430_), .A2(new_n9432_), .B(new_n9435_), .ZN(new_n9591_));
  NOR2_X1    g09399(.A1(new_n9590_), .A2(new_n9591_), .ZN(new_n9592_));
  XOR2_X1    g09400(.A1(new_n9592_), .A2(new_n9160_), .Z(new_n9593_));
  INV_X1     g09401(.I(new_n9593_), .ZN(new_n9594_));
  INV_X1     g09402(.I(new_n9180_), .ZN(new_n9595_));
  INV_X1     g09403(.I(new_n9572_), .ZN(new_n9596_));
  NOR2_X1    g09404(.A1(new_n9571_), .A2(new_n9565_), .ZN(new_n9597_));
  INV_X1     g09405(.I(new_n9575_), .ZN(new_n9598_));
  AOI21_X1   g09406(.A1(new_n9597_), .A2(new_n234_), .B(new_n9598_), .ZN(new_n9599_));
  OAI21_X1   g09407(.A1(new_n9599_), .A2(new_n9596_), .B(new_n9184_), .ZN(new_n9600_));
  OAI21_X1   g09408(.A1(new_n9600_), .A2(new_n9182_), .B(new_n193_), .ZN(new_n9601_));
  NOR2_X1    g09409(.A1(new_n9599_), .A2(new_n9596_), .ZN(new_n9602_));
  NAND2_X1   g09410(.A1(new_n9602_), .A2(new_n9182_), .ZN(new_n9603_));
  INV_X1     g09411(.I(new_n9589_), .ZN(new_n9604_));
  NAND4_X1   g09412(.A1(new_n9601_), .A2(new_n9595_), .A3(new_n9603_), .A4(new_n9604_), .ZN(\asqrt[21] ));
  NAND3_X1   g09413(.A1(\asqrt[21] ), .A2(new_n9449_), .A3(new_n9431_), .ZN(new_n9606_));
  XOR2_X1    g09414(.A1(new_n9606_), .A2(new_n9240_), .Z(new_n9607_));
  OAI21_X1   g09415(.A1(new_n9444_), .A2(new_n9445_), .B(new_n9448_), .ZN(new_n9608_));
  NOR2_X1    g09416(.A1(new_n9590_), .A2(new_n9608_), .ZN(new_n9609_));
  XOR2_X1    g09417(.A1(new_n9609_), .A2(new_n9242_), .Z(new_n9610_));
  INV_X1     g09418(.I(new_n9610_), .ZN(new_n9611_));
  NAND3_X1   g09419(.A1(\asqrt[21] ), .A2(new_n9408_), .A3(new_n9427_), .ZN(new_n9612_));
  XOR2_X1    g09420(.A1(new_n9612_), .A2(new_n9442_), .Z(new_n9613_));
  INV_X1     g09421(.I(new_n9613_), .ZN(new_n9614_));
  OAI21_X1   g09422(.A1(new_n9402_), .A2(new_n9404_), .B(new_n9407_), .ZN(new_n9615_));
  NOR2_X1    g09423(.A1(new_n9590_), .A2(new_n9615_), .ZN(new_n9616_));
  XOR2_X1    g09424(.A1(new_n9616_), .A2(new_n9248_), .Z(new_n9617_));
  NAND3_X1   g09425(.A1(\asqrt[21] ), .A2(new_n9421_), .A3(new_n9403_), .ZN(new_n9618_));
  XOR2_X1    g09426(.A1(new_n9618_), .A2(new_n9252_), .Z(new_n9619_));
  OAI21_X1   g09427(.A1(new_n9416_), .A2(new_n9417_), .B(new_n9420_), .ZN(new_n9620_));
  NOR2_X1    g09428(.A1(new_n9590_), .A2(new_n9620_), .ZN(new_n9621_));
  XOR2_X1    g09429(.A1(new_n9621_), .A2(new_n9254_), .Z(new_n9622_));
  INV_X1     g09430(.I(new_n9622_), .ZN(new_n9623_));
  NAND3_X1   g09431(.A1(\asqrt[21] ), .A2(new_n9380_), .A3(new_n9399_), .ZN(new_n9624_));
  XOR2_X1    g09432(.A1(new_n9624_), .A2(new_n9414_), .Z(new_n9625_));
  INV_X1     g09433(.I(new_n9625_), .ZN(new_n9626_));
  OAI21_X1   g09434(.A1(new_n9374_), .A2(new_n9376_), .B(new_n9379_), .ZN(new_n9627_));
  NOR2_X1    g09435(.A1(new_n9590_), .A2(new_n9627_), .ZN(new_n9628_));
  XOR2_X1    g09436(.A1(new_n9628_), .A2(new_n9260_), .Z(new_n9629_));
  NAND3_X1   g09437(.A1(\asqrt[21] ), .A2(new_n9393_), .A3(new_n9375_), .ZN(new_n9630_));
  XOR2_X1    g09438(.A1(new_n9630_), .A2(new_n9264_), .Z(new_n9631_));
  OAI21_X1   g09439(.A1(new_n9388_), .A2(new_n9389_), .B(new_n9392_), .ZN(new_n9632_));
  NOR2_X1    g09440(.A1(new_n9590_), .A2(new_n9632_), .ZN(new_n9633_));
  XOR2_X1    g09441(.A1(new_n9633_), .A2(new_n9266_), .Z(new_n9634_));
  INV_X1     g09442(.I(new_n9634_), .ZN(new_n9635_));
  NAND3_X1   g09443(.A1(\asqrt[21] ), .A2(new_n9352_), .A3(new_n9371_), .ZN(new_n9636_));
  XOR2_X1    g09444(.A1(new_n9636_), .A2(new_n9386_), .Z(new_n9637_));
  INV_X1     g09445(.I(new_n9637_), .ZN(new_n9638_));
  OAI21_X1   g09446(.A1(new_n9346_), .A2(new_n9348_), .B(new_n9351_), .ZN(new_n9639_));
  NOR2_X1    g09447(.A1(new_n9590_), .A2(new_n9639_), .ZN(new_n9640_));
  XOR2_X1    g09448(.A1(new_n9640_), .A2(new_n9272_), .Z(new_n9641_));
  NAND3_X1   g09449(.A1(\asqrt[21] ), .A2(new_n9365_), .A3(new_n9347_), .ZN(new_n9642_));
  XOR2_X1    g09450(.A1(new_n9642_), .A2(new_n9276_), .Z(new_n9643_));
  OAI21_X1   g09451(.A1(new_n9360_), .A2(new_n9361_), .B(new_n9364_), .ZN(new_n9644_));
  NOR2_X1    g09452(.A1(new_n9590_), .A2(new_n9644_), .ZN(new_n9645_));
  XOR2_X1    g09453(.A1(new_n9645_), .A2(new_n9278_), .Z(new_n9646_));
  INV_X1     g09454(.I(new_n9646_), .ZN(new_n9647_));
  NAND3_X1   g09455(.A1(\asqrt[21] ), .A2(new_n9317_), .A3(new_n9343_), .ZN(new_n9648_));
  XOR2_X1    g09456(.A1(new_n9648_), .A2(new_n9358_), .Z(new_n9649_));
  INV_X1     g09457(.I(new_n9649_), .ZN(new_n9650_));
  AOI21_X1   g09458(.A1(new_n9338_), .A2(new_n9339_), .B(new_n9342_), .ZN(new_n9651_));
  NAND2_X1   g09459(.A1(\asqrt[21] ), .A2(new_n9651_), .ZN(new_n9652_));
  XOR2_X1    g09460(.A1(new_n9652_), .A2(new_n9322_), .Z(new_n9653_));
  NOR2_X1    g09461(.A1(new_n9337_), .A2(\asqrt[26] ), .ZN(new_n9654_));
  NOR3_X1    g09462(.A1(new_n9590_), .A2(new_n9654_), .A3(new_n9315_), .ZN(new_n9655_));
  XOR2_X1    g09463(.A1(new_n9655_), .A2(new_n9287_), .Z(new_n9656_));
  NOR3_X1    g09464(.A1(new_n9590_), .A2(new_n9334_), .A3(new_n9310_), .ZN(new_n9657_));
  XOR2_X1    g09465(.A1(new_n9657_), .A2(new_n9309_), .Z(new_n9658_));
  INV_X1     g09466(.I(new_n9658_), .ZN(new_n9659_));
  NOR2_X1    g09467(.A1(new_n9304_), .A2(\asqrt[24] ), .ZN(new_n9660_));
  NOR3_X1    g09468(.A1(new_n9590_), .A2(new_n9660_), .A3(new_n9333_), .ZN(new_n9661_));
  XOR2_X1    g09469(.A1(new_n9661_), .A2(new_n9295_), .Z(new_n9662_));
  INV_X1     g09470(.I(new_n9662_), .ZN(new_n9663_));
  NAND3_X1   g09471(.A1(\asqrt[21] ), .A2(new_n9296_), .A3(new_n9297_), .ZN(new_n9664_));
  NOR4_X1    g09472(.A1(new_n9586_), .A2(new_n9177_), .A3(new_n9180_), .A4(new_n9588_), .ZN(new_n9665_));
  INV_X1     g09473(.I(new_n9665_), .ZN(new_n9666_));
  AOI21_X1   g09474(.A1(new_n9664_), .A2(new_n9666_), .B(\a[44] ), .ZN(new_n9667_));
  NOR3_X1    g09475(.A1(new_n9590_), .A2(\a[42] ), .A3(\a[43] ), .ZN(new_n9668_));
  NOR3_X1    g09476(.A1(new_n9668_), .A2(new_n8811_), .A3(new_n9665_), .ZN(new_n9669_));
  NOR2_X1    g09477(.A1(new_n9669_), .A2(new_n9667_), .ZN(new_n9670_));
  INV_X1     g09478(.I(\a[40] ), .ZN(new_n9671_));
  INV_X1     g09479(.I(\a[41] ), .ZN(new_n9672_));
  NAND3_X1   g09480(.A1(new_n9671_), .A2(new_n9672_), .A3(new_n9296_), .ZN(new_n9673_));
  OAI21_X1   g09481(.A1(new_n9590_), .A2(new_n9296_), .B(new_n9673_), .ZN(new_n9674_));
  NAND2_X1   g09482(.A1(new_n9674_), .A2(\asqrt[22] ), .ZN(new_n9675_));
  OAI21_X1   g09483(.A1(new_n9590_), .A2(\a[42] ), .B(\a[43] ), .ZN(new_n9676_));
  NAND2_X1   g09484(.A1(new_n9676_), .A2(new_n9664_), .ZN(new_n9677_));
  NOR2_X1    g09485(.A1(new_n9674_), .A2(\asqrt[22] ), .ZN(new_n9678_));
  OAI21_X1   g09486(.A1(new_n9677_), .A2(new_n9678_), .B(new_n9675_), .ZN(new_n9679_));
  OAI21_X1   g09487(.A1(\asqrt[23] ), .A2(new_n9679_), .B(new_n9670_), .ZN(new_n9680_));
  NAND2_X1   g09488(.A1(new_n9679_), .A2(\asqrt[23] ), .ZN(new_n9681_));
  NAND3_X1   g09489(.A1(new_n9680_), .A2(new_n8349_), .A3(new_n9681_), .ZN(new_n9682_));
  NOR3_X1    g09490(.A1(new_n9590_), .A2(new_n9327_), .A3(new_n9303_), .ZN(new_n9683_));
  XOR2_X1    g09491(.A1(new_n9683_), .A2(new_n9329_), .Z(new_n9684_));
  NAND2_X1   g09492(.A1(new_n9682_), .A2(new_n9684_), .ZN(new_n9685_));
  NAND2_X1   g09493(.A1(new_n9680_), .A2(new_n9681_), .ZN(new_n9686_));
  AOI21_X1   g09494(.A1(new_n9686_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n9687_));
  AOI21_X1   g09495(.A1(new_n9687_), .A2(new_n9685_), .B(new_n9663_), .ZN(new_n9688_));
  OAI21_X1   g09496(.A1(new_n9668_), .A2(new_n9665_), .B(new_n8811_), .ZN(new_n9689_));
  NAND3_X1   g09497(.A1(new_n9664_), .A2(\a[44] ), .A3(new_n9666_), .ZN(new_n9690_));
  NAND2_X1   g09498(.A1(new_n9689_), .A2(new_n9690_), .ZN(new_n9691_));
  NAND2_X1   g09499(.A1(\asqrt[21] ), .A2(\a[42] ), .ZN(new_n9692_));
  AOI21_X1   g09500(.A1(new_n9692_), .A2(new_n9673_), .B(new_n9177_), .ZN(new_n9693_));
  AOI21_X1   g09501(.A1(\asqrt[21] ), .A2(new_n9296_), .B(new_n9297_), .ZN(new_n9694_));
  NOR2_X1    g09502(.A1(new_n9694_), .A2(new_n9668_), .ZN(new_n9695_));
  NAND3_X1   g09503(.A1(new_n9692_), .A2(new_n9177_), .A3(new_n9673_), .ZN(new_n9696_));
  AOI21_X1   g09504(.A1(new_n9695_), .A2(new_n9696_), .B(new_n9693_), .ZN(new_n9697_));
  AOI21_X1   g09505(.A1(new_n9697_), .A2(new_n8742_), .B(new_n9691_), .ZN(new_n9698_));
  NOR2_X1    g09506(.A1(new_n9697_), .A2(new_n8742_), .ZN(new_n9699_));
  OAI21_X1   g09507(.A1(new_n9698_), .A2(new_n9699_), .B(\asqrt[24] ), .ZN(new_n9700_));
  AOI21_X1   g09508(.A1(new_n9685_), .A2(new_n9700_), .B(new_n7934_), .ZN(new_n9701_));
  NOR2_X1    g09509(.A1(new_n9688_), .A2(new_n9701_), .ZN(new_n9702_));
  AOI21_X1   g09510(.A1(new_n9702_), .A2(new_n7561_), .B(new_n9659_), .ZN(new_n9703_));
  OAI21_X1   g09511(.A1(new_n9688_), .A2(new_n9701_), .B(\asqrt[26] ), .ZN(new_n9704_));
  NAND2_X1   g09512(.A1(new_n9704_), .A2(new_n7166_), .ZN(new_n9705_));
  OAI21_X1   g09513(.A1(new_n9703_), .A2(new_n9705_), .B(new_n9656_), .ZN(new_n9706_));
  INV_X1     g09514(.I(new_n9704_), .ZN(new_n9707_));
  OAI21_X1   g09515(.A1(new_n9703_), .A2(new_n9707_), .B(\asqrt[27] ), .ZN(new_n9708_));
  NAND3_X1   g09516(.A1(new_n9706_), .A2(new_n9708_), .A3(new_n6813_), .ZN(new_n9709_));
  NAND2_X1   g09517(.A1(new_n9709_), .A2(new_n9653_), .ZN(new_n9710_));
  NAND2_X1   g09518(.A1(new_n9706_), .A2(new_n9708_), .ZN(new_n9711_));
  AOI21_X1   g09519(.A1(new_n9711_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n9712_));
  AOI21_X1   g09520(.A1(new_n9712_), .A2(new_n9710_), .B(new_n9650_), .ZN(new_n9713_));
  INV_X1     g09521(.I(new_n9656_), .ZN(new_n9714_));
  NOR2_X1    g09522(.A1(new_n9698_), .A2(new_n9699_), .ZN(new_n9715_));
  INV_X1     g09523(.I(new_n9684_), .ZN(new_n9716_));
  AOI21_X1   g09524(.A1(new_n9715_), .A2(new_n8349_), .B(new_n9716_), .ZN(new_n9717_));
  NAND2_X1   g09525(.A1(new_n9700_), .A2(new_n7934_), .ZN(new_n9718_));
  OAI21_X1   g09526(.A1(new_n9717_), .A2(new_n9718_), .B(new_n9662_), .ZN(new_n9719_));
  INV_X1     g09527(.I(new_n9700_), .ZN(new_n9720_));
  OAI21_X1   g09528(.A1(new_n9717_), .A2(new_n9720_), .B(\asqrt[25] ), .ZN(new_n9721_));
  NAND3_X1   g09529(.A1(new_n9719_), .A2(new_n9721_), .A3(new_n7561_), .ZN(new_n9722_));
  NAND2_X1   g09530(.A1(new_n9722_), .A2(new_n9658_), .ZN(new_n9723_));
  NAND2_X1   g09531(.A1(new_n9719_), .A2(new_n9721_), .ZN(new_n9724_));
  AOI21_X1   g09532(.A1(new_n9724_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n9725_));
  AOI21_X1   g09533(.A1(new_n9725_), .A2(new_n9723_), .B(new_n9714_), .ZN(new_n9726_));
  AOI21_X1   g09534(.A1(new_n9723_), .A2(new_n9704_), .B(new_n7166_), .ZN(new_n9727_));
  OAI21_X1   g09535(.A1(new_n9726_), .A2(new_n9727_), .B(\asqrt[28] ), .ZN(new_n9728_));
  AOI21_X1   g09536(.A1(new_n9710_), .A2(new_n9728_), .B(new_n6454_), .ZN(new_n9729_));
  NOR2_X1    g09537(.A1(new_n9713_), .A2(new_n9729_), .ZN(new_n9730_));
  AOI21_X1   g09538(.A1(new_n9730_), .A2(new_n6106_), .B(new_n9647_), .ZN(new_n9731_));
  OAI21_X1   g09539(.A1(new_n9713_), .A2(new_n9729_), .B(\asqrt[30] ), .ZN(new_n9732_));
  NAND2_X1   g09540(.A1(new_n9732_), .A2(new_n5750_), .ZN(new_n9733_));
  OAI21_X1   g09541(.A1(new_n9731_), .A2(new_n9733_), .B(new_n9643_), .ZN(new_n9734_));
  INV_X1     g09542(.I(new_n9732_), .ZN(new_n9735_));
  OAI21_X1   g09543(.A1(new_n9731_), .A2(new_n9735_), .B(\asqrt[31] ), .ZN(new_n9736_));
  NAND3_X1   g09544(.A1(new_n9734_), .A2(new_n9736_), .A3(new_n5435_), .ZN(new_n9737_));
  NAND2_X1   g09545(.A1(new_n9737_), .A2(new_n9641_), .ZN(new_n9738_));
  NAND2_X1   g09546(.A1(new_n9734_), .A2(new_n9736_), .ZN(new_n9739_));
  AOI21_X1   g09547(.A1(new_n9739_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n9740_));
  AOI21_X1   g09548(.A1(new_n9740_), .A2(new_n9738_), .B(new_n9638_), .ZN(new_n9741_));
  INV_X1     g09549(.I(new_n9643_), .ZN(new_n9742_));
  INV_X1     g09550(.I(new_n9653_), .ZN(new_n9743_));
  NOR2_X1    g09551(.A1(new_n9726_), .A2(new_n9727_), .ZN(new_n9744_));
  AOI21_X1   g09552(.A1(new_n9744_), .A2(new_n6813_), .B(new_n9743_), .ZN(new_n9745_));
  NAND2_X1   g09553(.A1(new_n9728_), .A2(new_n6454_), .ZN(new_n9746_));
  OAI21_X1   g09554(.A1(new_n9745_), .A2(new_n9746_), .B(new_n9649_), .ZN(new_n9747_));
  INV_X1     g09555(.I(new_n9728_), .ZN(new_n9748_));
  OAI21_X1   g09556(.A1(new_n9745_), .A2(new_n9748_), .B(\asqrt[29] ), .ZN(new_n9749_));
  NAND3_X1   g09557(.A1(new_n9747_), .A2(new_n9749_), .A3(new_n6106_), .ZN(new_n9750_));
  NAND2_X1   g09558(.A1(new_n9750_), .A2(new_n9646_), .ZN(new_n9751_));
  NAND2_X1   g09559(.A1(new_n9747_), .A2(new_n9749_), .ZN(new_n9752_));
  AOI21_X1   g09560(.A1(new_n9752_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n9753_));
  AOI21_X1   g09561(.A1(new_n9753_), .A2(new_n9751_), .B(new_n9742_), .ZN(new_n9754_));
  AOI21_X1   g09562(.A1(new_n9751_), .A2(new_n9732_), .B(new_n5750_), .ZN(new_n9755_));
  OAI21_X1   g09563(.A1(new_n9754_), .A2(new_n9755_), .B(\asqrt[32] ), .ZN(new_n9756_));
  AOI21_X1   g09564(.A1(new_n9738_), .A2(new_n9756_), .B(new_n5110_), .ZN(new_n9757_));
  NOR2_X1    g09565(.A1(new_n9741_), .A2(new_n9757_), .ZN(new_n9758_));
  AOI21_X1   g09566(.A1(new_n9758_), .A2(new_n4810_), .B(new_n9635_), .ZN(new_n9759_));
  OAI21_X1   g09567(.A1(new_n9741_), .A2(new_n9757_), .B(\asqrt[34] ), .ZN(new_n9760_));
  NAND2_X1   g09568(.A1(new_n9760_), .A2(new_n4510_), .ZN(new_n9761_));
  OAI21_X1   g09569(.A1(new_n9759_), .A2(new_n9761_), .B(new_n9631_), .ZN(new_n9762_));
  INV_X1     g09570(.I(new_n9760_), .ZN(new_n9763_));
  OAI21_X1   g09571(.A1(new_n9759_), .A2(new_n9763_), .B(\asqrt[35] ), .ZN(new_n9764_));
  NAND3_X1   g09572(.A1(new_n9762_), .A2(new_n9764_), .A3(new_n4224_), .ZN(new_n9765_));
  NAND2_X1   g09573(.A1(new_n9765_), .A2(new_n9629_), .ZN(new_n9766_));
  NAND2_X1   g09574(.A1(new_n9762_), .A2(new_n9764_), .ZN(new_n9767_));
  AOI21_X1   g09575(.A1(new_n9767_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n9768_));
  AOI21_X1   g09576(.A1(new_n9768_), .A2(new_n9766_), .B(new_n9626_), .ZN(new_n9769_));
  INV_X1     g09577(.I(new_n9631_), .ZN(new_n9770_));
  INV_X1     g09578(.I(new_n9641_), .ZN(new_n9771_));
  NOR2_X1    g09579(.A1(new_n9754_), .A2(new_n9755_), .ZN(new_n9772_));
  AOI21_X1   g09580(.A1(new_n9772_), .A2(new_n5435_), .B(new_n9771_), .ZN(new_n9773_));
  NAND2_X1   g09581(.A1(new_n9756_), .A2(new_n5110_), .ZN(new_n9774_));
  OAI21_X1   g09582(.A1(new_n9773_), .A2(new_n9774_), .B(new_n9637_), .ZN(new_n9775_));
  INV_X1     g09583(.I(new_n9756_), .ZN(new_n9776_));
  OAI21_X1   g09584(.A1(new_n9773_), .A2(new_n9776_), .B(\asqrt[33] ), .ZN(new_n9777_));
  NAND3_X1   g09585(.A1(new_n9775_), .A2(new_n9777_), .A3(new_n4810_), .ZN(new_n9778_));
  NAND2_X1   g09586(.A1(new_n9778_), .A2(new_n9634_), .ZN(new_n9779_));
  NAND2_X1   g09587(.A1(new_n9775_), .A2(new_n9777_), .ZN(new_n9780_));
  AOI21_X1   g09588(.A1(new_n9780_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n9781_));
  AOI21_X1   g09589(.A1(new_n9781_), .A2(new_n9779_), .B(new_n9770_), .ZN(new_n9782_));
  AOI21_X1   g09590(.A1(new_n9779_), .A2(new_n9760_), .B(new_n4510_), .ZN(new_n9783_));
  OAI21_X1   g09591(.A1(new_n9782_), .A2(new_n9783_), .B(\asqrt[36] ), .ZN(new_n9784_));
  AOI21_X1   g09592(.A1(new_n9766_), .A2(new_n9784_), .B(new_n3928_), .ZN(new_n9785_));
  NOR2_X1    g09593(.A1(new_n9769_), .A2(new_n9785_), .ZN(new_n9786_));
  AOI21_X1   g09594(.A1(new_n9786_), .A2(new_n3675_), .B(new_n9623_), .ZN(new_n9787_));
  OAI21_X1   g09595(.A1(new_n9769_), .A2(new_n9785_), .B(\asqrt[38] ), .ZN(new_n9788_));
  NAND2_X1   g09596(.A1(new_n9788_), .A2(new_n3400_), .ZN(new_n9789_));
  OAI21_X1   g09597(.A1(new_n9787_), .A2(new_n9789_), .B(new_n9619_), .ZN(new_n9790_));
  INV_X1     g09598(.I(new_n9788_), .ZN(new_n9791_));
  OAI21_X1   g09599(.A1(new_n9787_), .A2(new_n9791_), .B(\asqrt[39] ), .ZN(new_n9792_));
  NAND3_X1   g09600(.A1(new_n9790_), .A2(new_n9792_), .A3(new_n3167_), .ZN(new_n9793_));
  NAND2_X1   g09601(.A1(new_n9793_), .A2(new_n9617_), .ZN(new_n9794_));
  NAND2_X1   g09602(.A1(new_n9790_), .A2(new_n9792_), .ZN(new_n9795_));
  AOI21_X1   g09603(.A1(new_n9795_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n9796_));
  AOI21_X1   g09604(.A1(new_n9796_), .A2(new_n9794_), .B(new_n9614_), .ZN(new_n9797_));
  INV_X1     g09605(.I(new_n9619_), .ZN(new_n9798_));
  INV_X1     g09606(.I(new_n9629_), .ZN(new_n9799_));
  NOR2_X1    g09607(.A1(new_n9782_), .A2(new_n9783_), .ZN(new_n9800_));
  AOI21_X1   g09608(.A1(new_n9800_), .A2(new_n4224_), .B(new_n9799_), .ZN(new_n9801_));
  NAND2_X1   g09609(.A1(new_n9784_), .A2(new_n3928_), .ZN(new_n9802_));
  OAI21_X1   g09610(.A1(new_n9801_), .A2(new_n9802_), .B(new_n9625_), .ZN(new_n9803_));
  INV_X1     g09611(.I(new_n9784_), .ZN(new_n9804_));
  OAI21_X1   g09612(.A1(new_n9801_), .A2(new_n9804_), .B(\asqrt[37] ), .ZN(new_n9805_));
  NAND3_X1   g09613(.A1(new_n9803_), .A2(new_n9805_), .A3(new_n3675_), .ZN(new_n9806_));
  NAND2_X1   g09614(.A1(new_n9806_), .A2(new_n9622_), .ZN(new_n9807_));
  NAND2_X1   g09615(.A1(new_n9803_), .A2(new_n9805_), .ZN(new_n9808_));
  AOI21_X1   g09616(.A1(new_n9808_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n9809_));
  AOI21_X1   g09617(.A1(new_n9809_), .A2(new_n9807_), .B(new_n9798_), .ZN(new_n9810_));
  AOI21_X1   g09618(.A1(new_n9807_), .A2(new_n9788_), .B(new_n3400_), .ZN(new_n9811_));
  OAI21_X1   g09619(.A1(new_n9810_), .A2(new_n9811_), .B(\asqrt[40] ), .ZN(new_n9812_));
  AOI21_X1   g09620(.A1(new_n9794_), .A2(new_n9812_), .B(new_n2912_), .ZN(new_n9813_));
  NOR2_X1    g09621(.A1(new_n9797_), .A2(new_n9813_), .ZN(new_n9814_));
  AOI21_X1   g09622(.A1(new_n9814_), .A2(new_n2699_), .B(new_n9611_), .ZN(new_n9815_));
  OAI21_X1   g09623(.A1(new_n9797_), .A2(new_n9813_), .B(\asqrt[42] ), .ZN(new_n9816_));
  NAND2_X1   g09624(.A1(new_n9816_), .A2(new_n2464_), .ZN(new_n9817_));
  OAI21_X1   g09625(.A1(new_n9815_), .A2(new_n9817_), .B(new_n9607_), .ZN(new_n9818_));
  INV_X1     g09626(.I(new_n9816_), .ZN(new_n9819_));
  OAI21_X1   g09627(.A1(new_n9815_), .A2(new_n9819_), .B(\asqrt[43] ), .ZN(new_n9820_));
  NAND3_X1   g09628(.A1(new_n9818_), .A2(new_n9820_), .A3(new_n2271_), .ZN(new_n9821_));
  INV_X1     g09629(.I(new_n9607_), .ZN(new_n9822_));
  INV_X1     g09630(.I(new_n9617_), .ZN(new_n9823_));
  NOR2_X1    g09631(.A1(new_n9810_), .A2(new_n9811_), .ZN(new_n9824_));
  AOI21_X1   g09632(.A1(new_n9824_), .A2(new_n3167_), .B(new_n9823_), .ZN(new_n9825_));
  NAND2_X1   g09633(.A1(new_n9812_), .A2(new_n2912_), .ZN(new_n9826_));
  OAI21_X1   g09634(.A1(new_n9825_), .A2(new_n9826_), .B(new_n9613_), .ZN(new_n9827_));
  INV_X1     g09635(.I(new_n9812_), .ZN(new_n9828_));
  OAI21_X1   g09636(.A1(new_n9825_), .A2(new_n9828_), .B(\asqrt[41] ), .ZN(new_n9829_));
  NAND3_X1   g09637(.A1(new_n9827_), .A2(new_n9829_), .A3(new_n2699_), .ZN(new_n9830_));
  NAND2_X1   g09638(.A1(new_n9830_), .A2(new_n9610_), .ZN(new_n9831_));
  NAND2_X1   g09639(.A1(new_n9827_), .A2(new_n9829_), .ZN(new_n9832_));
  AOI21_X1   g09640(.A1(new_n9832_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n9833_));
  AOI21_X1   g09641(.A1(new_n9833_), .A2(new_n9831_), .B(new_n9822_), .ZN(new_n9834_));
  AOI21_X1   g09642(.A1(new_n9831_), .A2(new_n9816_), .B(new_n2464_), .ZN(new_n9835_));
  OAI21_X1   g09643(.A1(new_n9834_), .A2(new_n9835_), .B(\asqrt[44] ), .ZN(new_n9836_));
  NAND2_X1   g09644(.A1(new_n9587_), .A2(new_n9182_), .ZN(new_n9837_));
  NOR2_X1    g09645(.A1(new_n9590_), .A2(new_n9182_), .ZN(new_n9838_));
  NAND2_X1   g09646(.A1(new_n9838_), .A2(new_n9602_), .ZN(new_n9839_));
  AOI21_X1   g09647(.A1(new_n9839_), .A2(new_n9837_), .B(new_n193_), .ZN(new_n9840_));
  INV_X1     g09648(.I(new_n9840_), .ZN(new_n9841_));
  NAND3_X1   g09649(.A1(\asqrt[21] ), .A2(new_n9572_), .A3(new_n9583_), .ZN(new_n9842_));
  XOR2_X1    g09650(.A1(new_n9842_), .A2(new_n9575_), .Z(new_n9843_));
  AOI21_X1   g09651(.A1(new_n9838_), .A2(new_n9587_), .B(new_n9588_), .ZN(new_n9844_));
  OAI21_X1   g09652(.A1(new_n9542_), .A2(new_n9544_), .B(new_n9547_), .ZN(new_n9845_));
  NOR2_X1    g09653(.A1(new_n9590_), .A2(new_n9845_), .ZN(new_n9846_));
  XOR2_X1    g09654(.A1(new_n9846_), .A2(new_n9190_), .Z(new_n9847_));
  NAND3_X1   g09655(.A1(\asqrt[21] ), .A2(new_n9558_), .A3(new_n9543_), .ZN(new_n9848_));
  XOR2_X1    g09656(.A1(new_n9848_), .A2(new_n9194_), .Z(new_n9849_));
  OAI21_X1   g09657(.A1(new_n9553_), .A2(new_n9554_), .B(new_n9557_), .ZN(new_n9850_));
  NOR2_X1    g09658(.A1(new_n9590_), .A2(new_n9850_), .ZN(new_n9851_));
  XOR2_X1    g09659(.A1(new_n9851_), .A2(new_n9196_), .Z(new_n9852_));
  INV_X1     g09660(.I(new_n9852_), .ZN(new_n9853_));
  NAND3_X1   g09661(.A1(\asqrt[21] ), .A2(new_n9520_), .A3(new_n9539_), .ZN(new_n9854_));
  XOR2_X1    g09662(.A1(new_n9854_), .A2(new_n9551_), .Z(new_n9855_));
  INV_X1     g09663(.I(new_n9855_), .ZN(new_n9856_));
  OAI21_X1   g09664(.A1(new_n9514_), .A2(new_n9516_), .B(new_n9519_), .ZN(new_n9857_));
  NOR2_X1    g09665(.A1(new_n9590_), .A2(new_n9857_), .ZN(new_n9858_));
  XOR2_X1    g09666(.A1(new_n9858_), .A2(new_n9202_), .Z(new_n9859_));
  NAND3_X1   g09667(.A1(\asqrt[21] ), .A2(new_n9533_), .A3(new_n9515_), .ZN(new_n9860_));
  XOR2_X1    g09668(.A1(new_n9860_), .A2(new_n9206_), .Z(new_n9861_));
  OAI21_X1   g09669(.A1(new_n9528_), .A2(new_n9529_), .B(new_n9532_), .ZN(new_n9862_));
  NOR2_X1    g09670(.A1(new_n9590_), .A2(new_n9862_), .ZN(new_n9863_));
  XOR2_X1    g09671(.A1(new_n9863_), .A2(new_n9208_), .Z(new_n9864_));
  INV_X1     g09672(.I(new_n9864_), .ZN(new_n9865_));
  NAND3_X1   g09673(.A1(\asqrt[21] ), .A2(new_n9492_), .A3(new_n9511_), .ZN(new_n9866_));
  XOR2_X1    g09674(.A1(new_n9866_), .A2(new_n9526_), .Z(new_n9867_));
  INV_X1     g09675(.I(new_n9867_), .ZN(new_n9868_));
  OAI21_X1   g09676(.A1(new_n9486_), .A2(new_n9488_), .B(new_n9491_), .ZN(new_n9869_));
  NOR2_X1    g09677(.A1(new_n9590_), .A2(new_n9869_), .ZN(new_n9870_));
  XOR2_X1    g09678(.A1(new_n9870_), .A2(new_n9214_), .Z(new_n9871_));
  NAND3_X1   g09679(.A1(\asqrt[21] ), .A2(new_n9505_), .A3(new_n9487_), .ZN(new_n9872_));
  XOR2_X1    g09680(.A1(new_n9872_), .A2(new_n9218_), .Z(new_n9873_));
  OAI21_X1   g09681(.A1(new_n9500_), .A2(new_n9501_), .B(new_n9504_), .ZN(new_n9874_));
  NOR2_X1    g09682(.A1(new_n9590_), .A2(new_n9874_), .ZN(new_n9875_));
  XOR2_X1    g09683(.A1(new_n9875_), .A2(new_n9220_), .Z(new_n9876_));
  INV_X1     g09684(.I(new_n9876_), .ZN(new_n9877_));
  NAND3_X1   g09685(.A1(\asqrt[21] ), .A2(new_n9464_), .A3(new_n9483_), .ZN(new_n9878_));
  XOR2_X1    g09686(.A1(new_n9878_), .A2(new_n9498_), .Z(new_n9879_));
  INV_X1     g09687(.I(new_n9879_), .ZN(new_n9880_));
  OAI21_X1   g09688(.A1(new_n9458_), .A2(new_n9460_), .B(new_n9463_), .ZN(new_n9881_));
  NOR2_X1    g09689(.A1(new_n9590_), .A2(new_n9881_), .ZN(new_n9882_));
  XOR2_X1    g09690(.A1(new_n9882_), .A2(new_n9226_), .Z(new_n9883_));
  NAND3_X1   g09691(.A1(\asqrt[21] ), .A2(new_n9477_), .A3(new_n9459_), .ZN(new_n9884_));
  XOR2_X1    g09692(.A1(new_n9884_), .A2(new_n9230_), .Z(new_n9885_));
  OAI21_X1   g09693(.A1(new_n9472_), .A2(new_n9473_), .B(new_n9476_), .ZN(new_n9886_));
  NOR2_X1    g09694(.A1(new_n9590_), .A2(new_n9886_), .ZN(new_n9887_));
  XOR2_X1    g09695(.A1(new_n9887_), .A2(new_n9232_), .Z(new_n9888_));
  INV_X1     g09696(.I(new_n9888_), .ZN(new_n9889_));
  NAND3_X1   g09697(.A1(\asqrt[21] ), .A2(new_n9436_), .A3(new_n9455_), .ZN(new_n9890_));
  XOR2_X1    g09698(.A1(new_n9890_), .A2(new_n9470_), .Z(new_n9891_));
  INV_X1     g09699(.I(new_n9891_), .ZN(new_n9892_));
  NAND2_X1   g09700(.A1(new_n9821_), .A2(new_n9593_), .ZN(new_n9893_));
  NAND2_X1   g09701(.A1(new_n9818_), .A2(new_n9820_), .ZN(new_n9894_));
  AOI21_X1   g09702(.A1(new_n9894_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n9895_));
  AOI21_X1   g09703(.A1(new_n9895_), .A2(new_n9893_), .B(new_n9892_), .ZN(new_n9896_));
  AOI21_X1   g09704(.A1(new_n9893_), .A2(new_n9836_), .B(new_n2072_), .ZN(new_n9897_));
  NOR2_X1    g09705(.A1(new_n9896_), .A2(new_n9897_), .ZN(new_n9898_));
  AOI21_X1   g09706(.A1(new_n9898_), .A2(new_n1884_), .B(new_n9889_), .ZN(new_n9899_));
  OAI21_X1   g09707(.A1(new_n9896_), .A2(new_n9897_), .B(\asqrt[46] ), .ZN(new_n9900_));
  NAND2_X1   g09708(.A1(new_n9900_), .A2(new_n1688_), .ZN(new_n9901_));
  OAI21_X1   g09709(.A1(new_n9899_), .A2(new_n9901_), .B(new_n9885_), .ZN(new_n9902_));
  INV_X1     g09710(.I(new_n9900_), .ZN(new_n9903_));
  OAI21_X1   g09711(.A1(new_n9899_), .A2(new_n9903_), .B(\asqrt[47] ), .ZN(new_n9904_));
  NAND3_X1   g09712(.A1(new_n9902_), .A2(new_n9904_), .A3(new_n1533_), .ZN(new_n9905_));
  NAND2_X1   g09713(.A1(new_n9905_), .A2(new_n9883_), .ZN(new_n9906_));
  NAND2_X1   g09714(.A1(new_n9902_), .A2(new_n9904_), .ZN(new_n9907_));
  AOI21_X1   g09715(.A1(new_n9907_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n9908_));
  AOI21_X1   g09716(.A1(new_n9908_), .A2(new_n9906_), .B(new_n9880_), .ZN(new_n9909_));
  INV_X1     g09717(.I(new_n9885_), .ZN(new_n9910_));
  NOR2_X1    g09718(.A1(new_n9834_), .A2(new_n9835_), .ZN(new_n9911_));
  AOI21_X1   g09719(.A1(new_n9911_), .A2(new_n2271_), .B(new_n9594_), .ZN(new_n9912_));
  NAND2_X1   g09720(.A1(new_n9836_), .A2(new_n2072_), .ZN(new_n9913_));
  OAI21_X1   g09721(.A1(new_n9912_), .A2(new_n9913_), .B(new_n9891_), .ZN(new_n9914_));
  INV_X1     g09722(.I(new_n9836_), .ZN(new_n9915_));
  OAI21_X1   g09723(.A1(new_n9912_), .A2(new_n9915_), .B(\asqrt[45] ), .ZN(new_n9916_));
  NAND3_X1   g09724(.A1(new_n9914_), .A2(new_n9916_), .A3(new_n1884_), .ZN(new_n9917_));
  NAND2_X1   g09725(.A1(new_n9917_), .A2(new_n9888_), .ZN(new_n9918_));
  NAND2_X1   g09726(.A1(new_n9914_), .A2(new_n9916_), .ZN(new_n9919_));
  AOI21_X1   g09727(.A1(new_n9919_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n9920_));
  AOI21_X1   g09728(.A1(new_n9920_), .A2(new_n9918_), .B(new_n9910_), .ZN(new_n9921_));
  AOI21_X1   g09729(.A1(new_n9918_), .A2(new_n9900_), .B(new_n1688_), .ZN(new_n9922_));
  OAI21_X1   g09730(.A1(new_n9921_), .A2(new_n9922_), .B(\asqrt[48] ), .ZN(new_n9923_));
  AOI21_X1   g09731(.A1(new_n9906_), .A2(new_n9923_), .B(new_n1368_), .ZN(new_n9924_));
  NOR2_X1    g09732(.A1(new_n9909_), .A2(new_n9924_), .ZN(new_n9925_));
  AOI21_X1   g09733(.A1(new_n9925_), .A2(new_n1228_), .B(new_n9877_), .ZN(new_n9926_));
  OAI21_X1   g09734(.A1(new_n9909_), .A2(new_n9924_), .B(\asqrt[50] ), .ZN(new_n9927_));
  NAND2_X1   g09735(.A1(new_n9927_), .A2(new_n1088_), .ZN(new_n9928_));
  OAI21_X1   g09736(.A1(new_n9926_), .A2(new_n9928_), .B(new_n9873_), .ZN(new_n9929_));
  INV_X1     g09737(.I(new_n9927_), .ZN(new_n9930_));
  OAI21_X1   g09738(.A1(new_n9926_), .A2(new_n9930_), .B(\asqrt[51] ), .ZN(new_n9931_));
  NAND3_X1   g09739(.A1(new_n9929_), .A2(new_n9931_), .A3(new_n962_), .ZN(new_n9932_));
  NAND2_X1   g09740(.A1(new_n9932_), .A2(new_n9871_), .ZN(new_n9933_));
  NAND2_X1   g09741(.A1(new_n9929_), .A2(new_n9931_), .ZN(new_n9934_));
  AOI21_X1   g09742(.A1(new_n9934_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n9935_));
  AOI21_X1   g09743(.A1(new_n9935_), .A2(new_n9933_), .B(new_n9868_), .ZN(new_n9936_));
  INV_X1     g09744(.I(new_n9873_), .ZN(new_n9937_));
  INV_X1     g09745(.I(new_n9883_), .ZN(new_n9938_));
  NOR2_X1    g09746(.A1(new_n9921_), .A2(new_n9922_), .ZN(new_n9939_));
  AOI21_X1   g09747(.A1(new_n9939_), .A2(new_n1533_), .B(new_n9938_), .ZN(new_n9940_));
  NAND2_X1   g09748(.A1(new_n9923_), .A2(new_n1368_), .ZN(new_n9941_));
  OAI21_X1   g09749(.A1(new_n9940_), .A2(new_n9941_), .B(new_n9879_), .ZN(new_n9942_));
  INV_X1     g09750(.I(new_n9923_), .ZN(new_n9943_));
  OAI21_X1   g09751(.A1(new_n9940_), .A2(new_n9943_), .B(\asqrt[49] ), .ZN(new_n9944_));
  NAND3_X1   g09752(.A1(new_n9942_), .A2(new_n9944_), .A3(new_n1228_), .ZN(new_n9945_));
  NAND2_X1   g09753(.A1(new_n9945_), .A2(new_n9876_), .ZN(new_n9946_));
  NAND2_X1   g09754(.A1(new_n9942_), .A2(new_n9944_), .ZN(new_n9947_));
  AOI21_X1   g09755(.A1(new_n9947_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n9948_));
  AOI21_X1   g09756(.A1(new_n9948_), .A2(new_n9946_), .B(new_n9937_), .ZN(new_n9949_));
  AOI21_X1   g09757(.A1(new_n9946_), .A2(new_n9927_), .B(new_n1088_), .ZN(new_n9950_));
  OAI21_X1   g09758(.A1(new_n9949_), .A2(new_n9950_), .B(\asqrt[52] ), .ZN(new_n9951_));
  AOI21_X1   g09759(.A1(new_n9933_), .A2(new_n9951_), .B(new_n842_), .ZN(new_n9952_));
  NOR2_X1    g09760(.A1(new_n9936_), .A2(new_n9952_), .ZN(new_n9953_));
  AOI21_X1   g09761(.A1(new_n9953_), .A2(new_n720_), .B(new_n9865_), .ZN(new_n9954_));
  OAI21_X1   g09762(.A1(new_n9936_), .A2(new_n9952_), .B(\asqrt[54] ), .ZN(new_n9955_));
  NAND2_X1   g09763(.A1(new_n9955_), .A2(new_n630_), .ZN(new_n9956_));
  OAI21_X1   g09764(.A1(new_n9954_), .A2(new_n9956_), .B(new_n9861_), .ZN(new_n9957_));
  INV_X1     g09765(.I(new_n9955_), .ZN(new_n9958_));
  OAI21_X1   g09766(.A1(new_n9954_), .A2(new_n9958_), .B(\asqrt[55] ), .ZN(new_n9959_));
  NAND3_X1   g09767(.A1(new_n9957_), .A2(new_n9959_), .A3(new_n545_), .ZN(new_n9960_));
  NAND2_X1   g09768(.A1(new_n9960_), .A2(new_n9859_), .ZN(new_n9961_));
  NAND2_X1   g09769(.A1(new_n9957_), .A2(new_n9959_), .ZN(new_n9962_));
  AOI21_X1   g09770(.A1(new_n9962_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n9963_));
  AOI21_X1   g09771(.A1(new_n9963_), .A2(new_n9961_), .B(new_n9856_), .ZN(new_n9964_));
  INV_X1     g09772(.I(new_n9861_), .ZN(new_n9965_));
  INV_X1     g09773(.I(new_n9871_), .ZN(new_n9966_));
  NOR2_X1    g09774(.A1(new_n9949_), .A2(new_n9950_), .ZN(new_n9967_));
  AOI21_X1   g09775(.A1(new_n9967_), .A2(new_n962_), .B(new_n9966_), .ZN(new_n9968_));
  NAND2_X1   g09776(.A1(new_n9951_), .A2(new_n842_), .ZN(new_n9969_));
  OAI21_X1   g09777(.A1(new_n9968_), .A2(new_n9969_), .B(new_n9867_), .ZN(new_n9970_));
  INV_X1     g09778(.I(new_n9951_), .ZN(new_n9971_));
  OAI21_X1   g09779(.A1(new_n9968_), .A2(new_n9971_), .B(\asqrt[53] ), .ZN(new_n9972_));
  NAND3_X1   g09780(.A1(new_n9970_), .A2(new_n9972_), .A3(new_n720_), .ZN(new_n9973_));
  NAND2_X1   g09781(.A1(new_n9973_), .A2(new_n9864_), .ZN(new_n9974_));
  NAND2_X1   g09782(.A1(new_n9970_), .A2(new_n9972_), .ZN(new_n9975_));
  AOI21_X1   g09783(.A1(new_n9975_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n9976_));
  AOI21_X1   g09784(.A1(new_n9976_), .A2(new_n9974_), .B(new_n9965_), .ZN(new_n9977_));
  AOI21_X1   g09785(.A1(new_n9974_), .A2(new_n9955_), .B(new_n630_), .ZN(new_n9978_));
  OAI21_X1   g09786(.A1(new_n9977_), .A2(new_n9978_), .B(\asqrt[56] ), .ZN(new_n9979_));
  AOI21_X1   g09787(.A1(new_n9961_), .A2(new_n9979_), .B(new_n450_), .ZN(new_n9980_));
  NOR2_X1    g09788(.A1(new_n9964_), .A2(new_n9980_), .ZN(new_n9981_));
  AOI21_X1   g09789(.A1(new_n9981_), .A2(new_n403_), .B(new_n9853_), .ZN(new_n9982_));
  OAI21_X1   g09790(.A1(new_n9964_), .A2(new_n9980_), .B(\asqrt[58] ), .ZN(new_n9983_));
  NAND2_X1   g09791(.A1(new_n9983_), .A2(new_n339_), .ZN(new_n9984_));
  OAI21_X1   g09792(.A1(new_n9982_), .A2(new_n9984_), .B(new_n9849_), .ZN(new_n9985_));
  INV_X1     g09793(.I(new_n9983_), .ZN(new_n9986_));
  OAI21_X1   g09794(.A1(new_n9982_), .A2(new_n9986_), .B(\asqrt[59] ), .ZN(new_n9987_));
  NAND3_X1   g09795(.A1(new_n9985_), .A2(new_n9987_), .A3(new_n288_), .ZN(new_n9988_));
  NAND2_X1   g09796(.A1(new_n9988_), .A2(new_n9847_), .ZN(new_n9989_));
  INV_X1     g09797(.I(new_n9849_), .ZN(new_n9990_));
  INV_X1     g09798(.I(new_n9859_), .ZN(new_n9991_));
  NOR2_X1    g09799(.A1(new_n9977_), .A2(new_n9978_), .ZN(new_n9992_));
  AOI21_X1   g09800(.A1(new_n9992_), .A2(new_n545_), .B(new_n9991_), .ZN(new_n9993_));
  NAND2_X1   g09801(.A1(new_n9979_), .A2(new_n450_), .ZN(new_n9994_));
  OAI21_X1   g09802(.A1(new_n9993_), .A2(new_n9994_), .B(new_n9855_), .ZN(new_n9995_));
  INV_X1     g09803(.I(new_n9979_), .ZN(new_n9996_));
  OAI21_X1   g09804(.A1(new_n9993_), .A2(new_n9996_), .B(\asqrt[57] ), .ZN(new_n9997_));
  NAND3_X1   g09805(.A1(new_n9995_), .A2(new_n9997_), .A3(new_n403_), .ZN(new_n9998_));
  NAND2_X1   g09806(.A1(new_n9998_), .A2(new_n9852_), .ZN(new_n9999_));
  NAND2_X1   g09807(.A1(new_n9995_), .A2(new_n9997_), .ZN(new_n10000_));
  AOI21_X1   g09808(.A1(new_n10000_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n10001_));
  AOI21_X1   g09809(.A1(new_n10001_), .A2(new_n9999_), .B(new_n9990_), .ZN(new_n10002_));
  AOI21_X1   g09810(.A1(new_n9999_), .A2(new_n9983_), .B(new_n339_), .ZN(new_n10003_));
  OAI21_X1   g09811(.A1(new_n10002_), .A2(new_n10003_), .B(\asqrt[60] ), .ZN(new_n10004_));
  AOI21_X1   g09812(.A1(new_n9989_), .A2(new_n10004_), .B(new_n242_), .ZN(new_n10005_));
  NAND3_X1   g09813(.A1(\asqrt[21] ), .A2(new_n9548_), .A3(new_n9564_), .ZN(new_n10006_));
  XOR2_X1    g09814(.A1(new_n10006_), .A2(new_n9576_), .Z(new_n10007_));
  INV_X1     g09815(.I(new_n10007_), .ZN(new_n10008_));
  NAND2_X1   g09816(.A1(new_n9985_), .A2(new_n9987_), .ZN(new_n10009_));
  AOI21_X1   g09817(.A1(new_n10009_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n10010_));
  AOI21_X1   g09818(.A1(new_n10010_), .A2(new_n9989_), .B(new_n10008_), .ZN(new_n10011_));
  OAI21_X1   g09819(.A1(new_n10011_), .A2(new_n10005_), .B(\asqrt[62] ), .ZN(new_n10012_));
  INV_X1     g09820(.I(new_n10012_), .ZN(new_n10013_));
  NOR2_X1    g09821(.A1(new_n10011_), .A2(new_n10005_), .ZN(new_n10014_));
  AOI21_X1   g09822(.A1(new_n9549_), .A2(new_n9570_), .B(new_n9565_), .ZN(new_n10015_));
  NAND2_X1   g09823(.A1(\asqrt[21] ), .A2(new_n10015_), .ZN(new_n10016_));
  XOR2_X1    g09824(.A1(new_n10016_), .A2(new_n9568_), .Z(new_n10017_));
  INV_X1     g09825(.I(new_n10017_), .ZN(new_n10018_));
  AOI21_X1   g09826(.A1(new_n10014_), .A2(new_n234_), .B(new_n10018_), .ZN(new_n10019_));
  OAI21_X1   g09827(.A1(new_n10019_), .A2(new_n10013_), .B(new_n9844_), .ZN(new_n10020_));
  OAI21_X1   g09828(.A1(new_n10020_), .A2(new_n9843_), .B(new_n193_), .ZN(new_n10021_));
  NOR2_X1    g09829(.A1(new_n10019_), .A2(new_n10013_), .ZN(new_n10022_));
  NAND2_X1   g09830(.A1(new_n10022_), .A2(new_n9843_), .ZN(new_n10023_));
  NOR2_X1    g09831(.A1(\asqrt[21] ), .A2(new_n9183_), .ZN(new_n10024_));
  INV_X1     g09832(.I(new_n10024_), .ZN(new_n10025_));
  NAND4_X1   g09833(.A1(new_n10021_), .A2(new_n9841_), .A3(new_n10023_), .A4(new_n10025_), .ZN(\asqrt[20] ));
  NAND3_X1   g09834(.A1(\asqrt[20] ), .A2(new_n9821_), .A3(new_n9836_), .ZN(new_n10027_));
  XOR2_X1    g09835(.A1(new_n10027_), .A2(new_n9594_), .Z(new_n10028_));
  INV_X1     g09836(.I(new_n9847_), .ZN(new_n10029_));
  NOR2_X1    g09837(.A1(new_n10002_), .A2(new_n10003_), .ZN(new_n10030_));
  AOI21_X1   g09838(.A1(new_n10030_), .A2(new_n288_), .B(new_n10029_), .ZN(new_n10031_));
  INV_X1     g09839(.I(new_n10004_), .ZN(new_n10032_));
  OAI21_X1   g09840(.A1(new_n10031_), .A2(new_n10032_), .B(\asqrt[61] ), .ZN(new_n10033_));
  NAND2_X1   g09841(.A1(new_n10004_), .A2(new_n242_), .ZN(new_n10034_));
  OAI21_X1   g09842(.A1(new_n10031_), .A2(new_n10034_), .B(new_n10007_), .ZN(new_n10035_));
  NAND3_X1   g09843(.A1(new_n10035_), .A2(new_n10033_), .A3(new_n234_), .ZN(new_n10036_));
  NAND2_X1   g09844(.A1(new_n10036_), .A2(new_n10017_), .ZN(new_n10037_));
  NAND2_X1   g09845(.A1(new_n10037_), .A2(new_n10012_), .ZN(new_n10038_));
  NAND2_X1   g09846(.A1(new_n10038_), .A2(new_n9843_), .ZN(new_n10039_));
  INV_X1     g09847(.I(new_n9843_), .ZN(new_n10040_));
  INV_X1     g09848(.I(new_n9844_), .ZN(new_n10041_));
  AOI21_X1   g09849(.A1(new_n10037_), .A2(new_n10012_), .B(new_n10041_), .ZN(new_n10042_));
  AOI21_X1   g09850(.A1(new_n10042_), .A2(new_n10040_), .B(\asqrt[63] ), .ZN(new_n10043_));
  NOR2_X1    g09851(.A1(new_n10038_), .A2(new_n10040_), .ZN(new_n10044_));
  NOR4_X1    g09852(.A1(new_n10043_), .A2(new_n9840_), .A3(new_n10044_), .A4(new_n10024_), .ZN(new_n10045_));
  NOR2_X1    g09853(.A1(new_n10045_), .A2(new_n9843_), .ZN(new_n10046_));
  NAND2_X1   g09854(.A1(new_n10046_), .A2(new_n10022_), .ZN(new_n10047_));
  AOI21_X1   g09855(.A1(new_n10047_), .A2(new_n10039_), .B(new_n193_), .ZN(new_n10048_));
  NAND3_X1   g09856(.A1(\asqrt[20] ), .A2(new_n10012_), .A3(new_n10036_), .ZN(new_n10049_));
  XOR2_X1    g09857(.A1(new_n10049_), .A2(new_n10017_), .Z(new_n10050_));
  INV_X1     g09858(.I(new_n10050_), .ZN(new_n10051_));
  AOI21_X1   g09859(.A1(new_n10046_), .A2(new_n10038_), .B(new_n10044_), .ZN(new_n10052_));
  INV_X1     g09860(.I(new_n10052_), .ZN(new_n10053_));
  OAI21_X1   g09861(.A1(new_n9982_), .A2(new_n9984_), .B(new_n9987_), .ZN(new_n10054_));
  NOR2_X1    g09862(.A1(new_n10045_), .A2(new_n10054_), .ZN(new_n10055_));
  XOR2_X1    g09863(.A1(new_n10055_), .A2(new_n9849_), .Z(new_n10056_));
  NAND3_X1   g09864(.A1(\asqrt[20] ), .A2(new_n9998_), .A3(new_n9983_), .ZN(new_n10057_));
  XOR2_X1    g09865(.A1(new_n10057_), .A2(new_n9853_), .Z(new_n10058_));
  OAI21_X1   g09866(.A1(new_n9993_), .A2(new_n9994_), .B(new_n9997_), .ZN(new_n10059_));
  NOR2_X1    g09867(.A1(new_n10045_), .A2(new_n10059_), .ZN(new_n10060_));
  XOR2_X1    g09868(.A1(new_n10060_), .A2(new_n9855_), .Z(new_n10061_));
  INV_X1     g09869(.I(new_n10061_), .ZN(new_n10062_));
  NAND3_X1   g09870(.A1(\asqrt[20] ), .A2(new_n9960_), .A3(new_n9979_), .ZN(new_n10063_));
  XOR2_X1    g09871(.A1(new_n10063_), .A2(new_n9991_), .Z(new_n10064_));
  INV_X1     g09872(.I(new_n10064_), .ZN(new_n10065_));
  OAI21_X1   g09873(.A1(new_n9954_), .A2(new_n9956_), .B(new_n9959_), .ZN(new_n10066_));
  NOR2_X1    g09874(.A1(new_n10045_), .A2(new_n10066_), .ZN(new_n10067_));
  XOR2_X1    g09875(.A1(new_n10067_), .A2(new_n9861_), .Z(new_n10068_));
  NAND3_X1   g09876(.A1(\asqrt[20] ), .A2(new_n9973_), .A3(new_n9955_), .ZN(new_n10069_));
  XOR2_X1    g09877(.A1(new_n10069_), .A2(new_n9865_), .Z(new_n10070_));
  OAI21_X1   g09878(.A1(new_n9968_), .A2(new_n9969_), .B(new_n9972_), .ZN(new_n10071_));
  NOR2_X1    g09879(.A1(new_n10045_), .A2(new_n10071_), .ZN(new_n10072_));
  XOR2_X1    g09880(.A1(new_n10072_), .A2(new_n9867_), .Z(new_n10073_));
  INV_X1     g09881(.I(new_n10073_), .ZN(new_n10074_));
  NAND3_X1   g09882(.A1(\asqrt[20] ), .A2(new_n9932_), .A3(new_n9951_), .ZN(new_n10075_));
  XOR2_X1    g09883(.A1(new_n10075_), .A2(new_n9966_), .Z(new_n10076_));
  INV_X1     g09884(.I(new_n10076_), .ZN(new_n10077_));
  OAI21_X1   g09885(.A1(new_n9926_), .A2(new_n9928_), .B(new_n9931_), .ZN(new_n10078_));
  NOR2_X1    g09886(.A1(new_n10045_), .A2(new_n10078_), .ZN(new_n10079_));
  XOR2_X1    g09887(.A1(new_n10079_), .A2(new_n9873_), .Z(new_n10080_));
  NAND3_X1   g09888(.A1(\asqrt[20] ), .A2(new_n9945_), .A3(new_n9927_), .ZN(new_n10081_));
  XOR2_X1    g09889(.A1(new_n10081_), .A2(new_n9877_), .Z(new_n10082_));
  OAI21_X1   g09890(.A1(new_n9940_), .A2(new_n9941_), .B(new_n9944_), .ZN(new_n10083_));
  NOR2_X1    g09891(.A1(new_n10045_), .A2(new_n10083_), .ZN(new_n10084_));
  XOR2_X1    g09892(.A1(new_n10084_), .A2(new_n9879_), .Z(new_n10085_));
  INV_X1     g09893(.I(new_n10085_), .ZN(new_n10086_));
  NAND3_X1   g09894(.A1(\asqrt[20] ), .A2(new_n9905_), .A3(new_n9923_), .ZN(new_n10087_));
  XOR2_X1    g09895(.A1(new_n10087_), .A2(new_n9938_), .Z(new_n10088_));
  INV_X1     g09896(.I(new_n10088_), .ZN(new_n10089_));
  OAI21_X1   g09897(.A1(new_n9899_), .A2(new_n9901_), .B(new_n9904_), .ZN(new_n10090_));
  NOR2_X1    g09898(.A1(new_n10045_), .A2(new_n10090_), .ZN(new_n10091_));
  XOR2_X1    g09899(.A1(new_n10091_), .A2(new_n9885_), .Z(new_n10092_));
  NAND3_X1   g09900(.A1(\asqrt[20] ), .A2(new_n9917_), .A3(new_n9900_), .ZN(new_n10093_));
  XOR2_X1    g09901(.A1(new_n10093_), .A2(new_n9889_), .Z(new_n10094_));
  OAI21_X1   g09902(.A1(new_n9912_), .A2(new_n9913_), .B(new_n9916_), .ZN(new_n10095_));
  NOR2_X1    g09903(.A1(new_n10045_), .A2(new_n10095_), .ZN(new_n10096_));
  XOR2_X1    g09904(.A1(new_n10096_), .A2(new_n9891_), .Z(new_n10097_));
  INV_X1     g09905(.I(new_n10097_), .ZN(new_n10098_));
  INV_X1     g09906(.I(new_n10028_), .ZN(new_n10099_));
  OAI21_X1   g09907(.A1(new_n9815_), .A2(new_n9817_), .B(new_n9820_), .ZN(new_n10100_));
  NOR2_X1    g09908(.A1(new_n10045_), .A2(new_n10100_), .ZN(new_n10101_));
  XOR2_X1    g09909(.A1(new_n10101_), .A2(new_n9607_), .Z(new_n10102_));
  NAND3_X1   g09910(.A1(\asqrt[20] ), .A2(new_n9830_), .A3(new_n9816_), .ZN(new_n10103_));
  XOR2_X1    g09911(.A1(new_n10103_), .A2(new_n9611_), .Z(new_n10104_));
  OAI21_X1   g09912(.A1(new_n9825_), .A2(new_n9826_), .B(new_n9829_), .ZN(new_n10105_));
  NOR2_X1    g09913(.A1(new_n10045_), .A2(new_n10105_), .ZN(new_n10106_));
  XOR2_X1    g09914(.A1(new_n10106_), .A2(new_n9613_), .Z(new_n10107_));
  INV_X1     g09915(.I(new_n10107_), .ZN(new_n10108_));
  NAND3_X1   g09916(.A1(\asqrt[20] ), .A2(new_n9793_), .A3(new_n9812_), .ZN(new_n10109_));
  XOR2_X1    g09917(.A1(new_n10109_), .A2(new_n9823_), .Z(new_n10110_));
  INV_X1     g09918(.I(new_n10110_), .ZN(new_n10111_));
  OAI21_X1   g09919(.A1(new_n9787_), .A2(new_n9789_), .B(new_n9792_), .ZN(new_n10112_));
  NOR2_X1    g09920(.A1(new_n10045_), .A2(new_n10112_), .ZN(new_n10113_));
  XOR2_X1    g09921(.A1(new_n10113_), .A2(new_n9619_), .Z(new_n10114_));
  NAND3_X1   g09922(.A1(\asqrt[20] ), .A2(new_n9806_), .A3(new_n9788_), .ZN(new_n10115_));
  XOR2_X1    g09923(.A1(new_n10115_), .A2(new_n9623_), .Z(new_n10116_));
  OAI21_X1   g09924(.A1(new_n9801_), .A2(new_n9802_), .B(new_n9805_), .ZN(new_n10117_));
  NOR2_X1    g09925(.A1(new_n10045_), .A2(new_n10117_), .ZN(new_n10118_));
  XOR2_X1    g09926(.A1(new_n10118_), .A2(new_n9625_), .Z(new_n10119_));
  INV_X1     g09927(.I(new_n10119_), .ZN(new_n10120_));
  NAND3_X1   g09928(.A1(\asqrt[20] ), .A2(new_n9765_), .A3(new_n9784_), .ZN(new_n10121_));
  XOR2_X1    g09929(.A1(new_n10121_), .A2(new_n9799_), .Z(new_n10122_));
  INV_X1     g09930(.I(new_n10122_), .ZN(new_n10123_));
  OAI21_X1   g09931(.A1(new_n9759_), .A2(new_n9761_), .B(new_n9764_), .ZN(new_n10124_));
  NOR2_X1    g09932(.A1(new_n10045_), .A2(new_n10124_), .ZN(new_n10125_));
  XOR2_X1    g09933(.A1(new_n10125_), .A2(new_n9631_), .Z(new_n10126_));
  NAND3_X1   g09934(.A1(\asqrt[20] ), .A2(new_n9778_), .A3(new_n9760_), .ZN(new_n10127_));
  XOR2_X1    g09935(.A1(new_n10127_), .A2(new_n9635_), .Z(new_n10128_));
  OAI21_X1   g09936(.A1(new_n9773_), .A2(new_n9774_), .B(new_n9777_), .ZN(new_n10129_));
  NOR2_X1    g09937(.A1(new_n10045_), .A2(new_n10129_), .ZN(new_n10130_));
  XOR2_X1    g09938(.A1(new_n10130_), .A2(new_n9637_), .Z(new_n10131_));
  INV_X1     g09939(.I(new_n10131_), .ZN(new_n10132_));
  NAND3_X1   g09940(.A1(\asqrt[20] ), .A2(new_n9737_), .A3(new_n9756_), .ZN(new_n10133_));
  XOR2_X1    g09941(.A1(new_n10133_), .A2(new_n9771_), .Z(new_n10134_));
  INV_X1     g09942(.I(new_n10134_), .ZN(new_n10135_));
  OAI21_X1   g09943(.A1(new_n9731_), .A2(new_n9733_), .B(new_n9736_), .ZN(new_n10136_));
  NOR2_X1    g09944(.A1(new_n10045_), .A2(new_n10136_), .ZN(new_n10137_));
  XOR2_X1    g09945(.A1(new_n10137_), .A2(new_n9643_), .Z(new_n10138_));
  NAND3_X1   g09946(.A1(\asqrt[20] ), .A2(new_n9750_), .A3(new_n9732_), .ZN(new_n10139_));
  XOR2_X1    g09947(.A1(new_n10139_), .A2(new_n9647_), .Z(new_n10140_));
  OAI21_X1   g09948(.A1(new_n9745_), .A2(new_n9746_), .B(new_n9749_), .ZN(new_n10141_));
  NOR2_X1    g09949(.A1(new_n10045_), .A2(new_n10141_), .ZN(new_n10142_));
  XOR2_X1    g09950(.A1(new_n10142_), .A2(new_n9649_), .Z(new_n10143_));
  INV_X1     g09951(.I(new_n10143_), .ZN(new_n10144_));
  NAND3_X1   g09952(.A1(\asqrt[20] ), .A2(new_n9709_), .A3(new_n9728_), .ZN(new_n10145_));
  XOR2_X1    g09953(.A1(new_n10145_), .A2(new_n9743_), .Z(new_n10146_));
  INV_X1     g09954(.I(new_n10146_), .ZN(new_n10147_));
  OAI21_X1   g09955(.A1(new_n9703_), .A2(new_n9705_), .B(new_n9708_), .ZN(new_n10148_));
  NOR2_X1    g09956(.A1(new_n10045_), .A2(new_n10148_), .ZN(new_n10149_));
  XOR2_X1    g09957(.A1(new_n10149_), .A2(new_n9656_), .Z(new_n10150_));
  NAND3_X1   g09958(.A1(\asqrt[20] ), .A2(new_n9722_), .A3(new_n9704_), .ZN(new_n10151_));
  XOR2_X1    g09959(.A1(new_n10151_), .A2(new_n9659_), .Z(new_n10152_));
  OAI21_X1   g09960(.A1(new_n9717_), .A2(new_n9718_), .B(new_n9721_), .ZN(new_n10153_));
  NOR2_X1    g09961(.A1(new_n10045_), .A2(new_n10153_), .ZN(new_n10154_));
  XOR2_X1    g09962(.A1(new_n10154_), .A2(new_n9662_), .Z(new_n10155_));
  INV_X1     g09963(.I(new_n10155_), .ZN(new_n10156_));
  NAND3_X1   g09964(.A1(\asqrt[20] ), .A2(new_n9682_), .A3(new_n9700_), .ZN(new_n10157_));
  XOR2_X1    g09965(.A1(new_n10157_), .A2(new_n9716_), .Z(new_n10158_));
  INV_X1     g09966(.I(new_n10158_), .ZN(new_n10159_));
  NOR2_X1    g09967(.A1(new_n9679_), .A2(\asqrt[23] ), .ZN(new_n10160_));
  NOR3_X1    g09968(.A1(new_n10045_), .A2(new_n10160_), .A3(new_n9699_), .ZN(new_n10161_));
  XOR2_X1    g09969(.A1(new_n10161_), .A2(new_n9670_), .Z(new_n10162_));
  NOR3_X1    g09970(.A1(new_n10045_), .A2(\a[40] ), .A3(\a[41] ), .ZN(new_n10163_));
  NOR4_X1    g09971(.A1(new_n10043_), .A2(new_n9590_), .A3(new_n9840_), .A4(new_n10044_), .ZN(new_n10164_));
  OAI21_X1   g09972(.A1(new_n10163_), .A2(new_n10164_), .B(new_n9296_), .ZN(new_n10165_));
  NAND3_X1   g09973(.A1(\asqrt[20] ), .A2(new_n9671_), .A3(new_n9672_), .ZN(new_n10166_));
  INV_X1     g09974(.I(new_n10164_), .ZN(new_n10167_));
  NAND3_X1   g09975(.A1(new_n10166_), .A2(\a[42] ), .A3(new_n10167_), .ZN(new_n10168_));
  NAND2_X1   g09976(.A1(new_n10165_), .A2(new_n10168_), .ZN(new_n10169_));
  INV_X1     g09977(.I(\a[38] ), .ZN(new_n10170_));
  INV_X1     g09978(.I(\a[39] ), .ZN(new_n10171_));
  NAND3_X1   g09979(.A1(new_n10170_), .A2(new_n10171_), .A3(new_n9671_), .ZN(new_n10172_));
  NAND2_X1   g09980(.A1(\asqrt[20] ), .A2(\a[40] ), .ZN(new_n10173_));
  AOI21_X1   g09981(.A1(new_n10173_), .A2(new_n10172_), .B(new_n9590_), .ZN(new_n10174_));
  AOI21_X1   g09982(.A1(\asqrt[20] ), .A2(new_n9671_), .B(new_n9672_), .ZN(new_n10175_));
  NOR2_X1    g09983(.A1(new_n10163_), .A2(new_n10175_), .ZN(new_n10176_));
  NAND3_X1   g09984(.A1(new_n10173_), .A2(new_n9590_), .A3(new_n10172_), .ZN(new_n10177_));
  AOI21_X1   g09985(.A1(new_n10176_), .A2(new_n10177_), .B(new_n10174_), .ZN(new_n10178_));
  AOI21_X1   g09986(.A1(new_n10178_), .A2(new_n9177_), .B(new_n10169_), .ZN(new_n10179_));
  NOR2_X1    g09987(.A1(new_n10178_), .A2(new_n9177_), .ZN(new_n10180_));
  NOR3_X1    g09988(.A1(new_n10179_), .A2(\asqrt[23] ), .A3(new_n10180_), .ZN(new_n10181_));
  NOR3_X1    g09989(.A1(new_n10045_), .A2(new_n9693_), .A3(new_n9678_), .ZN(new_n10182_));
  XOR2_X1    g09990(.A1(new_n10182_), .A2(new_n9695_), .Z(new_n10183_));
  INV_X1     g09991(.I(new_n10183_), .ZN(new_n10184_));
  OAI21_X1   g09992(.A1(new_n10179_), .A2(new_n10180_), .B(\asqrt[23] ), .ZN(new_n10185_));
  OAI21_X1   g09993(.A1(new_n10181_), .A2(new_n10184_), .B(new_n10185_), .ZN(new_n10186_));
  OAI21_X1   g09994(.A1(new_n10186_), .A2(\asqrt[24] ), .B(new_n10162_), .ZN(new_n10187_));
  AOI21_X1   g09995(.A1(new_n10186_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n10188_));
  AOI21_X1   g09996(.A1(new_n10188_), .A2(new_n10187_), .B(new_n10159_), .ZN(new_n10189_));
  NAND2_X1   g09997(.A1(new_n10186_), .A2(\asqrt[24] ), .ZN(new_n10190_));
  AOI21_X1   g09998(.A1(new_n10187_), .A2(new_n10190_), .B(new_n7934_), .ZN(new_n10191_));
  NOR2_X1    g09999(.A1(new_n10189_), .A2(new_n10191_), .ZN(new_n10192_));
  AOI21_X1   g10000(.A1(new_n10192_), .A2(new_n7561_), .B(new_n10156_), .ZN(new_n10193_));
  OAI21_X1   g10001(.A1(new_n10189_), .A2(new_n10191_), .B(\asqrt[26] ), .ZN(new_n10194_));
  NAND2_X1   g10002(.A1(new_n10194_), .A2(new_n7166_), .ZN(new_n10195_));
  OAI21_X1   g10003(.A1(new_n10193_), .A2(new_n10195_), .B(new_n10152_), .ZN(new_n10196_));
  INV_X1     g10004(.I(new_n10194_), .ZN(new_n10197_));
  OAI21_X1   g10005(.A1(new_n10193_), .A2(new_n10197_), .B(\asqrt[27] ), .ZN(new_n10198_));
  NAND3_X1   g10006(.A1(new_n10196_), .A2(new_n10198_), .A3(new_n6813_), .ZN(new_n10199_));
  NAND2_X1   g10007(.A1(new_n10199_), .A2(new_n10150_), .ZN(new_n10200_));
  NAND2_X1   g10008(.A1(new_n10196_), .A2(new_n10198_), .ZN(new_n10201_));
  AOI21_X1   g10009(.A1(new_n10201_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n10202_));
  AOI21_X1   g10010(.A1(new_n10202_), .A2(new_n10200_), .B(new_n10147_), .ZN(new_n10203_));
  INV_X1     g10011(.I(new_n10152_), .ZN(new_n10204_));
  INV_X1     g10012(.I(new_n10162_), .ZN(new_n10205_));
  AOI21_X1   g10013(.A1(new_n10166_), .A2(new_n10167_), .B(\a[42] ), .ZN(new_n10206_));
  NOR3_X1    g10014(.A1(new_n10163_), .A2(new_n9296_), .A3(new_n10164_), .ZN(new_n10207_));
  NOR2_X1    g10015(.A1(new_n10207_), .A2(new_n10206_), .ZN(new_n10208_));
  OAI21_X1   g10016(.A1(new_n10045_), .A2(new_n9671_), .B(new_n10172_), .ZN(new_n10209_));
  NAND2_X1   g10017(.A1(new_n10209_), .A2(\asqrt[21] ), .ZN(new_n10210_));
  OAI21_X1   g10018(.A1(new_n10045_), .A2(\a[40] ), .B(\a[41] ), .ZN(new_n10211_));
  NAND2_X1   g10019(.A1(new_n10211_), .A2(new_n10166_), .ZN(new_n10212_));
  NOR2_X1    g10020(.A1(new_n10209_), .A2(\asqrt[21] ), .ZN(new_n10213_));
  OAI21_X1   g10021(.A1(new_n10212_), .A2(new_n10213_), .B(new_n10210_), .ZN(new_n10214_));
  OAI21_X1   g10022(.A1(\asqrt[22] ), .A2(new_n10214_), .B(new_n10208_), .ZN(new_n10215_));
  NAND2_X1   g10023(.A1(new_n10214_), .A2(\asqrt[22] ), .ZN(new_n10216_));
  NAND3_X1   g10024(.A1(new_n10215_), .A2(new_n8742_), .A3(new_n10216_), .ZN(new_n10217_));
  AOI21_X1   g10025(.A1(new_n10215_), .A2(new_n10216_), .B(new_n8742_), .ZN(new_n10218_));
  AOI21_X1   g10026(.A1(new_n10217_), .A2(new_n10183_), .B(new_n10218_), .ZN(new_n10219_));
  AOI21_X1   g10027(.A1(new_n10219_), .A2(new_n8349_), .B(new_n10205_), .ZN(new_n10220_));
  OAI21_X1   g10028(.A1(new_n10219_), .A2(new_n8349_), .B(new_n7934_), .ZN(new_n10221_));
  OAI21_X1   g10029(.A1(new_n10220_), .A2(new_n10221_), .B(new_n10158_), .ZN(new_n10222_));
  NOR2_X1    g10030(.A1(new_n10219_), .A2(new_n8349_), .ZN(new_n10223_));
  OAI21_X1   g10031(.A1(new_n10220_), .A2(new_n10223_), .B(\asqrt[25] ), .ZN(new_n10224_));
  NAND3_X1   g10032(.A1(new_n10222_), .A2(new_n10224_), .A3(new_n7561_), .ZN(new_n10225_));
  NAND2_X1   g10033(.A1(new_n10225_), .A2(new_n10155_), .ZN(new_n10226_));
  NAND2_X1   g10034(.A1(new_n10222_), .A2(new_n10224_), .ZN(new_n10227_));
  AOI21_X1   g10035(.A1(new_n10227_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n10228_));
  AOI21_X1   g10036(.A1(new_n10228_), .A2(new_n10226_), .B(new_n10204_), .ZN(new_n10229_));
  AOI21_X1   g10037(.A1(new_n10226_), .A2(new_n10194_), .B(new_n7166_), .ZN(new_n10230_));
  OAI21_X1   g10038(.A1(new_n10229_), .A2(new_n10230_), .B(\asqrt[28] ), .ZN(new_n10231_));
  AOI21_X1   g10039(.A1(new_n10200_), .A2(new_n10231_), .B(new_n6454_), .ZN(new_n10232_));
  NOR2_X1    g10040(.A1(new_n10203_), .A2(new_n10232_), .ZN(new_n10233_));
  AOI21_X1   g10041(.A1(new_n10233_), .A2(new_n6106_), .B(new_n10144_), .ZN(new_n10234_));
  OAI21_X1   g10042(.A1(new_n10203_), .A2(new_n10232_), .B(\asqrt[30] ), .ZN(new_n10235_));
  NAND2_X1   g10043(.A1(new_n10235_), .A2(new_n5750_), .ZN(new_n10236_));
  OAI21_X1   g10044(.A1(new_n10234_), .A2(new_n10236_), .B(new_n10140_), .ZN(new_n10237_));
  INV_X1     g10045(.I(new_n10235_), .ZN(new_n10238_));
  OAI21_X1   g10046(.A1(new_n10234_), .A2(new_n10238_), .B(\asqrt[31] ), .ZN(new_n10239_));
  NAND3_X1   g10047(.A1(new_n10237_), .A2(new_n10239_), .A3(new_n5435_), .ZN(new_n10240_));
  NAND2_X1   g10048(.A1(new_n10240_), .A2(new_n10138_), .ZN(new_n10241_));
  NAND2_X1   g10049(.A1(new_n10237_), .A2(new_n10239_), .ZN(new_n10242_));
  AOI21_X1   g10050(.A1(new_n10242_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n10243_));
  AOI21_X1   g10051(.A1(new_n10243_), .A2(new_n10241_), .B(new_n10135_), .ZN(new_n10244_));
  INV_X1     g10052(.I(new_n10140_), .ZN(new_n10245_));
  INV_X1     g10053(.I(new_n10150_), .ZN(new_n10246_));
  NOR2_X1    g10054(.A1(new_n10229_), .A2(new_n10230_), .ZN(new_n10247_));
  AOI21_X1   g10055(.A1(new_n10247_), .A2(new_n6813_), .B(new_n10246_), .ZN(new_n10248_));
  NAND2_X1   g10056(.A1(new_n10231_), .A2(new_n6454_), .ZN(new_n10249_));
  OAI21_X1   g10057(.A1(new_n10248_), .A2(new_n10249_), .B(new_n10146_), .ZN(new_n10250_));
  INV_X1     g10058(.I(new_n10231_), .ZN(new_n10251_));
  OAI21_X1   g10059(.A1(new_n10248_), .A2(new_n10251_), .B(\asqrt[29] ), .ZN(new_n10252_));
  NAND3_X1   g10060(.A1(new_n10250_), .A2(new_n10252_), .A3(new_n6106_), .ZN(new_n10253_));
  NAND2_X1   g10061(.A1(new_n10253_), .A2(new_n10143_), .ZN(new_n10254_));
  NAND2_X1   g10062(.A1(new_n10250_), .A2(new_n10252_), .ZN(new_n10255_));
  AOI21_X1   g10063(.A1(new_n10255_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n10256_));
  AOI21_X1   g10064(.A1(new_n10256_), .A2(new_n10254_), .B(new_n10245_), .ZN(new_n10257_));
  AOI21_X1   g10065(.A1(new_n10254_), .A2(new_n10235_), .B(new_n5750_), .ZN(new_n10258_));
  OAI21_X1   g10066(.A1(new_n10257_), .A2(new_n10258_), .B(\asqrt[32] ), .ZN(new_n10259_));
  AOI21_X1   g10067(.A1(new_n10241_), .A2(new_n10259_), .B(new_n5110_), .ZN(new_n10260_));
  NOR2_X1    g10068(.A1(new_n10244_), .A2(new_n10260_), .ZN(new_n10261_));
  AOI21_X1   g10069(.A1(new_n10261_), .A2(new_n4810_), .B(new_n10132_), .ZN(new_n10262_));
  OAI21_X1   g10070(.A1(new_n10244_), .A2(new_n10260_), .B(\asqrt[34] ), .ZN(new_n10263_));
  NAND2_X1   g10071(.A1(new_n10263_), .A2(new_n4510_), .ZN(new_n10264_));
  OAI21_X1   g10072(.A1(new_n10262_), .A2(new_n10264_), .B(new_n10128_), .ZN(new_n10265_));
  INV_X1     g10073(.I(new_n10263_), .ZN(new_n10266_));
  OAI21_X1   g10074(.A1(new_n10262_), .A2(new_n10266_), .B(\asqrt[35] ), .ZN(new_n10267_));
  NAND3_X1   g10075(.A1(new_n10265_), .A2(new_n10267_), .A3(new_n4224_), .ZN(new_n10268_));
  NAND2_X1   g10076(.A1(new_n10268_), .A2(new_n10126_), .ZN(new_n10269_));
  NAND2_X1   g10077(.A1(new_n10265_), .A2(new_n10267_), .ZN(new_n10270_));
  AOI21_X1   g10078(.A1(new_n10270_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n10271_));
  AOI21_X1   g10079(.A1(new_n10271_), .A2(new_n10269_), .B(new_n10123_), .ZN(new_n10272_));
  INV_X1     g10080(.I(new_n10128_), .ZN(new_n10273_));
  INV_X1     g10081(.I(new_n10138_), .ZN(new_n10274_));
  NOR2_X1    g10082(.A1(new_n10257_), .A2(new_n10258_), .ZN(new_n10275_));
  AOI21_X1   g10083(.A1(new_n10275_), .A2(new_n5435_), .B(new_n10274_), .ZN(new_n10276_));
  NAND2_X1   g10084(.A1(new_n10259_), .A2(new_n5110_), .ZN(new_n10277_));
  OAI21_X1   g10085(.A1(new_n10276_), .A2(new_n10277_), .B(new_n10134_), .ZN(new_n10278_));
  INV_X1     g10086(.I(new_n10259_), .ZN(new_n10279_));
  OAI21_X1   g10087(.A1(new_n10276_), .A2(new_n10279_), .B(\asqrt[33] ), .ZN(new_n10280_));
  NAND3_X1   g10088(.A1(new_n10278_), .A2(new_n10280_), .A3(new_n4810_), .ZN(new_n10281_));
  NAND2_X1   g10089(.A1(new_n10281_), .A2(new_n10131_), .ZN(new_n10282_));
  NAND2_X1   g10090(.A1(new_n10278_), .A2(new_n10280_), .ZN(new_n10283_));
  AOI21_X1   g10091(.A1(new_n10283_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n10284_));
  AOI21_X1   g10092(.A1(new_n10284_), .A2(new_n10282_), .B(new_n10273_), .ZN(new_n10285_));
  AOI21_X1   g10093(.A1(new_n10282_), .A2(new_n10263_), .B(new_n4510_), .ZN(new_n10286_));
  OAI21_X1   g10094(.A1(new_n10285_), .A2(new_n10286_), .B(\asqrt[36] ), .ZN(new_n10287_));
  AOI21_X1   g10095(.A1(new_n10269_), .A2(new_n10287_), .B(new_n3928_), .ZN(new_n10288_));
  NOR2_X1    g10096(.A1(new_n10272_), .A2(new_n10288_), .ZN(new_n10289_));
  AOI21_X1   g10097(.A1(new_n10289_), .A2(new_n3675_), .B(new_n10120_), .ZN(new_n10290_));
  OAI21_X1   g10098(.A1(new_n10272_), .A2(new_n10288_), .B(\asqrt[38] ), .ZN(new_n10291_));
  NAND2_X1   g10099(.A1(new_n10291_), .A2(new_n3400_), .ZN(new_n10292_));
  OAI21_X1   g10100(.A1(new_n10290_), .A2(new_n10292_), .B(new_n10116_), .ZN(new_n10293_));
  INV_X1     g10101(.I(new_n10291_), .ZN(new_n10294_));
  OAI21_X1   g10102(.A1(new_n10290_), .A2(new_n10294_), .B(\asqrt[39] ), .ZN(new_n10295_));
  NAND3_X1   g10103(.A1(new_n10293_), .A2(new_n10295_), .A3(new_n3167_), .ZN(new_n10296_));
  NAND2_X1   g10104(.A1(new_n10296_), .A2(new_n10114_), .ZN(new_n10297_));
  NAND2_X1   g10105(.A1(new_n10293_), .A2(new_n10295_), .ZN(new_n10298_));
  AOI21_X1   g10106(.A1(new_n10298_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n10299_));
  AOI21_X1   g10107(.A1(new_n10299_), .A2(new_n10297_), .B(new_n10111_), .ZN(new_n10300_));
  INV_X1     g10108(.I(new_n10116_), .ZN(new_n10301_));
  INV_X1     g10109(.I(new_n10126_), .ZN(new_n10302_));
  NOR2_X1    g10110(.A1(new_n10285_), .A2(new_n10286_), .ZN(new_n10303_));
  AOI21_X1   g10111(.A1(new_n10303_), .A2(new_n4224_), .B(new_n10302_), .ZN(new_n10304_));
  NAND2_X1   g10112(.A1(new_n10287_), .A2(new_n3928_), .ZN(new_n10305_));
  OAI21_X1   g10113(.A1(new_n10304_), .A2(new_n10305_), .B(new_n10122_), .ZN(new_n10306_));
  INV_X1     g10114(.I(new_n10287_), .ZN(new_n10307_));
  OAI21_X1   g10115(.A1(new_n10304_), .A2(new_n10307_), .B(\asqrt[37] ), .ZN(new_n10308_));
  NAND3_X1   g10116(.A1(new_n10306_), .A2(new_n10308_), .A3(new_n3675_), .ZN(new_n10309_));
  NAND2_X1   g10117(.A1(new_n10309_), .A2(new_n10119_), .ZN(new_n10310_));
  NAND2_X1   g10118(.A1(new_n10306_), .A2(new_n10308_), .ZN(new_n10311_));
  AOI21_X1   g10119(.A1(new_n10311_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n10312_));
  AOI21_X1   g10120(.A1(new_n10312_), .A2(new_n10310_), .B(new_n10301_), .ZN(new_n10313_));
  AOI21_X1   g10121(.A1(new_n10310_), .A2(new_n10291_), .B(new_n3400_), .ZN(new_n10314_));
  OAI21_X1   g10122(.A1(new_n10313_), .A2(new_n10314_), .B(\asqrt[40] ), .ZN(new_n10315_));
  AOI21_X1   g10123(.A1(new_n10297_), .A2(new_n10315_), .B(new_n2912_), .ZN(new_n10316_));
  NOR2_X1    g10124(.A1(new_n10300_), .A2(new_n10316_), .ZN(new_n10317_));
  AOI21_X1   g10125(.A1(new_n10317_), .A2(new_n2699_), .B(new_n10108_), .ZN(new_n10318_));
  OAI21_X1   g10126(.A1(new_n10300_), .A2(new_n10316_), .B(\asqrt[42] ), .ZN(new_n10319_));
  NAND2_X1   g10127(.A1(new_n10319_), .A2(new_n2464_), .ZN(new_n10320_));
  OAI21_X1   g10128(.A1(new_n10318_), .A2(new_n10320_), .B(new_n10104_), .ZN(new_n10321_));
  INV_X1     g10129(.I(new_n10319_), .ZN(new_n10322_));
  OAI21_X1   g10130(.A1(new_n10318_), .A2(new_n10322_), .B(\asqrt[43] ), .ZN(new_n10323_));
  NAND3_X1   g10131(.A1(new_n10321_), .A2(new_n10323_), .A3(new_n2271_), .ZN(new_n10324_));
  NAND2_X1   g10132(.A1(new_n10324_), .A2(new_n10102_), .ZN(new_n10325_));
  NAND2_X1   g10133(.A1(new_n10321_), .A2(new_n10323_), .ZN(new_n10326_));
  AOI21_X1   g10134(.A1(new_n10326_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n10327_));
  AOI21_X1   g10135(.A1(new_n10327_), .A2(new_n10325_), .B(new_n10099_), .ZN(new_n10328_));
  INV_X1     g10136(.I(new_n10104_), .ZN(new_n10329_));
  INV_X1     g10137(.I(new_n10114_), .ZN(new_n10330_));
  NOR2_X1    g10138(.A1(new_n10313_), .A2(new_n10314_), .ZN(new_n10331_));
  AOI21_X1   g10139(.A1(new_n10331_), .A2(new_n3167_), .B(new_n10330_), .ZN(new_n10332_));
  NAND2_X1   g10140(.A1(new_n10315_), .A2(new_n2912_), .ZN(new_n10333_));
  OAI21_X1   g10141(.A1(new_n10332_), .A2(new_n10333_), .B(new_n10110_), .ZN(new_n10334_));
  INV_X1     g10142(.I(new_n10315_), .ZN(new_n10335_));
  OAI21_X1   g10143(.A1(new_n10332_), .A2(new_n10335_), .B(\asqrt[41] ), .ZN(new_n10336_));
  NAND3_X1   g10144(.A1(new_n10334_), .A2(new_n10336_), .A3(new_n2699_), .ZN(new_n10337_));
  NAND2_X1   g10145(.A1(new_n10337_), .A2(new_n10107_), .ZN(new_n10338_));
  NAND2_X1   g10146(.A1(new_n10334_), .A2(new_n10336_), .ZN(new_n10339_));
  AOI21_X1   g10147(.A1(new_n10339_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n10340_));
  AOI21_X1   g10148(.A1(new_n10340_), .A2(new_n10338_), .B(new_n10329_), .ZN(new_n10341_));
  AOI21_X1   g10149(.A1(new_n10338_), .A2(new_n10319_), .B(new_n2464_), .ZN(new_n10342_));
  OAI21_X1   g10150(.A1(new_n10341_), .A2(new_n10342_), .B(\asqrt[44] ), .ZN(new_n10343_));
  AOI21_X1   g10151(.A1(new_n10325_), .A2(new_n10343_), .B(new_n2072_), .ZN(new_n10344_));
  NOR2_X1    g10152(.A1(new_n10328_), .A2(new_n10344_), .ZN(new_n10345_));
  AOI21_X1   g10153(.A1(new_n10345_), .A2(new_n1884_), .B(new_n10098_), .ZN(new_n10346_));
  OAI21_X1   g10154(.A1(new_n10328_), .A2(new_n10344_), .B(\asqrt[46] ), .ZN(new_n10347_));
  NAND2_X1   g10155(.A1(new_n10347_), .A2(new_n1688_), .ZN(new_n10348_));
  OAI21_X1   g10156(.A1(new_n10346_), .A2(new_n10348_), .B(new_n10094_), .ZN(new_n10349_));
  INV_X1     g10157(.I(new_n10347_), .ZN(new_n10350_));
  OAI21_X1   g10158(.A1(new_n10346_), .A2(new_n10350_), .B(\asqrt[47] ), .ZN(new_n10351_));
  NAND3_X1   g10159(.A1(new_n10349_), .A2(new_n10351_), .A3(new_n1533_), .ZN(new_n10352_));
  NAND2_X1   g10160(.A1(new_n10352_), .A2(new_n10092_), .ZN(new_n10353_));
  NAND2_X1   g10161(.A1(new_n10349_), .A2(new_n10351_), .ZN(new_n10354_));
  AOI21_X1   g10162(.A1(new_n10354_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n10355_));
  AOI21_X1   g10163(.A1(new_n10355_), .A2(new_n10353_), .B(new_n10089_), .ZN(new_n10356_));
  INV_X1     g10164(.I(new_n10094_), .ZN(new_n10357_));
  INV_X1     g10165(.I(new_n10102_), .ZN(new_n10358_));
  NOR2_X1    g10166(.A1(new_n10341_), .A2(new_n10342_), .ZN(new_n10359_));
  AOI21_X1   g10167(.A1(new_n10359_), .A2(new_n2271_), .B(new_n10358_), .ZN(new_n10360_));
  NAND2_X1   g10168(.A1(new_n10343_), .A2(new_n2072_), .ZN(new_n10361_));
  OAI21_X1   g10169(.A1(new_n10360_), .A2(new_n10361_), .B(new_n10028_), .ZN(new_n10362_));
  INV_X1     g10170(.I(new_n10343_), .ZN(new_n10363_));
  OAI21_X1   g10171(.A1(new_n10360_), .A2(new_n10363_), .B(\asqrt[45] ), .ZN(new_n10364_));
  NAND3_X1   g10172(.A1(new_n10362_), .A2(new_n10364_), .A3(new_n1884_), .ZN(new_n10365_));
  NAND2_X1   g10173(.A1(new_n10365_), .A2(new_n10097_), .ZN(new_n10366_));
  NAND2_X1   g10174(.A1(new_n10362_), .A2(new_n10364_), .ZN(new_n10367_));
  AOI21_X1   g10175(.A1(new_n10367_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n10368_));
  AOI21_X1   g10176(.A1(new_n10368_), .A2(new_n10366_), .B(new_n10357_), .ZN(new_n10369_));
  AOI21_X1   g10177(.A1(new_n10366_), .A2(new_n10347_), .B(new_n1688_), .ZN(new_n10370_));
  OAI21_X1   g10178(.A1(new_n10369_), .A2(new_n10370_), .B(\asqrt[48] ), .ZN(new_n10371_));
  AOI21_X1   g10179(.A1(new_n10353_), .A2(new_n10371_), .B(new_n1368_), .ZN(new_n10372_));
  NOR2_X1    g10180(.A1(new_n10356_), .A2(new_n10372_), .ZN(new_n10373_));
  AOI21_X1   g10181(.A1(new_n10373_), .A2(new_n1228_), .B(new_n10086_), .ZN(new_n10374_));
  OAI21_X1   g10182(.A1(new_n10356_), .A2(new_n10372_), .B(\asqrt[50] ), .ZN(new_n10375_));
  NAND2_X1   g10183(.A1(new_n10375_), .A2(new_n1088_), .ZN(new_n10376_));
  OAI21_X1   g10184(.A1(new_n10374_), .A2(new_n10376_), .B(new_n10082_), .ZN(new_n10377_));
  INV_X1     g10185(.I(new_n10375_), .ZN(new_n10378_));
  OAI21_X1   g10186(.A1(new_n10374_), .A2(new_n10378_), .B(\asqrt[51] ), .ZN(new_n10379_));
  NAND3_X1   g10187(.A1(new_n10377_), .A2(new_n10379_), .A3(new_n962_), .ZN(new_n10380_));
  NAND2_X1   g10188(.A1(new_n10380_), .A2(new_n10080_), .ZN(new_n10381_));
  NAND2_X1   g10189(.A1(new_n10377_), .A2(new_n10379_), .ZN(new_n10382_));
  AOI21_X1   g10190(.A1(new_n10382_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n10383_));
  AOI21_X1   g10191(.A1(new_n10383_), .A2(new_n10381_), .B(new_n10077_), .ZN(new_n10384_));
  INV_X1     g10192(.I(new_n10082_), .ZN(new_n10385_));
  INV_X1     g10193(.I(new_n10092_), .ZN(new_n10386_));
  NOR2_X1    g10194(.A1(new_n10369_), .A2(new_n10370_), .ZN(new_n10387_));
  AOI21_X1   g10195(.A1(new_n10387_), .A2(new_n1533_), .B(new_n10386_), .ZN(new_n10388_));
  NAND2_X1   g10196(.A1(new_n10371_), .A2(new_n1368_), .ZN(new_n10389_));
  OAI21_X1   g10197(.A1(new_n10388_), .A2(new_n10389_), .B(new_n10088_), .ZN(new_n10390_));
  INV_X1     g10198(.I(new_n10371_), .ZN(new_n10391_));
  OAI21_X1   g10199(.A1(new_n10388_), .A2(new_n10391_), .B(\asqrt[49] ), .ZN(new_n10392_));
  NAND3_X1   g10200(.A1(new_n10390_), .A2(new_n10392_), .A3(new_n1228_), .ZN(new_n10393_));
  NAND2_X1   g10201(.A1(new_n10393_), .A2(new_n10085_), .ZN(new_n10394_));
  NAND2_X1   g10202(.A1(new_n10390_), .A2(new_n10392_), .ZN(new_n10395_));
  AOI21_X1   g10203(.A1(new_n10395_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n10396_));
  AOI21_X1   g10204(.A1(new_n10396_), .A2(new_n10394_), .B(new_n10385_), .ZN(new_n10397_));
  AOI21_X1   g10205(.A1(new_n10394_), .A2(new_n10375_), .B(new_n1088_), .ZN(new_n10398_));
  OAI21_X1   g10206(.A1(new_n10397_), .A2(new_n10398_), .B(\asqrt[52] ), .ZN(new_n10399_));
  AOI21_X1   g10207(.A1(new_n10381_), .A2(new_n10399_), .B(new_n842_), .ZN(new_n10400_));
  NOR2_X1    g10208(.A1(new_n10384_), .A2(new_n10400_), .ZN(new_n10401_));
  AOI21_X1   g10209(.A1(new_n10401_), .A2(new_n720_), .B(new_n10074_), .ZN(new_n10402_));
  OAI21_X1   g10210(.A1(new_n10384_), .A2(new_n10400_), .B(\asqrt[54] ), .ZN(new_n10403_));
  NAND2_X1   g10211(.A1(new_n10403_), .A2(new_n630_), .ZN(new_n10404_));
  OAI21_X1   g10212(.A1(new_n10402_), .A2(new_n10404_), .B(new_n10070_), .ZN(new_n10405_));
  INV_X1     g10213(.I(new_n10403_), .ZN(new_n10406_));
  OAI21_X1   g10214(.A1(new_n10402_), .A2(new_n10406_), .B(\asqrt[55] ), .ZN(new_n10407_));
  NAND3_X1   g10215(.A1(new_n10405_), .A2(new_n10407_), .A3(new_n545_), .ZN(new_n10408_));
  NAND2_X1   g10216(.A1(new_n10408_), .A2(new_n10068_), .ZN(new_n10409_));
  NAND2_X1   g10217(.A1(new_n10405_), .A2(new_n10407_), .ZN(new_n10410_));
  AOI21_X1   g10218(.A1(new_n10410_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n10411_));
  AOI21_X1   g10219(.A1(new_n10411_), .A2(new_n10409_), .B(new_n10065_), .ZN(new_n10412_));
  INV_X1     g10220(.I(new_n10070_), .ZN(new_n10413_));
  INV_X1     g10221(.I(new_n10080_), .ZN(new_n10414_));
  NOR2_X1    g10222(.A1(new_n10397_), .A2(new_n10398_), .ZN(new_n10415_));
  AOI21_X1   g10223(.A1(new_n10415_), .A2(new_n962_), .B(new_n10414_), .ZN(new_n10416_));
  NAND2_X1   g10224(.A1(new_n10399_), .A2(new_n842_), .ZN(new_n10417_));
  OAI21_X1   g10225(.A1(new_n10416_), .A2(new_n10417_), .B(new_n10076_), .ZN(new_n10418_));
  INV_X1     g10226(.I(new_n10399_), .ZN(new_n10419_));
  OAI21_X1   g10227(.A1(new_n10416_), .A2(new_n10419_), .B(\asqrt[53] ), .ZN(new_n10420_));
  NAND3_X1   g10228(.A1(new_n10418_), .A2(new_n10420_), .A3(new_n720_), .ZN(new_n10421_));
  NAND2_X1   g10229(.A1(new_n10421_), .A2(new_n10073_), .ZN(new_n10422_));
  NAND2_X1   g10230(.A1(new_n10418_), .A2(new_n10420_), .ZN(new_n10423_));
  AOI21_X1   g10231(.A1(new_n10423_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n10424_));
  AOI21_X1   g10232(.A1(new_n10424_), .A2(new_n10422_), .B(new_n10413_), .ZN(new_n10425_));
  AOI21_X1   g10233(.A1(new_n10422_), .A2(new_n10403_), .B(new_n630_), .ZN(new_n10426_));
  OAI21_X1   g10234(.A1(new_n10425_), .A2(new_n10426_), .B(\asqrt[56] ), .ZN(new_n10427_));
  AOI21_X1   g10235(.A1(new_n10409_), .A2(new_n10427_), .B(new_n450_), .ZN(new_n10428_));
  NOR2_X1    g10236(.A1(new_n10412_), .A2(new_n10428_), .ZN(new_n10429_));
  AOI21_X1   g10237(.A1(new_n10429_), .A2(new_n403_), .B(new_n10062_), .ZN(new_n10430_));
  OAI21_X1   g10238(.A1(new_n10412_), .A2(new_n10428_), .B(\asqrt[58] ), .ZN(new_n10431_));
  NAND2_X1   g10239(.A1(new_n10431_), .A2(new_n339_), .ZN(new_n10432_));
  OAI21_X1   g10240(.A1(new_n10430_), .A2(new_n10432_), .B(new_n10058_), .ZN(new_n10433_));
  INV_X1     g10241(.I(new_n10431_), .ZN(new_n10434_));
  OAI21_X1   g10242(.A1(new_n10430_), .A2(new_n10434_), .B(\asqrt[59] ), .ZN(new_n10435_));
  NAND3_X1   g10243(.A1(new_n10433_), .A2(new_n10435_), .A3(new_n288_), .ZN(new_n10436_));
  NAND2_X1   g10244(.A1(new_n10436_), .A2(new_n10056_), .ZN(new_n10437_));
  INV_X1     g10245(.I(new_n10058_), .ZN(new_n10438_));
  INV_X1     g10246(.I(new_n10068_), .ZN(new_n10439_));
  NOR2_X1    g10247(.A1(new_n10425_), .A2(new_n10426_), .ZN(new_n10440_));
  AOI21_X1   g10248(.A1(new_n10440_), .A2(new_n545_), .B(new_n10439_), .ZN(new_n10441_));
  NAND2_X1   g10249(.A1(new_n10427_), .A2(new_n450_), .ZN(new_n10442_));
  OAI21_X1   g10250(.A1(new_n10441_), .A2(new_n10442_), .B(new_n10064_), .ZN(new_n10443_));
  INV_X1     g10251(.I(new_n10427_), .ZN(new_n10444_));
  OAI21_X1   g10252(.A1(new_n10441_), .A2(new_n10444_), .B(\asqrt[57] ), .ZN(new_n10445_));
  NAND3_X1   g10253(.A1(new_n10443_), .A2(new_n10445_), .A3(new_n403_), .ZN(new_n10446_));
  NAND2_X1   g10254(.A1(new_n10446_), .A2(new_n10061_), .ZN(new_n10447_));
  NAND2_X1   g10255(.A1(new_n10443_), .A2(new_n10445_), .ZN(new_n10448_));
  AOI21_X1   g10256(.A1(new_n10448_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n10449_));
  AOI21_X1   g10257(.A1(new_n10449_), .A2(new_n10447_), .B(new_n10438_), .ZN(new_n10450_));
  AOI21_X1   g10258(.A1(new_n10447_), .A2(new_n10431_), .B(new_n339_), .ZN(new_n10451_));
  OAI21_X1   g10259(.A1(new_n10450_), .A2(new_n10451_), .B(\asqrt[60] ), .ZN(new_n10452_));
  AOI21_X1   g10260(.A1(new_n10437_), .A2(new_n10452_), .B(new_n242_), .ZN(new_n10453_));
  NAND3_X1   g10261(.A1(\asqrt[20] ), .A2(new_n9988_), .A3(new_n10004_), .ZN(new_n10454_));
  XOR2_X1    g10262(.A1(new_n10454_), .A2(new_n10029_), .Z(new_n10455_));
  INV_X1     g10263(.I(new_n10455_), .ZN(new_n10456_));
  NAND2_X1   g10264(.A1(new_n10433_), .A2(new_n10435_), .ZN(new_n10457_));
  AOI21_X1   g10265(.A1(new_n10457_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n10458_));
  AOI21_X1   g10266(.A1(new_n10458_), .A2(new_n10437_), .B(new_n10456_), .ZN(new_n10459_));
  OAI21_X1   g10267(.A1(new_n10459_), .A2(new_n10453_), .B(\asqrt[62] ), .ZN(new_n10460_));
  AOI21_X1   g10268(.A1(new_n9989_), .A2(new_n10010_), .B(new_n10005_), .ZN(new_n10461_));
  NAND2_X1   g10269(.A1(\asqrt[20] ), .A2(new_n10461_), .ZN(new_n10462_));
  XOR2_X1    g10270(.A1(new_n10462_), .A2(new_n10008_), .Z(new_n10463_));
  INV_X1     g10271(.I(new_n10056_), .ZN(new_n10464_));
  NOR2_X1    g10272(.A1(new_n10450_), .A2(new_n10451_), .ZN(new_n10465_));
  AOI21_X1   g10273(.A1(new_n10465_), .A2(new_n288_), .B(new_n10464_), .ZN(new_n10466_));
  INV_X1     g10274(.I(new_n10452_), .ZN(new_n10467_));
  OAI21_X1   g10275(.A1(new_n10466_), .A2(new_n10467_), .B(\asqrt[61] ), .ZN(new_n10468_));
  NAND2_X1   g10276(.A1(new_n10452_), .A2(new_n242_), .ZN(new_n10469_));
  OAI21_X1   g10277(.A1(new_n10466_), .A2(new_n10469_), .B(new_n10455_), .ZN(new_n10470_));
  NAND3_X1   g10278(.A1(new_n10470_), .A2(new_n10468_), .A3(new_n234_), .ZN(new_n10471_));
  NAND2_X1   g10279(.A1(new_n10471_), .A2(new_n10463_), .ZN(new_n10472_));
  AOI21_X1   g10280(.A1(new_n10472_), .A2(new_n10460_), .B(new_n10053_), .ZN(new_n10473_));
  AOI21_X1   g10281(.A1(new_n10473_), .A2(new_n10051_), .B(\asqrt[63] ), .ZN(new_n10474_));
  NAND2_X1   g10282(.A1(new_n10472_), .A2(new_n10460_), .ZN(new_n10475_));
  NOR2_X1    g10283(.A1(new_n10475_), .A2(new_n10051_), .ZN(new_n10476_));
  NOR2_X1    g10284(.A1(\asqrt[20] ), .A2(new_n10040_), .ZN(new_n10477_));
  NOR4_X1    g10285(.A1(new_n10474_), .A2(new_n10048_), .A3(new_n10476_), .A4(new_n10477_), .ZN(new_n10478_));
  OAI21_X1   g10286(.A1(new_n10360_), .A2(new_n10361_), .B(new_n10364_), .ZN(new_n10479_));
  NOR2_X1    g10287(.A1(new_n10478_), .A2(new_n10479_), .ZN(new_n10480_));
  XOR2_X1    g10288(.A1(new_n10480_), .A2(new_n10028_), .Z(new_n10481_));
  INV_X1     g10289(.I(new_n10481_), .ZN(new_n10482_));
  INV_X1     g10290(.I(new_n10048_), .ZN(new_n10483_));
  INV_X1     g10291(.I(new_n10460_), .ZN(new_n10484_));
  NOR2_X1    g10292(.A1(new_n10459_), .A2(new_n10453_), .ZN(new_n10485_));
  INV_X1     g10293(.I(new_n10463_), .ZN(new_n10486_));
  AOI21_X1   g10294(.A1(new_n10485_), .A2(new_n234_), .B(new_n10486_), .ZN(new_n10487_));
  OAI21_X1   g10295(.A1(new_n10487_), .A2(new_n10484_), .B(new_n10052_), .ZN(new_n10488_));
  OAI21_X1   g10296(.A1(new_n10488_), .A2(new_n10050_), .B(new_n193_), .ZN(new_n10489_));
  NOR2_X1    g10297(.A1(new_n10487_), .A2(new_n10484_), .ZN(new_n10490_));
  NAND2_X1   g10298(.A1(new_n10490_), .A2(new_n10050_), .ZN(new_n10491_));
  INV_X1     g10299(.I(new_n10477_), .ZN(new_n10492_));
  NAND4_X1   g10300(.A1(new_n10489_), .A2(new_n10483_), .A3(new_n10491_), .A4(new_n10492_), .ZN(\asqrt[19] ));
  NAND3_X1   g10301(.A1(\asqrt[19] ), .A2(new_n10324_), .A3(new_n10343_), .ZN(new_n10494_));
  XOR2_X1    g10302(.A1(new_n10494_), .A2(new_n10358_), .Z(new_n10495_));
  OAI21_X1   g10303(.A1(new_n10318_), .A2(new_n10320_), .B(new_n10323_), .ZN(new_n10496_));
  NOR2_X1    g10304(.A1(new_n10478_), .A2(new_n10496_), .ZN(new_n10497_));
  XOR2_X1    g10305(.A1(new_n10497_), .A2(new_n10104_), .Z(new_n10498_));
  INV_X1     g10306(.I(new_n10498_), .ZN(new_n10499_));
  NAND3_X1   g10307(.A1(\asqrt[19] ), .A2(new_n10337_), .A3(new_n10319_), .ZN(new_n10500_));
  XOR2_X1    g10308(.A1(new_n10500_), .A2(new_n10108_), .Z(new_n10501_));
  INV_X1     g10309(.I(new_n10501_), .ZN(new_n10502_));
  OAI21_X1   g10310(.A1(new_n10332_), .A2(new_n10333_), .B(new_n10336_), .ZN(new_n10503_));
  NOR2_X1    g10311(.A1(new_n10478_), .A2(new_n10503_), .ZN(new_n10504_));
  XOR2_X1    g10312(.A1(new_n10504_), .A2(new_n10110_), .Z(new_n10505_));
  NAND3_X1   g10313(.A1(\asqrt[19] ), .A2(new_n10296_), .A3(new_n10315_), .ZN(new_n10506_));
  XOR2_X1    g10314(.A1(new_n10506_), .A2(new_n10330_), .Z(new_n10507_));
  OAI21_X1   g10315(.A1(new_n10290_), .A2(new_n10292_), .B(new_n10295_), .ZN(new_n10508_));
  NOR2_X1    g10316(.A1(new_n10478_), .A2(new_n10508_), .ZN(new_n10509_));
  XOR2_X1    g10317(.A1(new_n10509_), .A2(new_n10116_), .Z(new_n10510_));
  INV_X1     g10318(.I(new_n10510_), .ZN(new_n10511_));
  NAND3_X1   g10319(.A1(\asqrt[19] ), .A2(new_n10309_), .A3(new_n10291_), .ZN(new_n10512_));
  XOR2_X1    g10320(.A1(new_n10512_), .A2(new_n10120_), .Z(new_n10513_));
  INV_X1     g10321(.I(new_n10513_), .ZN(new_n10514_));
  OAI21_X1   g10322(.A1(new_n10304_), .A2(new_n10305_), .B(new_n10308_), .ZN(new_n10515_));
  NOR2_X1    g10323(.A1(new_n10478_), .A2(new_n10515_), .ZN(new_n10516_));
  XOR2_X1    g10324(.A1(new_n10516_), .A2(new_n10122_), .Z(new_n10517_));
  NAND3_X1   g10325(.A1(\asqrt[19] ), .A2(new_n10268_), .A3(new_n10287_), .ZN(new_n10518_));
  XOR2_X1    g10326(.A1(new_n10518_), .A2(new_n10302_), .Z(new_n10519_));
  OAI21_X1   g10327(.A1(new_n10262_), .A2(new_n10264_), .B(new_n10267_), .ZN(new_n10520_));
  NOR2_X1    g10328(.A1(new_n10478_), .A2(new_n10520_), .ZN(new_n10521_));
  XOR2_X1    g10329(.A1(new_n10521_), .A2(new_n10128_), .Z(new_n10522_));
  INV_X1     g10330(.I(new_n10522_), .ZN(new_n10523_));
  NAND3_X1   g10331(.A1(\asqrt[19] ), .A2(new_n10281_), .A3(new_n10263_), .ZN(new_n10524_));
  XOR2_X1    g10332(.A1(new_n10524_), .A2(new_n10132_), .Z(new_n10525_));
  INV_X1     g10333(.I(new_n10525_), .ZN(new_n10526_));
  OAI21_X1   g10334(.A1(new_n10276_), .A2(new_n10277_), .B(new_n10280_), .ZN(new_n10527_));
  NOR2_X1    g10335(.A1(new_n10478_), .A2(new_n10527_), .ZN(new_n10528_));
  XOR2_X1    g10336(.A1(new_n10528_), .A2(new_n10134_), .Z(new_n10529_));
  NAND3_X1   g10337(.A1(\asqrt[19] ), .A2(new_n10240_), .A3(new_n10259_), .ZN(new_n10530_));
  XOR2_X1    g10338(.A1(new_n10530_), .A2(new_n10274_), .Z(new_n10531_));
  OAI21_X1   g10339(.A1(new_n10234_), .A2(new_n10236_), .B(new_n10239_), .ZN(new_n10532_));
  NOR2_X1    g10340(.A1(new_n10478_), .A2(new_n10532_), .ZN(new_n10533_));
  XOR2_X1    g10341(.A1(new_n10533_), .A2(new_n10140_), .Z(new_n10534_));
  INV_X1     g10342(.I(new_n10534_), .ZN(new_n10535_));
  NAND3_X1   g10343(.A1(\asqrt[19] ), .A2(new_n10253_), .A3(new_n10235_), .ZN(new_n10536_));
  XOR2_X1    g10344(.A1(new_n10536_), .A2(new_n10144_), .Z(new_n10537_));
  INV_X1     g10345(.I(new_n10537_), .ZN(new_n10538_));
  OAI21_X1   g10346(.A1(new_n10248_), .A2(new_n10249_), .B(new_n10252_), .ZN(new_n10539_));
  NOR2_X1    g10347(.A1(new_n10478_), .A2(new_n10539_), .ZN(new_n10540_));
  XOR2_X1    g10348(.A1(new_n10540_), .A2(new_n10146_), .Z(new_n10541_));
  NAND3_X1   g10349(.A1(\asqrt[19] ), .A2(new_n10199_), .A3(new_n10231_), .ZN(new_n10542_));
  XOR2_X1    g10350(.A1(new_n10542_), .A2(new_n10246_), .Z(new_n10543_));
  OAI21_X1   g10351(.A1(new_n10193_), .A2(new_n10195_), .B(new_n10198_), .ZN(new_n10544_));
  NOR2_X1    g10352(.A1(new_n10478_), .A2(new_n10544_), .ZN(new_n10545_));
  XOR2_X1    g10353(.A1(new_n10545_), .A2(new_n10152_), .Z(new_n10546_));
  INV_X1     g10354(.I(new_n10546_), .ZN(new_n10547_));
  NAND3_X1   g10355(.A1(\asqrt[19] ), .A2(new_n10225_), .A3(new_n10194_), .ZN(new_n10548_));
  XOR2_X1    g10356(.A1(new_n10548_), .A2(new_n10156_), .Z(new_n10549_));
  INV_X1     g10357(.I(new_n10549_), .ZN(new_n10550_));
  AOI21_X1   g10358(.A1(new_n10187_), .A2(new_n10188_), .B(new_n10191_), .ZN(new_n10551_));
  NAND2_X1   g10359(.A1(\asqrt[19] ), .A2(new_n10551_), .ZN(new_n10552_));
  XOR2_X1    g10360(.A1(new_n10552_), .A2(new_n10159_), .Z(new_n10553_));
  NOR2_X1    g10361(.A1(new_n10186_), .A2(\asqrt[24] ), .ZN(new_n10554_));
  NOR3_X1    g10362(.A1(new_n10478_), .A2(new_n10554_), .A3(new_n10223_), .ZN(new_n10555_));
  XOR2_X1    g10363(.A1(new_n10555_), .A2(new_n10162_), .Z(new_n10556_));
  NOR3_X1    g10364(.A1(new_n10478_), .A2(new_n10181_), .A3(new_n10218_), .ZN(new_n10557_));
  XOR2_X1    g10365(.A1(new_n10557_), .A2(new_n10183_), .Z(new_n10558_));
  INV_X1     g10366(.I(new_n10558_), .ZN(new_n10559_));
  NOR2_X1    g10367(.A1(new_n10214_), .A2(\asqrt[22] ), .ZN(new_n10560_));
  NOR3_X1    g10368(.A1(new_n10478_), .A2(new_n10560_), .A3(new_n10180_), .ZN(new_n10561_));
  XOR2_X1    g10369(.A1(new_n10561_), .A2(new_n10208_), .Z(new_n10562_));
  INV_X1     g10370(.I(new_n10562_), .ZN(new_n10563_));
  NAND3_X1   g10371(.A1(\asqrt[19] ), .A2(new_n10170_), .A3(new_n10171_), .ZN(new_n10564_));
  NAND4_X1   g10372(.A1(new_n10489_), .A2(\asqrt[20] ), .A3(new_n10491_), .A4(new_n10483_), .ZN(new_n10565_));
  AOI21_X1   g10373(.A1(new_n10564_), .A2(new_n10565_), .B(\a[40] ), .ZN(new_n10566_));
  NOR3_X1    g10374(.A1(new_n10478_), .A2(\a[38] ), .A3(\a[39] ), .ZN(new_n10567_));
  INV_X1     g10375(.I(new_n10565_), .ZN(new_n10568_));
  NOR3_X1    g10376(.A1(new_n10567_), .A2(new_n9671_), .A3(new_n10568_), .ZN(new_n10569_));
  NOR2_X1    g10377(.A1(new_n10569_), .A2(new_n10566_), .ZN(new_n10570_));
  INV_X1     g10378(.I(\a[36] ), .ZN(new_n10571_));
  INV_X1     g10379(.I(\a[37] ), .ZN(new_n10572_));
  NAND3_X1   g10380(.A1(new_n10571_), .A2(new_n10572_), .A3(new_n10170_), .ZN(new_n10573_));
  OAI21_X1   g10381(.A1(new_n10478_), .A2(new_n10170_), .B(new_n10573_), .ZN(new_n10574_));
  NAND2_X1   g10382(.A1(new_n10574_), .A2(\asqrt[20] ), .ZN(new_n10575_));
  OAI21_X1   g10383(.A1(new_n10478_), .A2(\a[38] ), .B(\a[39] ), .ZN(new_n10576_));
  NAND2_X1   g10384(.A1(new_n10576_), .A2(new_n10564_), .ZN(new_n10577_));
  NOR2_X1    g10385(.A1(new_n10574_), .A2(\asqrt[20] ), .ZN(new_n10578_));
  OAI21_X1   g10386(.A1(new_n10577_), .A2(new_n10578_), .B(new_n10575_), .ZN(new_n10579_));
  OAI21_X1   g10387(.A1(new_n10579_), .A2(\asqrt[21] ), .B(new_n10570_), .ZN(new_n10580_));
  NAND2_X1   g10388(.A1(new_n10579_), .A2(\asqrt[21] ), .ZN(new_n10581_));
  NAND3_X1   g10389(.A1(new_n10580_), .A2(new_n9177_), .A3(new_n10581_), .ZN(new_n10582_));
  NOR3_X1    g10390(.A1(new_n10478_), .A2(new_n10174_), .A3(new_n10213_), .ZN(new_n10583_));
  XOR2_X1    g10391(.A1(new_n10583_), .A2(new_n10176_), .Z(new_n10584_));
  NAND2_X1   g10392(.A1(new_n10582_), .A2(new_n10584_), .ZN(new_n10585_));
  NAND2_X1   g10393(.A1(new_n10580_), .A2(new_n10581_), .ZN(new_n10586_));
  AOI21_X1   g10394(.A1(new_n10586_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n10587_));
  AOI21_X1   g10395(.A1(new_n10587_), .A2(new_n10585_), .B(new_n10563_), .ZN(new_n10588_));
  OAI21_X1   g10396(.A1(new_n10567_), .A2(new_n10568_), .B(new_n9671_), .ZN(new_n10589_));
  NAND3_X1   g10397(.A1(new_n10564_), .A2(\a[40] ), .A3(new_n10565_), .ZN(new_n10590_));
  NAND2_X1   g10398(.A1(new_n10589_), .A2(new_n10590_), .ZN(new_n10591_));
  NAND2_X1   g10399(.A1(\asqrt[19] ), .A2(\a[38] ), .ZN(new_n10592_));
  AOI21_X1   g10400(.A1(new_n10592_), .A2(new_n10573_), .B(new_n10045_), .ZN(new_n10593_));
  AOI21_X1   g10401(.A1(\asqrt[19] ), .A2(new_n10170_), .B(new_n10171_), .ZN(new_n10594_));
  NOR2_X1    g10402(.A1(new_n10567_), .A2(new_n10594_), .ZN(new_n10595_));
  NAND3_X1   g10403(.A1(new_n10592_), .A2(new_n10045_), .A3(new_n10573_), .ZN(new_n10596_));
  AOI21_X1   g10404(.A1(new_n10595_), .A2(new_n10596_), .B(new_n10593_), .ZN(new_n10597_));
  AOI21_X1   g10405(.A1(new_n10597_), .A2(new_n9590_), .B(new_n10591_), .ZN(new_n10598_));
  NOR2_X1    g10406(.A1(new_n10597_), .A2(new_n9590_), .ZN(new_n10599_));
  OAI21_X1   g10407(.A1(new_n10598_), .A2(new_n10599_), .B(\asqrt[22] ), .ZN(new_n10600_));
  AOI21_X1   g10408(.A1(new_n10585_), .A2(new_n10600_), .B(new_n8742_), .ZN(new_n10601_));
  NOR2_X1    g10409(.A1(new_n10588_), .A2(new_n10601_), .ZN(new_n10602_));
  AOI21_X1   g10410(.A1(new_n10602_), .A2(new_n8349_), .B(new_n10559_), .ZN(new_n10603_));
  OAI21_X1   g10411(.A1(new_n10588_), .A2(new_n10601_), .B(\asqrt[24] ), .ZN(new_n10604_));
  NAND2_X1   g10412(.A1(new_n10604_), .A2(new_n7934_), .ZN(new_n10605_));
  OAI21_X1   g10413(.A1(new_n10603_), .A2(new_n10605_), .B(new_n10556_), .ZN(new_n10606_));
  INV_X1     g10414(.I(new_n10604_), .ZN(new_n10607_));
  OAI21_X1   g10415(.A1(new_n10603_), .A2(new_n10607_), .B(\asqrt[25] ), .ZN(new_n10608_));
  NAND3_X1   g10416(.A1(new_n10606_), .A2(new_n10608_), .A3(new_n7561_), .ZN(new_n10609_));
  NAND2_X1   g10417(.A1(new_n10609_), .A2(new_n10553_), .ZN(new_n10610_));
  NAND2_X1   g10418(.A1(new_n10606_), .A2(new_n10608_), .ZN(new_n10611_));
  AOI21_X1   g10419(.A1(new_n10611_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n10612_));
  AOI21_X1   g10420(.A1(new_n10612_), .A2(new_n10610_), .B(new_n10550_), .ZN(new_n10613_));
  INV_X1     g10421(.I(new_n10556_), .ZN(new_n10614_));
  NOR2_X1    g10422(.A1(new_n10598_), .A2(new_n10599_), .ZN(new_n10615_));
  INV_X1     g10423(.I(new_n10584_), .ZN(new_n10616_));
  AOI21_X1   g10424(.A1(new_n10615_), .A2(new_n9177_), .B(new_n10616_), .ZN(new_n10617_));
  NAND2_X1   g10425(.A1(new_n10600_), .A2(new_n8742_), .ZN(new_n10618_));
  OAI21_X1   g10426(.A1(new_n10617_), .A2(new_n10618_), .B(new_n10562_), .ZN(new_n10619_));
  INV_X1     g10427(.I(new_n10600_), .ZN(new_n10620_));
  OAI21_X1   g10428(.A1(new_n10617_), .A2(new_n10620_), .B(\asqrt[23] ), .ZN(new_n10621_));
  NAND3_X1   g10429(.A1(new_n10619_), .A2(new_n10621_), .A3(new_n8349_), .ZN(new_n10622_));
  NAND2_X1   g10430(.A1(new_n10622_), .A2(new_n10558_), .ZN(new_n10623_));
  NAND2_X1   g10431(.A1(new_n10619_), .A2(new_n10621_), .ZN(new_n10624_));
  AOI21_X1   g10432(.A1(new_n10624_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n10625_));
  AOI21_X1   g10433(.A1(new_n10625_), .A2(new_n10623_), .B(new_n10614_), .ZN(new_n10626_));
  AOI21_X1   g10434(.A1(new_n10623_), .A2(new_n10604_), .B(new_n7934_), .ZN(new_n10627_));
  OAI21_X1   g10435(.A1(new_n10626_), .A2(new_n10627_), .B(\asqrt[26] ), .ZN(new_n10628_));
  AOI21_X1   g10436(.A1(new_n10610_), .A2(new_n10628_), .B(new_n7166_), .ZN(new_n10629_));
  NOR2_X1    g10437(.A1(new_n10613_), .A2(new_n10629_), .ZN(new_n10630_));
  AOI21_X1   g10438(.A1(new_n10630_), .A2(new_n6813_), .B(new_n10547_), .ZN(new_n10631_));
  OAI21_X1   g10439(.A1(new_n10613_), .A2(new_n10629_), .B(\asqrt[28] ), .ZN(new_n10632_));
  NAND2_X1   g10440(.A1(new_n10632_), .A2(new_n6454_), .ZN(new_n10633_));
  OAI21_X1   g10441(.A1(new_n10631_), .A2(new_n10633_), .B(new_n10543_), .ZN(new_n10634_));
  INV_X1     g10442(.I(new_n10632_), .ZN(new_n10635_));
  OAI21_X1   g10443(.A1(new_n10631_), .A2(new_n10635_), .B(\asqrt[29] ), .ZN(new_n10636_));
  NAND3_X1   g10444(.A1(new_n10634_), .A2(new_n10636_), .A3(new_n6106_), .ZN(new_n10637_));
  NAND2_X1   g10445(.A1(new_n10637_), .A2(new_n10541_), .ZN(new_n10638_));
  NAND2_X1   g10446(.A1(new_n10634_), .A2(new_n10636_), .ZN(new_n10639_));
  AOI21_X1   g10447(.A1(new_n10639_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n10640_));
  AOI21_X1   g10448(.A1(new_n10640_), .A2(new_n10638_), .B(new_n10538_), .ZN(new_n10641_));
  INV_X1     g10449(.I(new_n10543_), .ZN(new_n10642_));
  INV_X1     g10450(.I(new_n10553_), .ZN(new_n10643_));
  NOR2_X1    g10451(.A1(new_n10626_), .A2(new_n10627_), .ZN(new_n10644_));
  AOI21_X1   g10452(.A1(new_n10644_), .A2(new_n7561_), .B(new_n10643_), .ZN(new_n10645_));
  NAND2_X1   g10453(.A1(new_n10628_), .A2(new_n7166_), .ZN(new_n10646_));
  OAI21_X1   g10454(.A1(new_n10645_), .A2(new_n10646_), .B(new_n10549_), .ZN(new_n10647_));
  INV_X1     g10455(.I(new_n10628_), .ZN(new_n10648_));
  OAI21_X1   g10456(.A1(new_n10645_), .A2(new_n10648_), .B(\asqrt[27] ), .ZN(new_n10649_));
  NAND3_X1   g10457(.A1(new_n10647_), .A2(new_n10649_), .A3(new_n6813_), .ZN(new_n10650_));
  NAND2_X1   g10458(.A1(new_n10650_), .A2(new_n10546_), .ZN(new_n10651_));
  NAND2_X1   g10459(.A1(new_n10647_), .A2(new_n10649_), .ZN(new_n10652_));
  AOI21_X1   g10460(.A1(new_n10652_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n10653_));
  AOI21_X1   g10461(.A1(new_n10653_), .A2(new_n10651_), .B(new_n10642_), .ZN(new_n10654_));
  AOI21_X1   g10462(.A1(new_n10651_), .A2(new_n10632_), .B(new_n6454_), .ZN(new_n10655_));
  OAI21_X1   g10463(.A1(new_n10654_), .A2(new_n10655_), .B(\asqrt[30] ), .ZN(new_n10656_));
  AOI21_X1   g10464(.A1(new_n10638_), .A2(new_n10656_), .B(new_n5750_), .ZN(new_n10657_));
  NOR2_X1    g10465(.A1(new_n10641_), .A2(new_n10657_), .ZN(new_n10658_));
  AOI21_X1   g10466(.A1(new_n10658_), .A2(new_n5435_), .B(new_n10535_), .ZN(new_n10659_));
  OAI21_X1   g10467(.A1(new_n10641_), .A2(new_n10657_), .B(\asqrt[32] ), .ZN(new_n10660_));
  NAND2_X1   g10468(.A1(new_n10660_), .A2(new_n5110_), .ZN(new_n10661_));
  OAI21_X1   g10469(.A1(new_n10659_), .A2(new_n10661_), .B(new_n10531_), .ZN(new_n10662_));
  INV_X1     g10470(.I(new_n10660_), .ZN(new_n10663_));
  OAI21_X1   g10471(.A1(new_n10659_), .A2(new_n10663_), .B(\asqrt[33] ), .ZN(new_n10664_));
  NAND3_X1   g10472(.A1(new_n10662_), .A2(new_n10664_), .A3(new_n4810_), .ZN(new_n10665_));
  NAND2_X1   g10473(.A1(new_n10665_), .A2(new_n10529_), .ZN(new_n10666_));
  NAND2_X1   g10474(.A1(new_n10662_), .A2(new_n10664_), .ZN(new_n10667_));
  AOI21_X1   g10475(.A1(new_n10667_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n10668_));
  AOI21_X1   g10476(.A1(new_n10668_), .A2(new_n10666_), .B(new_n10526_), .ZN(new_n10669_));
  INV_X1     g10477(.I(new_n10531_), .ZN(new_n10670_));
  INV_X1     g10478(.I(new_n10541_), .ZN(new_n10671_));
  NOR2_X1    g10479(.A1(new_n10654_), .A2(new_n10655_), .ZN(new_n10672_));
  AOI21_X1   g10480(.A1(new_n10672_), .A2(new_n6106_), .B(new_n10671_), .ZN(new_n10673_));
  NAND2_X1   g10481(.A1(new_n10656_), .A2(new_n5750_), .ZN(new_n10674_));
  OAI21_X1   g10482(.A1(new_n10673_), .A2(new_n10674_), .B(new_n10537_), .ZN(new_n10675_));
  INV_X1     g10483(.I(new_n10656_), .ZN(new_n10676_));
  OAI21_X1   g10484(.A1(new_n10673_), .A2(new_n10676_), .B(\asqrt[31] ), .ZN(new_n10677_));
  NAND3_X1   g10485(.A1(new_n10675_), .A2(new_n10677_), .A3(new_n5435_), .ZN(new_n10678_));
  NAND2_X1   g10486(.A1(new_n10678_), .A2(new_n10534_), .ZN(new_n10679_));
  NAND2_X1   g10487(.A1(new_n10675_), .A2(new_n10677_), .ZN(new_n10680_));
  AOI21_X1   g10488(.A1(new_n10680_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n10681_));
  AOI21_X1   g10489(.A1(new_n10681_), .A2(new_n10679_), .B(new_n10670_), .ZN(new_n10682_));
  AOI21_X1   g10490(.A1(new_n10679_), .A2(new_n10660_), .B(new_n5110_), .ZN(new_n10683_));
  OAI21_X1   g10491(.A1(new_n10682_), .A2(new_n10683_), .B(\asqrt[34] ), .ZN(new_n10684_));
  AOI21_X1   g10492(.A1(new_n10666_), .A2(new_n10684_), .B(new_n4510_), .ZN(new_n10685_));
  NOR2_X1    g10493(.A1(new_n10669_), .A2(new_n10685_), .ZN(new_n10686_));
  AOI21_X1   g10494(.A1(new_n10686_), .A2(new_n4224_), .B(new_n10523_), .ZN(new_n10687_));
  OAI21_X1   g10495(.A1(new_n10669_), .A2(new_n10685_), .B(\asqrt[36] ), .ZN(new_n10688_));
  NAND2_X1   g10496(.A1(new_n10688_), .A2(new_n3928_), .ZN(new_n10689_));
  OAI21_X1   g10497(.A1(new_n10687_), .A2(new_n10689_), .B(new_n10519_), .ZN(new_n10690_));
  INV_X1     g10498(.I(new_n10688_), .ZN(new_n10691_));
  OAI21_X1   g10499(.A1(new_n10687_), .A2(new_n10691_), .B(\asqrt[37] ), .ZN(new_n10692_));
  NAND3_X1   g10500(.A1(new_n10690_), .A2(new_n10692_), .A3(new_n3675_), .ZN(new_n10693_));
  NAND2_X1   g10501(.A1(new_n10693_), .A2(new_n10517_), .ZN(new_n10694_));
  NAND2_X1   g10502(.A1(new_n10690_), .A2(new_n10692_), .ZN(new_n10695_));
  AOI21_X1   g10503(.A1(new_n10695_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n10696_));
  AOI21_X1   g10504(.A1(new_n10696_), .A2(new_n10694_), .B(new_n10514_), .ZN(new_n10697_));
  INV_X1     g10505(.I(new_n10519_), .ZN(new_n10698_));
  INV_X1     g10506(.I(new_n10529_), .ZN(new_n10699_));
  NOR2_X1    g10507(.A1(new_n10682_), .A2(new_n10683_), .ZN(new_n10700_));
  AOI21_X1   g10508(.A1(new_n10700_), .A2(new_n4810_), .B(new_n10699_), .ZN(new_n10701_));
  NAND2_X1   g10509(.A1(new_n10684_), .A2(new_n4510_), .ZN(new_n10702_));
  OAI21_X1   g10510(.A1(new_n10701_), .A2(new_n10702_), .B(new_n10525_), .ZN(new_n10703_));
  INV_X1     g10511(.I(new_n10684_), .ZN(new_n10704_));
  OAI21_X1   g10512(.A1(new_n10701_), .A2(new_n10704_), .B(\asqrt[35] ), .ZN(new_n10705_));
  NAND3_X1   g10513(.A1(new_n10703_), .A2(new_n10705_), .A3(new_n4224_), .ZN(new_n10706_));
  NAND2_X1   g10514(.A1(new_n10706_), .A2(new_n10522_), .ZN(new_n10707_));
  NAND2_X1   g10515(.A1(new_n10703_), .A2(new_n10705_), .ZN(new_n10708_));
  AOI21_X1   g10516(.A1(new_n10708_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n10709_));
  AOI21_X1   g10517(.A1(new_n10709_), .A2(new_n10707_), .B(new_n10698_), .ZN(new_n10710_));
  AOI21_X1   g10518(.A1(new_n10707_), .A2(new_n10688_), .B(new_n3928_), .ZN(new_n10711_));
  OAI21_X1   g10519(.A1(new_n10710_), .A2(new_n10711_), .B(\asqrt[38] ), .ZN(new_n10712_));
  AOI21_X1   g10520(.A1(new_n10694_), .A2(new_n10712_), .B(new_n3400_), .ZN(new_n10713_));
  NOR2_X1    g10521(.A1(new_n10697_), .A2(new_n10713_), .ZN(new_n10714_));
  AOI21_X1   g10522(.A1(new_n10714_), .A2(new_n3167_), .B(new_n10511_), .ZN(new_n10715_));
  OAI21_X1   g10523(.A1(new_n10697_), .A2(new_n10713_), .B(\asqrt[40] ), .ZN(new_n10716_));
  NAND2_X1   g10524(.A1(new_n10716_), .A2(new_n2912_), .ZN(new_n10717_));
  OAI21_X1   g10525(.A1(new_n10715_), .A2(new_n10717_), .B(new_n10507_), .ZN(new_n10718_));
  INV_X1     g10526(.I(new_n10716_), .ZN(new_n10719_));
  OAI21_X1   g10527(.A1(new_n10715_), .A2(new_n10719_), .B(\asqrt[41] ), .ZN(new_n10720_));
  NAND3_X1   g10528(.A1(new_n10718_), .A2(new_n10720_), .A3(new_n2699_), .ZN(new_n10721_));
  NAND2_X1   g10529(.A1(new_n10721_), .A2(new_n10505_), .ZN(new_n10722_));
  NAND2_X1   g10530(.A1(new_n10718_), .A2(new_n10720_), .ZN(new_n10723_));
  AOI21_X1   g10531(.A1(new_n10723_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n10724_));
  AOI21_X1   g10532(.A1(new_n10724_), .A2(new_n10722_), .B(new_n10502_), .ZN(new_n10725_));
  INV_X1     g10533(.I(new_n10507_), .ZN(new_n10726_));
  INV_X1     g10534(.I(new_n10517_), .ZN(new_n10727_));
  NOR2_X1    g10535(.A1(new_n10710_), .A2(new_n10711_), .ZN(new_n10728_));
  AOI21_X1   g10536(.A1(new_n10728_), .A2(new_n3675_), .B(new_n10727_), .ZN(new_n10729_));
  NAND2_X1   g10537(.A1(new_n10712_), .A2(new_n3400_), .ZN(new_n10730_));
  OAI21_X1   g10538(.A1(new_n10729_), .A2(new_n10730_), .B(new_n10513_), .ZN(new_n10731_));
  INV_X1     g10539(.I(new_n10712_), .ZN(new_n10732_));
  OAI21_X1   g10540(.A1(new_n10729_), .A2(new_n10732_), .B(\asqrt[39] ), .ZN(new_n10733_));
  NAND3_X1   g10541(.A1(new_n10731_), .A2(new_n10733_), .A3(new_n3167_), .ZN(new_n10734_));
  NAND2_X1   g10542(.A1(new_n10734_), .A2(new_n10510_), .ZN(new_n10735_));
  NAND2_X1   g10543(.A1(new_n10731_), .A2(new_n10733_), .ZN(new_n10736_));
  AOI21_X1   g10544(.A1(new_n10736_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n10737_));
  AOI21_X1   g10545(.A1(new_n10737_), .A2(new_n10735_), .B(new_n10726_), .ZN(new_n10738_));
  AOI21_X1   g10546(.A1(new_n10735_), .A2(new_n10716_), .B(new_n2912_), .ZN(new_n10739_));
  OAI21_X1   g10547(.A1(new_n10738_), .A2(new_n10739_), .B(\asqrt[42] ), .ZN(new_n10740_));
  AOI21_X1   g10548(.A1(new_n10722_), .A2(new_n10740_), .B(new_n2464_), .ZN(new_n10741_));
  NOR2_X1    g10549(.A1(new_n10725_), .A2(new_n10741_), .ZN(new_n10742_));
  AOI21_X1   g10550(.A1(new_n10742_), .A2(new_n2271_), .B(new_n10499_), .ZN(new_n10743_));
  OAI21_X1   g10551(.A1(new_n10725_), .A2(new_n10741_), .B(\asqrt[44] ), .ZN(new_n10744_));
  NAND2_X1   g10552(.A1(new_n10744_), .A2(new_n2072_), .ZN(new_n10745_));
  OAI21_X1   g10553(.A1(new_n10743_), .A2(new_n10745_), .B(new_n10495_), .ZN(new_n10746_));
  INV_X1     g10554(.I(new_n10744_), .ZN(new_n10747_));
  OAI21_X1   g10555(.A1(new_n10743_), .A2(new_n10747_), .B(\asqrt[45] ), .ZN(new_n10748_));
  NAND3_X1   g10556(.A1(new_n10746_), .A2(new_n10748_), .A3(new_n1884_), .ZN(new_n10749_));
  INV_X1     g10557(.I(new_n10495_), .ZN(new_n10750_));
  INV_X1     g10558(.I(new_n10505_), .ZN(new_n10751_));
  NOR2_X1    g10559(.A1(new_n10738_), .A2(new_n10739_), .ZN(new_n10752_));
  AOI21_X1   g10560(.A1(new_n10752_), .A2(new_n2699_), .B(new_n10751_), .ZN(new_n10753_));
  NAND2_X1   g10561(.A1(new_n10740_), .A2(new_n2464_), .ZN(new_n10754_));
  OAI21_X1   g10562(.A1(new_n10753_), .A2(new_n10754_), .B(new_n10501_), .ZN(new_n10755_));
  INV_X1     g10563(.I(new_n10740_), .ZN(new_n10756_));
  OAI21_X1   g10564(.A1(new_n10753_), .A2(new_n10756_), .B(\asqrt[43] ), .ZN(new_n10757_));
  NAND3_X1   g10565(.A1(new_n10755_), .A2(new_n10757_), .A3(new_n2271_), .ZN(new_n10758_));
  NAND2_X1   g10566(.A1(new_n10758_), .A2(new_n10498_), .ZN(new_n10759_));
  NAND2_X1   g10567(.A1(new_n10755_), .A2(new_n10757_), .ZN(new_n10760_));
  AOI21_X1   g10568(.A1(new_n10760_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n10761_));
  AOI21_X1   g10569(.A1(new_n10761_), .A2(new_n10759_), .B(new_n10750_), .ZN(new_n10762_));
  AOI21_X1   g10570(.A1(new_n10759_), .A2(new_n10744_), .B(new_n2072_), .ZN(new_n10763_));
  OAI21_X1   g10571(.A1(new_n10762_), .A2(new_n10763_), .B(\asqrt[46] ), .ZN(new_n10764_));
  NAND2_X1   g10572(.A1(new_n10475_), .A2(new_n10050_), .ZN(new_n10765_));
  NOR2_X1    g10573(.A1(new_n10478_), .A2(new_n10050_), .ZN(new_n10766_));
  NAND2_X1   g10574(.A1(new_n10766_), .A2(new_n10490_), .ZN(new_n10767_));
  AOI21_X1   g10575(.A1(new_n10767_), .A2(new_n10765_), .B(new_n193_), .ZN(new_n10768_));
  INV_X1     g10576(.I(new_n10768_), .ZN(new_n10769_));
  NAND3_X1   g10577(.A1(\asqrt[19] ), .A2(new_n10460_), .A3(new_n10471_), .ZN(new_n10770_));
  XOR2_X1    g10578(.A1(new_n10770_), .A2(new_n10463_), .Z(new_n10771_));
  AOI21_X1   g10579(.A1(new_n10766_), .A2(new_n10475_), .B(new_n10476_), .ZN(new_n10772_));
  OAI21_X1   g10580(.A1(new_n10430_), .A2(new_n10432_), .B(new_n10435_), .ZN(new_n10773_));
  NOR2_X1    g10581(.A1(new_n10478_), .A2(new_n10773_), .ZN(new_n10774_));
  XOR2_X1    g10582(.A1(new_n10774_), .A2(new_n10058_), .Z(new_n10775_));
  NAND3_X1   g10583(.A1(\asqrt[19] ), .A2(new_n10446_), .A3(new_n10431_), .ZN(new_n10776_));
  XOR2_X1    g10584(.A1(new_n10776_), .A2(new_n10062_), .Z(new_n10777_));
  OAI21_X1   g10585(.A1(new_n10441_), .A2(new_n10442_), .B(new_n10445_), .ZN(new_n10778_));
  NOR2_X1    g10586(.A1(new_n10478_), .A2(new_n10778_), .ZN(new_n10779_));
  XOR2_X1    g10587(.A1(new_n10779_), .A2(new_n10064_), .Z(new_n10780_));
  INV_X1     g10588(.I(new_n10780_), .ZN(new_n10781_));
  NAND3_X1   g10589(.A1(\asqrt[19] ), .A2(new_n10408_), .A3(new_n10427_), .ZN(new_n10782_));
  XOR2_X1    g10590(.A1(new_n10782_), .A2(new_n10439_), .Z(new_n10783_));
  INV_X1     g10591(.I(new_n10783_), .ZN(new_n10784_));
  OAI21_X1   g10592(.A1(new_n10402_), .A2(new_n10404_), .B(new_n10407_), .ZN(new_n10785_));
  NOR2_X1    g10593(.A1(new_n10478_), .A2(new_n10785_), .ZN(new_n10786_));
  XOR2_X1    g10594(.A1(new_n10786_), .A2(new_n10070_), .Z(new_n10787_));
  NAND3_X1   g10595(.A1(\asqrt[19] ), .A2(new_n10421_), .A3(new_n10403_), .ZN(new_n10788_));
  XOR2_X1    g10596(.A1(new_n10788_), .A2(new_n10074_), .Z(new_n10789_));
  OAI21_X1   g10597(.A1(new_n10416_), .A2(new_n10417_), .B(new_n10420_), .ZN(new_n10790_));
  NOR2_X1    g10598(.A1(new_n10478_), .A2(new_n10790_), .ZN(new_n10791_));
  XOR2_X1    g10599(.A1(new_n10791_), .A2(new_n10076_), .Z(new_n10792_));
  INV_X1     g10600(.I(new_n10792_), .ZN(new_n10793_));
  NAND3_X1   g10601(.A1(\asqrt[19] ), .A2(new_n10380_), .A3(new_n10399_), .ZN(new_n10794_));
  XOR2_X1    g10602(.A1(new_n10794_), .A2(new_n10414_), .Z(new_n10795_));
  INV_X1     g10603(.I(new_n10795_), .ZN(new_n10796_));
  OAI21_X1   g10604(.A1(new_n10374_), .A2(new_n10376_), .B(new_n10379_), .ZN(new_n10797_));
  NOR2_X1    g10605(.A1(new_n10478_), .A2(new_n10797_), .ZN(new_n10798_));
  XOR2_X1    g10606(.A1(new_n10798_), .A2(new_n10082_), .Z(new_n10799_));
  NAND3_X1   g10607(.A1(\asqrt[19] ), .A2(new_n10393_), .A3(new_n10375_), .ZN(new_n10800_));
  XOR2_X1    g10608(.A1(new_n10800_), .A2(new_n10086_), .Z(new_n10801_));
  OAI21_X1   g10609(.A1(new_n10388_), .A2(new_n10389_), .B(new_n10392_), .ZN(new_n10802_));
  NOR2_X1    g10610(.A1(new_n10478_), .A2(new_n10802_), .ZN(new_n10803_));
  XOR2_X1    g10611(.A1(new_n10803_), .A2(new_n10088_), .Z(new_n10804_));
  INV_X1     g10612(.I(new_n10804_), .ZN(new_n10805_));
  NAND3_X1   g10613(.A1(\asqrt[19] ), .A2(new_n10352_), .A3(new_n10371_), .ZN(new_n10806_));
  XOR2_X1    g10614(.A1(new_n10806_), .A2(new_n10386_), .Z(new_n10807_));
  INV_X1     g10615(.I(new_n10807_), .ZN(new_n10808_));
  OAI21_X1   g10616(.A1(new_n10346_), .A2(new_n10348_), .B(new_n10351_), .ZN(new_n10809_));
  NOR2_X1    g10617(.A1(new_n10478_), .A2(new_n10809_), .ZN(new_n10810_));
  XOR2_X1    g10618(.A1(new_n10810_), .A2(new_n10094_), .Z(new_n10811_));
  NAND3_X1   g10619(.A1(\asqrt[19] ), .A2(new_n10365_), .A3(new_n10347_), .ZN(new_n10812_));
  XOR2_X1    g10620(.A1(new_n10812_), .A2(new_n10098_), .Z(new_n10813_));
  NOR2_X1    g10621(.A1(new_n10762_), .A2(new_n10763_), .ZN(new_n10814_));
  AOI21_X1   g10622(.A1(new_n10814_), .A2(new_n1884_), .B(new_n10482_), .ZN(new_n10815_));
  NAND2_X1   g10623(.A1(new_n10764_), .A2(new_n1688_), .ZN(new_n10816_));
  OAI21_X1   g10624(.A1(new_n10815_), .A2(new_n10816_), .B(new_n10813_), .ZN(new_n10817_));
  INV_X1     g10625(.I(new_n10764_), .ZN(new_n10818_));
  OAI21_X1   g10626(.A1(new_n10815_), .A2(new_n10818_), .B(\asqrt[47] ), .ZN(new_n10819_));
  NAND3_X1   g10627(.A1(new_n10817_), .A2(new_n10819_), .A3(new_n1533_), .ZN(new_n10820_));
  NAND2_X1   g10628(.A1(new_n10820_), .A2(new_n10811_), .ZN(new_n10821_));
  NAND2_X1   g10629(.A1(new_n10817_), .A2(new_n10819_), .ZN(new_n10822_));
  AOI21_X1   g10630(.A1(new_n10822_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n10823_));
  AOI21_X1   g10631(.A1(new_n10823_), .A2(new_n10821_), .B(new_n10808_), .ZN(new_n10824_));
  INV_X1     g10632(.I(new_n10813_), .ZN(new_n10825_));
  NAND2_X1   g10633(.A1(new_n10749_), .A2(new_n10481_), .ZN(new_n10826_));
  NAND2_X1   g10634(.A1(new_n10746_), .A2(new_n10748_), .ZN(new_n10827_));
  AOI21_X1   g10635(.A1(new_n10827_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n10828_));
  AOI21_X1   g10636(.A1(new_n10828_), .A2(new_n10826_), .B(new_n10825_), .ZN(new_n10829_));
  AOI21_X1   g10637(.A1(new_n10826_), .A2(new_n10764_), .B(new_n1688_), .ZN(new_n10830_));
  OAI21_X1   g10638(.A1(new_n10829_), .A2(new_n10830_), .B(\asqrt[48] ), .ZN(new_n10831_));
  AOI21_X1   g10639(.A1(new_n10821_), .A2(new_n10831_), .B(new_n1368_), .ZN(new_n10832_));
  NOR2_X1    g10640(.A1(new_n10824_), .A2(new_n10832_), .ZN(new_n10833_));
  AOI21_X1   g10641(.A1(new_n10833_), .A2(new_n1228_), .B(new_n10805_), .ZN(new_n10834_));
  OAI21_X1   g10642(.A1(new_n10824_), .A2(new_n10832_), .B(\asqrt[50] ), .ZN(new_n10835_));
  NAND2_X1   g10643(.A1(new_n10835_), .A2(new_n1088_), .ZN(new_n10836_));
  OAI21_X1   g10644(.A1(new_n10834_), .A2(new_n10836_), .B(new_n10801_), .ZN(new_n10837_));
  INV_X1     g10645(.I(new_n10835_), .ZN(new_n10838_));
  OAI21_X1   g10646(.A1(new_n10834_), .A2(new_n10838_), .B(\asqrt[51] ), .ZN(new_n10839_));
  NAND3_X1   g10647(.A1(new_n10837_), .A2(new_n10839_), .A3(new_n962_), .ZN(new_n10840_));
  NAND2_X1   g10648(.A1(new_n10840_), .A2(new_n10799_), .ZN(new_n10841_));
  NAND2_X1   g10649(.A1(new_n10837_), .A2(new_n10839_), .ZN(new_n10842_));
  AOI21_X1   g10650(.A1(new_n10842_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n10843_));
  AOI21_X1   g10651(.A1(new_n10843_), .A2(new_n10841_), .B(new_n10796_), .ZN(new_n10844_));
  INV_X1     g10652(.I(new_n10801_), .ZN(new_n10845_));
  INV_X1     g10653(.I(new_n10811_), .ZN(new_n10846_));
  NOR2_X1    g10654(.A1(new_n10829_), .A2(new_n10830_), .ZN(new_n10847_));
  AOI21_X1   g10655(.A1(new_n10847_), .A2(new_n1533_), .B(new_n10846_), .ZN(new_n10848_));
  NAND2_X1   g10656(.A1(new_n10831_), .A2(new_n1368_), .ZN(new_n10849_));
  OAI21_X1   g10657(.A1(new_n10848_), .A2(new_n10849_), .B(new_n10807_), .ZN(new_n10850_));
  INV_X1     g10658(.I(new_n10831_), .ZN(new_n10851_));
  OAI21_X1   g10659(.A1(new_n10848_), .A2(new_n10851_), .B(\asqrt[49] ), .ZN(new_n10852_));
  NAND3_X1   g10660(.A1(new_n10850_), .A2(new_n10852_), .A3(new_n1228_), .ZN(new_n10853_));
  NAND2_X1   g10661(.A1(new_n10853_), .A2(new_n10804_), .ZN(new_n10854_));
  NAND2_X1   g10662(.A1(new_n10850_), .A2(new_n10852_), .ZN(new_n10855_));
  AOI21_X1   g10663(.A1(new_n10855_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n10856_));
  AOI21_X1   g10664(.A1(new_n10856_), .A2(new_n10854_), .B(new_n10845_), .ZN(new_n10857_));
  AOI21_X1   g10665(.A1(new_n10854_), .A2(new_n10835_), .B(new_n1088_), .ZN(new_n10858_));
  OAI21_X1   g10666(.A1(new_n10857_), .A2(new_n10858_), .B(\asqrt[52] ), .ZN(new_n10859_));
  AOI21_X1   g10667(.A1(new_n10841_), .A2(new_n10859_), .B(new_n842_), .ZN(new_n10860_));
  NOR2_X1    g10668(.A1(new_n10844_), .A2(new_n10860_), .ZN(new_n10861_));
  AOI21_X1   g10669(.A1(new_n10861_), .A2(new_n720_), .B(new_n10793_), .ZN(new_n10862_));
  OAI21_X1   g10670(.A1(new_n10844_), .A2(new_n10860_), .B(\asqrt[54] ), .ZN(new_n10863_));
  NAND2_X1   g10671(.A1(new_n10863_), .A2(new_n630_), .ZN(new_n10864_));
  OAI21_X1   g10672(.A1(new_n10862_), .A2(new_n10864_), .B(new_n10789_), .ZN(new_n10865_));
  INV_X1     g10673(.I(new_n10863_), .ZN(new_n10866_));
  OAI21_X1   g10674(.A1(new_n10862_), .A2(new_n10866_), .B(\asqrt[55] ), .ZN(new_n10867_));
  NAND3_X1   g10675(.A1(new_n10865_), .A2(new_n10867_), .A3(new_n545_), .ZN(new_n10868_));
  NAND2_X1   g10676(.A1(new_n10868_), .A2(new_n10787_), .ZN(new_n10869_));
  NAND2_X1   g10677(.A1(new_n10865_), .A2(new_n10867_), .ZN(new_n10870_));
  AOI21_X1   g10678(.A1(new_n10870_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n10871_));
  AOI21_X1   g10679(.A1(new_n10871_), .A2(new_n10869_), .B(new_n10784_), .ZN(new_n10872_));
  INV_X1     g10680(.I(new_n10789_), .ZN(new_n10873_));
  INV_X1     g10681(.I(new_n10799_), .ZN(new_n10874_));
  NOR2_X1    g10682(.A1(new_n10857_), .A2(new_n10858_), .ZN(new_n10875_));
  AOI21_X1   g10683(.A1(new_n10875_), .A2(new_n962_), .B(new_n10874_), .ZN(new_n10876_));
  NAND2_X1   g10684(.A1(new_n10859_), .A2(new_n842_), .ZN(new_n10877_));
  OAI21_X1   g10685(.A1(new_n10876_), .A2(new_n10877_), .B(new_n10795_), .ZN(new_n10878_));
  INV_X1     g10686(.I(new_n10859_), .ZN(new_n10879_));
  OAI21_X1   g10687(.A1(new_n10876_), .A2(new_n10879_), .B(\asqrt[53] ), .ZN(new_n10880_));
  NAND3_X1   g10688(.A1(new_n10878_), .A2(new_n10880_), .A3(new_n720_), .ZN(new_n10881_));
  NAND2_X1   g10689(.A1(new_n10881_), .A2(new_n10792_), .ZN(new_n10882_));
  NAND2_X1   g10690(.A1(new_n10878_), .A2(new_n10880_), .ZN(new_n10883_));
  AOI21_X1   g10691(.A1(new_n10883_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n10884_));
  AOI21_X1   g10692(.A1(new_n10884_), .A2(new_n10882_), .B(new_n10873_), .ZN(new_n10885_));
  AOI21_X1   g10693(.A1(new_n10882_), .A2(new_n10863_), .B(new_n630_), .ZN(new_n10886_));
  OAI21_X1   g10694(.A1(new_n10885_), .A2(new_n10886_), .B(\asqrt[56] ), .ZN(new_n10887_));
  AOI21_X1   g10695(.A1(new_n10869_), .A2(new_n10887_), .B(new_n450_), .ZN(new_n10888_));
  NOR2_X1    g10696(.A1(new_n10872_), .A2(new_n10888_), .ZN(new_n10889_));
  AOI21_X1   g10697(.A1(new_n10889_), .A2(new_n403_), .B(new_n10781_), .ZN(new_n10890_));
  OAI21_X1   g10698(.A1(new_n10872_), .A2(new_n10888_), .B(\asqrt[58] ), .ZN(new_n10891_));
  NAND2_X1   g10699(.A1(new_n10891_), .A2(new_n339_), .ZN(new_n10892_));
  OAI21_X1   g10700(.A1(new_n10890_), .A2(new_n10892_), .B(new_n10777_), .ZN(new_n10893_));
  INV_X1     g10701(.I(new_n10891_), .ZN(new_n10894_));
  OAI21_X1   g10702(.A1(new_n10890_), .A2(new_n10894_), .B(\asqrt[59] ), .ZN(new_n10895_));
  NAND3_X1   g10703(.A1(new_n10893_), .A2(new_n10895_), .A3(new_n288_), .ZN(new_n10896_));
  NAND2_X1   g10704(.A1(new_n10896_), .A2(new_n10775_), .ZN(new_n10897_));
  INV_X1     g10705(.I(new_n10777_), .ZN(new_n10898_));
  INV_X1     g10706(.I(new_n10787_), .ZN(new_n10899_));
  NOR2_X1    g10707(.A1(new_n10885_), .A2(new_n10886_), .ZN(new_n10900_));
  AOI21_X1   g10708(.A1(new_n10900_), .A2(new_n545_), .B(new_n10899_), .ZN(new_n10901_));
  NAND2_X1   g10709(.A1(new_n10887_), .A2(new_n450_), .ZN(new_n10902_));
  OAI21_X1   g10710(.A1(new_n10901_), .A2(new_n10902_), .B(new_n10783_), .ZN(new_n10903_));
  INV_X1     g10711(.I(new_n10887_), .ZN(new_n10904_));
  OAI21_X1   g10712(.A1(new_n10901_), .A2(new_n10904_), .B(\asqrt[57] ), .ZN(new_n10905_));
  NAND3_X1   g10713(.A1(new_n10903_), .A2(new_n10905_), .A3(new_n403_), .ZN(new_n10906_));
  NAND2_X1   g10714(.A1(new_n10906_), .A2(new_n10780_), .ZN(new_n10907_));
  NAND2_X1   g10715(.A1(new_n10903_), .A2(new_n10905_), .ZN(new_n10908_));
  AOI21_X1   g10716(.A1(new_n10908_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n10909_));
  AOI21_X1   g10717(.A1(new_n10909_), .A2(new_n10907_), .B(new_n10898_), .ZN(new_n10910_));
  AOI21_X1   g10718(.A1(new_n10907_), .A2(new_n10891_), .B(new_n339_), .ZN(new_n10911_));
  OAI21_X1   g10719(.A1(new_n10910_), .A2(new_n10911_), .B(\asqrt[60] ), .ZN(new_n10912_));
  AOI21_X1   g10720(.A1(new_n10897_), .A2(new_n10912_), .B(new_n242_), .ZN(new_n10913_));
  NAND3_X1   g10721(.A1(\asqrt[19] ), .A2(new_n10436_), .A3(new_n10452_), .ZN(new_n10914_));
  XOR2_X1    g10722(.A1(new_n10914_), .A2(new_n10464_), .Z(new_n10915_));
  INV_X1     g10723(.I(new_n10915_), .ZN(new_n10916_));
  NAND2_X1   g10724(.A1(new_n10893_), .A2(new_n10895_), .ZN(new_n10917_));
  AOI21_X1   g10725(.A1(new_n10917_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n10918_));
  AOI21_X1   g10726(.A1(new_n10918_), .A2(new_n10897_), .B(new_n10916_), .ZN(new_n10919_));
  OAI21_X1   g10727(.A1(new_n10919_), .A2(new_n10913_), .B(\asqrt[62] ), .ZN(new_n10920_));
  INV_X1     g10728(.I(new_n10920_), .ZN(new_n10921_));
  NOR2_X1    g10729(.A1(new_n10919_), .A2(new_n10913_), .ZN(new_n10922_));
  AOI21_X1   g10730(.A1(new_n10437_), .A2(new_n10458_), .B(new_n10453_), .ZN(new_n10923_));
  NAND2_X1   g10731(.A1(\asqrt[19] ), .A2(new_n10923_), .ZN(new_n10924_));
  XOR2_X1    g10732(.A1(new_n10924_), .A2(new_n10456_), .Z(new_n10925_));
  INV_X1     g10733(.I(new_n10925_), .ZN(new_n10926_));
  AOI21_X1   g10734(.A1(new_n10922_), .A2(new_n234_), .B(new_n10926_), .ZN(new_n10927_));
  OAI21_X1   g10735(.A1(new_n10927_), .A2(new_n10921_), .B(new_n10772_), .ZN(new_n10928_));
  OAI21_X1   g10736(.A1(new_n10928_), .A2(new_n10771_), .B(new_n193_), .ZN(new_n10929_));
  NOR2_X1    g10737(.A1(new_n10927_), .A2(new_n10921_), .ZN(new_n10930_));
  NAND2_X1   g10738(.A1(new_n10930_), .A2(new_n10771_), .ZN(new_n10931_));
  NOR2_X1    g10739(.A1(\asqrt[19] ), .A2(new_n10051_), .ZN(new_n10932_));
  INV_X1     g10740(.I(new_n10932_), .ZN(new_n10933_));
  NAND4_X1   g10741(.A1(new_n10929_), .A2(new_n10769_), .A3(new_n10931_), .A4(new_n10933_), .ZN(\asqrt[18] ));
  NAND3_X1   g10742(.A1(\asqrt[18] ), .A2(new_n10749_), .A3(new_n10764_), .ZN(new_n10935_));
  XOR2_X1    g10743(.A1(new_n10935_), .A2(new_n10482_), .Z(new_n10936_));
  INV_X1     g10744(.I(new_n10775_), .ZN(new_n10937_));
  NOR2_X1    g10745(.A1(new_n10910_), .A2(new_n10911_), .ZN(new_n10938_));
  AOI21_X1   g10746(.A1(new_n10938_), .A2(new_n288_), .B(new_n10937_), .ZN(new_n10939_));
  INV_X1     g10747(.I(new_n10912_), .ZN(new_n10940_));
  OAI21_X1   g10748(.A1(new_n10939_), .A2(new_n10940_), .B(\asqrt[61] ), .ZN(new_n10941_));
  NAND2_X1   g10749(.A1(new_n10912_), .A2(new_n242_), .ZN(new_n10942_));
  OAI21_X1   g10750(.A1(new_n10939_), .A2(new_n10942_), .B(new_n10915_), .ZN(new_n10943_));
  NAND3_X1   g10751(.A1(new_n10943_), .A2(new_n10941_), .A3(new_n234_), .ZN(new_n10944_));
  NAND2_X1   g10752(.A1(new_n10944_), .A2(new_n10925_), .ZN(new_n10945_));
  NAND2_X1   g10753(.A1(new_n10945_), .A2(new_n10920_), .ZN(new_n10946_));
  NAND2_X1   g10754(.A1(new_n10946_), .A2(new_n10771_), .ZN(new_n10947_));
  INV_X1     g10755(.I(new_n10771_), .ZN(new_n10948_));
  INV_X1     g10756(.I(new_n10772_), .ZN(new_n10949_));
  AOI21_X1   g10757(.A1(new_n10945_), .A2(new_n10920_), .B(new_n10949_), .ZN(new_n10950_));
  AOI21_X1   g10758(.A1(new_n10950_), .A2(new_n10948_), .B(\asqrt[63] ), .ZN(new_n10951_));
  NOR2_X1    g10759(.A1(new_n10946_), .A2(new_n10948_), .ZN(new_n10952_));
  NOR4_X1    g10760(.A1(new_n10951_), .A2(new_n10768_), .A3(new_n10952_), .A4(new_n10932_), .ZN(new_n10953_));
  NOR2_X1    g10761(.A1(new_n10953_), .A2(new_n10771_), .ZN(new_n10954_));
  NAND2_X1   g10762(.A1(new_n10954_), .A2(new_n10930_), .ZN(new_n10955_));
  AOI21_X1   g10763(.A1(new_n10955_), .A2(new_n10947_), .B(new_n193_), .ZN(new_n10956_));
  NAND3_X1   g10764(.A1(\asqrt[18] ), .A2(new_n10920_), .A3(new_n10944_), .ZN(new_n10957_));
  XOR2_X1    g10765(.A1(new_n10957_), .A2(new_n10925_), .Z(new_n10958_));
  INV_X1     g10766(.I(new_n10958_), .ZN(new_n10959_));
  AOI21_X1   g10767(.A1(new_n10954_), .A2(new_n10946_), .B(new_n10952_), .ZN(new_n10960_));
  INV_X1     g10768(.I(new_n10960_), .ZN(new_n10961_));
  OAI21_X1   g10769(.A1(new_n10890_), .A2(new_n10892_), .B(new_n10895_), .ZN(new_n10962_));
  NOR2_X1    g10770(.A1(new_n10953_), .A2(new_n10962_), .ZN(new_n10963_));
  XOR2_X1    g10771(.A1(new_n10963_), .A2(new_n10777_), .Z(new_n10964_));
  NAND3_X1   g10772(.A1(\asqrt[18] ), .A2(new_n10906_), .A3(new_n10891_), .ZN(new_n10965_));
  XOR2_X1    g10773(.A1(new_n10965_), .A2(new_n10781_), .Z(new_n10966_));
  OAI21_X1   g10774(.A1(new_n10901_), .A2(new_n10902_), .B(new_n10905_), .ZN(new_n10967_));
  NOR2_X1    g10775(.A1(new_n10953_), .A2(new_n10967_), .ZN(new_n10968_));
  XOR2_X1    g10776(.A1(new_n10968_), .A2(new_n10783_), .Z(new_n10969_));
  INV_X1     g10777(.I(new_n10969_), .ZN(new_n10970_));
  NAND3_X1   g10778(.A1(\asqrt[18] ), .A2(new_n10868_), .A3(new_n10887_), .ZN(new_n10971_));
  XOR2_X1    g10779(.A1(new_n10971_), .A2(new_n10899_), .Z(new_n10972_));
  INV_X1     g10780(.I(new_n10972_), .ZN(new_n10973_));
  OAI21_X1   g10781(.A1(new_n10862_), .A2(new_n10864_), .B(new_n10867_), .ZN(new_n10974_));
  NOR2_X1    g10782(.A1(new_n10953_), .A2(new_n10974_), .ZN(new_n10975_));
  XOR2_X1    g10783(.A1(new_n10975_), .A2(new_n10789_), .Z(new_n10976_));
  NAND3_X1   g10784(.A1(\asqrt[18] ), .A2(new_n10881_), .A3(new_n10863_), .ZN(new_n10977_));
  XOR2_X1    g10785(.A1(new_n10977_), .A2(new_n10793_), .Z(new_n10978_));
  OAI21_X1   g10786(.A1(new_n10876_), .A2(new_n10877_), .B(new_n10880_), .ZN(new_n10979_));
  NOR2_X1    g10787(.A1(new_n10953_), .A2(new_n10979_), .ZN(new_n10980_));
  XOR2_X1    g10788(.A1(new_n10980_), .A2(new_n10795_), .Z(new_n10981_));
  INV_X1     g10789(.I(new_n10981_), .ZN(new_n10982_));
  NAND3_X1   g10790(.A1(\asqrt[18] ), .A2(new_n10840_), .A3(new_n10859_), .ZN(new_n10983_));
  XOR2_X1    g10791(.A1(new_n10983_), .A2(new_n10874_), .Z(new_n10984_));
  INV_X1     g10792(.I(new_n10984_), .ZN(new_n10985_));
  OAI21_X1   g10793(.A1(new_n10834_), .A2(new_n10836_), .B(new_n10839_), .ZN(new_n10986_));
  NOR2_X1    g10794(.A1(new_n10953_), .A2(new_n10986_), .ZN(new_n10987_));
  XOR2_X1    g10795(.A1(new_n10987_), .A2(new_n10801_), .Z(new_n10988_));
  NAND3_X1   g10796(.A1(\asqrt[18] ), .A2(new_n10853_), .A3(new_n10835_), .ZN(new_n10989_));
  XOR2_X1    g10797(.A1(new_n10989_), .A2(new_n10805_), .Z(new_n10990_));
  OAI21_X1   g10798(.A1(new_n10848_), .A2(new_n10849_), .B(new_n10852_), .ZN(new_n10991_));
  NOR2_X1    g10799(.A1(new_n10953_), .A2(new_n10991_), .ZN(new_n10992_));
  XOR2_X1    g10800(.A1(new_n10992_), .A2(new_n10807_), .Z(new_n10993_));
  INV_X1     g10801(.I(new_n10993_), .ZN(new_n10994_));
  NAND3_X1   g10802(.A1(\asqrt[18] ), .A2(new_n10820_), .A3(new_n10831_), .ZN(new_n10995_));
  XOR2_X1    g10803(.A1(new_n10995_), .A2(new_n10846_), .Z(new_n10996_));
  INV_X1     g10804(.I(new_n10996_), .ZN(new_n10997_));
  OAI21_X1   g10805(.A1(new_n10815_), .A2(new_n10816_), .B(new_n10819_), .ZN(new_n10998_));
  NOR2_X1    g10806(.A1(new_n10953_), .A2(new_n10998_), .ZN(new_n10999_));
  XOR2_X1    g10807(.A1(new_n10999_), .A2(new_n10813_), .Z(new_n11000_));
  OAI21_X1   g10808(.A1(new_n10743_), .A2(new_n10745_), .B(new_n10748_), .ZN(new_n11001_));
  NOR2_X1    g10809(.A1(new_n10953_), .A2(new_n11001_), .ZN(new_n11002_));
  XOR2_X1    g10810(.A1(new_n11002_), .A2(new_n10495_), .Z(new_n11003_));
  INV_X1     g10811(.I(new_n11003_), .ZN(new_n11004_));
  NAND3_X1   g10812(.A1(\asqrt[18] ), .A2(new_n10758_), .A3(new_n10744_), .ZN(new_n11005_));
  XOR2_X1    g10813(.A1(new_n11005_), .A2(new_n10499_), .Z(new_n11006_));
  INV_X1     g10814(.I(new_n11006_), .ZN(new_n11007_));
  OAI21_X1   g10815(.A1(new_n10753_), .A2(new_n10754_), .B(new_n10757_), .ZN(new_n11008_));
  NOR2_X1    g10816(.A1(new_n10953_), .A2(new_n11008_), .ZN(new_n11009_));
  XOR2_X1    g10817(.A1(new_n11009_), .A2(new_n10501_), .Z(new_n11010_));
  NAND3_X1   g10818(.A1(\asqrt[18] ), .A2(new_n10721_), .A3(new_n10740_), .ZN(new_n11011_));
  XOR2_X1    g10819(.A1(new_n11011_), .A2(new_n10751_), .Z(new_n11012_));
  OAI21_X1   g10820(.A1(new_n10715_), .A2(new_n10717_), .B(new_n10720_), .ZN(new_n11013_));
  NOR2_X1    g10821(.A1(new_n10953_), .A2(new_n11013_), .ZN(new_n11014_));
  XOR2_X1    g10822(.A1(new_n11014_), .A2(new_n10507_), .Z(new_n11015_));
  INV_X1     g10823(.I(new_n11015_), .ZN(new_n11016_));
  NAND3_X1   g10824(.A1(\asqrt[18] ), .A2(new_n10734_), .A3(new_n10716_), .ZN(new_n11017_));
  XOR2_X1    g10825(.A1(new_n11017_), .A2(new_n10511_), .Z(new_n11018_));
  INV_X1     g10826(.I(new_n11018_), .ZN(new_n11019_));
  OAI21_X1   g10827(.A1(new_n10729_), .A2(new_n10730_), .B(new_n10733_), .ZN(new_n11020_));
  NOR2_X1    g10828(.A1(new_n10953_), .A2(new_n11020_), .ZN(new_n11021_));
  XOR2_X1    g10829(.A1(new_n11021_), .A2(new_n10513_), .Z(new_n11022_));
  NAND3_X1   g10830(.A1(\asqrt[18] ), .A2(new_n10693_), .A3(new_n10712_), .ZN(new_n11023_));
  XOR2_X1    g10831(.A1(new_n11023_), .A2(new_n10727_), .Z(new_n11024_));
  OAI21_X1   g10832(.A1(new_n10687_), .A2(new_n10689_), .B(new_n10692_), .ZN(new_n11025_));
  NOR2_X1    g10833(.A1(new_n10953_), .A2(new_n11025_), .ZN(new_n11026_));
  XOR2_X1    g10834(.A1(new_n11026_), .A2(new_n10519_), .Z(new_n11027_));
  INV_X1     g10835(.I(new_n11027_), .ZN(new_n11028_));
  NAND3_X1   g10836(.A1(\asqrt[18] ), .A2(new_n10706_), .A3(new_n10688_), .ZN(new_n11029_));
  XOR2_X1    g10837(.A1(new_n11029_), .A2(new_n10523_), .Z(new_n11030_));
  INV_X1     g10838(.I(new_n11030_), .ZN(new_n11031_));
  OAI21_X1   g10839(.A1(new_n10701_), .A2(new_n10702_), .B(new_n10705_), .ZN(new_n11032_));
  NOR2_X1    g10840(.A1(new_n10953_), .A2(new_n11032_), .ZN(new_n11033_));
  XOR2_X1    g10841(.A1(new_n11033_), .A2(new_n10525_), .Z(new_n11034_));
  NAND3_X1   g10842(.A1(\asqrt[18] ), .A2(new_n10665_), .A3(new_n10684_), .ZN(new_n11035_));
  XOR2_X1    g10843(.A1(new_n11035_), .A2(new_n10699_), .Z(new_n11036_));
  OAI21_X1   g10844(.A1(new_n10659_), .A2(new_n10661_), .B(new_n10664_), .ZN(new_n11037_));
  NOR2_X1    g10845(.A1(new_n10953_), .A2(new_n11037_), .ZN(new_n11038_));
  XOR2_X1    g10846(.A1(new_n11038_), .A2(new_n10531_), .Z(new_n11039_));
  INV_X1     g10847(.I(new_n11039_), .ZN(new_n11040_));
  NAND3_X1   g10848(.A1(\asqrt[18] ), .A2(new_n10678_), .A3(new_n10660_), .ZN(new_n11041_));
  XOR2_X1    g10849(.A1(new_n11041_), .A2(new_n10535_), .Z(new_n11042_));
  INV_X1     g10850(.I(new_n11042_), .ZN(new_n11043_));
  OAI21_X1   g10851(.A1(new_n10673_), .A2(new_n10674_), .B(new_n10677_), .ZN(new_n11044_));
  NOR2_X1    g10852(.A1(new_n10953_), .A2(new_n11044_), .ZN(new_n11045_));
  XOR2_X1    g10853(.A1(new_n11045_), .A2(new_n10537_), .Z(new_n11046_));
  NAND3_X1   g10854(.A1(\asqrt[18] ), .A2(new_n10637_), .A3(new_n10656_), .ZN(new_n11047_));
  XOR2_X1    g10855(.A1(new_n11047_), .A2(new_n10671_), .Z(new_n11048_));
  OAI21_X1   g10856(.A1(new_n10631_), .A2(new_n10633_), .B(new_n10636_), .ZN(new_n11049_));
  NOR2_X1    g10857(.A1(new_n10953_), .A2(new_n11049_), .ZN(new_n11050_));
  XOR2_X1    g10858(.A1(new_n11050_), .A2(new_n10543_), .Z(new_n11051_));
  INV_X1     g10859(.I(new_n11051_), .ZN(new_n11052_));
  NAND3_X1   g10860(.A1(\asqrt[18] ), .A2(new_n10650_), .A3(new_n10632_), .ZN(new_n11053_));
  XOR2_X1    g10861(.A1(new_n11053_), .A2(new_n10547_), .Z(new_n11054_));
  INV_X1     g10862(.I(new_n11054_), .ZN(new_n11055_));
  OAI21_X1   g10863(.A1(new_n10645_), .A2(new_n10646_), .B(new_n10649_), .ZN(new_n11056_));
  NOR2_X1    g10864(.A1(new_n10953_), .A2(new_n11056_), .ZN(new_n11057_));
  XOR2_X1    g10865(.A1(new_n11057_), .A2(new_n10549_), .Z(new_n11058_));
  NAND3_X1   g10866(.A1(\asqrt[18] ), .A2(new_n10609_), .A3(new_n10628_), .ZN(new_n11059_));
  XOR2_X1    g10867(.A1(new_n11059_), .A2(new_n10643_), .Z(new_n11060_));
  OAI21_X1   g10868(.A1(new_n10603_), .A2(new_n10605_), .B(new_n10608_), .ZN(new_n11061_));
  NOR2_X1    g10869(.A1(new_n10953_), .A2(new_n11061_), .ZN(new_n11062_));
  XOR2_X1    g10870(.A1(new_n11062_), .A2(new_n10556_), .Z(new_n11063_));
  INV_X1     g10871(.I(new_n11063_), .ZN(new_n11064_));
  NAND3_X1   g10872(.A1(\asqrt[18] ), .A2(new_n10622_), .A3(new_n10604_), .ZN(new_n11065_));
  XOR2_X1    g10873(.A1(new_n11065_), .A2(new_n10559_), .Z(new_n11066_));
  INV_X1     g10874(.I(new_n11066_), .ZN(new_n11067_));
  OAI21_X1   g10875(.A1(new_n10617_), .A2(new_n10618_), .B(new_n10621_), .ZN(new_n11068_));
  NOR2_X1    g10876(.A1(new_n10953_), .A2(new_n11068_), .ZN(new_n11069_));
  XOR2_X1    g10877(.A1(new_n11069_), .A2(new_n10562_), .Z(new_n11070_));
  NAND3_X1   g10878(.A1(\asqrt[18] ), .A2(new_n10582_), .A3(new_n10600_), .ZN(new_n11071_));
  XOR2_X1    g10879(.A1(new_n11071_), .A2(new_n10616_), .Z(new_n11072_));
  NOR2_X1    g10880(.A1(new_n10579_), .A2(\asqrt[21] ), .ZN(new_n11073_));
  NOR3_X1    g10881(.A1(new_n10953_), .A2(new_n11073_), .A3(new_n10599_), .ZN(new_n11074_));
  XOR2_X1    g10882(.A1(new_n11074_), .A2(new_n10570_), .Z(new_n11075_));
  INV_X1     g10883(.I(new_n11075_), .ZN(new_n11076_));
  NAND3_X1   g10884(.A1(\asqrt[18] ), .A2(new_n10571_), .A3(new_n10572_), .ZN(new_n11077_));
  NOR4_X1    g10885(.A1(new_n10951_), .A2(new_n10478_), .A3(new_n10768_), .A4(new_n10952_), .ZN(new_n11078_));
  INV_X1     g10886(.I(new_n11078_), .ZN(new_n11079_));
  AOI21_X1   g10887(.A1(new_n11077_), .A2(new_n11079_), .B(\a[38] ), .ZN(new_n11080_));
  NOR3_X1    g10888(.A1(new_n10953_), .A2(\a[36] ), .A3(\a[37] ), .ZN(new_n11081_));
  NOR3_X1    g10889(.A1(new_n11081_), .A2(new_n10170_), .A3(new_n11078_), .ZN(new_n11082_));
  NOR2_X1    g10890(.A1(new_n11082_), .A2(new_n11080_), .ZN(new_n11083_));
  INV_X1     g10891(.I(\a[34] ), .ZN(new_n11084_));
  INV_X1     g10892(.I(\a[35] ), .ZN(new_n11085_));
  NAND3_X1   g10893(.A1(new_n11084_), .A2(new_n11085_), .A3(new_n10571_), .ZN(new_n11086_));
  OAI21_X1   g10894(.A1(new_n10953_), .A2(new_n10571_), .B(new_n11086_), .ZN(new_n11087_));
  NAND2_X1   g10895(.A1(new_n11087_), .A2(\asqrt[19] ), .ZN(new_n11088_));
  OAI21_X1   g10896(.A1(new_n10953_), .A2(\a[36] ), .B(\a[37] ), .ZN(new_n11089_));
  NAND2_X1   g10897(.A1(new_n11089_), .A2(new_n11077_), .ZN(new_n11090_));
  NOR2_X1    g10898(.A1(new_n11087_), .A2(\asqrt[19] ), .ZN(new_n11091_));
  OAI21_X1   g10899(.A1(new_n11090_), .A2(new_n11091_), .B(new_n11088_), .ZN(new_n11092_));
  OAI21_X1   g10900(.A1(new_n11092_), .A2(\asqrt[20] ), .B(new_n11083_), .ZN(new_n11093_));
  NAND2_X1   g10901(.A1(new_n11092_), .A2(\asqrt[20] ), .ZN(new_n11094_));
  NAND3_X1   g10902(.A1(new_n11093_), .A2(new_n9590_), .A3(new_n11094_), .ZN(new_n11095_));
  NOR3_X1    g10903(.A1(new_n10953_), .A2(new_n10593_), .A3(new_n10578_), .ZN(new_n11096_));
  XOR2_X1    g10904(.A1(new_n11096_), .A2(new_n10595_), .Z(new_n11097_));
  AOI21_X1   g10905(.A1(new_n11093_), .A2(new_n11094_), .B(new_n9590_), .ZN(new_n11098_));
  AOI21_X1   g10906(.A1(new_n11095_), .A2(new_n11097_), .B(new_n11098_), .ZN(new_n11099_));
  AOI21_X1   g10907(.A1(new_n11099_), .A2(new_n9177_), .B(new_n11076_), .ZN(new_n11100_));
  OAI21_X1   g10908(.A1(new_n11099_), .A2(new_n9177_), .B(new_n8742_), .ZN(new_n11101_));
  OAI21_X1   g10909(.A1(new_n11100_), .A2(new_n11101_), .B(new_n11072_), .ZN(new_n11102_));
  NOR2_X1    g10910(.A1(new_n11099_), .A2(new_n9177_), .ZN(new_n11103_));
  OAI21_X1   g10911(.A1(new_n11100_), .A2(new_n11103_), .B(\asqrt[23] ), .ZN(new_n11104_));
  NAND3_X1   g10912(.A1(new_n11102_), .A2(new_n11104_), .A3(new_n8349_), .ZN(new_n11105_));
  NAND2_X1   g10913(.A1(new_n11105_), .A2(new_n11070_), .ZN(new_n11106_));
  NAND2_X1   g10914(.A1(new_n11102_), .A2(new_n11104_), .ZN(new_n11107_));
  AOI21_X1   g10915(.A1(new_n11107_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n11108_));
  AOI21_X1   g10916(.A1(new_n11108_), .A2(new_n11106_), .B(new_n11067_), .ZN(new_n11109_));
  INV_X1     g10917(.I(new_n11072_), .ZN(new_n11110_));
  OAI21_X1   g10918(.A1(new_n11081_), .A2(new_n11078_), .B(new_n10170_), .ZN(new_n11111_));
  NAND3_X1   g10919(.A1(new_n11077_), .A2(new_n11079_), .A3(\a[38] ), .ZN(new_n11112_));
  NAND2_X1   g10920(.A1(new_n11111_), .A2(new_n11112_), .ZN(new_n11113_));
  NAND2_X1   g10921(.A1(\asqrt[18] ), .A2(\a[36] ), .ZN(new_n11114_));
  AOI21_X1   g10922(.A1(new_n11114_), .A2(new_n11086_), .B(new_n10478_), .ZN(new_n11115_));
  AOI21_X1   g10923(.A1(\asqrt[18] ), .A2(new_n10571_), .B(new_n10572_), .ZN(new_n11116_));
  NOR2_X1    g10924(.A1(new_n11081_), .A2(new_n11116_), .ZN(new_n11117_));
  NAND3_X1   g10925(.A1(new_n11114_), .A2(new_n10478_), .A3(new_n11086_), .ZN(new_n11118_));
  AOI21_X1   g10926(.A1(new_n11117_), .A2(new_n11118_), .B(new_n11115_), .ZN(new_n11119_));
  AOI21_X1   g10927(.A1(new_n11119_), .A2(new_n10045_), .B(new_n11113_), .ZN(new_n11120_));
  NOR2_X1    g10928(.A1(new_n11119_), .A2(new_n10045_), .ZN(new_n11121_));
  NOR3_X1    g10929(.A1(new_n11120_), .A2(\asqrt[21] ), .A3(new_n11121_), .ZN(new_n11122_));
  INV_X1     g10930(.I(new_n11097_), .ZN(new_n11123_));
  OAI21_X1   g10931(.A1(new_n11120_), .A2(new_n11121_), .B(\asqrt[21] ), .ZN(new_n11124_));
  OAI21_X1   g10932(.A1(new_n11122_), .A2(new_n11123_), .B(new_n11124_), .ZN(new_n11125_));
  OAI21_X1   g10933(.A1(new_n11125_), .A2(\asqrt[22] ), .B(new_n11075_), .ZN(new_n11126_));
  AOI21_X1   g10934(.A1(new_n11125_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n11127_));
  AOI21_X1   g10935(.A1(new_n11127_), .A2(new_n11126_), .B(new_n11110_), .ZN(new_n11128_));
  NAND2_X1   g10936(.A1(new_n11125_), .A2(\asqrt[22] ), .ZN(new_n11129_));
  AOI21_X1   g10937(.A1(new_n11126_), .A2(new_n11129_), .B(new_n8742_), .ZN(new_n11130_));
  OAI21_X1   g10938(.A1(new_n11128_), .A2(new_n11130_), .B(\asqrt[24] ), .ZN(new_n11131_));
  AOI21_X1   g10939(.A1(new_n11106_), .A2(new_n11131_), .B(new_n7934_), .ZN(new_n11132_));
  NOR2_X1    g10940(.A1(new_n11109_), .A2(new_n11132_), .ZN(new_n11133_));
  AOI21_X1   g10941(.A1(new_n11133_), .A2(new_n7561_), .B(new_n11064_), .ZN(new_n11134_));
  OAI21_X1   g10942(.A1(new_n11109_), .A2(new_n11132_), .B(\asqrt[26] ), .ZN(new_n11135_));
  NAND2_X1   g10943(.A1(new_n11135_), .A2(new_n7166_), .ZN(new_n11136_));
  OAI21_X1   g10944(.A1(new_n11134_), .A2(new_n11136_), .B(new_n11060_), .ZN(new_n11137_));
  INV_X1     g10945(.I(new_n11135_), .ZN(new_n11138_));
  OAI21_X1   g10946(.A1(new_n11134_), .A2(new_n11138_), .B(\asqrt[27] ), .ZN(new_n11139_));
  NAND3_X1   g10947(.A1(new_n11137_), .A2(new_n11139_), .A3(new_n6813_), .ZN(new_n11140_));
  NAND2_X1   g10948(.A1(new_n11140_), .A2(new_n11058_), .ZN(new_n11141_));
  NAND2_X1   g10949(.A1(new_n11137_), .A2(new_n11139_), .ZN(new_n11142_));
  AOI21_X1   g10950(.A1(new_n11142_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n11143_));
  AOI21_X1   g10951(.A1(new_n11143_), .A2(new_n11141_), .B(new_n11055_), .ZN(new_n11144_));
  INV_X1     g10952(.I(new_n11060_), .ZN(new_n11145_));
  INV_X1     g10953(.I(new_n11070_), .ZN(new_n11146_));
  NOR2_X1    g10954(.A1(new_n11128_), .A2(new_n11130_), .ZN(new_n11147_));
  AOI21_X1   g10955(.A1(new_n11147_), .A2(new_n8349_), .B(new_n11146_), .ZN(new_n11148_));
  NAND2_X1   g10956(.A1(new_n11131_), .A2(new_n7934_), .ZN(new_n11149_));
  OAI21_X1   g10957(.A1(new_n11148_), .A2(new_n11149_), .B(new_n11066_), .ZN(new_n11150_));
  INV_X1     g10958(.I(new_n11131_), .ZN(new_n11151_));
  OAI21_X1   g10959(.A1(new_n11148_), .A2(new_n11151_), .B(\asqrt[25] ), .ZN(new_n11152_));
  NAND3_X1   g10960(.A1(new_n11150_), .A2(new_n11152_), .A3(new_n7561_), .ZN(new_n11153_));
  NAND2_X1   g10961(.A1(new_n11153_), .A2(new_n11063_), .ZN(new_n11154_));
  NAND2_X1   g10962(.A1(new_n11150_), .A2(new_n11152_), .ZN(new_n11155_));
  AOI21_X1   g10963(.A1(new_n11155_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n11156_));
  AOI21_X1   g10964(.A1(new_n11156_), .A2(new_n11154_), .B(new_n11145_), .ZN(new_n11157_));
  AOI21_X1   g10965(.A1(new_n11154_), .A2(new_n11135_), .B(new_n7166_), .ZN(new_n11158_));
  OAI21_X1   g10966(.A1(new_n11157_), .A2(new_n11158_), .B(\asqrt[28] ), .ZN(new_n11159_));
  AOI21_X1   g10967(.A1(new_n11141_), .A2(new_n11159_), .B(new_n6454_), .ZN(new_n11160_));
  NOR2_X1    g10968(.A1(new_n11144_), .A2(new_n11160_), .ZN(new_n11161_));
  AOI21_X1   g10969(.A1(new_n11161_), .A2(new_n6106_), .B(new_n11052_), .ZN(new_n11162_));
  OAI21_X1   g10970(.A1(new_n11144_), .A2(new_n11160_), .B(\asqrt[30] ), .ZN(new_n11163_));
  NAND2_X1   g10971(.A1(new_n11163_), .A2(new_n5750_), .ZN(new_n11164_));
  OAI21_X1   g10972(.A1(new_n11162_), .A2(new_n11164_), .B(new_n11048_), .ZN(new_n11165_));
  INV_X1     g10973(.I(new_n11163_), .ZN(new_n11166_));
  OAI21_X1   g10974(.A1(new_n11162_), .A2(new_n11166_), .B(\asqrt[31] ), .ZN(new_n11167_));
  NAND3_X1   g10975(.A1(new_n11165_), .A2(new_n11167_), .A3(new_n5435_), .ZN(new_n11168_));
  NAND2_X1   g10976(.A1(new_n11168_), .A2(new_n11046_), .ZN(new_n11169_));
  NAND2_X1   g10977(.A1(new_n11165_), .A2(new_n11167_), .ZN(new_n11170_));
  AOI21_X1   g10978(.A1(new_n11170_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n11171_));
  AOI21_X1   g10979(.A1(new_n11171_), .A2(new_n11169_), .B(new_n11043_), .ZN(new_n11172_));
  INV_X1     g10980(.I(new_n11048_), .ZN(new_n11173_));
  INV_X1     g10981(.I(new_n11058_), .ZN(new_n11174_));
  NOR2_X1    g10982(.A1(new_n11157_), .A2(new_n11158_), .ZN(new_n11175_));
  AOI21_X1   g10983(.A1(new_n11175_), .A2(new_n6813_), .B(new_n11174_), .ZN(new_n11176_));
  NAND2_X1   g10984(.A1(new_n11159_), .A2(new_n6454_), .ZN(new_n11177_));
  OAI21_X1   g10985(.A1(new_n11176_), .A2(new_n11177_), .B(new_n11054_), .ZN(new_n11178_));
  INV_X1     g10986(.I(new_n11159_), .ZN(new_n11179_));
  OAI21_X1   g10987(.A1(new_n11176_), .A2(new_n11179_), .B(\asqrt[29] ), .ZN(new_n11180_));
  NAND3_X1   g10988(.A1(new_n11178_), .A2(new_n11180_), .A3(new_n6106_), .ZN(new_n11181_));
  NAND2_X1   g10989(.A1(new_n11181_), .A2(new_n11051_), .ZN(new_n11182_));
  NAND2_X1   g10990(.A1(new_n11178_), .A2(new_n11180_), .ZN(new_n11183_));
  AOI21_X1   g10991(.A1(new_n11183_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n11184_));
  AOI21_X1   g10992(.A1(new_n11184_), .A2(new_n11182_), .B(new_n11173_), .ZN(new_n11185_));
  AOI21_X1   g10993(.A1(new_n11182_), .A2(new_n11163_), .B(new_n5750_), .ZN(new_n11186_));
  OAI21_X1   g10994(.A1(new_n11185_), .A2(new_n11186_), .B(\asqrt[32] ), .ZN(new_n11187_));
  AOI21_X1   g10995(.A1(new_n11169_), .A2(new_n11187_), .B(new_n5110_), .ZN(new_n11188_));
  NOR2_X1    g10996(.A1(new_n11172_), .A2(new_n11188_), .ZN(new_n11189_));
  AOI21_X1   g10997(.A1(new_n11189_), .A2(new_n4810_), .B(new_n11040_), .ZN(new_n11190_));
  OAI21_X1   g10998(.A1(new_n11172_), .A2(new_n11188_), .B(\asqrt[34] ), .ZN(new_n11191_));
  NAND2_X1   g10999(.A1(new_n11191_), .A2(new_n4510_), .ZN(new_n11192_));
  OAI21_X1   g11000(.A1(new_n11190_), .A2(new_n11192_), .B(new_n11036_), .ZN(new_n11193_));
  INV_X1     g11001(.I(new_n11191_), .ZN(new_n11194_));
  OAI21_X1   g11002(.A1(new_n11190_), .A2(new_n11194_), .B(\asqrt[35] ), .ZN(new_n11195_));
  NAND3_X1   g11003(.A1(new_n11193_), .A2(new_n11195_), .A3(new_n4224_), .ZN(new_n11196_));
  NAND2_X1   g11004(.A1(new_n11196_), .A2(new_n11034_), .ZN(new_n11197_));
  NAND2_X1   g11005(.A1(new_n11193_), .A2(new_n11195_), .ZN(new_n11198_));
  AOI21_X1   g11006(.A1(new_n11198_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n11199_));
  AOI21_X1   g11007(.A1(new_n11199_), .A2(new_n11197_), .B(new_n11031_), .ZN(new_n11200_));
  INV_X1     g11008(.I(new_n11036_), .ZN(new_n11201_));
  INV_X1     g11009(.I(new_n11046_), .ZN(new_n11202_));
  NOR2_X1    g11010(.A1(new_n11185_), .A2(new_n11186_), .ZN(new_n11203_));
  AOI21_X1   g11011(.A1(new_n11203_), .A2(new_n5435_), .B(new_n11202_), .ZN(new_n11204_));
  NAND2_X1   g11012(.A1(new_n11187_), .A2(new_n5110_), .ZN(new_n11205_));
  OAI21_X1   g11013(.A1(new_n11204_), .A2(new_n11205_), .B(new_n11042_), .ZN(new_n11206_));
  INV_X1     g11014(.I(new_n11187_), .ZN(new_n11207_));
  OAI21_X1   g11015(.A1(new_n11204_), .A2(new_n11207_), .B(\asqrt[33] ), .ZN(new_n11208_));
  NAND3_X1   g11016(.A1(new_n11206_), .A2(new_n11208_), .A3(new_n4810_), .ZN(new_n11209_));
  NAND2_X1   g11017(.A1(new_n11209_), .A2(new_n11039_), .ZN(new_n11210_));
  NAND2_X1   g11018(.A1(new_n11206_), .A2(new_n11208_), .ZN(new_n11211_));
  AOI21_X1   g11019(.A1(new_n11211_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n11212_));
  AOI21_X1   g11020(.A1(new_n11212_), .A2(new_n11210_), .B(new_n11201_), .ZN(new_n11213_));
  AOI21_X1   g11021(.A1(new_n11210_), .A2(new_n11191_), .B(new_n4510_), .ZN(new_n11214_));
  OAI21_X1   g11022(.A1(new_n11213_), .A2(new_n11214_), .B(\asqrt[36] ), .ZN(new_n11215_));
  AOI21_X1   g11023(.A1(new_n11197_), .A2(new_n11215_), .B(new_n3928_), .ZN(new_n11216_));
  NOR2_X1    g11024(.A1(new_n11200_), .A2(new_n11216_), .ZN(new_n11217_));
  AOI21_X1   g11025(.A1(new_n11217_), .A2(new_n3675_), .B(new_n11028_), .ZN(new_n11218_));
  OAI21_X1   g11026(.A1(new_n11200_), .A2(new_n11216_), .B(\asqrt[38] ), .ZN(new_n11219_));
  NAND2_X1   g11027(.A1(new_n11219_), .A2(new_n3400_), .ZN(new_n11220_));
  OAI21_X1   g11028(.A1(new_n11218_), .A2(new_n11220_), .B(new_n11024_), .ZN(new_n11221_));
  INV_X1     g11029(.I(new_n11219_), .ZN(new_n11222_));
  OAI21_X1   g11030(.A1(new_n11218_), .A2(new_n11222_), .B(\asqrt[39] ), .ZN(new_n11223_));
  NAND3_X1   g11031(.A1(new_n11221_), .A2(new_n11223_), .A3(new_n3167_), .ZN(new_n11224_));
  NAND2_X1   g11032(.A1(new_n11224_), .A2(new_n11022_), .ZN(new_n11225_));
  NAND2_X1   g11033(.A1(new_n11221_), .A2(new_n11223_), .ZN(new_n11226_));
  AOI21_X1   g11034(.A1(new_n11226_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n11227_));
  AOI21_X1   g11035(.A1(new_n11227_), .A2(new_n11225_), .B(new_n11019_), .ZN(new_n11228_));
  INV_X1     g11036(.I(new_n11024_), .ZN(new_n11229_));
  INV_X1     g11037(.I(new_n11034_), .ZN(new_n11230_));
  NOR2_X1    g11038(.A1(new_n11213_), .A2(new_n11214_), .ZN(new_n11231_));
  AOI21_X1   g11039(.A1(new_n11231_), .A2(new_n4224_), .B(new_n11230_), .ZN(new_n11232_));
  NAND2_X1   g11040(.A1(new_n11215_), .A2(new_n3928_), .ZN(new_n11233_));
  OAI21_X1   g11041(.A1(new_n11232_), .A2(new_n11233_), .B(new_n11030_), .ZN(new_n11234_));
  INV_X1     g11042(.I(new_n11215_), .ZN(new_n11235_));
  OAI21_X1   g11043(.A1(new_n11232_), .A2(new_n11235_), .B(\asqrt[37] ), .ZN(new_n11236_));
  NAND3_X1   g11044(.A1(new_n11234_), .A2(new_n11236_), .A3(new_n3675_), .ZN(new_n11237_));
  NAND2_X1   g11045(.A1(new_n11237_), .A2(new_n11027_), .ZN(new_n11238_));
  NAND2_X1   g11046(.A1(new_n11234_), .A2(new_n11236_), .ZN(new_n11239_));
  AOI21_X1   g11047(.A1(new_n11239_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n11240_));
  AOI21_X1   g11048(.A1(new_n11240_), .A2(new_n11238_), .B(new_n11229_), .ZN(new_n11241_));
  AOI21_X1   g11049(.A1(new_n11238_), .A2(new_n11219_), .B(new_n3400_), .ZN(new_n11242_));
  OAI21_X1   g11050(.A1(new_n11241_), .A2(new_n11242_), .B(\asqrt[40] ), .ZN(new_n11243_));
  AOI21_X1   g11051(.A1(new_n11225_), .A2(new_n11243_), .B(new_n2912_), .ZN(new_n11244_));
  NOR2_X1    g11052(.A1(new_n11228_), .A2(new_n11244_), .ZN(new_n11245_));
  AOI21_X1   g11053(.A1(new_n11245_), .A2(new_n2699_), .B(new_n11016_), .ZN(new_n11246_));
  OAI21_X1   g11054(.A1(new_n11228_), .A2(new_n11244_), .B(\asqrt[42] ), .ZN(new_n11247_));
  NAND2_X1   g11055(.A1(new_n11247_), .A2(new_n2464_), .ZN(new_n11248_));
  OAI21_X1   g11056(.A1(new_n11246_), .A2(new_n11248_), .B(new_n11012_), .ZN(new_n11249_));
  INV_X1     g11057(.I(new_n11247_), .ZN(new_n11250_));
  OAI21_X1   g11058(.A1(new_n11246_), .A2(new_n11250_), .B(\asqrt[43] ), .ZN(new_n11251_));
  NAND3_X1   g11059(.A1(new_n11249_), .A2(new_n11251_), .A3(new_n2271_), .ZN(new_n11252_));
  NAND2_X1   g11060(.A1(new_n11252_), .A2(new_n11010_), .ZN(new_n11253_));
  NAND2_X1   g11061(.A1(new_n11249_), .A2(new_n11251_), .ZN(new_n11254_));
  AOI21_X1   g11062(.A1(new_n11254_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n11255_));
  AOI21_X1   g11063(.A1(new_n11255_), .A2(new_n11253_), .B(new_n11007_), .ZN(new_n11256_));
  INV_X1     g11064(.I(new_n11012_), .ZN(new_n11257_));
  INV_X1     g11065(.I(new_n11022_), .ZN(new_n11258_));
  NOR2_X1    g11066(.A1(new_n11241_), .A2(new_n11242_), .ZN(new_n11259_));
  AOI21_X1   g11067(.A1(new_n11259_), .A2(new_n3167_), .B(new_n11258_), .ZN(new_n11260_));
  NAND2_X1   g11068(.A1(new_n11243_), .A2(new_n2912_), .ZN(new_n11261_));
  OAI21_X1   g11069(.A1(new_n11260_), .A2(new_n11261_), .B(new_n11018_), .ZN(new_n11262_));
  INV_X1     g11070(.I(new_n11243_), .ZN(new_n11263_));
  OAI21_X1   g11071(.A1(new_n11260_), .A2(new_n11263_), .B(\asqrt[41] ), .ZN(new_n11264_));
  NAND3_X1   g11072(.A1(new_n11262_), .A2(new_n11264_), .A3(new_n2699_), .ZN(new_n11265_));
  NAND2_X1   g11073(.A1(new_n11265_), .A2(new_n11015_), .ZN(new_n11266_));
  NAND2_X1   g11074(.A1(new_n11262_), .A2(new_n11264_), .ZN(new_n11267_));
  AOI21_X1   g11075(.A1(new_n11267_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n11268_));
  AOI21_X1   g11076(.A1(new_n11268_), .A2(new_n11266_), .B(new_n11257_), .ZN(new_n11269_));
  AOI21_X1   g11077(.A1(new_n11266_), .A2(new_n11247_), .B(new_n2464_), .ZN(new_n11270_));
  OAI21_X1   g11078(.A1(new_n11269_), .A2(new_n11270_), .B(\asqrt[44] ), .ZN(new_n11271_));
  AOI21_X1   g11079(.A1(new_n11253_), .A2(new_n11271_), .B(new_n2072_), .ZN(new_n11272_));
  NOR2_X1    g11080(.A1(new_n11256_), .A2(new_n11272_), .ZN(new_n11273_));
  AOI21_X1   g11081(.A1(new_n11273_), .A2(new_n1884_), .B(new_n11004_), .ZN(new_n11274_));
  OAI21_X1   g11082(.A1(new_n11256_), .A2(new_n11272_), .B(\asqrt[46] ), .ZN(new_n11275_));
  NAND2_X1   g11083(.A1(new_n11275_), .A2(new_n1688_), .ZN(new_n11276_));
  OAI21_X1   g11084(.A1(new_n11274_), .A2(new_n11276_), .B(new_n10936_), .ZN(new_n11277_));
  INV_X1     g11085(.I(new_n11275_), .ZN(new_n11278_));
  OAI21_X1   g11086(.A1(new_n11274_), .A2(new_n11278_), .B(\asqrt[47] ), .ZN(new_n11279_));
  NAND3_X1   g11087(.A1(new_n11277_), .A2(new_n11279_), .A3(new_n1533_), .ZN(new_n11280_));
  NAND2_X1   g11088(.A1(new_n11280_), .A2(new_n11000_), .ZN(new_n11281_));
  NAND2_X1   g11089(.A1(new_n11277_), .A2(new_n11279_), .ZN(new_n11282_));
  AOI21_X1   g11090(.A1(new_n11282_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n11283_));
  AOI21_X1   g11091(.A1(new_n11283_), .A2(new_n11281_), .B(new_n10997_), .ZN(new_n11284_));
  INV_X1     g11092(.I(new_n10936_), .ZN(new_n11285_));
  INV_X1     g11093(.I(new_n11010_), .ZN(new_n11286_));
  NOR2_X1    g11094(.A1(new_n11269_), .A2(new_n11270_), .ZN(new_n11287_));
  AOI21_X1   g11095(.A1(new_n11287_), .A2(new_n2271_), .B(new_n11286_), .ZN(new_n11288_));
  NAND2_X1   g11096(.A1(new_n11271_), .A2(new_n2072_), .ZN(new_n11289_));
  OAI21_X1   g11097(.A1(new_n11288_), .A2(new_n11289_), .B(new_n11006_), .ZN(new_n11290_));
  INV_X1     g11098(.I(new_n11271_), .ZN(new_n11291_));
  OAI21_X1   g11099(.A1(new_n11288_), .A2(new_n11291_), .B(\asqrt[45] ), .ZN(new_n11292_));
  NAND3_X1   g11100(.A1(new_n11290_), .A2(new_n11292_), .A3(new_n1884_), .ZN(new_n11293_));
  NAND2_X1   g11101(.A1(new_n11293_), .A2(new_n11003_), .ZN(new_n11294_));
  NAND2_X1   g11102(.A1(new_n11290_), .A2(new_n11292_), .ZN(new_n11295_));
  AOI21_X1   g11103(.A1(new_n11295_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n11296_));
  AOI21_X1   g11104(.A1(new_n11296_), .A2(new_n11294_), .B(new_n11285_), .ZN(new_n11297_));
  AOI21_X1   g11105(.A1(new_n11294_), .A2(new_n11275_), .B(new_n1688_), .ZN(new_n11298_));
  OAI21_X1   g11106(.A1(new_n11297_), .A2(new_n11298_), .B(\asqrt[48] ), .ZN(new_n11299_));
  AOI21_X1   g11107(.A1(new_n11281_), .A2(new_n11299_), .B(new_n1368_), .ZN(new_n11300_));
  NOR2_X1    g11108(.A1(new_n11284_), .A2(new_n11300_), .ZN(new_n11301_));
  AOI21_X1   g11109(.A1(new_n11301_), .A2(new_n1228_), .B(new_n10994_), .ZN(new_n11302_));
  OAI21_X1   g11110(.A1(new_n11284_), .A2(new_n11300_), .B(\asqrt[50] ), .ZN(new_n11303_));
  NAND2_X1   g11111(.A1(new_n11303_), .A2(new_n1088_), .ZN(new_n11304_));
  OAI21_X1   g11112(.A1(new_n11302_), .A2(new_n11304_), .B(new_n10990_), .ZN(new_n11305_));
  INV_X1     g11113(.I(new_n11303_), .ZN(new_n11306_));
  OAI21_X1   g11114(.A1(new_n11302_), .A2(new_n11306_), .B(\asqrt[51] ), .ZN(new_n11307_));
  NAND3_X1   g11115(.A1(new_n11305_), .A2(new_n11307_), .A3(new_n962_), .ZN(new_n11308_));
  NAND2_X1   g11116(.A1(new_n11308_), .A2(new_n10988_), .ZN(new_n11309_));
  NAND2_X1   g11117(.A1(new_n11305_), .A2(new_n11307_), .ZN(new_n11310_));
  AOI21_X1   g11118(.A1(new_n11310_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n11311_));
  AOI21_X1   g11119(.A1(new_n11311_), .A2(new_n11309_), .B(new_n10985_), .ZN(new_n11312_));
  INV_X1     g11120(.I(new_n10990_), .ZN(new_n11313_));
  INV_X1     g11121(.I(new_n11000_), .ZN(new_n11314_));
  NOR2_X1    g11122(.A1(new_n11297_), .A2(new_n11298_), .ZN(new_n11315_));
  AOI21_X1   g11123(.A1(new_n11315_), .A2(new_n1533_), .B(new_n11314_), .ZN(new_n11316_));
  NAND2_X1   g11124(.A1(new_n11299_), .A2(new_n1368_), .ZN(new_n11317_));
  OAI21_X1   g11125(.A1(new_n11316_), .A2(new_n11317_), .B(new_n10996_), .ZN(new_n11318_));
  INV_X1     g11126(.I(new_n11299_), .ZN(new_n11319_));
  OAI21_X1   g11127(.A1(new_n11316_), .A2(new_n11319_), .B(\asqrt[49] ), .ZN(new_n11320_));
  NAND3_X1   g11128(.A1(new_n11318_), .A2(new_n11320_), .A3(new_n1228_), .ZN(new_n11321_));
  NAND2_X1   g11129(.A1(new_n11321_), .A2(new_n10993_), .ZN(new_n11322_));
  NAND2_X1   g11130(.A1(new_n11318_), .A2(new_n11320_), .ZN(new_n11323_));
  AOI21_X1   g11131(.A1(new_n11323_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n11324_));
  AOI21_X1   g11132(.A1(new_n11324_), .A2(new_n11322_), .B(new_n11313_), .ZN(new_n11325_));
  AOI21_X1   g11133(.A1(new_n11322_), .A2(new_n11303_), .B(new_n1088_), .ZN(new_n11326_));
  OAI21_X1   g11134(.A1(new_n11325_), .A2(new_n11326_), .B(\asqrt[52] ), .ZN(new_n11327_));
  AOI21_X1   g11135(.A1(new_n11309_), .A2(new_n11327_), .B(new_n842_), .ZN(new_n11328_));
  NOR2_X1    g11136(.A1(new_n11312_), .A2(new_n11328_), .ZN(new_n11329_));
  AOI21_X1   g11137(.A1(new_n11329_), .A2(new_n720_), .B(new_n10982_), .ZN(new_n11330_));
  OAI21_X1   g11138(.A1(new_n11312_), .A2(new_n11328_), .B(\asqrt[54] ), .ZN(new_n11331_));
  NAND2_X1   g11139(.A1(new_n11331_), .A2(new_n630_), .ZN(new_n11332_));
  OAI21_X1   g11140(.A1(new_n11330_), .A2(new_n11332_), .B(new_n10978_), .ZN(new_n11333_));
  INV_X1     g11141(.I(new_n11331_), .ZN(new_n11334_));
  OAI21_X1   g11142(.A1(new_n11330_), .A2(new_n11334_), .B(\asqrt[55] ), .ZN(new_n11335_));
  NAND3_X1   g11143(.A1(new_n11333_), .A2(new_n11335_), .A3(new_n545_), .ZN(new_n11336_));
  NAND2_X1   g11144(.A1(new_n11336_), .A2(new_n10976_), .ZN(new_n11337_));
  NAND2_X1   g11145(.A1(new_n11333_), .A2(new_n11335_), .ZN(new_n11338_));
  AOI21_X1   g11146(.A1(new_n11338_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n11339_));
  AOI21_X1   g11147(.A1(new_n11339_), .A2(new_n11337_), .B(new_n10973_), .ZN(new_n11340_));
  INV_X1     g11148(.I(new_n10978_), .ZN(new_n11341_));
  INV_X1     g11149(.I(new_n10988_), .ZN(new_n11342_));
  NOR2_X1    g11150(.A1(new_n11325_), .A2(new_n11326_), .ZN(new_n11343_));
  AOI21_X1   g11151(.A1(new_n11343_), .A2(new_n962_), .B(new_n11342_), .ZN(new_n11344_));
  NAND2_X1   g11152(.A1(new_n11327_), .A2(new_n842_), .ZN(new_n11345_));
  OAI21_X1   g11153(.A1(new_n11344_), .A2(new_n11345_), .B(new_n10984_), .ZN(new_n11346_));
  INV_X1     g11154(.I(new_n11327_), .ZN(new_n11347_));
  OAI21_X1   g11155(.A1(new_n11344_), .A2(new_n11347_), .B(\asqrt[53] ), .ZN(new_n11348_));
  NAND3_X1   g11156(.A1(new_n11346_), .A2(new_n11348_), .A3(new_n720_), .ZN(new_n11349_));
  NAND2_X1   g11157(.A1(new_n11349_), .A2(new_n10981_), .ZN(new_n11350_));
  NAND2_X1   g11158(.A1(new_n11346_), .A2(new_n11348_), .ZN(new_n11351_));
  AOI21_X1   g11159(.A1(new_n11351_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n11352_));
  AOI21_X1   g11160(.A1(new_n11352_), .A2(new_n11350_), .B(new_n11341_), .ZN(new_n11353_));
  AOI21_X1   g11161(.A1(new_n11350_), .A2(new_n11331_), .B(new_n630_), .ZN(new_n11354_));
  OAI21_X1   g11162(.A1(new_n11353_), .A2(new_n11354_), .B(\asqrt[56] ), .ZN(new_n11355_));
  AOI21_X1   g11163(.A1(new_n11337_), .A2(new_n11355_), .B(new_n450_), .ZN(new_n11356_));
  NOR2_X1    g11164(.A1(new_n11340_), .A2(new_n11356_), .ZN(new_n11357_));
  AOI21_X1   g11165(.A1(new_n11357_), .A2(new_n403_), .B(new_n10970_), .ZN(new_n11358_));
  OAI21_X1   g11166(.A1(new_n11340_), .A2(new_n11356_), .B(\asqrt[58] ), .ZN(new_n11359_));
  NAND2_X1   g11167(.A1(new_n11359_), .A2(new_n339_), .ZN(new_n11360_));
  OAI21_X1   g11168(.A1(new_n11358_), .A2(new_n11360_), .B(new_n10966_), .ZN(new_n11361_));
  INV_X1     g11169(.I(new_n11359_), .ZN(new_n11362_));
  OAI21_X1   g11170(.A1(new_n11358_), .A2(new_n11362_), .B(\asqrt[59] ), .ZN(new_n11363_));
  NAND3_X1   g11171(.A1(new_n11361_), .A2(new_n11363_), .A3(new_n288_), .ZN(new_n11364_));
  NAND2_X1   g11172(.A1(new_n11364_), .A2(new_n10964_), .ZN(new_n11365_));
  INV_X1     g11173(.I(new_n10966_), .ZN(new_n11366_));
  INV_X1     g11174(.I(new_n10976_), .ZN(new_n11367_));
  NOR2_X1    g11175(.A1(new_n11353_), .A2(new_n11354_), .ZN(new_n11368_));
  AOI21_X1   g11176(.A1(new_n11368_), .A2(new_n545_), .B(new_n11367_), .ZN(new_n11369_));
  NAND2_X1   g11177(.A1(new_n11355_), .A2(new_n450_), .ZN(new_n11370_));
  OAI21_X1   g11178(.A1(new_n11369_), .A2(new_n11370_), .B(new_n10972_), .ZN(new_n11371_));
  INV_X1     g11179(.I(new_n11355_), .ZN(new_n11372_));
  OAI21_X1   g11180(.A1(new_n11369_), .A2(new_n11372_), .B(\asqrt[57] ), .ZN(new_n11373_));
  NAND3_X1   g11181(.A1(new_n11371_), .A2(new_n11373_), .A3(new_n403_), .ZN(new_n11374_));
  NAND2_X1   g11182(.A1(new_n11374_), .A2(new_n10969_), .ZN(new_n11375_));
  NAND2_X1   g11183(.A1(new_n11371_), .A2(new_n11373_), .ZN(new_n11376_));
  AOI21_X1   g11184(.A1(new_n11376_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n11377_));
  AOI21_X1   g11185(.A1(new_n11377_), .A2(new_n11375_), .B(new_n11366_), .ZN(new_n11378_));
  AOI21_X1   g11186(.A1(new_n11375_), .A2(new_n11359_), .B(new_n339_), .ZN(new_n11379_));
  OAI21_X1   g11187(.A1(new_n11378_), .A2(new_n11379_), .B(\asqrt[60] ), .ZN(new_n11380_));
  AOI21_X1   g11188(.A1(new_n11365_), .A2(new_n11380_), .B(new_n242_), .ZN(new_n11381_));
  NAND3_X1   g11189(.A1(\asqrt[18] ), .A2(new_n10896_), .A3(new_n10912_), .ZN(new_n11382_));
  XOR2_X1    g11190(.A1(new_n11382_), .A2(new_n10937_), .Z(new_n11383_));
  INV_X1     g11191(.I(new_n11383_), .ZN(new_n11384_));
  NAND2_X1   g11192(.A1(new_n11361_), .A2(new_n11363_), .ZN(new_n11385_));
  AOI21_X1   g11193(.A1(new_n11385_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n11386_));
  AOI21_X1   g11194(.A1(new_n11386_), .A2(new_n11365_), .B(new_n11384_), .ZN(new_n11387_));
  OAI21_X1   g11195(.A1(new_n11387_), .A2(new_n11381_), .B(\asqrt[62] ), .ZN(new_n11388_));
  AOI21_X1   g11196(.A1(new_n10897_), .A2(new_n10918_), .B(new_n10913_), .ZN(new_n11389_));
  NAND2_X1   g11197(.A1(\asqrt[18] ), .A2(new_n11389_), .ZN(new_n11390_));
  XOR2_X1    g11198(.A1(new_n11390_), .A2(new_n10916_), .Z(new_n11391_));
  INV_X1     g11199(.I(new_n10964_), .ZN(new_n11392_));
  NOR2_X1    g11200(.A1(new_n11378_), .A2(new_n11379_), .ZN(new_n11393_));
  AOI21_X1   g11201(.A1(new_n11393_), .A2(new_n288_), .B(new_n11392_), .ZN(new_n11394_));
  INV_X1     g11202(.I(new_n11380_), .ZN(new_n11395_));
  OAI21_X1   g11203(.A1(new_n11394_), .A2(new_n11395_), .B(\asqrt[61] ), .ZN(new_n11396_));
  NAND2_X1   g11204(.A1(new_n11380_), .A2(new_n242_), .ZN(new_n11397_));
  OAI21_X1   g11205(.A1(new_n11394_), .A2(new_n11397_), .B(new_n11383_), .ZN(new_n11398_));
  NAND3_X1   g11206(.A1(new_n11398_), .A2(new_n11396_), .A3(new_n234_), .ZN(new_n11399_));
  NAND2_X1   g11207(.A1(new_n11399_), .A2(new_n11391_), .ZN(new_n11400_));
  AOI21_X1   g11208(.A1(new_n11400_), .A2(new_n11388_), .B(new_n10961_), .ZN(new_n11401_));
  AOI21_X1   g11209(.A1(new_n11401_), .A2(new_n10959_), .B(\asqrt[63] ), .ZN(new_n11402_));
  NAND2_X1   g11210(.A1(new_n11400_), .A2(new_n11388_), .ZN(new_n11403_));
  NOR2_X1    g11211(.A1(new_n11403_), .A2(new_n10959_), .ZN(new_n11404_));
  NOR2_X1    g11212(.A1(\asqrt[18] ), .A2(new_n10948_), .ZN(new_n11405_));
  NOR4_X1    g11213(.A1(new_n11402_), .A2(new_n10956_), .A3(new_n11404_), .A4(new_n11405_), .ZN(new_n11406_));
  OAI21_X1   g11214(.A1(new_n11274_), .A2(new_n11276_), .B(new_n11279_), .ZN(new_n11407_));
  NOR2_X1    g11215(.A1(new_n11406_), .A2(new_n11407_), .ZN(new_n11408_));
  XOR2_X1    g11216(.A1(new_n11408_), .A2(new_n10936_), .Z(new_n11409_));
  INV_X1     g11217(.I(new_n11409_), .ZN(new_n11410_));
  INV_X1     g11218(.I(new_n10956_), .ZN(new_n11411_));
  INV_X1     g11219(.I(new_n11388_), .ZN(new_n11412_));
  NOR2_X1    g11220(.A1(new_n11387_), .A2(new_n11381_), .ZN(new_n11413_));
  INV_X1     g11221(.I(new_n11391_), .ZN(new_n11414_));
  AOI21_X1   g11222(.A1(new_n11413_), .A2(new_n234_), .B(new_n11414_), .ZN(new_n11415_));
  OAI21_X1   g11223(.A1(new_n11415_), .A2(new_n11412_), .B(new_n10960_), .ZN(new_n11416_));
  OAI21_X1   g11224(.A1(new_n11416_), .A2(new_n10958_), .B(new_n193_), .ZN(new_n11417_));
  NOR2_X1    g11225(.A1(new_n11415_), .A2(new_n11412_), .ZN(new_n11418_));
  NAND2_X1   g11226(.A1(new_n11418_), .A2(new_n10958_), .ZN(new_n11419_));
  INV_X1     g11227(.I(new_n11405_), .ZN(new_n11420_));
  NAND4_X1   g11228(.A1(new_n11417_), .A2(new_n11411_), .A3(new_n11419_), .A4(new_n11420_), .ZN(\asqrt[17] ));
  NAND3_X1   g11229(.A1(\asqrt[17] ), .A2(new_n11293_), .A3(new_n11275_), .ZN(new_n11422_));
  XOR2_X1    g11230(.A1(new_n11422_), .A2(new_n11004_), .Z(new_n11423_));
  OAI21_X1   g11231(.A1(new_n11288_), .A2(new_n11289_), .B(new_n11292_), .ZN(new_n11424_));
  NOR2_X1    g11232(.A1(new_n11406_), .A2(new_n11424_), .ZN(new_n11425_));
  XOR2_X1    g11233(.A1(new_n11425_), .A2(new_n11006_), .Z(new_n11426_));
  INV_X1     g11234(.I(new_n11426_), .ZN(new_n11427_));
  NAND3_X1   g11235(.A1(\asqrt[17] ), .A2(new_n11252_), .A3(new_n11271_), .ZN(new_n11428_));
  XOR2_X1    g11236(.A1(new_n11428_), .A2(new_n11286_), .Z(new_n11429_));
  INV_X1     g11237(.I(new_n11429_), .ZN(new_n11430_));
  OAI21_X1   g11238(.A1(new_n11246_), .A2(new_n11248_), .B(new_n11251_), .ZN(new_n11431_));
  NOR2_X1    g11239(.A1(new_n11406_), .A2(new_n11431_), .ZN(new_n11432_));
  XOR2_X1    g11240(.A1(new_n11432_), .A2(new_n11012_), .Z(new_n11433_));
  NAND3_X1   g11241(.A1(\asqrt[17] ), .A2(new_n11265_), .A3(new_n11247_), .ZN(new_n11434_));
  XOR2_X1    g11242(.A1(new_n11434_), .A2(new_n11016_), .Z(new_n11435_));
  OAI21_X1   g11243(.A1(new_n11260_), .A2(new_n11261_), .B(new_n11264_), .ZN(new_n11436_));
  NOR2_X1    g11244(.A1(new_n11406_), .A2(new_n11436_), .ZN(new_n11437_));
  XOR2_X1    g11245(.A1(new_n11437_), .A2(new_n11018_), .Z(new_n11438_));
  INV_X1     g11246(.I(new_n11438_), .ZN(new_n11439_));
  NAND3_X1   g11247(.A1(\asqrt[17] ), .A2(new_n11224_), .A3(new_n11243_), .ZN(new_n11440_));
  XOR2_X1    g11248(.A1(new_n11440_), .A2(new_n11258_), .Z(new_n11441_));
  INV_X1     g11249(.I(new_n11441_), .ZN(new_n11442_));
  OAI21_X1   g11250(.A1(new_n11218_), .A2(new_n11220_), .B(new_n11223_), .ZN(new_n11443_));
  NOR2_X1    g11251(.A1(new_n11406_), .A2(new_n11443_), .ZN(new_n11444_));
  XOR2_X1    g11252(.A1(new_n11444_), .A2(new_n11024_), .Z(new_n11445_));
  NAND3_X1   g11253(.A1(\asqrt[17] ), .A2(new_n11237_), .A3(new_n11219_), .ZN(new_n11446_));
  XOR2_X1    g11254(.A1(new_n11446_), .A2(new_n11028_), .Z(new_n11447_));
  OAI21_X1   g11255(.A1(new_n11232_), .A2(new_n11233_), .B(new_n11236_), .ZN(new_n11448_));
  NOR2_X1    g11256(.A1(new_n11406_), .A2(new_n11448_), .ZN(new_n11449_));
  XOR2_X1    g11257(.A1(new_n11449_), .A2(new_n11030_), .Z(new_n11450_));
  INV_X1     g11258(.I(new_n11450_), .ZN(new_n11451_));
  NAND3_X1   g11259(.A1(\asqrt[17] ), .A2(new_n11196_), .A3(new_n11215_), .ZN(new_n11452_));
  XOR2_X1    g11260(.A1(new_n11452_), .A2(new_n11230_), .Z(new_n11453_));
  INV_X1     g11261(.I(new_n11453_), .ZN(new_n11454_));
  OAI21_X1   g11262(.A1(new_n11190_), .A2(new_n11192_), .B(new_n11195_), .ZN(new_n11455_));
  NOR2_X1    g11263(.A1(new_n11406_), .A2(new_n11455_), .ZN(new_n11456_));
  XOR2_X1    g11264(.A1(new_n11456_), .A2(new_n11036_), .Z(new_n11457_));
  NAND3_X1   g11265(.A1(\asqrt[17] ), .A2(new_n11209_), .A3(new_n11191_), .ZN(new_n11458_));
  XOR2_X1    g11266(.A1(new_n11458_), .A2(new_n11040_), .Z(new_n11459_));
  OAI21_X1   g11267(.A1(new_n11204_), .A2(new_n11205_), .B(new_n11208_), .ZN(new_n11460_));
  NOR2_X1    g11268(.A1(new_n11406_), .A2(new_n11460_), .ZN(new_n11461_));
  XOR2_X1    g11269(.A1(new_n11461_), .A2(new_n11042_), .Z(new_n11462_));
  INV_X1     g11270(.I(new_n11462_), .ZN(new_n11463_));
  NAND3_X1   g11271(.A1(\asqrt[17] ), .A2(new_n11168_), .A3(new_n11187_), .ZN(new_n11464_));
  XOR2_X1    g11272(.A1(new_n11464_), .A2(new_n11202_), .Z(new_n11465_));
  INV_X1     g11273(.I(new_n11465_), .ZN(new_n11466_));
  OAI21_X1   g11274(.A1(new_n11162_), .A2(new_n11164_), .B(new_n11167_), .ZN(new_n11467_));
  NOR2_X1    g11275(.A1(new_n11406_), .A2(new_n11467_), .ZN(new_n11468_));
  XOR2_X1    g11276(.A1(new_n11468_), .A2(new_n11048_), .Z(new_n11469_));
  NAND3_X1   g11277(.A1(\asqrt[17] ), .A2(new_n11181_), .A3(new_n11163_), .ZN(new_n11470_));
  XOR2_X1    g11278(.A1(new_n11470_), .A2(new_n11052_), .Z(new_n11471_));
  OAI21_X1   g11279(.A1(new_n11176_), .A2(new_n11177_), .B(new_n11180_), .ZN(new_n11472_));
  NOR2_X1    g11280(.A1(new_n11406_), .A2(new_n11472_), .ZN(new_n11473_));
  XOR2_X1    g11281(.A1(new_n11473_), .A2(new_n11054_), .Z(new_n11474_));
  INV_X1     g11282(.I(new_n11474_), .ZN(new_n11475_));
  NAND3_X1   g11283(.A1(\asqrt[17] ), .A2(new_n11140_), .A3(new_n11159_), .ZN(new_n11476_));
  XOR2_X1    g11284(.A1(new_n11476_), .A2(new_n11174_), .Z(new_n11477_));
  INV_X1     g11285(.I(new_n11477_), .ZN(new_n11478_));
  OAI21_X1   g11286(.A1(new_n11134_), .A2(new_n11136_), .B(new_n11139_), .ZN(new_n11479_));
  NOR2_X1    g11287(.A1(new_n11406_), .A2(new_n11479_), .ZN(new_n11480_));
  XOR2_X1    g11288(.A1(new_n11480_), .A2(new_n11060_), .Z(new_n11481_));
  NAND3_X1   g11289(.A1(\asqrt[17] ), .A2(new_n11153_), .A3(new_n11135_), .ZN(new_n11482_));
  XOR2_X1    g11290(.A1(new_n11482_), .A2(new_n11064_), .Z(new_n11483_));
  OAI21_X1   g11291(.A1(new_n11148_), .A2(new_n11149_), .B(new_n11152_), .ZN(new_n11484_));
  NOR2_X1    g11292(.A1(new_n11406_), .A2(new_n11484_), .ZN(new_n11485_));
  XOR2_X1    g11293(.A1(new_n11485_), .A2(new_n11066_), .Z(new_n11486_));
  INV_X1     g11294(.I(new_n11486_), .ZN(new_n11487_));
  NAND3_X1   g11295(.A1(\asqrt[17] ), .A2(new_n11105_), .A3(new_n11131_), .ZN(new_n11488_));
  XOR2_X1    g11296(.A1(new_n11488_), .A2(new_n11146_), .Z(new_n11489_));
  INV_X1     g11297(.I(new_n11489_), .ZN(new_n11490_));
  AOI21_X1   g11298(.A1(new_n11126_), .A2(new_n11127_), .B(new_n11130_), .ZN(new_n11491_));
  NAND2_X1   g11299(.A1(\asqrt[17] ), .A2(new_n11491_), .ZN(new_n11492_));
  XOR2_X1    g11300(.A1(new_n11492_), .A2(new_n11110_), .Z(new_n11493_));
  NOR2_X1    g11301(.A1(new_n11125_), .A2(\asqrt[22] ), .ZN(new_n11494_));
  NOR3_X1    g11302(.A1(new_n11406_), .A2(new_n11494_), .A3(new_n11103_), .ZN(new_n11495_));
  XOR2_X1    g11303(.A1(new_n11495_), .A2(new_n11075_), .Z(new_n11496_));
  NOR3_X1    g11304(.A1(new_n11406_), .A2(new_n11122_), .A3(new_n11098_), .ZN(new_n11497_));
  XOR2_X1    g11305(.A1(new_n11497_), .A2(new_n11097_), .Z(new_n11498_));
  INV_X1     g11306(.I(new_n11498_), .ZN(new_n11499_));
  NOR2_X1    g11307(.A1(new_n11092_), .A2(\asqrt[20] ), .ZN(new_n11500_));
  NOR3_X1    g11308(.A1(new_n11406_), .A2(new_n11500_), .A3(new_n11121_), .ZN(new_n11501_));
  XOR2_X1    g11309(.A1(new_n11501_), .A2(new_n11083_), .Z(new_n11502_));
  INV_X1     g11310(.I(new_n11502_), .ZN(new_n11503_));
  NAND3_X1   g11311(.A1(\asqrt[17] ), .A2(new_n11084_), .A3(new_n11085_), .ZN(new_n11504_));
  NOR4_X1    g11312(.A1(new_n11402_), .A2(new_n10953_), .A3(new_n10956_), .A4(new_n11404_), .ZN(new_n11505_));
  INV_X1     g11313(.I(new_n11505_), .ZN(new_n11506_));
  AOI21_X1   g11314(.A1(new_n11504_), .A2(new_n11506_), .B(\a[36] ), .ZN(new_n11507_));
  NOR3_X1    g11315(.A1(new_n11406_), .A2(\a[34] ), .A3(\a[35] ), .ZN(new_n11508_));
  NOR3_X1    g11316(.A1(new_n11508_), .A2(new_n10571_), .A3(new_n11505_), .ZN(new_n11509_));
  NOR2_X1    g11317(.A1(new_n11509_), .A2(new_n11507_), .ZN(new_n11510_));
  INV_X1     g11318(.I(\a[32] ), .ZN(new_n11511_));
  INV_X1     g11319(.I(\a[33] ), .ZN(new_n11512_));
  NAND3_X1   g11320(.A1(new_n11511_), .A2(new_n11512_), .A3(new_n11084_), .ZN(new_n11513_));
  OAI21_X1   g11321(.A1(new_n11406_), .A2(new_n11084_), .B(new_n11513_), .ZN(new_n11514_));
  NAND2_X1   g11322(.A1(new_n11514_), .A2(\asqrt[18] ), .ZN(new_n11515_));
  OAI21_X1   g11323(.A1(new_n11406_), .A2(\a[34] ), .B(\a[35] ), .ZN(new_n11516_));
  NAND2_X1   g11324(.A1(new_n11516_), .A2(new_n11504_), .ZN(new_n11517_));
  NOR2_X1    g11325(.A1(new_n11514_), .A2(\asqrt[18] ), .ZN(new_n11518_));
  OAI21_X1   g11326(.A1(new_n11517_), .A2(new_n11518_), .B(new_n11515_), .ZN(new_n11519_));
  OAI21_X1   g11327(.A1(\asqrt[19] ), .A2(new_n11519_), .B(new_n11510_), .ZN(new_n11520_));
  NAND2_X1   g11328(.A1(new_n11519_), .A2(\asqrt[19] ), .ZN(new_n11521_));
  NAND3_X1   g11329(.A1(new_n11520_), .A2(new_n10045_), .A3(new_n11521_), .ZN(new_n11522_));
  NOR3_X1    g11330(.A1(new_n11406_), .A2(new_n11115_), .A3(new_n11091_), .ZN(new_n11523_));
  XOR2_X1    g11331(.A1(new_n11523_), .A2(new_n11117_), .Z(new_n11524_));
  NAND2_X1   g11332(.A1(new_n11522_), .A2(new_n11524_), .ZN(new_n11525_));
  NAND2_X1   g11333(.A1(new_n11520_), .A2(new_n11521_), .ZN(new_n11526_));
  AOI21_X1   g11334(.A1(new_n11526_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n11527_));
  AOI21_X1   g11335(.A1(new_n11527_), .A2(new_n11525_), .B(new_n11503_), .ZN(new_n11528_));
  OAI21_X1   g11336(.A1(new_n11508_), .A2(new_n11505_), .B(new_n10571_), .ZN(new_n11529_));
  NAND3_X1   g11337(.A1(new_n11504_), .A2(\a[36] ), .A3(new_n11506_), .ZN(new_n11530_));
  NAND2_X1   g11338(.A1(new_n11529_), .A2(new_n11530_), .ZN(new_n11531_));
  NAND2_X1   g11339(.A1(\asqrt[17] ), .A2(\a[34] ), .ZN(new_n11532_));
  AOI21_X1   g11340(.A1(new_n11532_), .A2(new_n11513_), .B(new_n10953_), .ZN(new_n11533_));
  AOI21_X1   g11341(.A1(\asqrt[17] ), .A2(new_n11084_), .B(new_n11085_), .ZN(new_n11534_));
  NOR2_X1    g11342(.A1(new_n11534_), .A2(new_n11508_), .ZN(new_n11535_));
  NAND3_X1   g11343(.A1(new_n11532_), .A2(new_n10953_), .A3(new_n11513_), .ZN(new_n11536_));
  AOI21_X1   g11344(.A1(new_n11535_), .A2(new_n11536_), .B(new_n11533_), .ZN(new_n11537_));
  AOI21_X1   g11345(.A1(new_n11537_), .A2(new_n10478_), .B(new_n11531_), .ZN(new_n11538_));
  NOR2_X1    g11346(.A1(new_n11537_), .A2(new_n10478_), .ZN(new_n11539_));
  OAI21_X1   g11347(.A1(new_n11538_), .A2(new_n11539_), .B(\asqrt[20] ), .ZN(new_n11540_));
  AOI21_X1   g11348(.A1(new_n11525_), .A2(new_n11540_), .B(new_n9590_), .ZN(new_n11541_));
  NOR2_X1    g11349(.A1(new_n11528_), .A2(new_n11541_), .ZN(new_n11542_));
  AOI21_X1   g11350(.A1(new_n11542_), .A2(new_n9177_), .B(new_n11499_), .ZN(new_n11543_));
  OAI21_X1   g11351(.A1(new_n11528_), .A2(new_n11541_), .B(\asqrt[22] ), .ZN(new_n11544_));
  NAND2_X1   g11352(.A1(new_n11544_), .A2(new_n8742_), .ZN(new_n11545_));
  OAI21_X1   g11353(.A1(new_n11543_), .A2(new_n11545_), .B(new_n11496_), .ZN(new_n11546_));
  INV_X1     g11354(.I(new_n11544_), .ZN(new_n11547_));
  OAI21_X1   g11355(.A1(new_n11543_), .A2(new_n11547_), .B(\asqrt[23] ), .ZN(new_n11548_));
  NAND3_X1   g11356(.A1(new_n11546_), .A2(new_n11548_), .A3(new_n8349_), .ZN(new_n11549_));
  NAND2_X1   g11357(.A1(new_n11549_), .A2(new_n11493_), .ZN(new_n11550_));
  NAND2_X1   g11358(.A1(new_n11546_), .A2(new_n11548_), .ZN(new_n11551_));
  AOI21_X1   g11359(.A1(new_n11551_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n11552_));
  AOI21_X1   g11360(.A1(new_n11552_), .A2(new_n11550_), .B(new_n11490_), .ZN(new_n11553_));
  INV_X1     g11361(.I(new_n11496_), .ZN(new_n11554_));
  NOR2_X1    g11362(.A1(new_n11538_), .A2(new_n11539_), .ZN(new_n11555_));
  INV_X1     g11363(.I(new_n11524_), .ZN(new_n11556_));
  AOI21_X1   g11364(.A1(new_n11555_), .A2(new_n10045_), .B(new_n11556_), .ZN(new_n11557_));
  NAND2_X1   g11365(.A1(new_n11540_), .A2(new_n9590_), .ZN(new_n11558_));
  OAI21_X1   g11366(.A1(new_n11557_), .A2(new_n11558_), .B(new_n11502_), .ZN(new_n11559_));
  INV_X1     g11367(.I(new_n11540_), .ZN(new_n11560_));
  OAI21_X1   g11368(.A1(new_n11557_), .A2(new_n11560_), .B(\asqrt[21] ), .ZN(new_n11561_));
  NAND3_X1   g11369(.A1(new_n11559_), .A2(new_n11561_), .A3(new_n9177_), .ZN(new_n11562_));
  NAND2_X1   g11370(.A1(new_n11562_), .A2(new_n11498_), .ZN(new_n11563_));
  NAND2_X1   g11371(.A1(new_n11559_), .A2(new_n11561_), .ZN(new_n11564_));
  AOI21_X1   g11372(.A1(new_n11564_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n11565_));
  AOI21_X1   g11373(.A1(new_n11565_), .A2(new_n11563_), .B(new_n11554_), .ZN(new_n11566_));
  AOI21_X1   g11374(.A1(new_n11563_), .A2(new_n11544_), .B(new_n8742_), .ZN(new_n11567_));
  OAI21_X1   g11375(.A1(new_n11566_), .A2(new_n11567_), .B(\asqrt[24] ), .ZN(new_n11568_));
  AOI21_X1   g11376(.A1(new_n11550_), .A2(new_n11568_), .B(new_n7934_), .ZN(new_n11569_));
  NOR2_X1    g11377(.A1(new_n11553_), .A2(new_n11569_), .ZN(new_n11570_));
  AOI21_X1   g11378(.A1(new_n11570_), .A2(new_n7561_), .B(new_n11487_), .ZN(new_n11571_));
  OAI21_X1   g11379(.A1(new_n11553_), .A2(new_n11569_), .B(\asqrt[26] ), .ZN(new_n11572_));
  NAND2_X1   g11380(.A1(new_n11572_), .A2(new_n7166_), .ZN(new_n11573_));
  OAI21_X1   g11381(.A1(new_n11571_), .A2(new_n11573_), .B(new_n11483_), .ZN(new_n11574_));
  INV_X1     g11382(.I(new_n11572_), .ZN(new_n11575_));
  OAI21_X1   g11383(.A1(new_n11571_), .A2(new_n11575_), .B(\asqrt[27] ), .ZN(new_n11576_));
  NAND3_X1   g11384(.A1(new_n11574_), .A2(new_n11576_), .A3(new_n6813_), .ZN(new_n11577_));
  NAND2_X1   g11385(.A1(new_n11577_), .A2(new_n11481_), .ZN(new_n11578_));
  NAND2_X1   g11386(.A1(new_n11574_), .A2(new_n11576_), .ZN(new_n11579_));
  AOI21_X1   g11387(.A1(new_n11579_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n11580_));
  AOI21_X1   g11388(.A1(new_n11580_), .A2(new_n11578_), .B(new_n11478_), .ZN(new_n11581_));
  INV_X1     g11389(.I(new_n11483_), .ZN(new_n11582_));
  INV_X1     g11390(.I(new_n11493_), .ZN(new_n11583_));
  NOR2_X1    g11391(.A1(new_n11566_), .A2(new_n11567_), .ZN(new_n11584_));
  AOI21_X1   g11392(.A1(new_n11584_), .A2(new_n8349_), .B(new_n11583_), .ZN(new_n11585_));
  NAND2_X1   g11393(.A1(new_n11568_), .A2(new_n7934_), .ZN(new_n11586_));
  OAI21_X1   g11394(.A1(new_n11585_), .A2(new_n11586_), .B(new_n11489_), .ZN(new_n11587_));
  INV_X1     g11395(.I(new_n11568_), .ZN(new_n11588_));
  OAI21_X1   g11396(.A1(new_n11585_), .A2(new_n11588_), .B(\asqrt[25] ), .ZN(new_n11589_));
  NAND3_X1   g11397(.A1(new_n11587_), .A2(new_n11589_), .A3(new_n7561_), .ZN(new_n11590_));
  NAND2_X1   g11398(.A1(new_n11590_), .A2(new_n11486_), .ZN(new_n11591_));
  NAND2_X1   g11399(.A1(new_n11587_), .A2(new_n11589_), .ZN(new_n11592_));
  AOI21_X1   g11400(.A1(new_n11592_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n11593_));
  AOI21_X1   g11401(.A1(new_n11593_), .A2(new_n11591_), .B(new_n11582_), .ZN(new_n11594_));
  AOI21_X1   g11402(.A1(new_n11591_), .A2(new_n11572_), .B(new_n7166_), .ZN(new_n11595_));
  OAI21_X1   g11403(.A1(new_n11594_), .A2(new_n11595_), .B(\asqrt[28] ), .ZN(new_n11596_));
  AOI21_X1   g11404(.A1(new_n11578_), .A2(new_n11596_), .B(new_n6454_), .ZN(new_n11597_));
  NOR2_X1    g11405(.A1(new_n11581_), .A2(new_n11597_), .ZN(new_n11598_));
  AOI21_X1   g11406(.A1(new_n11598_), .A2(new_n6106_), .B(new_n11475_), .ZN(new_n11599_));
  OAI21_X1   g11407(.A1(new_n11581_), .A2(new_n11597_), .B(\asqrt[30] ), .ZN(new_n11600_));
  NAND2_X1   g11408(.A1(new_n11600_), .A2(new_n5750_), .ZN(new_n11601_));
  OAI21_X1   g11409(.A1(new_n11599_), .A2(new_n11601_), .B(new_n11471_), .ZN(new_n11602_));
  INV_X1     g11410(.I(new_n11600_), .ZN(new_n11603_));
  OAI21_X1   g11411(.A1(new_n11599_), .A2(new_n11603_), .B(\asqrt[31] ), .ZN(new_n11604_));
  NAND3_X1   g11412(.A1(new_n11602_), .A2(new_n11604_), .A3(new_n5435_), .ZN(new_n11605_));
  NAND2_X1   g11413(.A1(new_n11605_), .A2(new_n11469_), .ZN(new_n11606_));
  NAND2_X1   g11414(.A1(new_n11602_), .A2(new_n11604_), .ZN(new_n11607_));
  AOI21_X1   g11415(.A1(new_n11607_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n11608_));
  AOI21_X1   g11416(.A1(new_n11608_), .A2(new_n11606_), .B(new_n11466_), .ZN(new_n11609_));
  INV_X1     g11417(.I(new_n11471_), .ZN(new_n11610_));
  INV_X1     g11418(.I(new_n11481_), .ZN(new_n11611_));
  NOR2_X1    g11419(.A1(new_n11594_), .A2(new_n11595_), .ZN(new_n11612_));
  AOI21_X1   g11420(.A1(new_n11612_), .A2(new_n6813_), .B(new_n11611_), .ZN(new_n11613_));
  NAND2_X1   g11421(.A1(new_n11596_), .A2(new_n6454_), .ZN(new_n11614_));
  OAI21_X1   g11422(.A1(new_n11613_), .A2(new_n11614_), .B(new_n11477_), .ZN(new_n11615_));
  INV_X1     g11423(.I(new_n11596_), .ZN(new_n11616_));
  OAI21_X1   g11424(.A1(new_n11613_), .A2(new_n11616_), .B(\asqrt[29] ), .ZN(new_n11617_));
  NAND3_X1   g11425(.A1(new_n11615_), .A2(new_n11617_), .A3(new_n6106_), .ZN(new_n11618_));
  NAND2_X1   g11426(.A1(new_n11618_), .A2(new_n11474_), .ZN(new_n11619_));
  NAND2_X1   g11427(.A1(new_n11615_), .A2(new_n11617_), .ZN(new_n11620_));
  AOI21_X1   g11428(.A1(new_n11620_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n11621_));
  AOI21_X1   g11429(.A1(new_n11621_), .A2(new_n11619_), .B(new_n11610_), .ZN(new_n11622_));
  AOI21_X1   g11430(.A1(new_n11619_), .A2(new_n11600_), .B(new_n5750_), .ZN(new_n11623_));
  OAI21_X1   g11431(.A1(new_n11622_), .A2(new_n11623_), .B(\asqrt[32] ), .ZN(new_n11624_));
  AOI21_X1   g11432(.A1(new_n11606_), .A2(new_n11624_), .B(new_n5110_), .ZN(new_n11625_));
  NOR2_X1    g11433(.A1(new_n11609_), .A2(new_n11625_), .ZN(new_n11626_));
  AOI21_X1   g11434(.A1(new_n11626_), .A2(new_n4810_), .B(new_n11463_), .ZN(new_n11627_));
  OAI21_X1   g11435(.A1(new_n11609_), .A2(new_n11625_), .B(\asqrt[34] ), .ZN(new_n11628_));
  NAND2_X1   g11436(.A1(new_n11628_), .A2(new_n4510_), .ZN(new_n11629_));
  OAI21_X1   g11437(.A1(new_n11627_), .A2(new_n11629_), .B(new_n11459_), .ZN(new_n11630_));
  INV_X1     g11438(.I(new_n11628_), .ZN(new_n11631_));
  OAI21_X1   g11439(.A1(new_n11627_), .A2(new_n11631_), .B(\asqrt[35] ), .ZN(new_n11632_));
  NAND3_X1   g11440(.A1(new_n11630_), .A2(new_n11632_), .A3(new_n4224_), .ZN(new_n11633_));
  NAND2_X1   g11441(.A1(new_n11633_), .A2(new_n11457_), .ZN(new_n11634_));
  NAND2_X1   g11442(.A1(new_n11630_), .A2(new_n11632_), .ZN(new_n11635_));
  AOI21_X1   g11443(.A1(new_n11635_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n11636_));
  AOI21_X1   g11444(.A1(new_n11636_), .A2(new_n11634_), .B(new_n11454_), .ZN(new_n11637_));
  INV_X1     g11445(.I(new_n11459_), .ZN(new_n11638_));
  INV_X1     g11446(.I(new_n11469_), .ZN(new_n11639_));
  NOR2_X1    g11447(.A1(new_n11622_), .A2(new_n11623_), .ZN(new_n11640_));
  AOI21_X1   g11448(.A1(new_n11640_), .A2(new_n5435_), .B(new_n11639_), .ZN(new_n11641_));
  NAND2_X1   g11449(.A1(new_n11624_), .A2(new_n5110_), .ZN(new_n11642_));
  OAI21_X1   g11450(.A1(new_n11641_), .A2(new_n11642_), .B(new_n11465_), .ZN(new_n11643_));
  INV_X1     g11451(.I(new_n11624_), .ZN(new_n11644_));
  OAI21_X1   g11452(.A1(new_n11641_), .A2(new_n11644_), .B(\asqrt[33] ), .ZN(new_n11645_));
  NAND3_X1   g11453(.A1(new_n11643_), .A2(new_n11645_), .A3(new_n4810_), .ZN(new_n11646_));
  NAND2_X1   g11454(.A1(new_n11646_), .A2(new_n11462_), .ZN(new_n11647_));
  NAND2_X1   g11455(.A1(new_n11643_), .A2(new_n11645_), .ZN(new_n11648_));
  AOI21_X1   g11456(.A1(new_n11648_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n11649_));
  AOI21_X1   g11457(.A1(new_n11649_), .A2(new_n11647_), .B(new_n11638_), .ZN(new_n11650_));
  AOI21_X1   g11458(.A1(new_n11647_), .A2(new_n11628_), .B(new_n4510_), .ZN(new_n11651_));
  OAI21_X1   g11459(.A1(new_n11650_), .A2(new_n11651_), .B(\asqrt[36] ), .ZN(new_n11652_));
  AOI21_X1   g11460(.A1(new_n11634_), .A2(new_n11652_), .B(new_n3928_), .ZN(new_n11653_));
  NOR2_X1    g11461(.A1(new_n11637_), .A2(new_n11653_), .ZN(new_n11654_));
  AOI21_X1   g11462(.A1(new_n11654_), .A2(new_n3675_), .B(new_n11451_), .ZN(new_n11655_));
  OAI21_X1   g11463(.A1(new_n11637_), .A2(new_n11653_), .B(\asqrt[38] ), .ZN(new_n11656_));
  NAND2_X1   g11464(.A1(new_n11656_), .A2(new_n3400_), .ZN(new_n11657_));
  OAI21_X1   g11465(.A1(new_n11655_), .A2(new_n11657_), .B(new_n11447_), .ZN(new_n11658_));
  INV_X1     g11466(.I(new_n11656_), .ZN(new_n11659_));
  OAI21_X1   g11467(.A1(new_n11655_), .A2(new_n11659_), .B(\asqrt[39] ), .ZN(new_n11660_));
  NAND3_X1   g11468(.A1(new_n11658_), .A2(new_n11660_), .A3(new_n3167_), .ZN(new_n11661_));
  NAND2_X1   g11469(.A1(new_n11661_), .A2(new_n11445_), .ZN(new_n11662_));
  NAND2_X1   g11470(.A1(new_n11658_), .A2(new_n11660_), .ZN(new_n11663_));
  AOI21_X1   g11471(.A1(new_n11663_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n11664_));
  AOI21_X1   g11472(.A1(new_n11664_), .A2(new_n11662_), .B(new_n11442_), .ZN(new_n11665_));
  INV_X1     g11473(.I(new_n11447_), .ZN(new_n11666_));
  INV_X1     g11474(.I(new_n11457_), .ZN(new_n11667_));
  NOR2_X1    g11475(.A1(new_n11650_), .A2(new_n11651_), .ZN(new_n11668_));
  AOI21_X1   g11476(.A1(new_n11668_), .A2(new_n4224_), .B(new_n11667_), .ZN(new_n11669_));
  NAND2_X1   g11477(.A1(new_n11652_), .A2(new_n3928_), .ZN(new_n11670_));
  OAI21_X1   g11478(.A1(new_n11669_), .A2(new_n11670_), .B(new_n11453_), .ZN(new_n11671_));
  INV_X1     g11479(.I(new_n11652_), .ZN(new_n11672_));
  OAI21_X1   g11480(.A1(new_n11669_), .A2(new_n11672_), .B(\asqrt[37] ), .ZN(new_n11673_));
  NAND3_X1   g11481(.A1(new_n11671_), .A2(new_n11673_), .A3(new_n3675_), .ZN(new_n11674_));
  NAND2_X1   g11482(.A1(new_n11674_), .A2(new_n11450_), .ZN(new_n11675_));
  NAND2_X1   g11483(.A1(new_n11671_), .A2(new_n11673_), .ZN(new_n11676_));
  AOI21_X1   g11484(.A1(new_n11676_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n11677_));
  AOI21_X1   g11485(.A1(new_n11677_), .A2(new_n11675_), .B(new_n11666_), .ZN(new_n11678_));
  AOI21_X1   g11486(.A1(new_n11675_), .A2(new_n11656_), .B(new_n3400_), .ZN(new_n11679_));
  OAI21_X1   g11487(.A1(new_n11678_), .A2(new_n11679_), .B(\asqrt[40] ), .ZN(new_n11680_));
  AOI21_X1   g11488(.A1(new_n11662_), .A2(new_n11680_), .B(new_n2912_), .ZN(new_n11681_));
  NOR2_X1    g11489(.A1(new_n11665_), .A2(new_n11681_), .ZN(new_n11682_));
  AOI21_X1   g11490(.A1(new_n11682_), .A2(new_n2699_), .B(new_n11439_), .ZN(new_n11683_));
  OAI21_X1   g11491(.A1(new_n11665_), .A2(new_n11681_), .B(\asqrt[42] ), .ZN(new_n11684_));
  NAND2_X1   g11492(.A1(new_n11684_), .A2(new_n2464_), .ZN(new_n11685_));
  OAI21_X1   g11493(.A1(new_n11683_), .A2(new_n11685_), .B(new_n11435_), .ZN(new_n11686_));
  INV_X1     g11494(.I(new_n11684_), .ZN(new_n11687_));
  OAI21_X1   g11495(.A1(new_n11683_), .A2(new_n11687_), .B(\asqrt[43] ), .ZN(new_n11688_));
  NAND3_X1   g11496(.A1(new_n11686_), .A2(new_n11688_), .A3(new_n2271_), .ZN(new_n11689_));
  NAND2_X1   g11497(.A1(new_n11689_), .A2(new_n11433_), .ZN(new_n11690_));
  NAND2_X1   g11498(.A1(new_n11686_), .A2(new_n11688_), .ZN(new_n11691_));
  AOI21_X1   g11499(.A1(new_n11691_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n11692_));
  AOI21_X1   g11500(.A1(new_n11692_), .A2(new_n11690_), .B(new_n11430_), .ZN(new_n11693_));
  INV_X1     g11501(.I(new_n11435_), .ZN(new_n11694_));
  INV_X1     g11502(.I(new_n11445_), .ZN(new_n11695_));
  NOR2_X1    g11503(.A1(new_n11678_), .A2(new_n11679_), .ZN(new_n11696_));
  AOI21_X1   g11504(.A1(new_n11696_), .A2(new_n3167_), .B(new_n11695_), .ZN(new_n11697_));
  NAND2_X1   g11505(.A1(new_n11680_), .A2(new_n2912_), .ZN(new_n11698_));
  OAI21_X1   g11506(.A1(new_n11697_), .A2(new_n11698_), .B(new_n11441_), .ZN(new_n11699_));
  INV_X1     g11507(.I(new_n11680_), .ZN(new_n11700_));
  OAI21_X1   g11508(.A1(new_n11697_), .A2(new_n11700_), .B(\asqrt[41] ), .ZN(new_n11701_));
  NAND3_X1   g11509(.A1(new_n11699_), .A2(new_n11701_), .A3(new_n2699_), .ZN(new_n11702_));
  NAND2_X1   g11510(.A1(new_n11702_), .A2(new_n11438_), .ZN(new_n11703_));
  NAND2_X1   g11511(.A1(new_n11699_), .A2(new_n11701_), .ZN(new_n11704_));
  AOI21_X1   g11512(.A1(new_n11704_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n11705_));
  AOI21_X1   g11513(.A1(new_n11705_), .A2(new_n11703_), .B(new_n11694_), .ZN(new_n11706_));
  AOI21_X1   g11514(.A1(new_n11703_), .A2(new_n11684_), .B(new_n2464_), .ZN(new_n11707_));
  OAI21_X1   g11515(.A1(new_n11706_), .A2(new_n11707_), .B(\asqrt[44] ), .ZN(new_n11708_));
  AOI21_X1   g11516(.A1(new_n11690_), .A2(new_n11708_), .B(new_n2072_), .ZN(new_n11709_));
  NOR2_X1    g11517(.A1(new_n11693_), .A2(new_n11709_), .ZN(new_n11710_));
  AOI21_X1   g11518(.A1(new_n11710_), .A2(new_n1884_), .B(new_n11427_), .ZN(new_n11711_));
  OAI21_X1   g11519(.A1(new_n11693_), .A2(new_n11709_), .B(\asqrt[46] ), .ZN(new_n11712_));
  NAND2_X1   g11520(.A1(new_n11712_), .A2(new_n1688_), .ZN(new_n11713_));
  OAI21_X1   g11521(.A1(new_n11711_), .A2(new_n11713_), .B(new_n11423_), .ZN(new_n11714_));
  INV_X1     g11522(.I(new_n11712_), .ZN(new_n11715_));
  OAI21_X1   g11523(.A1(new_n11711_), .A2(new_n11715_), .B(\asqrt[47] ), .ZN(new_n11716_));
  NAND3_X1   g11524(.A1(new_n11714_), .A2(new_n11716_), .A3(new_n1533_), .ZN(new_n11717_));
  INV_X1     g11525(.I(new_n11423_), .ZN(new_n11718_));
  INV_X1     g11526(.I(new_n11433_), .ZN(new_n11719_));
  NOR2_X1    g11527(.A1(new_n11706_), .A2(new_n11707_), .ZN(new_n11720_));
  AOI21_X1   g11528(.A1(new_n11720_), .A2(new_n2271_), .B(new_n11719_), .ZN(new_n11721_));
  NAND2_X1   g11529(.A1(new_n11708_), .A2(new_n2072_), .ZN(new_n11722_));
  OAI21_X1   g11530(.A1(new_n11721_), .A2(new_n11722_), .B(new_n11429_), .ZN(new_n11723_));
  INV_X1     g11531(.I(new_n11708_), .ZN(new_n11724_));
  OAI21_X1   g11532(.A1(new_n11721_), .A2(new_n11724_), .B(\asqrt[45] ), .ZN(new_n11725_));
  NAND3_X1   g11533(.A1(new_n11723_), .A2(new_n11725_), .A3(new_n1884_), .ZN(new_n11726_));
  NAND2_X1   g11534(.A1(new_n11726_), .A2(new_n11426_), .ZN(new_n11727_));
  NAND2_X1   g11535(.A1(new_n11723_), .A2(new_n11725_), .ZN(new_n11728_));
  AOI21_X1   g11536(.A1(new_n11728_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n11729_));
  AOI21_X1   g11537(.A1(new_n11729_), .A2(new_n11727_), .B(new_n11718_), .ZN(new_n11730_));
  AOI21_X1   g11538(.A1(new_n11727_), .A2(new_n11712_), .B(new_n1688_), .ZN(new_n11731_));
  OAI21_X1   g11539(.A1(new_n11730_), .A2(new_n11731_), .B(\asqrt[48] ), .ZN(new_n11732_));
  NAND2_X1   g11540(.A1(new_n11403_), .A2(new_n10958_), .ZN(new_n11733_));
  NOR2_X1    g11541(.A1(new_n11406_), .A2(new_n10958_), .ZN(new_n11734_));
  NAND2_X1   g11542(.A1(new_n11734_), .A2(new_n11418_), .ZN(new_n11735_));
  AOI21_X1   g11543(.A1(new_n11735_), .A2(new_n11733_), .B(new_n193_), .ZN(new_n11736_));
  INV_X1     g11544(.I(new_n11736_), .ZN(new_n11737_));
  NAND3_X1   g11545(.A1(\asqrt[17] ), .A2(new_n11388_), .A3(new_n11399_), .ZN(new_n11738_));
  XOR2_X1    g11546(.A1(new_n11738_), .A2(new_n11391_), .Z(new_n11739_));
  AOI21_X1   g11547(.A1(new_n11734_), .A2(new_n11403_), .B(new_n11404_), .ZN(new_n11740_));
  OAI21_X1   g11548(.A1(new_n11358_), .A2(new_n11360_), .B(new_n11363_), .ZN(new_n11741_));
  NOR2_X1    g11549(.A1(new_n11406_), .A2(new_n11741_), .ZN(new_n11742_));
  XOR2_X1    g11550(.A1(new_n11742_), .A2(new_n10966_), .Z(new_n11743_));
  NAND3_X1   g11551(.A1(\asqrt[17] ), .A2(new_n11374_), .A3(new_n11359_), .ZN(new_n11744_));
  XOR2_X1    g11552(.A1(new_n11744_), .A2(new_n10970_), .Z(new_n11745_));
  OAI21_X1   g11553(.A1(new_n11369_), .A2(new_n11370_), .B(new_n11373_), .ZN(new_n11746_));
  NOR2_X1    g11554(.A1(new_n11406_), .A2(new_n11746_), .ZN(new_n11747_));
  XOR2_X1    g11555(.A1(new_n11747_), .A2(new_n10972_), .Z(new_n11748_));
  INV_X1     g11556(.I(new_n11748_), .ZN(new_n11749_));
  NAND3_X1   g11557(.A1(\asqrt[17] ), .A2(new_n11336_), .A3(new_n11355_), .ZN(new_n11750_));
  XOR2_X1    g11558(.A1(new_n11750_), .A2(new_n11367_), .Z(new_n11751_));
  INV_X1     g11559(.I(new_n11751_), .ZN(new_n11752_));
  OAI21_X1   g11560(.A1(new_n11330_), .A2(new_n11332_), .B(new_n11335_), .ZN(new_n11753_));
  NOR2_X1    g11561(.A1(new_n11406_), .A2(new_n11753_), .ZN(new_n11754_));
  XOR2_X1    g11562(.A1(new_n11754_), .A2(new_n10978_), .Z(new_n11755_));
  NAND3_X1   g11563(.A1(\asqrt[17] ), .A2(new_n11349_), .A3(new_n11331_), .ZN(new_n11756_));
  XOR2_X1    g11564(.A1(new_n11756_), .A2(new_n10982_), .Z(new_n11757_));
  OAI21_X1   g11565(.A1(new_n11344_), .A2(new_n11345_), .B(new_n11348_), .ZN(new_n11758_));
  NOR2_X1    g11566(.A1(new_n11406_), .A2(new_n11758_), .ZN(new_n11759_));
  XOR2_X1    g11567(.A1(new_n11759_), .A2(new_n10984_), .Z(new_n11760_));
  INV_X1     g11568(.I(new_n11760_), .ZN(new_n11761_));
  NAND3_X1   g11569(.A1(\asqrt[17] ), .A2(new_n11308_), .A3(new_n11327_), .ZN(new_n11762_));
  XOR2_X1    g11570(.A1(new_n11762_), .A2(new_n11342_), .Z(new_n11763_));
  INV_X1     g11571(.I(new_n11763_), .ZN(new_n11764_));
  OAI21_X1   g11572(.A1(new_n11302_), .A2(new_n11304_), .B(new_n11307_), .ZN(new_n11765_));
  NOR2_X1    g11573(.A1(new_n11406_), .A2(new_n11765_), .ZN(new_n11766_));
  XOR2_X1    g11574(.A1(new_n11766_), .A2(new_n10990_), .Z(new_n11767_));
  NAND3_X1   g11575(.A1(\asqrt[17] ), .A2(new_n11321_), .A3(new_n11303_), .ZN(new_n11768_));
  XOR2_X1    g11576(.A1(new_n11768_), .A2(new_n10994_), .Z(new_n11769_));
  OAI21_X1   g11577(.A1(new_n11316_), .A2(new_n11317_), .B(new_n11320_), .ZN(new_n11770_));
  NOR2_X1    g11578(.A1(new_n11406_), .A2(new_n11770_), .ZN(new_n11771_));
  XOR2_X1    g11579(.A1(new_n11771_), .A2(new_n10996_), .Z(new_n11772_));
  INV_X1     g11580(.I(new_n11772_), .ZN(new_n11773_));
  NAND3_X1   g11581(.A1(\asqrt[17] ), .A2(new_n11280_), .A3(new_n11299_), .ZN(new_n11774_));
  XOR2_X1    g11582(.A1(new_n11774_), .A2(new_n11314_), .Z(new_n11775_));
  INV_X1     g11583(.I(new_n11775_), .ZN(new_n11776_));
  NAND2_X1   g11584(.A1(new_n11717_), .A2(new_n11409_), .ZN(new_n11777_));
  NAND2_X1   g11585(.A1(new_n11714_), .A2(new_n11716_), .ZN(new_n11778_));
  AOI21_X1   g11586(.A1(new_n11778_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n11779_));
  AOI21_X1   g11587(.A1(new_n11779_), .A2(new_n11777_), .B(new_n11776_), .ZN(new_n11780_));
  AOI21_X1   g11588(.A1(new_n11777_), .A2(new_n11732_), .B(new_n1368_), .ZN(new_n11781_));
  NOR2_X1    g11589(.A1(new_n11780_), .A2(new_n11781_), .ZN(new_n11782_));
  AOI21_X1   g11590(.A1(new_n11782_), .A2(new_n1228_), .B(new_n11773_), .ZN(new_n11783_));
  OAI21_X1   g11591(.A1(new_n11780_), .A2(new_n11781_), .B(\asqrt[50] ), .ZN(new_n11784_));
  NAND2_X1   g11592(.A1(new_n11784_), .A2(new_n1088_), .ZN(new_n11785_));
  OAI21_X1   g11593(.A1(new_n11783_), .A2(new_n11785_), .B(new_n11769_), .ZN(new_n11786_));
  INV_X1     g11594(.I(new_n11784_), .ZN(new_n11787_));
  OAI21_X1   g11595(.A1(new_n11783_), .A2(new_n11787_), .B(\asqrt[51] ), .ZN(new_n11788_));
  NAND3_X1   g11596(.A1(new_n11786_), .A2(new_n11788_), .A3(new_n962_), .ZN(new_n11789_));
  NAND2_X1   g11597(.A1(new_n11789_), .A2(new_n11767_), .ZN(new_n11790_));
  NAND2_X1   g11598(.A1(new_n11786_), .A2(new_n11788_), .ZN(new_n11791_));
  AOI21_X1   g11599(.A1(new_n11791_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n11792_));
  AOI21_X1   g11600(.A1(new_n11792_), .A2(new_n11790_), .B(new_n11764_), .ZN(new_n11793_));
  INV_X1     g11601(.I(new_n11769_), .ZN(new_n11794_));
  NOR2_X1    g11602(.A1(new_n11730_), .A2(new_n11731_), .ZN(new_n11795_));
  AOI21_X1   g11603(.A1(new_n11795_), .A2(new_n1533_), .B(new_n11410_), .ZN(new_n11796_));
  NAND2_X1   g11604(.A1(new_n11732_), .A2(new_n1368_), .ZN(new_n11797_));
  OAI21_X1   g11605(.A1(new_n11796_), .A2(new_n11797_), .B(new_n11775_), .ZN(new_n11798_));
  INV_X1     g11606(.I(new_n11732_), .ZN(new_n11799_));
  OAI21_X1   g11607(.A1(new_n11796_), .A2(new_n11799_), .B(\asqrt[49] ), .ZN(new_n11800_));
  NAND3_X1   g11608(.A1(new_n11798_), .A2(new_n11800_), .A3(new_n1228_), .ZN(new_n11801_));
  NAND2_X1   g11609(.A1(new_n11801_), .A2(new_n11772_), .ZN(new_n11802_));
  NAND2_X1   g11610(.A1(new_n11798_), .A2(new_n11800_), .ZN(new_n11803_));
  AOI21_X1   g11611(.A1(new_n11803_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n11804_));
  AOI21_X1   g11612(.A1(new_n11804_), .A2(new_n11802_), .B(new_n11794_), .ZN(new_n11805_));
  AOI21_X1   g11613(.A1(new_n11802_), .A2(new_n11784_), .B(new_n1088_), .ZN(new_n11806_));
  OAI21_X1   g11614(.A1(new_n11805_), .A2(new_n11806_), .B(\asqrt[52] ), .ZN(new_n11807_));
  AOI21_X1   g11615(.A1(new_n11790_), .A2(new_n11807_), .B(new_n842_), .ZN(new_n11808_));
  NOR2_X1    g11616(.A1(new_n11793_), .A2(new_n11808_), .ZN(new_n11809_));
  AOI21_X1   g11617(.A1(new_n11809_), .A2(new_n720_), .B(new_n11761_), .ZN(new_n11810_));
  OAI21_X1   g11618(.A1(new_n11793_), .A2(new_n11808_), .B(\asqrt[54] ), .ZN(new_n11811_));
  NAND2_X1   g11619(.A1(new_n11811_), .A2(new_n630_), .ZN(new_n11812_));
  OAI21_X1   g11620(.A1(new_n11810_), .A2(new_n11812_), .B(new_n11757_), .ZN(new_n11813_));
  INV_X1     g11621(.I(new_n11811_), .ZN(new_n11814_));
  OAI21_X1   g11622(.A1(new_n11810_), .A2(new_n11814_), .B(\asqrt[55] ), .ZN(new_n11815_));
  NAND3_X1   g11623(.A1(new_n11813_), .A2(new_n11815_), .A3(new_n545_), .ZN(new_n11816_));
  NAND2_X1   g11624(.A1(new_n11816_), .A2(new_n11755_), .ZN(new_n11817_));
  NAND2_X1   g11625(.A1(new_n11813_), .A2(new_n11815_), .ZN(new_n11818_));
  AOI21_X1   g11626(.A1(new_n11818_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n11819_));
  AOI21_X1   g11627(.A1(new_n11819_), .A2(new_n11817_), .B(new_n11752_), .ZN(new_n11820_));
  INV_X1     g11628(.I(new_n11757_), .ZN(new_n11821_));
  INV_X1     g11629(.I(new_n11767_), .ZN(new_n11822_));
  NOR2_X1    g11630(.A1(new_n11805_), .A2(new_n11806_), .ZN(new_n11823_));
  AOI21_X1   g11631(.A1(new_n11823_), .A2(new_n962_), .B(new_n11822_), .ZN(new_n11824_));
  NAND2_X1   g11632(.A1(new_n11807_), .A2(new_n842_), .ZN(new_n11825_));
  OAI21_X1   g11633(.A1(new_n11824_), .A2(new_n11825_), .B(new_n11763_), .ZN(new_n11826_));
  INV_X1     g11634(.I(new_n11807_), .ZN(new_n11827_));
  OAI21_X1   g11635(.A1(new_n11824_), .A2(new_n11827_), .B(\asqrt[53] ), .ZN(new_n11828_));
  NAND3_X1   g11636(.A1(new_n11826_), .A2(new_n11828_), .A3(new_n720_), .ZN(new_n11829_));
  NAND2_X1   g11637(.A1(new_n11829_), .A2(new_n11760_), .ZN(new_n11830_));
  NAND2_X1   g11638(.A1(new_n11826_), .A2(new_n11828_), .ZN(new_n11831_));
  AOI21_X1   g11639(.A1(new_n11831_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n11832_));
  AOI21_X1   g11640(.A1(new_n11832_), .A2(new_n11830_), .B(new_n11821_), .ZN(new_n11833_));
  AOI21_X1   g11641(.A1(new_n11830_), .A2(new_n11811_), .B(new_n630_), .ZN(new_n11834_));
  OAI21_X1   g11642(.A1(new_n11833_), .A2(new_n11834_), .B(\asqrt[56] ), .ZN(new_n11835_));
  AOI21_X1   g11643(.A1(new_n11817_), .A2(new_n11835_), .B(new_n450_), .ZN(new_n11836_));
  NOR2_X1    g11644(.A1(new_n11820_), .A2(new_n11836_), .ZN(new_n11837_));
  AOI21_X1   g11645(.A1(new_n11837_), .A2(new_n403_), .B(new_n11749_), .ZN(new_n11838_));
  OAI21_X1   g11646(.A1(new_n11820_), .A2(new_n11836_), .B(\asqrt[58] ), .ZN(new_n11839_));
  NAND2_X1   g11647(.A1(new_n11839_), .A2(new_n339_), .ZN(new_n11840_));
  OAI21_X1   g11648(.A1(new_n11838_), .A2(new_n11840_), .B(new_n11745_), .ZN(new_n11841_));
  INV_X1     g11649(.I(new_n11839_), .ZN(new_n11842_));
  OAI21_X1   g11650(.A1(new_n11838_), .A2(new_n11842_), .B(\asqrt[59] ), .ZN(new_n11843_));
  NAND3_X1   g11651(.A1(new_n11841_), .A2(new_n11843_), .A3(new_n288_), .ZN(new_n11844_));
  NAND2_X1   g11652(.A1(new_n11844_), .A2(new_n11743_), .ZN(new_n11845_));
  INV_X1     g11653(.I(new_n11745_), .ZN(new_n11846_));
  INV_X1     g11654(.I(new_n11755_), .ZN(new_n11847_));
  NOR2_X1    g11655(.A1(new_n11833_), .A2(new_n11834_), .ZN(new_n11848_));
  AOI21_X1   g11656(.A1(new_n11848_), .A2(new_n545_), .B(new_n11847_), .ZN(new_n11849_));
  NAND2_X1   g11657(.A1(new_n11835_), .A2(new_n450_), .ZN(new_n11850_));
  OAI21_X1   g11658(.A1(new_n11849_), .A2(new_n11850_), .B(new_n11751_), .ZN(new_n11851_));
  INV_X1     g11659(.I(new_n11835_), .ZN(new_n11852_));
  OAI21_X1   g11660(.A1(new_n11849_), .A2(new_n11852_), .B(\asqrt[57] ), .ZN(new_n11853_));
  NAND3_X1   g11661(.A1(new_n11851_), .A2(new_n11853_), .A3(new_n403_), .ZN(new_n11854_));
  NAND2_X1   g11662(.A1(new_n11854_), .A2(new_n11748_), .ZN(new_n11855_));
  NAND2_X1   g11663(.A1(new_n11851_), .A2(new_n11853_), .ZN(new_n11856_));
  AOI21_X1   g11664(.A1(new_n11856_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n11857_));
  AOI21_X1   g11665(.A1(new_n11857_), .A2(new_n11855_), .B(new_n11846_), .ZN(new_n11858_));
  AOI21_X1   g11666(.A1(new_n11855_), .A2(new_n11839_), .B(new_n339_), .ZN(new_n11859_));
  OAI21_X1   g11667(.A1(new_n11858_), .A2(new_n11859_), .B(\asqrt[60] ), .ZN(new_n11860_));
  AOI21_X1   g11668(.A1(new_n11845_), .A2(new_n11860_), .B(new_n242_), .ZN(new_n11861_));
  NAND3_X1   g11669(.A1(\asqrt[17] ), .A2(new_n11364_), .A3(new_n11380_), .ZN(new_n11862_));
  XOR2_X1    g11670(.A1(new_n11862_), .A2(new_n11392_), .Z(new_n11863_));
  INV_X1     g11671(.I(new_n11863_), .ZN(new_n11864_));
  NAND2_X1   g11672(.A1(new_n11841_), .A2(new_n11843_), .ZN(new_n11865_));
  AOI21_X1   g11673(.A1(new_n11865_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n11866_));
  AOI21_X1   g11674(.A1(new_n11866_), .A2(new_n11845_), .B(new_n11864_), .ZN(new_n11867_));
  OAI21_X1   g11675(.A1(new_n11867_), .A2(new_n11861_), .B(\asqrt[62] ), .ZN(new_n11868_));
  INV_X1     g11676(.I(new_n11868_), .ZN(new_n11869_));
  NOR2_X1    g11677(.A1(new_n11867_), .A2(new_n11861_), .ZN(new_n11870_));
  AOI21_X1   g11678(.A1(new_n11365_), .A2(new_n11386_), .B(new_n11381_), .ZN(new_n11871_));
  NAND2_X1   g11679(.A1(\asqrt[17] ), .A2(new_n11871_), .ZN(new_n11872_));
  XOR2_X1    g11680(.A1(new_n11872_), .A2(new_n11384_), .Z(new_n11873_));
  INV_X1     g11681(.I(new_n11873_), .ZN(new_n11874_));
  AOI21_X1   g11682(.A1(new_n11870_), .A2(new_n234_), .B(new_n11874_), .ZN(new_n11875_));
  OAI21_X1   g11683(.A1(new_n11875_), .A2(new_n11869_), .B(new_n11740_), .ZN(new_n11876_));
  OAI21_X1   g11684(.A1(new_n11876_), .A2(new_n11739_), .B(new_n193_), .ZN(new_n11877_));
  NOR2_X1    g11685(.A1(new_n11875_), .A2(new_n11869_), .ZN(new_n11878_));
  NAND2_X1   g11686(.A1(new_n11878_), .A2(new_n11739_), .ZN(new_n11879_));
  NOR2_X1    g11687(.A1(\asqrt[17] ), .A2(new_n10959_), .ZN(new_n11880_));
  INV_X1     g11688(.I(new_n11880_), .ZN(new_n11881_));
  NAND4_X1   g11689(.A1(new_n11877_), .A2(new_n11737_), .A3(new_n11879_), .A4(new_n11881_), .ZN(\asqrt[16] ));
  NAND3_X1   g11690(.A1(\asqrt[16] ), .A2(new_n11717_), .A3(new_n11732_), .ZN(new_n11883_));
  XOR2_X1    g11691(.A1(new_n11883_), .A2(new_n11410_), .Z(new_n11884_));
  INV_X1     g11692(.I(new_n11743_), .ZN(new_n11885_));
  NOR2_X1    g11693(.A1(new_n11858_), .A2(new_n11859_), .ZN(new_n11886_));
  AOI21_X1   g11694(.A1(new_n11886_), .A2(new_n288_), .B(new_n11885_), .ZN(new_n11887_));
  INV_X1     g11695(.I(new_n11860_), .ZN(new_n11888_));
  OAI21_X1   g11696(.A1(new_n11887_), .A2(new_n11888_), .B(\asqrt[61] ), .ZN(new_n11889_));
  NAND2_X1   g11697(.A1(new_n11860_), .A2(new_n242_), .ZN(new_n11890_));
  OAI21_X1   g11698(.A1(new_n11887_), .A2(new_n11890_), .B(new_n11863_), .ZN(new_n11891_));
  NAND3_X1   g11699(.A1(new_n11891_), .A2(new_n11889_), .A3(new_n234_), .ZN(new_n11892_));
  NAND2_X1   g11700(.A1(new_n11892_), .A2(new_n11873_), .ZN(new_n11893_));
  NAND2_X1   g11701(.A1(new_n11893_), .A2(new_n11868_), .ZN(new_n11894_));
  NAND2_X1   g11702(.A1(new_n11894_), .A2(new_n11739_), .ZN(new_n11895_));
  INV_X1     g11703(.I(new_n11739_), .ZN(new_n11896_));
  INV_X1     g11704(.I(new_n11740_), .ZN(new_n11897_));
  AOI21_X1   g11705(.A1(new_n11893_), .A2(new_n11868_), .B(new_n11897_), .ZN(new_n11898_));
  AOI21_X1   g11706(.A1(new_n11898_), .A2(new_n11896_), .B(\asqrt[63] ), .ZN(new_n11899_));
  NOR2_X1    g11707(.A1(new_n11894_), .A2(new_n11896_), .ZN(new_n11900_));
  NOR4_X1    g11708(.A1(new_n11899_), .A2(new_n11736_), .A3(new_n11900_), .A4(new_n11880_), .ZN(new_n11901_));
  NOR2_X1    g11709(.A1(new_n11901_), .A2(new_n11739_), .ZN(new_n11902_));
  NAND2_X1   g11710(.A1(new_n11902_), .A2(new_n11878_), .ZN(new_n11903_));
  AOI21_X1   g11711(.A1(new_n11903_), .A2(new_n11895_), .B(new_n193_), .ZN(new_n11904_));
  NAND3_X1   g11712(.A1(\asqrt[16] ), .A2(new_n11868_), .A3(new_n11892_), .ZN(new_n11905_));
  XOR2_X1    g11713(.A1(new_n11905_), .A2(new_n11873_), .Z(new_n11906_));
  INV_X1     g11714(.I(new_n11906_), .ZN(new_n11907_));
  AOI21_X1   g11715(.A1(new_n11902_), .A2(new_n11894_), .B(new_n11900_), .ZN(new_n11908_));
  INV_X1     g11716(.I(new_n11908_), .ZN(new_n11909_));
  OAI21_X1   g11717(.A1(new_n11838_), .A2(new_n11840_), .B(new_n11843_), .ZN(new_n11910_));
  NOR2_X1    g11718(.A1(new_n11901_), .A2(new_n11910_), .ZN(new_n11911_));
  XOR2_X1    g11719(.A1(new_n11911_), .A2(new_n11745_), .Z(new_n11912_));
  NAND3_X1   g11720(.A1(\asqrt[16] ), .A2(new_n11854_), .A3(new_n11839_), .ZN(new_n11913_));
  XOR2_X1    g11721(.A1(new_n11913_), .A2(new_n11749_), .Z(new_n11914_));
  OAI21_X1   g11722(.A1(new_n11849_), .A2(new_n11850_), .B(new_n11853_), .ZN(new_n11915_));
  NOR2_X1    g11723(.A1(new_n11901_), .A2(new_n11915_), .ZN(new_n11916_));
  XOR2_X1    g11724(.A1(new_n11916_), .A2(new_n11751_), .Z(new_n11917_));
  INV_X1     g11725(.I(new_n11917_), .ZN(new_n11918_));
  NAND3_X1   g11726(.A1(\asqrt[16] ), .A2(new_n11816_), .A3(new_n11835_), .ZN(new_n11919_));
  XOR2_X1    g11727(.A1(new_n11919_), .A2(new_n11847_), .Z(new_n11920_));
  INV_X1     g11728(.I(new_n11920_), .ZN(new_n11921_));
  OAI21_X1   g11729(.A1(new_n11810_), .A2(new_n11812_), .B(new_n11815_), .ZN(new_n11922_));
  NOR2_X1    g11730(.A1(new_n11901_), .A2(new_n11922_), .ZN(new_n11923_));
  XOR2_X1    g11731(.A1(new_n11923_), .A2(new_n11757_), .Z(new_n11924_));
  NAND3_X1   g11732(.A1(\asqrt[16] ), .A2(new_n11829_), .A3(new_n11811_), .ZN(new_n11925_));
  XOR2_X1    g11733(.A1(new_n11925_), .A2(new_n11761_), .Z(new_n11926_));
  OAI21_X1   g11734(.A1(new_n11824_), .A2(new_n11825_), .B(new_n11828_), .ZN(new_n11927_));
  NOR2_X1    g11735(.A1(new_n11901_), .A2(new_n11927_), .ZN(new_n11928_));
  XOR2_X1    g11736(.A1(new_n11928_), .A2(new_n11763_), .Z(new_n11929_));
  INV_X1     g11737(.I(new_n11929_), .ZN(new_n11930_));
  NAND3_X1   g11738(.A1(\asqrt[16] ), .A2(new_n11789_), .A3(new_n11807_), .ZN(new_n11931_));
  XOR2_X1    g11739(.A1(new_n11931_), .A2(new_n11822_), .Z(new_n11932_));
  INV_X1     g11740(.I(new_n11932_), .ZN(new_n11933_));
  OAI21_X1   g11741(.A1(new_n11783_), .A2(new_n11785_), .B(new_n11788_), .ZN(new_n11934_));
  NOR2_X1    g11742(.A1(new_n11901_), .A2(new_n11934_), .ZN(new_n11935_));
  XOR2_X1    g11743(.A1(new_n11935_), .A2(new_n11769_), .Z(new_n11936_));
  NAND3_X1   g11744(.A1(\asqrt[16] ), .A2(new_n11801_), .A3(new_n11784_), .ZN(new_n11937_));
  XOR2_X1    g11745(.A1(new_n11937_), .A2(new_n11773_), .Z(new_n11938_));
  OAI21_X1   g11746(.A1(new_n11796_), .A2(new_n11797_), .B(new_n11800_), .ZN(new_n11939_));
  NOR2_X1    g11747(.A1(new_n11901_), .A2(new_n11939_), .ZN(new_n11940_));
  XOR2_X1    g11748(.A1(new_n11940_), .A2(new_n11775_), .Z(new_n11941_));
  INV_X1     g11749(.I(new_n11941_), .ZN(new_n11942_));
  INV_X1     g11750(.I(new_n11884_), .ZN(new_n11943_));
  OAI21_X1   g11751(.A1(new_n11711_), .A2(new_n11713_), .B(new_n11716_), .ZN(new_n11944_));
  NOR2_X1    g11752(.A1(new_n11901_), .A2(new_n11944_), .ZN(new_n11945_));
  XOR2_X1    g11753(.A1(new_n11945_), .A2(new_n11423_), .Z(new_n11946_));
  NAND3_X1   g11754(.A1(\asqrt[16] ), .A2(new_n11726_), .A3(new_n11712_), .ZN(new_n11947_));
  XOR2_X1    g11755(.A1(new_n11947_), .A2(new_n11427_), .Z(new_n11948_));
  OAI21_X1   g11756(.A1(new_n11721_), .A2(new_n11722_), .B(new_n11725_), .ZN(new_n11949_));
  NOR2_X1    g11757(.A1(new_n11901_), .A2(new_n11949_), .ZN(new_n11950_));
  XOR2_X1    g11758(.A1(new_n11950_), .A2(new_n11429_), .Z(new_n11951_));
  INV_X1     g11759(.I(new_n11951_), .ZN(new_n11952_));
  NAND3_X1   g11760(.A1(\asqrt[16] ), .A2(new_n11689_), .A3(new_n11708_), .ZN(new_n11953_));
  XOR2_X1    g11761(.A1(new_n11953_), .A2(new_n11719_), .Z(new_n11954_));
  INV_X1     g11762(.I(new_n11954_), .ZN(new_n11955_));
  OAI21_X1   g11763(.A1(new_n11683_), .A2(new_n11685_), .B(new_n11688_), .ZN(new_n11956_));
  NOR2_X1    g11764(.A1(new_n11901_), .A2(new_n11956_), .ZN(new_n11957_));
  XOR2_X1    g11765(.A1(new_n11957_), .A2(new_n11435_), .Z(new_n11958_));
  NAND3_X1   g11766(.A1(\asqrt[16] ), .A2(new_n11702_), .A3(new_n11684_), .ZN(new_n11959_));
  XOR2_X1    g11767(.A1(new_n11959_), .A2(new_n11439_), .Z(new_n11960_));
  OAI21_X1   g11768(.A1(new_n11697_), .A2(new_n11698_), .B(new_n11701_), .ZN(new_n11961_));
  NOR2_X1    g11769(.A1(new_n11901_), .A2(new_n11961_), .ZN(new_n11962_));
  XOR2_X1    g11770(.A1(new_n11962_), .A2(new_n11441_), .Z(new_n11963_));
  INV_X1     g11771(.I(new_n11963_), .ZN(new_n11964_));
  NAND3_X1   g11772(.A1(\asqrt[16] ), .A2(new_n11661_), .A3(new_n11680_), .ZN(new_n11965_));
  XOR2_X1    g11773(.A1(new_n11965_), .A2(new_n11695_), .Z(new_n11966_));
  INV_X1     g11774(.I(new_n11966_), .ZN(new_n11967_));
  OAI21_X1   g11775(.A1(new_n11655_), .A2(new_n11657_), .B(new_n11660_), .ZN(new_n11968_));
  NOR2_X1    g11776(.A1(new_n11901_), .A2(new_n11968_), .ZN(new_n11969_));
  XOR2_X1    g11777(.A1(new_n11969_), .A2(new_n11447_), .Z(new_n11970_));
  NAND3_X1   g11778(.A1(\asqrt[16] ), .A2(new_n11674_), .A3(new_n11656_), .ZN(new_n11971_));
  XOR2_X1    g11779(.A1(new_n11971_), .A2(new_n11451_), .Z(new_n11972_));
  OAI21_X1   g11780(.A1(new_n11669_), .A2(new_n11670_), .B(new_n11673_), .ZN(new_n11973_));
  NOR2_X1    g11781(.A1(new_n11901_), .A2(new_n11973_), .ZN(new_n11974_));
  XOR2_X1    g11782(.A1(new_n11974_), .A2(new_n11453_), .Z(new_n11975_));
  INV_X1     g11783(.I(new_n11975_), .ZN(new_n11976_));
  NAND3_X1   g11784(.A1(\asqrt[16] ), .A2(new_n11633_), .A3(new_n11652_), .ZN(new_n11977_));
  XOR2_X1    g11785(.A1(new_n11977_), .A2(new_n11667_), .Z(new_n11978_));
  INV_X1     g11786(.I(new_n11978_), .ZN(new_n11979_));
  OAI21_X1   g11787(.A1(new_n11627_), .A2(new_n11629_), .B(new_n11632_), .ZN(new_n11980_));
  NOR2_X1    g11788(.A1(new_n11901_), .A2(new_n11980_), .ZN(new_n11981_));
  XOR2_X1    g11789(.A1(new_n11981_), .A2(new_n11459_), .Z(new_n11982_));
  NAND3_X1   g11790(.A1(\asqrt[16] ), .A2(new_n11646_), .A3(new_n11628_), .ZN(new_n11983_));
  XOR2_X1    g11791(.A1(new_n11983_), .A2(new_n11463_), .Z(new_n11984_));
  OAI21_X1   g11792(.A1(new_n11641_), .A2(new_n11642_), .B(new_n11645_), .ZN(new_n11985_));
  NOR2_X1    g11793(.A1(new_n11901_), .A2(new_n11985_), .ZN(new_n11986_));
  XOR2_X1    g11794(.A1(new_n11986_), .A2(new_n11465_), .Z(new_n11987_));
  INV_X1     g11795(.I(new_n11987_), .ZN(new_n11988_));
  NAND3_X1   g11796(.A1(\asqrt[16] ), .A2(new_n11605_), .A3(new_n11624_), .ZN(new_n11989_));
  XOR2_X1    g11797(.A1(new_n11989_), .A2(new_n11639_), .Z(new_n11990_));
  INV_X1     g11798(.I(new_n11990_), .ZN(new_n11991_));
  OAI21_X1   g11799(.A1(new_n11599_), .A2(new_n11601_), .B(new_n11604_), .ZN(new_n11992_));
  NOR2_X1    g11800(.A1(new_n11901_), .A2(new_n11992_), .ZN(new_n11993_));
  XOR2_X1    g11801(.A1(new_n11993_), .A2(new_n11471_), .Z(new_n11994_));
  NAND3_X1   g11802(.A1(\asqrt[16] ), .A2(new_n11618_), .A3(new_n11600_), .ZN(new_n11995_));
  XOR2_X1    g11803(.A1(new_n11995_), .A2(new_n11475_), .Z(new_n11996_));
  OAI21_X1   g11804(.A1(new_n11613_), .A2(new_n11614_), .B(new_n11617_), .ZN(new_n11997_));
  NOR2_X1    g11805(.A1(new_n11901_), .A2(new_n11997_), .ZN(new_n11998_));
  XOR2_X1    g11806(.A1(new_n11998_), .A2(new_n11477_), .Z(new_n11999_));
  INV_X1     g11807(.I(new_n11999_), .ZN(new_n12000_));
  NAND3_X1   g11808(.A1(\asqrt[16] ), .A2(new_n11577_), .A3(new_n11596_), .ZN(new_n12001_));
  XOR2_X1    g11809(.A1(new_n12001_), .A2(new_n11611_), .Z(new_n12002_));
  INV_X1     g11810(.I(new_n12002_), .ZN(new_n12003_));
  OAI21_X1   g11811(.A1(new_n11571_), .A2(new_n11573_), .B(new_n11576_), .ZN(new_n12004_));
  NOR2_X1    g11812(.A1(new_n11901_), .A2(new_n12004_), .ZN(new_n12005_));
  XOR2_X1    g11813(.A1(new_n12005_), .A2(new_n11483_), .Z(new_n12006_));
  NAND3_X1   g11814(.A1(\asqrt[16] ), .A2(new_n11590_), .A3(new_n11572_), .ZN(new_n12007_));
  XOR2_X1    g11815(.A1(new_n12007_), .A2(new_n11487_), .Z(new_n12008_));
  OAI21_X1   g11816(.A1(new_n11585_), .A2(new_n11586_), .B(new_n11589_), .ZN(new_n12009_));
  NOR2_X1    g11817(.A1(new_n11901_), .A2(new_n12009_), .ZN(new_n12010_));
  XOR2_X1    g11818(.A1(new_n12010_), .A2(new_n11489_), .Z(new_n12011_));
  INV_X1     g11819(.I(new_n12011_), .ZN(new_n12012_));
  NAND3_X1   g11820(.A1(\asqrt[16] ), .A2(new_n11549_), .A3(new_n11568_), .ZN(new_n12013_));
  XOR2_X1    g11821(.A1(new_n12013_), .A2(new_n11583_), .Z(new_n12014_));
  INV_X1     g11822(.I(new_n12014_), .ZN(new_n12015_));
  OAI21_X1   g11823(.A1(new_n11543_), .A2(new_n11545_), .B(new_n11548_), .ZN(new_n12016_));
  NOR2_X1    g11824(.A1(new_n11901_), .A2(new_n12016_), .ZN(new_n12017_));
  XOR2_X1    g11825(.A1(new_n12017_), .A2(new_n11496_), .Z(new_n12018_));
  NAND3_X1   g11826(.A1(\asqrt[16] ), .A2(new_n11562_), .A3(new_n11544_), .ZN(new_n12019_));
  XOR2_X1    g11827(.A1(new_n12019_), .A2(new_n11499_), .Z(new_n12020_));
  OAI21_X1   g11828(.A1(new_n11557_), .A2(new_n11558_), .B(new_n11561_), .ZN(new_n12021_));
  NOR2_X1    g11829(.A1(new_n11901_), .A2(new_n12021_), .ZN(new_n12022_));
  XOR2_X1    g11830(.A1(new_n12022_), .A2(new_n11502_), .Z(new_n12023_));
  INV_X1     g11831(.I(new_n12023_), .ZN(new_n12024_));
  NAND3_X1   g11832(.A1(\asqrt[16] ), .A2(new_n11522_), .A3(new_n11540_), .ZN(new_n12025_));
  XOR2_X1    g11833(.A1(new_n12025_), .A2(new_n11556_), .Z(new_n12026_));
  INV_X1     g11834(.I(new_n12026_), .ZN(new_n12027_));
  NOR2_X1    g11835(.A1(new_n11519_), .A2(\asqrt[19] ), .ZN(new_n12028_));
  NOR3_X1    g11836(.A1(new_n11901_), .A2(new_n12028_), .A3(new_n11539_), .ZN(new_n12029_));
  XOR2_X1    g11837(.A1(new_n12029_), .A2(new_n11510_), .Z(new_n12030_));
  NOR3_X1    g11838(.A1(new_n11901_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n12031_));
  NOR4_X1    g11839(.A1(new_n11899_), .A2(new_n11406_), .A3(new_n11736_), .A4(new_n11900_), .ZN(new_n12032_));
  OAI21_X1   g11840(.A1(new_n12031_), .A2(new_n12032_), .B(new_n11084_), .ZN(new_n12033_));
  NAND3_X1   g11841(.A1(\asqrt[16] ), .A2(new_n11511_), .A3(new_n11512_), .ZN(new_n12034_));
  INV_X1     g11842(.I(new_n12032_), .ZN(new_n12035_));
  NAND3_X1   g11843(.A1(new_n12034_), .A2(\a[34] ), .A3(new_n12035_), .ZN(new_n12036_));
  NAND2_X1   g11844(.A1(new_n12033_), .A2(new_n12036_), .ZN(new_n12037_));
  INV_X1     g11845(.I(\a[30] ), .ZN(new_n12038_));
  INV_X1     g11846(.I(\a[31] ), .ZN(new_n12039_));
  NAND3_X1   g11847(.A1(new_n12038_), .A2(new_n12039_), .A3(new_n11511_), .ZN(new_n12040_));
  NAND2_X1   g11848(.A1(\asqrt[16] ), .A2(\a[32] ), .ZN(new_n12041_));
  AOI21_X1   g11849(.A1(new_n12041_), .A2(new_n12040_), .B(new_n11406_), .ZN(new_n12042_));
  AOI21_X1   g11850(.A1(\asqrt[16] ), .A2(new_n11511_), .B(new_n11512_), .ZN(new_n12043_));
  NOR2_X1    g11851(.A1(new_n12031_), .A2(new_n12043_), .ZN(new_n12044_));
  NAND3_X1   g11852(.A1(new_n12041_), .A2(new_n11406_), .A3(new_n12040_), .ZN(new_n12045_));
  AOI21_X1   g11853(.A1(new_n12044_), .A2(new_n12045_), .B(new_n12042_), .ZN(new_n12046_));
  AOI21_X1   g11854(.A1(new_n12046_), .A2(new_n10953_), .B(new_n12037_), .ZN(new_n12047_));
  NOR2_X1    g11855(.A1(new_n12046_), .A2(new_n10953_), .ZN(new_n12048_));
  NOR3_X1    g11856(.A1(new_n12047_), .A2(\asqrt[19] ), .A3(new_n12048_), .ZN(new_n12049_));
  NOR3_X1    g11857(.A1(new_n11901_), .A2(new_n11533_), .A3(new_n11518_), .ZN(new_n12050_));
  XOR2_X1    g11858(.A1(new_n12050_), .A2(new_n11535_), .Z(new_n12051_));
  INV_X1     g11859(.I(new_n12051_), .ZN(new_n12052_));
  OAI21_X1   g11860(.A1(new_n12047_), .A2(new_n12048_), .B(\asqrt[19] ), .ZN(new_n12053_));
  OAI21_X1   g11861(.A1(new_n12049_), .A2(new_n12052_), .B(new_n12053_), .ZN(new_n12054_));
  OAI21_X1   g11862(.A1(new_n12054_), .A2(\asqrt[20] ), .B(new_n12030_), .ZN(new_n12055_));
  AOI21_X1   g11863(.A1(new_n12054_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n12056_));
  AOI21_X1   g11864(.A1(new_n12056_), .A2(new_n12055_), .B(new_n12027_), .ZN(new_n12057_));
  NAND2_X1   g11865(.A1(new_n12054_), .A2(\asqrt[20] ), .ZN(new_n12058_));
  AOI21_X1   g11866(.A1(new_n12055_), .A2(new_n12058_), .B(new_n9590_), .ZN(new_n12059_));
  NOR2_X1    g11867(.A1(new_n12057_), .A2(new_n12059_), .ZN(new_n12060_));
  AOI21_X1   g11868(.A1(new_n12060_), .A2(new_n9177_), .B(new_n12024_), .ZN(new_n12061_));
  OAI21_X1   g11869(.A1(new_n12057_), .A2(new_n12059_), .B(\asqrt[22] ), .ZN(new_n12062_));
  NAND2_X1   g11870(.A1(new_n12062_), .A2(new_n8742_), .ZN(new_n12063_));
  OAI21_X1   g11871(.A1(new_n12061_), .A2(new_n12063_), .B(new_n12020_), .ZN(new_n12064_));
  INV_X1     g11872(.I(new_n12062_), .ZN(new_n12065_));
  OAI21_X1   g11873(.A1(new_n12061_), .A2(new_n12065_), .B(\asqrt[23] ), .ZN(new_n12066_));
  NAND3_X1   g11874(.A1(new_n12064_), .A2(new_n12066_), .A3(new_n8349_), .ZN(new_n12067_));
  NAND2_X1   g11875(.A1(new_n12067_), .A2(new_n12018_), .ZN(new_n12068_));
  NAND2_X1   g11876(.A1(new_n12064_), .A2(new_n12066_), .ZN(new_n12069_));
  AOI21_X1   g11877(.A1(new_n12069_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n12070_));
  AOI21_X1   g11878(.A1(new_n12070_), .A2(new_n12068_), .B(new_n12015_), .ZN(new_n12071_));
  INV_X1     g11879(.I(new_n12020_), .ZN(new_n12072_));
  INV_X1     g11880(.I(new_n12030_), .ZN(new_n12073_));
  AOI21_X1   g11881(.A1(new_n12034_), .A2(new_n12035_), .B(\a[34] ), .ZN(new_n12074_));
  NOR3_X1    g11882(.A1(new_n12031_), .A2(new_n11084_), .A3(new_n12032_), .ZN(new_n12075_));
  NOR2_X1    g11883(.A1(new_n12075_), .A2(new_n12074_), .ZN(new_n12076_));
  OAI21_X1   g11884(.A1(new_n11901_), .A2(new_n11511_), .B(new_n12040_), .ZN(new_n12077_));
  NAND2_X1   g11885(.A1(new_n12077_), .A2(\asqrt[17] ), .ZN(new_n12078_));
  OAI21_X1   g11886(.A1(new_n11901_), .A2(\a[32] ), .B(\a[33] ), .ZN(new_n12079_));
  NAND2_X1   g11887(.A1(new_n12079_), .A2(new_n12034_), .ZN(new_n12080_));
  NOR2_X1    g11888(.A1(new_n12077_), .A2(\asqrt[17] ), .ZN(new_n12081_));
  OAI21_X1   g11889(.A1(new_n12080_), .A2(new_n12081_), .B(new_n12078_), .ZN(new_n12082_));
  OAI21_X1   g11890(.A1(\asqrt[18] ), .A2(new_n12082_), .B(new_n12076_), .ZN(new_n12083_));
  NAND2_X1   g11891(.A1(new_n12082_), .A2(\asqrt[18] ), .ZN(new_n12084_));
  NAND3_X1   g11892(.A1(new_n12083_), .A2(new_n10478_), .A3(new_n12084_), .ZN(new_n12085_));
  AOI21_X1   g11893(.A1(new_n12083_), .A2(new_n12084_), .B(new_n10478_), .ZN(new_n12086_));
  AOI21_X1   g11894(.A1(new_n12085_), .A2(new_n12051_), .B(new_n12086_), .ZN(new_n12087_));
  AOI21_X1   g11895(.A1(new_n12087_), .A2(new_n10045_), .B(new_n12073_), .ZN(new_n12088_));
  OAI21_X1   g11896(.A1(new_n12087_), .A2(new_n10045_), .B(new_n9590_), .ZN(new_n12089_));
  OAI21_X1   g11897(.A1(new_n12088_), .A2(new_n12089_), .B(new_n12026_), .ZN(new_n12090_));
  NOR2_X1    g11898(.A1(new_n12087_), .A2(new_n10045_), .ZN(new_n12091_));
  OAI21_X1   g11899(.A1(new_n12088_), .A2(new_n12091_), .B(\asqrt[21] ), .ZN(new_n12092_));
  NAND3_X1   g11900(.A1(new_n12090_), .A2(new_n12092_), .A3(new_n9177_), .ZN(new_n12093_));
  NAND2_X1   g11901(.A1(new_n12093_), .A2(new_n12023_), .ZN(new_n12094_));
  NAND2_X1   g11902(.A1(new_n12090_), .A2(new_n12092_), .ZN(new_n12095_));
  AOI21_X1   g11903(.A1(new_n12095_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n12096_));
  AOI21_X1   g11904(.A1(new_n12096_), .A2(new_n12094_), .B(new_n12072_), .ZN(new_n12097_));
  AOI21_X1   g11905(.A1(new_n12094_), .A2(new_n12062_), .B(new_n8742_), .ZN(new_n12098_));
  OAI21_X1   g11906(.A1(new_n12097_), .A2(new_n12098_), .B(\asqrt[24] ), .ZN(new_n12099_));
  AOI21_X1   g11907(.A1(new_n12068_), .A2(new_n12099_), .B(new_n7934_), .ZN(new_n12100_));
  NOR2_X1    g11908(.A1(new_n12071_), .A2(new_n12100_), .ZN(new_n12101_));
  AOI21_X1   g11909(.A1(new_n12101_), .A2(new_n7561_), .B(new_n12012_), .ZN(new_n12102_));
  OAI21_X1   g11910(.A1(new_n12071_), .A2(new_n12100_), .B(\asqrt[26] ), .ZN(new_n12103_));
  NAND2_X1   g11911(.A1(new_n12103_), .A2(new_n7166_), .ZN(new_n12104_));
  OAI21_X1   g11912(.A1(new_n12102_), .A2(new_n12104_), .B(new_n12008_), .ZN(new_n12105_));
  INV_X1     g11913(.I(new_n12103_), .ZN(new_n12106_));
  OAI21_X1   g11914(.A1(new_n12102_), .A2(new_n12106_), .B(\asqrt[27] ), .ZN(new_n12107_));
  NAND3_X1   g11915(.A1(new_n12105_), .A2(new_n12107_), .A3(new_n6813_), .ZN(new_n12108_));
  NAND2_X1   g11916(.A1(new_n12108_), .A2(new_n12006_), .ZN(new_n12109_));
  NAND2_X1   g11917(.A1(new_n12105_), .A2(new_n12107_), .ZN(new_n12110_));
  AOI21_X1   g11918(.A1(new_n12110_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n12111_));
  AOI21_X1   g11919(.A1(new_n12111_), .A2(new_n12109_), .B(new_n12003_), .ZN(new_n12112_));
  INV_X1     g11920(.I(new_n12008_), .ZN(new_n12113_));
  INV_X1     g11921(.I(new_n12018_), .ZN(new_n12114_));
  NOR2_X1    g11922(.A1(new_n12097_), .A2(new_n12098_), .ZN(new_n12115_));
  AOI21_X1   g11923(.A1(new_n12115_), .A2(new_n8349_), .B(new_n12114_), .ZN(new_n12116_));
  NAND2_X1   g11924(.A1(new_n12099_), .A2(new_n7934_), .ZN(new_n12117_));
  OAI21_X1   g11925(.A1(new_n12116_), .A2(new_n12117_), .B(new_n12014_), .ZN(new_n12118_));
  INV_X1     g11926(.I(new_n12099_), .ZN(new_n12119_));
  OAI21_X1   g11927(.A1(new_n12116_), .A2(new_n12119_), .B(\asqrt[25] ), .ZN(new_n12120_));
  NAND3_X1   g11928(.A1(new_n12118_), .A2(new_n12120_), .A3(new_n7561_), .ZN(new_n12121_));
  NAND2_X1   g11929(.A1(new_n12121_), .A2(new_n12011_), .ZN(new_n12122_));
  NAND2_X1   g11930(.A1(new_n12118_), .A2(new_n12120_), .ZN(new_n12123_));
  AOI21_X1   g11931(.A1(new_n12123_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n12124_));
  AOI21_X1   g11932(.A1(new_n12124_), .A2(new_n12122_), .B(new_n12113_), .ZN(new_n12125_));
  AOI21_X1   g11933(.A1(new_n12122_), .A2(new_n12103_), .B(new_n7166_), .ZN(new_n12126_));
  OAI21_X1   g11934(.A1(new_n12125_), .A2(new_n12126_), .B(\asqrt[28] ), .ZN(new_n12127_));
  AOI21_X1   g11935(.A1(new_n12109_), .A2(new_n12127_), .B(new_n6454_), .ZN(new_n12128_));
  NOR2_X1    g11936(.A1(new_n12112_), .A2(new_n12128_), .ZN(new_n12129_));
  AOI21_X1   g11937(.A1(new_n12129_), .A2(new_n6106_), .B(new_n12000_), .ZN(new_n12130_));
  OAI21_X1   g11938(.A1(new_n12112_), .A2(new_n12128_), .B(\asqrt[30] ), .ZN(new_n12131_));
  NAND2_X1   g11939(.A1(new_n12131_), .A2(new_n5750_), .ZN(new_n12132_));
  OAI21_X1   g11940(.A1(new_n12130_), .A2(new_n12132_), .B(new_n11996_), .ZN(new_n12133_));
  INV_X1     g11941(.I(new_n12131_), .ZN(new_n12134_));
  OAI21_X1   g11942(.A1(new_n12130_), .A2(new_n12134_), .B(\asqrt[31] ), .ZN(new_n12135_));
  NAND3_X1   g11943(.A1(new_n12133_), .A2(new_n12135_), .A3(new_n5435_), .ZN(new_n12136_));
  NAND2_X1   g11944(.A1(new_n12136_), .A2(new_n11994_), .ZN(new_n12137_));
  NAND2_X1   g11945(.A1(new_n12133_), .A2(new_n12135_), .ZN(new_n12138_));
  AOI21_X1   g11946(.A1(new_n12138_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n12139_));
  AOI21_X1   g11947(.A1(new_n12139_), .A2(new_n12137_), .B(new_n11991_), .ZN(new_n12140_));
  INV_X1     g11948(.I(new_n11996_), .ZN(new_n12141_));
  INV_X1     g11949(.I(new_n12006_), .ZN(new_n12142_));
  NOR2_X1    g11950(.A1(new_n12125_), .A2(new_n12126_), .ZN(new_n12143_));
  AOI21_X1   g11951(.A1(new_n12143_), .A2(new_n6813_), .B(new_n12142_), .ZN(new_n12144_));
  NAND2_X1   g11952(.A1(new_n12127_), .A2(new_n6454_), .ZN(new_n12145_));
  OAI21_X1   g11953(.A1(new_n12144_), .A2(new_n12145_), .B(new_n12002_), .ZN(new_n12146_));
  INV_X1     g11954(.I(new_n12127_), .ZN(new_n12147_));
  OAI21_X1   g11955(.A1(new_n12144_), .A2(new_n12147_), .B(\asqrt[29] ), .ZN(new_n12148_));
  NAND3_X1   g11956(.A1(new_n12146_), .A2(new_n12148_), .A3(new_n6106_), .ZN(new_n12149_));
  NAND2_X1   g11957(.A1(new_n12149_), .A2(new_n11999_), .ZN(new_n12150_));
  NAND2_X1   g11958(.A1(new_n12146_), .A2(new_n12148_), .ZN(new_n12151_));
  AOI21_X1   g11959(.A1(new_n12151_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n12152_));
  AOI21_X1   g11960(.A1(new_n12152_), .A2(new_n12150_), .B(new_n12141_), .ZN(new_n12153_));
  AOI21_X1   g11961(.A1(new_n12150_), .A2(new_n12131_), .B(new_n5750_), .ZN(new_n12154_));
  OAI21_X1   g11962(.A1(new_n12153_), .A2(new_n12154_), .B(\asqrt[32] ), .ZN(new_n12155_));
  AOI21_X1   g11963(.A1(new_n12137_), .A2(new_n12155_), .B(new_n5110_), .ZN(new_n12156_));
  NOR2_X1    g11964(.A1(new_n12140_), .A2(new_n12156_), .ZN(new_n12157_));
  AOI21_X1   g11965(.A1(new_n12157_), .A2(new_n4810_), .B(new_n11988_), .ZN(new_n12158_));
  OAI21_X1   g11966(.A1(new_n12140_), .A2(new_n12156_), .B(\asqrt[34] ), .ZN(new_n12159_));
  NAND2_X1   g11967(.A1(new_n12159_), .A2(new_n4510_), .ZN(new_n12160_));
  OAI21_X1   g11968(.A1(new_n12158_), .A2(new_n12160_), .B(new_n11984_), .ZN(new_n12161_));
  INV_X1     g11969(.I(new_n12159_), .ZN(new_n12162_));
  OAI21_X1   g11970(.A1(new_n12158_), .A2(new_n12162_), .B(\asqrt[35] ), .ZN(new_n12163_));
  NAND3_X1   g11971(.A1(new_n12161_), .A2(new_n12163_), .A3(new_n4224_), .ZN(new_n12164_));
  NAND2_X1   g11972(.A1(new_n12164_), .A2(new_n11982_), .ZN(new_n12165_));
  NAND2_X1   g11973(.A1(new_n12161_), .A2(new_n12163_), .ZN(new_n12166_));
  AOI21_X1   g11974(.A1(new_n12166_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n12167_));
  AOI21_X1   g11975(.A1(new_n12167_), .A2(new_n12165_), .B(new_n11979_), .ZN(new_n12168_));
  INV_X1     g11976(.I(new_n11984_), .ZN(new_n12169_));
  INV_X1     g11977(.I(new_n11994_), .ZN(new_n12170_));
  NOR2_X1    g11978(.A1(new_n12153_), .A2(new_n12154_), .ZN(new_n12171_));
  AOI21_X1   g11979(.A1(new_n12171_), .A2(new_n5435_), .B(new_n12170_), .ZN(new_n12172_));
  NAND2_X1   g11980(.A1(new_n12155_), .A2(new_n5110_), .ZN(new_n12173_));
  OAI21_X1   g11981(.A1(new_n12172_), .A2(new_n12173_), .B(new_n11990_), .ZN(new_n12174_));
  INV_X1     g11982(.I(new_n12155_), .ZN(new_n12175_));
  OAI21_X1   g11983(.A1(new_n12172_), .A2(new_n12175_), .B(\asqrt[33] ), .ZN(new_n12176_));
  NAND3_X1   g11984(.A1(new_n12174_), .A2(new_n12176_), .A3(new_n4810_), .ZN(new_n12177_));
  NAND2_X1   g11985(.A1(new_n12177_), .A2(new_n11987_), .ZN(new_n12178_));
  NAND2_X1   g11986(.A1(new_n12174_), .A2(new_n12176_), .ZN(new_n12179_));
  AOI21_X1   g11987(.A1(new_n12179_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n12180_));
  AOI21_X1   g11988(.A1(new_n12180_), .A2(new_n12178_), .B(new_n12169_), .ZN(new_n12181_));
  AOI21_X1   g11989(.A1(new_n12178_), .A2(new_n12159_), .B(new_n4510_), .ZN(new_n12182_));
  OAI21_X1   g11990(.A1(new_n12181_), .A2(new_n12182_), .B(\asqrt[36] ), .ZN(new_n12183_));
  AOI21_X1   g11991(.A1(new_n12165_), .A2(new_n12183_), .B(new_n3928_), .ZN(new_n12184_));
  NOR2_X1    g11992(.A1(new_n12168_), .A2(new_n12184_), .ZN(new_n12185_));
  AOI21_X1   g11993(.A1(new_n12185_), .A2(new_n3675_), .B(new_n11976_), .ZN(new_n12186_));
  OAI21_X1   g11994(.A1(new_n12168_), .A2(new_n12184_), .B(\asqrt[38] ), .ZN(new_n12187_));
  NAND2_X1   g11995(.A1(new_n12187_), .A2(new_n3400_), .ZN(new_n12188_));
  OAI21_X1   g11996(.A1(new_n12186_), .A2(new_n12188_), .B(new_n11972_), .ZN(new_n12189_));
  INV_X1     g11997(.I(new_n12187_), .ZN(new_n12190_));
  OAI21_X1   g11998(.A1(new_n12186_), .A2(new_n12190_), .B(\asqrt[39] ), .ZN(new_n12191_));
  NAND3_X1   g11999(.A1(new_n12189_), .A2(new_n12191_), .A3(new_n3167_), .ZN(new_n12192_));
  NAND2_X1   g12000(.A1(new_n12192_), .A2(new_n11970_), .ZN(new_n12193_));
  NAND2_X1   g12001(.A1(new_n12189_), .A2(new_n12191_), .ZN(new_n12194_));
  AOI21_X1   g12002(.A1(new_n12194_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n12195_));
  AOI21_X1   g12003(.A1(new_n12195_), .A2(new_n12193_), .B(new_n11967_), .ZN(new_n12196_));
  INV_X1     g12004(.I(new_n11972_), .ZN(new_n12197_));
  INV_X1     g12005(.I(new_n11982_), .ZN(new_n12198_));
  NOR2_X1    g12006(.A1(new_n12181_), .A2(new_n12182_), .ZN(new_n12199_));
  AOI21_X1   g12007(.A1(new_n12199_), .A2(new_n4224_), .B(new_n12198_), .ZN(new_n12200_));
  NAND2_X1   g12008(.A1(new_n12183_), .A2(new_n3928_), .ZN(new_n12201_));
  OAI21_X1   g12009(.A1(new_n12200_), .A2(new_n12201_), .B(new_n11978_), .ZN(new_n12202_));
  INV_X1     g12010(.I(new_n12183_), .ZN(new_n12203_));
  OAI21_X1   g12011(.A1(new_n12200_), .A2(new_n12203_), .B(\asqrt[37] ), .ZN(new_n12204_));
  NAND3_X1   g12012(.A1(new_n12202_), .A2(new_n12204_), .A3(new_n3675_), .ZN(new_n12205_));
  NAND2_X1   g12013(.A1(new_n12205_), .A2(new_n11975_), .ZN(new_n12206_));
  NAND2_X1   g12014(.A1(new_n12202_), .A2(new_n12204_), .ZN(new_n12207_));
  AOI21_X1   g12015(.A1(new_n12207_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n12208_));
  AOI21_X1   g12016(.A1(new_n12208_), .A2(new_n12206_), .B(new_n12197_), .ZN(new_n12209_));
  AOI21_X1   g12017(.A1(new_n12206_), .A2(new_n12187_), .B(new_n3400_), .ZN(new_n12210_));
  OAI21_X1   g12018(.A1(new_n12209_), .A2(new_n12210_), .B(\asqrt[40] ), .ZN(new_n12211_));
  AOI21_X1   g12019(.A1(new_n12193_), .A2(new_n12211_), .B(new_n2912_), .ZN(new_n12212_));
  NOR2_X1    g12020(.A1(new_n12196_), .A2(new_n12212_), .ZN(new_n12213_));
  AOI21_X1   g12021(.A1(new_n12213_), .A2(new_n2699_), .B(new_n11964_), .ZN(new_n12214_));
  OAI21_X1   g12022(.A1(new_n12196_), .A2(new_n12212_), .B(\asqrt[42] ), .ZN(new_n12215_));
  NAND2_X1   g12023(.A1(new_n12215_), .A2(new_n2464_), .ZN(new_n12216_));
  OAI21_X1   g12024(.A1(new_n12214_), .A2(new_n12216_), .B(new_n11960_), .ZN(new_n12217_));
  INV_X1     g12025(.I(new_n12215_), .ZN(new_n12218_));
  OAI21_X1   g12026(.A1(new_n12214_), .A2(new_n12218_), .B(\asqrt[43] ), .ZN(new_n12219_));
  NAND3_X1   g12027(.A1(new_n12217_), .A2(new_n12219_), .A3(new_n2271_), .ZN(new_n12220_));
  NAND2_X1   g12028(.A1(new_n12220_), .A2(new_n11958_), .ZN(new_n12221_));
  NAND2_X1   g12029(.A1(new_n12217_), .A2(new_n12219_), .ZN(new_n12222_));
  AOI21_X1   g12030(.A1(new_n12222_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n12223_));
  AOI21_X1   g12031(.A1(new_n12223_), .A2(new_n12221_), .B(new_n11955_), .ZN(new_n12224_));
  INV_X1     g12032(.I(new_n11960_), .ZN(new_n12225_));
  INV_X1     g12033(.I(new_n11970_), .ZN(new_n12226_));
  NOR2_X1    g12034(.A1(new_n12209_), .A2(new_n12210_), .ZN(new_n12227_));
  AOI21_X1   g12035(.A1(new_n12227_), .A2(new_n3167_), .B(new_n12226_), .ZN(new_n12228_));
  NAND2_X1   g12036(.A1(new_n12211_), .A2(new_n2912_), .ZN(new_n12229_));
  OAI21_X1   g12037(.A1(new_n12228_), .A2(new_n12229_), .B(new_n11966_), .ZN(new_n12230_));
  INV_X1     g12038(.I(new_n12211_), .ZN(new_n12231_));
  OAI21_X1   g12039(.A1(new_n12228_), .A2(new_n12231_), .B(\asqrt[41] ), .ZN(new_n12232_));
  NAND3_X1   g12040(.A1(new_n12230_), .A2(new_n12232_), .A3(new_n2699_), .ZN(new_n12233_));
  NAND2_X1   g12041(.A1(new_n12233_), .A2(new_n11963_), .ZN(new_n12234_));
  NAND2_X1   g12042(.A1(new_n12230_), .A2(new_n12232_), .ZN(new_n12235_));
  AOI21_X1   g12043(.A1(new_n12235_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n12236_));
  AOI21_X1   g12044(.A1(new_n12236_), .A2(new_n12234_), .B(new_n12225_), .ZN(new_n12237_));
  AOI21_X1   g12045(.A1(new_n12234_), .A2(new_n12215_), .B(new_n2464_), .ZN(new_n12238_));
  OAI21_X1   g12046(.A1(new_n12237_), .A2(new_n12238_), .B(\asqrt[44] ), .ZN(new_n12239_));
  AOI21_X1   g12047(.A1(new_n12221_), .A2(new_n12239_), .B(new_n2072_), .ZN(new_n12240_));
  NOR2_X1    g12048(.A1(new_n12224_), .A2(new_n12240_), .ZN(new_n12241_));
  AOI21_X1   g12049(.A1(new_n12241_), .A2(new_n1884_), .B(new_n11952_), .ZN(new_n12242_));
  OAI21_X1   g12050(.A1(new_n12224_), .A2(new_n12240_), .B(\asqrt[46] ), .ZN(new_n12243_));
  NAND2_X1   g12051(.A1(new_n12243_), .A2(new_n1688_), .ZN(new_n12244_));
  OAI21_X1   g12052(.A1(new_n12242_), .A2(new_n12244_), .B(new_n11948_), .ZN(new_n12245_));
  INV_X1     g12053(.I(new_n12243_), .ZN(new_n12246_));
  OAI21_X1   g12054(.A1(new_n12242_), .A2(new_n12246_), .B(\asqrt[47] ), .ZN(new_n12247_));
  NAND3_X1   g12055(.A1(new_n12245_), .A2(new_n12247_), .A3(new_n1533_), .ZN(new_n12248_));
  NAND2_X1   g12056(.A1(new_n12248_), .A2(new_n11946_), .ZN(new_n12249_));
  NAND2_X1   g12057(.A1(new_n12245_), .A2(new_n12247_), .ZN(new_n12250_));
  AOI21_X1   g12058(.A1(new_n12250_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n12251_));
  AOI21_X1   g12059(.A1(new_n12251_), .A2(new_n12249_), .B(new_n11943_), .ZN(new_n12252_));
  INV_X1     g12060(.I(new_n11948_), .ZN(new_n12253_));
  INV_X1     g12061(.I(new_n11958_), .ZN(new_n12254_));
  NOR2_X1    g12062(.A1(new_n12237_), .A2(new_n12238_), .ZN(new_n12255_));
  AOI21_X1   g12063(.A1(new_n12255_), .A2(new_n2271_), .B(new_n12254_), .ZN(new_n12256_));
  NAND2_X1   g12064(.A1(new_n12239_), .A2(new_n2072_), .ZN(new_n12257_));
  OAI21_X1   g12065(.A1(new_n12256_), .A2(new_n12257_), .B(new_n11954_), .ZN(new_n12258_));
  INV_X1     g12066(.I(new_n12239_), .ZN(new_n12259_));
  OAI21_X1   g12067(.A1(new_n12256_), .A2(new_n12259_), .B(\asqrt[45] ), .ZN(new_n12260_));
  NAND3_X1   g12068(.A1(new_n12258_), .A2(new_n12260_), .A3(new_n1884_), .ZN(new_n12261_));
  NAND2_X1   g12069(.A1(new_n12261_), .A2(new_n11951_), .ZN(new_n12262_));
  NAND2_X1   g12070(.A1(new_n12258_), .A2(new_n12260_), .ZN(new_n12263_));
  AOI21_X1   g12071(.A1(new_n12263_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n12264_));
  AOI21_X1   g12072(.A1(new_n12264_), .A2(new_n12262_), .B(new_n12253_), .ZN(new_n12265_));
  AOI21_X1   g12073(.A1(new_n12262_), .A2(new_n12243_), .B(new_n1688_), .ZN(new_n12266_));
  OAI21_X1   g12074(.A1(new_n12265_), .A2(new_n12266_), .B(\asqrt[48] ), .ZN(new_n12267_));
  AOI21_X1   g12075(.A1(new_n12249_), .A2(new_n12267_), .B(new_n1368_), .ZN(new_n12268_));
  NOR2_X1    g12076(.A1(new_n12252_), .A2(new_n12268_), .ZN(new_n12269_));
  AOI21_X1   g12077(.A1(new_n12269_), .A2(new_n1228_), .B(new_n11942_), .ZN(new_n12270_));
  OAI21_X1   g12078(.A1(new_n12252_), .A2(new_n12268_), .B(\asqrt[50] ), .ZN(new_n12271_));
  NAND2_X1   g12079(.A1(new_n12271_), .A2(new_n1088_), .ZN(new_n12272_));
  OAI21_X1   g12080(.A1(new_n12270_), .A2(new_n12272_), .B(new_n11938_), .ZN(new_n12273_));
  INV_X1     g12081(.I(new_n12271_), .ZN(new_n12274_));
  OAI21_X1   g12082(.A1(new_n12270_), .A2(new_n12274_), .B(\asqrt[51] ), .ZN(new_n12275_));
  NAND3_X1   g12083(.A1(new_n12273_), .A2(new_n12275_), .A3(new_n962_), .ZN(new_n12276_));
  NAND2_X1   g12084(.A1(new_n12276_), .A2(new_n11936_), .ZN(new_n12277_));
  NAND2_X1   g12085(.A1(new_n12273_), .A2(new_n12275_), .ZN(new_n12278_));
  AOI21_X1   g12086(.A1(new_n12278_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n12279_));
  AOI21_X1   g12087(.A1(new_n12279_), .A2(new_n12277_), .B(new_n11933_), .ZN(new_n12280_));
  INV_X1     g12088(.I(new_n11938_), .ZN(new_n12281_));
  INV_X1     g12089(.I(new_n11946_), .ZN(new_n12282_));
  NOR2_X1    g12090(.A1(new_n12265_), .A2(new_n12266_), .ZN(new_n12283_));
  AOI21_X1   g12091(.A1(new_n12283_), .A2(new_n1533_), .B(new_n12282_), .ZN(new_n12284_));
  NAND2_X1   g12092(.A1(new_n12267_), .A2(new_n1368_), .ZN(new_n12285_));
  OAI21_X1   g12093(.A1(new_n12284_), .A2(new_n12285_), .B(new_n11884_), .ZN(new_n12286_));
  INV_X1     g12094(.I(new_n12267_), .ZN(new_n12287_));
  OAI21_X1   g12095(.A1(new_n12284_), .A2(new_n12287_), .B(\asqrt[49] ), .ZN(new_n12288_));
  NAND3_X1   g12096(.A1(new_n12286_), .A2(new_n12288_), .A3(new_n1228_), .ZN(new_n12289_));
  NAND2_X1   g12097(.A1(new_n12289_), .A2(new_n11941_), .ZN(new_n12290_));
  NAND2_X1   g12098(.A1(new_n12286_), .A2(new_n12288_), .ZN(new_n12291_));
  AOI21_X1   g12099(.A1(new_n12291_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n12292_));
  AOI21_X1   g12100(.A1(new_n12292_), .A2(new_n12290_), .B(new_n12281_), .ZN(new_n12293_));
  AOI21_X1   g12101(.A1(new_n12290_), .A2(new_n12271_), .B(new_n1088_), .ZN(new_n12294_));
  OAI21_X1   g12102(.A1(new_n12293_), .A2(new_n12294_), .B(\asqrt[52] ), .ZN(new_n12295_));
  AOI21_X1   g12103(.A1(new_n12277_), .A2(new_n12295_), .B(new_n842_), .ZN(new_n12296_));
  NOR2_X1    g12104(.A1(new_n12280_), .A2(new_n12296_), .ZN(new_n12297_));
  AOI21_X1   g12105(.A1(new_n12297_), .A2(new_n720_), .B(new_n11930_), .ZN(new_n12298_));
  OAI21_X1   g12106(.A1(new_n12280_), .A2(new_n12296_), .B(\asqrt[54] ), .ZN(new_n12299_));
  NAND2_X1   g12107(.A1(new_n12299_), .A2(new_n630_), .ZN(new_n12300_));
  OAI21_X1   g12108(.A1(new_n12298_), .A2(new_n12300_), .B(new_n11926_), .ZN(new_n12301_));
  INV_X1     g12109(.I(new_n12299_), .ZN(new_n12302_));
  OAI21_X1   g12110(.A1(new_n12298_), .A2(new_n12302_), .B(\asqrt[55] ), .ZN(new_n12303_));
  NAND3_X1   g12111(.A1(new_n12301_), .A2(new_n12303_), .A3(new_n545_), .ZN(new_n12304_));
  NAND2_X1   g12112(.A1(new_n12304_), .A2(new_n11924_), .ZN(new_n12305_));
  NAND2_X1   g12113(.A1(new_n12301_), .A2(new_n12303_), .ZN(new_n12306_));
  AOI21_X1   g12114(.A1(new_n12306_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n12307_));
  AOI21_X1   g12115(.A1(new_n12307_), .A2(new_n12305_), .B(new_n11921_), .ZN(new_n12308_));
  INV_X1     g12116(.I(new_n11926_), .ZN(new_n12309_));
  INV_X1     g12117(.I(new_n11936_), .ZN(new_n12310_));
  NOR2_X1    g12118(.A1(new_n12293_), .A2(new_n12294_), .ZN(new_n12311_));
  AOI21_X1   g12119(.A1(new_n12311_), .A2(new_n962_), .B(new_n12310_), .ZN(new_n12312_));
  NAND2_X1   g12120(.A1(new_n12295_), .A2(new_n842_), .ZN(new_n12313_));
  OAI21_X1   g12121(.A1(new_n12312_), .A2(new_n12313_), .B(new_n11932_), .ZN(new_n12314_));
  INV_X1     g12122(.I(new_n12295_), .ZN(new_n12315_));
  OAI21_X1   g12123(.A1(new_n12312_), .A2(new_n12315_), .B(\asqrt[53] ), .ZN(new_n12316_));
  NAND3_X1   g12124(.A1(new_n12314_), .A2(new_n12316_), .A3(new_n720_), .ZN(new_n12317_));
  NAND2_X1   g12125(.A1(new_n12317_), .A2(new_n11929_), .ZN(new_n12318_));
  NAND2_X1   g12126(.A1(new_n12314_), .A2(new_n12316_), .ZN(new_n12319_));
  AOI21_X1   g12127(.A1(new_n12319_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n12320_));
  AOI21_X1   g12128(.A1(new_n12320_), .A2(new_n12318_), .B(new_n12309_), .ZN(new_n12321_));
  AOI21_X1   g12129(.A1(new_n12318_), .A2(new_n12299_), .B(new_n630_), .ZN(new_n12322_));
  OAI21_X1   g12130(.A1(new_n12321_), .A2(new_n12322_), .B(\asqrt[56] ), .ZN(new_n12323_));
  AOI21_X1   g12131(.A1(new_n12305_), .A2(new_n12323_), .B(new_n450_), .ZN(new_n12324_));
  NOR2_X1    g12132(.A1(new_n12308_), .A2(new_n12324_), .ZN(new_n12325_));
  AOI21_X1   g12133(.A1(new_n12325_), .A2(new_n403_), .B(new_n11918_), .ZN(new_n12326_));
  OAI21_X1   g12134(.A1(new_n12308_), .A2(new_n12324_), .B(\asqrt[58] ), .ZN(new_n12327_));
  NAND2_X1   g12135(.A1(new_n12327_), .A2(new_n339_), .ZN(new_n12328_));
  OAI21_X1   g12136(.A1(new_n12326_), .A2(new_n12328_), .B(new_n11914_), .ZN(new_n12329_));
  INV_X1     g12137(.I(new_n12327_), .ZN(new_n12330_));
  OAI21_X1   g12138(.A1(new_n12326_), .A2(new_n12330_), .B(\asqrt[59] ), .ZN(new_n12331_));
  NAND3_X1   g12139(.A1(new_n12329_), .A2(new_n12331_), .A3(new_n288_), .ZN(new_n12332_));
  NAND2_X1   g12140(.A1(new_n12332_), .A2(new_n11912_), .ZN(new_n12333_));
  INV_X1     g12141(.I(new_n11914_), .ZN(new_n12334_));
  INV_X1     g12142(.I(new_n11924_), .ZN(new_n12335_));
  NOR2_X1    g12143(.A1(new_n12321_), .A2(new_n12322_), .ZN(new_n12336_));
  AOI21_X1   g12144(.A1(new_n12336_), .A2(new_n545_), .B(new_n12335_), .ZN(new_n12337_));
  NAND2_X1   g12145(.A1(new_n12323_), .A2(new_n450_), .ZN(new_n12338_));
  OAI21_X1   g12146(.A1(new_n12337_), .A2(new_n12338_), .B(new_n11920_), .ZN(new_n12339_));
  INV_X1     g12147(.I(new_n12323_), .ZN(new_n12340_));
  OAI21_X1   g12148(.A1(new_n12337_), .A2(new_n12340_), .B(\asqrt[57] ), .ZN(new_n12341_));
  NAND3_X1   g12149(.A1(new_n12339_), .A2(new_n12341_), .A3(new_n403_), .ZN(new_n12342_));
  NAND2_X1   g12150(.A1(new_n12342_), .A2(new_n11917_), .ZN(new_n12343_));
  NAND2_X1   g12151(.A1(new_n12339_), .A2(new_n12341_), .ZN(new_n12344_));
  AOI21_X1   g12152(.A1(new_n12344_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n12345_));
  AOI21_X1   g12153(.A1(new_n12345_), .A2(new_n12343_), .B(new_n12334_), .ZN(new_n12346_));
  AOI21_X1   g12154(.A1(new_n12343_), .A2(new_n12327_), .B(new_n339_), .ZN(new_n12347_));
  OAI21_X1   g12155(.A1(new_n12346_), .A2(new_n12347_), .B(\asqrt[60] ), .ZN(new_n12348_));
  AOI21_X1   g12156(.A1(new_n12333_), .A2(new_n12348_), .B(new_n242_), .ZN(new_n12349_));
  NAND3_X1   g12157(.A1(\asqrt[16] ), .A2(new_n11844_), .A3(new_n11860_), .ZN(new_n12350_));
  XOR2_X1    g12158(.A1(new_n12350_), .A2(new_n11885_), .Z(new_n12351_));
  INV_X1     g12159(.I(new_n12351_), .ZN(new_n12352_));
  NAND2_X1   g12160(.A1(new_n12329_), .A2(new_n12331_), .ZN(new_n12353_));
  AOI21_X1   g12161(.A1(new_n12353_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n12354_));
  AOI21_X1   g12162(.A1(new_n12354_), .A2(new_n12333_), .B(new_n12352_), .ZN(new_n12355_));
  OAI21_X1   g12163(.A1(new_n12355_), .A2(new_n12349_), .B(\asqrt[62] ), .ZN(new_n12356_));
  AOI21_X1   g12164(.A1(new_n11845_), .A2(new_n11866_), .B(new_n11861_), .ZN(new_n12357_));
  NAND2_X1   g12165(.A1(\asqrt[16] ), .A2(new_n12357_), .ZN(new_n12358_));
  XOR2_X1    g12166(.A1(new_n12358_), .A2(new_n11864_), .Z(new_n12359_));
  INV_X1     g12167(.I(new_n11912_), .ZN(new_n12360_));
  NOR2_X1    g12168(.A1(new_n12346_), .A2(new_n12347_), .ZN(new_n12361_));
  AOI21_X1   g12169(.A1(new_n12361_), .A2(new_n288_), .B(new_n12360_), .ZN(new_n12362_));
  INV_X1     g12170(.I(new_n12348_), .ZN(new_n12363_));
  OAI21_X1   g12171(.A1(new_n12362_), .A2(new_n12363_), .B(\asqrt[61] ), .ZN(new_n12364_));
  NAND2_X1   g12172(.A1(new_n12348_), .A2(new_n242_), .ZN(new_n12365_));
  OAI21_X1   g12173(.A1(new_n12362_), .A2(new_n12365_), .B(new_n12351_), .ZN(new_n12366_));
  NAND3_X1   g12174(.A1(new_n12366_), .A2(new_n12364_), .A3(new_n234_), .ZN(new_n12367_));
  NAND2_X1   g12175(.A1(new_n12367_), .A2(new_n12359_), .ZN(new_n12368_));
  AOI21_X1   g12176(.A1(new_n12368_), .A2(new_n12356_), .B(new_n11909_), .ZN(new_n12369_));
  AOI21_X1   g12177(.A1(new_n12369_), .A2(new_n11907_), .B(\asqrt[63] ), .ZN(new_n12370_));
  NAND2_X1   g12178(.A1(new_n12368_), .A2(new_n12356_), .ZN(new_n12371_));
  NOR2_X1    g12179(.A1(new_n12371_), .A2(new_n11907_), .ZN(new_n12372_));
  NOR2_X1    g12180(.A1(\asqrt[16] ), .A2(new_n11896_), .ZN(new_n12373_));
  NOR4_X1    g12181(.A1(new_n12370_), .A2(new_n11904_), .A3(new_n12372_), .A4(new_n12373_), .ZN(new_n12374_));
  OAI21_X1   g12182(.A1(new_n12284_), .A2(new_n12285_), .B(new_n12288_), .ZN(new_n12375_));
  NOR2_X1    g12183(.A1(new_n12374_), .A2(new_n12375_), .ZN(new_n12376_));
  XOR2_X1    g12184(.A1(new_n12376_), .A2(new_n11884_), .Z(new_n12377_));
  INV_X1     g12185(.I(new_n12377_), .ZN(new_n12378_));
  INV_X1     g12186(.I(new_n11904_), .ZN(new_n12379_));
  INV_X1     g12187(.I(new_n12356_), .ZN(new_n12380_));
  NOR2_X1    g12188(.A1(new_n12355_), .A2(new_n12349_), .ZN(new_n12381_));
  INV_X1     g12189(.I(new_n12359_), .ZN(new_n12382_));
  AOI21_X1   g12190(.A1(new_n12381_), .A2(new_n234_), .B(new_n12382_), .ZN(new_n12383_));
  OAI21_X1   g12191(.A1(new_n12383_), .A2(new_n12380_), .B(new_n11908_), .ZN(new_n12384_));
  OAI21_X1   g12192(.A1(new_n12384_), .A2(new_n11906_), .B(new_n193_), .ZN(new_n12385_));
  NOR2_X1    g12193(.A1(new_n12383_), .A2(new_n12380_), .ZN(new_n12386_));
  NAND2_X1   g12194(.A1(new_n12386_), .A2(new_n11906_), .ZN(new_n12387_));
  INV_X1     g12195(.I(new_n12373_), .ZN(new_n12388_));
  NAND4_X1   g12196(.A1(new_n12385_), .A2(new_n12379_), .A3(new_n12387_), .A4(new_n12388_), .ZN(\asqrt[15] ));
  NAND3_X1   g12197(.A1(\asqrt[15] ), .A2(new_n12248_), .A3(new_n12267_), .ZN(new_n12390_));
  XOR2_X1    g12198(.A1(new_n12390_), .A2(new_n12282_), .Z(new_n12391_));
  OAI21_X1   g12199(.A1(new_n12242_), .A2(new_n12244_), .B(new_n12247_), .ZN(new_n12392_));
  NOR2_X1    g12200(.A1(new_n12374_), .A2(new_n12392_), .ZN(new_n12393_));
  XOR2_X1    g12201(.A1(new_n12393_), .A2(new_n11948_), .Z(new_n12394_));
  INV_X1     g12202(.I(new_n12394_), .ZN(new_n12395_));
  NAND3_X1   g12203(.A1(\asqrt[15] ), .A2(new_n12261_), .A3(new_n12243_), .ZN(new_n12396_));
  XOR2_X1    g12204(.A1(new_n12396_), .A2(new_n11952_), .Z(new_n12397_));
  INV_X1     g12205(.I(new_n12397_), .ZN(new_n12398_));
  OAI21_X1   g12206(.A1(new_n12256_), .A2(new_n12257_), .B(new_n12260_), .ZN(new_n12399_));
  NOR2_X1    g12207(.A1(new_n12374_), .A2(new_n12399_), .ZN(new_n12400_));
  XOR2_X1    g12208(.A1(new_n12400_), .A2(new_n11954_), .Z(new_n12401_));
  NAND3_X1   g12209(.A1(\asqrt[15] ), .A2(new_n12220_), .A3(new_n12239_), .ZN(new_n12402_));
  XOR2_X1    g12210(.A1(new_n12402_), .A2(new_n12254_), .Z(new_n12403_));
  OAI21_X1   g12211(.A1(new_n12214_), .A2(new_n12216_), .B(new_n12219_), .ZN(new_n12404_));
  NOR2_X1    g12212(.A1(new_n12374_), .A2(new_n12404_), .ZN(new_n12405_));
  XOR2_X1    g12213(.A1(new_n12405_), .A2(new_n11960_), .Z(new_n12406_));
  INV_X1     g12214(.I(new_n12406_), .ZN(new_n12407_));
  NAND3_X1   g12215(.A1(\asqrt[15] ), .A2(new_n12233_), .A3(new_n12215_), .ZN(new_n12408_));
  XOR2_X1    g12216(.A1(new_n12408_), .A2(new_n11964_), .Z(new_n12409_));
  INV_X1     g12217(.I(new_n12409_), .ZN(new_n12410_));
  OAI21_X1   g12218(.A1(new_n12228_), .A2(new_n12229_), .B(new_n12232_), .ZN(new_n12411_));
  NOR2_X1    g12219(.A1(new_n12374_), .A2(new_n12411_), .ZN(new_n12412_));
  XOR2_X1    g12220(.A1(new_n12412_), .A2(new_n11966_), .Z(new_n12413_));
  NAND3_X1   g12221(.A1(\asqrt[15] ), .A2(new_n12192_), .A3(new_n12211_), .ZN(new_n12414_));
  XOR2_X1    g12222(.A1(new_n12414_), .A2(new_n12226_), .Z(new_n12415_));
  OAI21_X1   g12223(.A1(new_n12186_), .A2(new_n12188_), .B(new_n12191_), .ZN(new_n12416_));
  NOR2_X1    g12224(.A1(new_n12374_), .A2(new_n12416_), .ZN(new_n12417_));
  XOR2_X1    g12225(.A1(new_n12417_), .A2(new_n11972_), .Z(new_n12418_));
  INV_X1     g12226(.I(new_n12418_), .ZN(new_n12419_));
  NAND3_X1   g12227(.A1(\asqrt[15] ), .A2(new_n12205_), .A3(new_n12187_), .ZN(new_n12420_));
  XOR2_X1    g12228(.A1(new_n12420_), .A2(new_n11976_), .Z(new_n12421_));
  INV_X1     g12229(.I(new_n12421_), .ZN(new_n12422_));
  OAI21_X1   g12230(.A1(new_n12200_), .A2(new_n12201_), .B(new_n12204_), .ZN(new_n12423_));
  NOR2_X1    g12231(.A1(new_n12374_), .A2(new_n12423_), .ZN(new_n12424_));
  XOR2_X1    g12232(.A1(new_n12424_), .A2(new_n11978_), .Z(new_n12425_));
  NAND3_X1   g12233(.A1(\asqrt[15] ), .A2(new_n12164_), .A3(new_n12183_), .ZN(new_n12426_));
  XOR2_X1    g12234(.A1(new_n12426_), .A2(new_n12198_), .Z(new_n12427_));
  OAI21_X1   g12235(.A1(new_n12158_), .A2(new_n12160_), .B(new_n12163_), .ZN(new_n12428_));
  NOR2_X1    g12236(.A1(new_n12374_), .A2(new_n12428_), .ZN(new_n12429_));
  XOR2_X1    g12237(.A1(new_n12429_), .A2(new_n11984_), .Z(new_n12430_));
  INV_X1     g12238(.I(new_n12430_), .ZN(new_n12431_));
  NAND3_X1   g12239(.A1(\asqrt[15] ), .A2(new_n12177_), .A3(new_n12159_), .ZN(new_n12432_));
  XOR2_X1    g12240(.A1(new_n12432_), .A2(new_n11988_), .Z(new_n12433_));
  INV_X1     g12241(.I(new_n12433_), .ZN(new_n12434_));
  OAI21_X1   g12242(.A1(new_n12172_), .A2(new_n12173_), .B(new_n12176_), .ZN(new_n12435_));
  NOR2_X1    g12243(.A1(new_n12374_), .A2(new_n12435_), .ZN(new_n12436_));
  XOR2_X1    g12244(.A1(new_n12436_), .A2(new_n11990_), .Z(new_n12437_));
  NAND3_X1   g12245(.A1(\asqrt[15] ), .A2(new_n12136_), .A3(new_n12155_), .ZN(new_n12438_));
  XOR2_X1    g12246(.A1(new_n12438_), .A2(new_n12170_), .Z(new_n12439_));
  OAI21_X1   g12247(.A1(new_n12130_), .A2(new_n12132_), .B(new_n12135_), .ZN(new_n12440_));
  NOR2_X1    g12248(.A1(new_n12374_), .A2(new_n12440_), .ZN(new_n12441_));
  XOR2_X1    g12249(.A1(new_n12441_), .A2(new_n11996_), .Z(new_n12442_));
  INV_X1     g12250(.I(new_n12442_), .ZN(new_n12443_));
  NAND3_X1   g12251(.A1(\asqrt[15] ), .A2(new_n12149_), .A3(new_n12131_), .ZN(new_n12444_));
  XOR2_X1    g12252(.A1(new_n12444_), .A2(new_n12000_), .Z(new_n12445_));
  INV_X1     g12253(.I(new_n12445_), .ZN(new_n12446_));
  OAI21_X1   g12254(.A1(new_n12144_), .A2(new_n12145_), .B(new_n12148_), .ZN(new_n12447_));
  NOR2_X1    g12255(.A1(new_n12374_), .A2(new_n12447_), .ZN(new_n12448_));
  XOR2_X1    g12256(.A1(new_n12448_), .A2(new_n12002_), .Z(new_n12449_));
  NAND3_X1   g12257(.A1(\asqrt[15] ), .A2(new_n12108_), .A3(new_n12127_), .ZN(new_n12450_));
  XOR2_X1    g12258(.A1(new_n12450_), .A2(new_n12142_), .Z(new_n12451_));
  OAI21_X1   g12259(.A1(new_n12102_), .A2(new_n12104_), .B(new_n12107_), .ZN(new_n12452_));
  NOR2_X1    g12260(.A1(new_n12374_), .A2(new_n12452_), .ZN(new_n12453_));
  XOR2_X1    g12261(.A1(new_n12453_), .A2(new_n12008_), .Z(new_n12454_));
  INV_X1     g12262(.I(new_n12454_), .ZN(new_n12455_));
  NAND3_X1   g12263(.A1(\asqrt[15] ), .A2(new_n12121_), .A3(new_n12103_), .ZN(new_n12456_));
  XOR2_X1    g12264(.A1(new_n12456_), .A2(new_n12012_), .Z(new_n12457_));
  INV_X1     g12265(.I(new_n12457_), .ZN(new_n12458_));
  OAI21_X1   g12266(.A1(new_n12116_), .A2(new_n12117_), .B(new_n12120_), .ZN(new_n12459_));
  NOR2_X1    g12267(.A1(new_n12374_), .A2(new_n12459_), .ZN(new_n12460_));
  XOR2_X1    g12268(.A1(new_n12460_), .A2(new_n12014_), .Z(new_n12461_));
  NAND3_X1   g12269(.A1(\asqrt[15] ), .A2(new_n12067_), .A3(new_n12099_), .ZN(new_n12462_));
  XOR2_X1    g12270(.A1(new_n12462_), .A2(new_n12114_), .Z(new_n12463_));
  OAI21_X1   g12271(.A1(new_n12061_), .A2(new_n12063_), .B(new_n12066_), .ZN(new_n12464_));
  NOR2_X1    g12272(.A1(new_n12374_), .A2(new_n12464_), .ZN(new_n12465_));
  XOR2_X1    g12273(.A1(new_n12465_), .A2(new_n12020_), .Z(new_n12466_));
  INV_X1     g12274(.I(new_n12466_), .ZN(new_n12467_));
  NAND3_X1   g12275(.A1(\asqrt[15] ), .A2(new_n12093_), .A3(new_n12062_), .ZN(new_n12468_));
  XOR2_X1    g12276(.A1(new_n12468_), .A2(new_n12024_), .Z(new_n12469_));
  INV_X1     g12277(.I(new_n12469_), .ZN(new_n12470_));
  AOI21_X1   g12278(.A1(new_n12055_), .A2(new_n12056_), .B(new_n12059_), .ZN(new_n12471_));
  NAND2_X1   g12279(.A1(\asqrt[15] ), .A2(new_n12471_), .ZN(new_n12472_));
  XOR2_X1    g12280(.A1(new_n12472_), .A2(new_n12027_), .Z(new_n12473_));
  NOR2_X1    g12281(.A1(new_n12054_), .A2(\asqrt[20] ), .ZN(new_n12474_));
  NOR3_X1    g12282(.A1(new_n12374_), .A2(new_n12474_), .A3(new_n12091_), .ZN(new_n12475_));
  XOR2_X1    g12283(.A1(new_n12475_), .A2(new_n12030_), .Z(new_n12476_));
  NOR3_X1    g12284(.A1(new_n12374_), .A2(new_n12049_), .A3(new_n12086_), .ZN(new_n12477_));
  XOR2_X1    g12285(.A1(new_n12477_), .A2(new_n12051_), .Z(new_n12478_));
  INV_X1     g12286(.I(new_n12478_), .ZN(new_n12479_));
  NOR2_X1    g12287(.A1(new_n12082_), .A2(\asqrt[18] ), .ZN(new_n12480_));
  NOR3_X1    g12288(.A1(new_n12374_), .A2(new_n12480_), .A3(new_n12048_), .ZN(new_n12481_));
  XOR2_X1    g12289(.A1(new_n12481_), .A2(new_n12076_), .Z(new_n12482_));
  INV_X1     g12290(.I(new_n12482_), .ZN(new_n12483_));
  NAND3_X1   g12291(.A1(\asqrt[15] ), .A2(new_n12038_), .A3(new_n12039_), .ZN(new_n12484_));
  NAND4_X1   g12292(.A1(new_n12385_), .A2(\asqrt[16] ), .A3(new_n12387_), .A4(new_n12379_), .ZN(new_n12485_));
  AOI21_X1   g12293(.A1(new_n12484_), .A2(new_n12485_), .B(\a[32] ), .ZN(new_n12486_));
  NOR3_X1    g12294(.A1(new_n12374_), .A2(\a[30] ), .A3(\a[31] ), .ZN(new_n12487_));
  INV_X1     g12295(.I(new_n12485_), .ZN(new_n12488_));
  NOR3_X1    g12296(.A1(new_n12487_), .A2(new_n11511_), .A3(new_n12488_), .ZN(new_n12489_));
  NOR2_X1    g12297(.A1(new_n12489_), .A2(new_n12486_), .ZN(new_n12490_));
  INV_X1     g12298(.I(\a[28] ), .ZN(new_n12491_));
  INV_X1     g12299(.I(\a[29] ), .ZN(new_n12492_));
  NAND3_X1   g12300(.A1(new_n12491_), .A2(new_n12492_), .A3(new_n12038_), .ZN(new_n12493_));
  OAI21_X1   g12301(.A1(new_n12374_), .A2(new_n12038_), .B(new_n12493_), .ZN(new_n12494_));
  NAND2_X1   g12302(.A1(new_n12494_), .A2(\asqrt[16] ), .ZN(new_n12495_));
  OAI21_X1   g12303(.A1(new_n12374_), .A2(\a[30] ), .B(\a[31] ), .ZN(new_n12496_));
  NAND2_X1   g12304(.A1(new_n12496_), .A2(new_n12484_), .ZN(new_n12497_));
  NOR2_X1    g12305(.A1(new_n12494_), .A2(\asqrt[16] ), .ZN(new_n12498_));
  OAI21_X1   g12306(.A1(new_n12497_), .A2(new_n12498_), .B(new_n12495_), .ZN(new_n12499_));
  OAI21_X1   g12307(.A1(new_n12499_), .A2(\asqrt[17] ), .B(new_n12490_), .ZN(new_n12500_));
  NAND2_X1   g12308(.A1(new_n12499_), .A2(\asqrt[17] ), .ZN(new_n12501_));
  NAND3_X1   g12309(.A1(new_n12500_), .A2(new_n10953_), .A3(new_n12501_), .ZN(new_n12502_));
  NOR3_X1    g12310(.A1(new_n12374_), .A2(new_n12042_), .A3(new_n12081_), .ZN(new_n12503_));
  XOR2_X1    g12311(.A1(new_n12503_), .A2(new_n12044_), .Z(new_n12504_));
  NAND2_X1   g12312(.A1(new_n12502_), .A2(new_n12504_), .ZN(new_n12505_));
  NAND2_X1   g12313(.A1(new_n12500_), .A2(new_n12501_), .ZN(new_n12506_));
  AOI21_X1   g12314(.A1(new_n12506_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n12507_));
  AOI21_X1   g12315(.A1(new_n12507_), .A2(new_n12505_), .B(new_n12483_), .ZN(new_n12508_));
  OAI21_X1   g12316(.A1(new_n12487_), .A2(new_n12488_), .B(new_n11511_), .ZN(new_n12509_));
  NAND3_X1   g12317(.A1(new_n12484_), .A2(\a[32] ), .A3(new_n12485_), .ZN(new_n12510_));
  NAND2_X1   g12318(.A1(new_n12509_), .A2(new_n12510_), .ZN(new_n12511_));
  NAND2_X1   g12319(.A1(\asqrt[15] ), .A2(\a[30] ), .ZN(new_n12512_));
  AOI21_X1   g12320(.A1(new_n12512_), .A2(new_n12493_), .B(new_n11901_), .ZN(new_n12513_));
  AOI21_X1   g12321(.A1(\asqrt[15] ), .A2(new_n12038_), .B(new_n12039_), .ZN(new_n12514_));
  NOR2_X1    g12322(.A1(new_n12487_), .A2(new_n12514_), .ZN(new_n12515_));
  NAND3_X1   g12323(.A1(new_n12512_), .A2(new_n11901_), .A3(new_n12493_), .ZN(new_n12516_));
  AOI21_X1   g12324(.A1(new_n12515_), .A2(new_n12516_), .B(new_n12513_), .ZN(new_n12517_));
  AOI21_X1   g12325(.A1(new_n12517_), .A2(new_n11406_), .B(new_n12511_), .ZN(new_n12518_));
  NOR2_X1    g12326(.A1(new_n12517_), .A2(new_n11406_), .ZN(new_n12519_));
  OAI21_X1   g12327(.A1(new_n12518_), .A2(new_n12519_), .B(\asqrt[18] ), .ZN(new_n12520_));
  AOI21_X1   g12328(.A1(new_n12505_), .A2(new_n12520_), .B(new_n10478_), .ZN(new_n12521_));
  NOR2_X1    g12329(.A1(new_n12508_), .A2(new_n12521_), .ZN(new_n12522_));
  AOI21_X1   g12330(.A1(new_n12522_), .A2(new_n10045_), .B(new_n12479_), .ZN(new_n12523_));
  OAI21_X1   g12331(.A1(new_n12508_), .A2(new_n12521_), .B(\asqrt[20] ), .ZN(new_n12524_));
  NAND2_X1   g12332(.A1(new_n12524_), .A2(new_n9590_), .ZN(new_n12525_));
  OAI21_X1   g12333(.A1(new_n12523_), .A2(new_n12525_), .B(new_n12476_), .ZN(new_n12526_));
  INV_X1     g12334(.I(new_n12524_), .ZN(new_n12527_));
  OAI21_X1   g12335(.A1(new_n12523_), .A2(new_n12527_), .B(\asqrt[21] ), .ZN(new_n12528_));
  NAND3_X1   g12336(.A1(new_n12526_), .A2(new_n12528_), .A3(new_n9177_), .ZN(new_n12529_));
  NAND2_X1   g12337(.A1(new_n12529_), .A2(new_n12473_), .ZN(new_n12530_));
  NAND2_X1   g12338(.A1(new_n12526_), .A2(new_n12528_), .ZN(new_n12531_));
  AOI21_X1   g12339(.A1(new_n12531_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n12532_));
  AOI21_X1   g12340(.A1(new_n12532_), .A2(new_n12530_), .B(new_n12470_), .ZN(new_n12533_));
  INV_X1     g12341(.I(new_n12476_), .ZN(new_n12534_));
  NOR2_X1    g12342(.A1(new_n12518_), .A2(new_n12519_), .ZN(new_n12535_));
  INV_X1     g12343(.I(new_n12504_), .ZN(new_n12536_));
  AOI21_X1   g12344(.A1(new_n12535_), .A2(new_n10953_), .B(new_n12536_), .ZN(new_n12537_));
  NAND2_X1   g12345(.A1(new_n12520_), .A2(new_n10478_), .ZN(new_n12538_));
  OAI21_X1   g12346(.A1(new_n12537_), .A2(new_n12538_), .B(new_n12482_), .ZN(new_n12539_));
  INV_X1     g12347(.I(new_n12520_), .ZN(new_n12540_));
  OAI21_X1   g12348(.A1(new_n12537_), .A2(new_n12540_), .B(\asqrt[19] ), .ZN(new_n12541_));
  NAND3_X1   g12349(.A1(new_n12539_), .A2(new_n12541_), .A3(new_n10045_), .ZN(new_n12542_));
  NAND2_X1   g12350(.A1(new_n12542_), .A2(new_n12478_), .ZN(new_n12543_));
  NAND2_X1   g12351(.A1(new_n12539_), .A2(new_n12541_), .ZN(new_n12544_));
  AOI21_X1   g12352(.A1(new_n12544_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n12545_));
  AOI21_X1   g12353(.A1(new_n12545_), .A2(new_n12543_), .B(new_n12534_), .ZN(new_n12546_));
  AOI21_X1   g12354(.A1(new_n12543_), .A2(new_n12524_), .B(new_n9590_), .ZN(new_n12547_));
  OAI21_X1   g12355(.A1(new_n12546_), .A2(new_n12547_), .B(\asqrt[22] ), .ZN(new_n12548_));
  AOI21_X1   g12356(.A1(new_n12530_), .A2(new_n12548_), .B(new_n8742_), .ZN(new_n12549_));
  NOR2_X1    g12357(.A1(new_n12533_), .A2(new_n12549_), .ZN(new_n12550_));
  AOI21_X1   g12358(.A1(new_n12550_), .A2(new_n8349_), .B(new_n12467_), .ZN(new_n12551_));
  OAI21_X1   g12359(.A1(new_n12533_), .A2(new_n12549_), .B(\asqrt[24] ), .ZN(new_n12552_));
  NAND2_X1   g12360(.A1(new_n12552_), .A2(new_n7934_), .ZN(new_n12553_));
  OAI21_X1   g12361(.A1(new_n12551_), .A2(new_n12553_), .B(new_n12463_), .ZN(new_n12554_));
  INV_X1     g12362(.I(new_n12552_), .ZN(new_n12555_));
  OAI21_X1   g12363(.A1(new_n12551_), .A2(new_n12555_), .B(\asqrt[25] ), .ZN(new_n12556_));
  NAND3_X1   g12364(.A1(new_n12554_), .A2(new_n12556_), .A3(new_n7561_), .ZN(new_n12557_));
  NAND2_X1   g12365(.A1(new_n12557_), .A2(new_n12461_), .ZN(new_n12558_));
  NAND2_X1   g12366(.A1(new_n12554_), .A2(new_n12556_), .ZN(new_n12559_));
  AOI21_X1   g12367(.A1(new_n12559_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n12560_));
  AOI21_X1   g12368(.A1(new_n12560_), .A2(new_n12558_), .B(new_n12458_), .ZN(new_n12561_));
  INV_X1     g12369(.I(new_n12463_), .ZN(new_n12562_));
  INV_X1     g12370(.I(new_n12473_), .ZN(new_n12563_));
  NOR2_X1    g12371(.A1(new_n12546_), .A2(new_n12547_), .ZN(new_n12564_));
  AOI21_X1   g12372(.A1(new_n12564_), .A2(new_n9177_), .B(new_n12563_), .ZN(new_n12565_));
  NAND2_X1   g12373(.A1(new_n12548_), .A2(new_n8742_), .ZN(new_n12566_));
  OAI21_X1   g12374(.A1(new_n12565_), .A2(new_n12566_), .B(new_n12469_), .ZN(new_n12567_));
  INV_X1     g12375(.I(new_n12548_), .ZN(new_n12568_));
  OAI21_X1   g12376(.A1(new_n12565_), .A2(new_n12568_), .B(\asqrt[23] ), .ZN(new_n12569_));
  NAND3_X1   g12377(.A1(new_n12567_), .A2(new_n12569_), .A3(new_n8349_), .ZN(new_n12570_));
  NAND2_X1   g12378(.A1(new_n12570_), .A2(new_n12466_), .ZN(new_n12571_));
  NAND2_X1   g12379(.A1(new_n12567_), .A2(new_n12569_), .ZN(new_n12572_));
  AOI21_X1   g12380(.A1(new_n12572_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n12573_));
  AOI21_X1   g12381(.A1(new_n12573_), .A2(new_n12571_), .B(new_n12562_), .ZN(new_n12574_));
  AOI21_X1   g12382(.A1(new_n12571_), .A2(new_n12552_), .B(new_n7934_), .ZN(new_n12575_));
  OAI21_X1   g12383(.A1(new_n12574_), .A2(new_n12575_), .B(\asqrt[26] ), .ZN(new_n12576_));
  AOI21_X1   g12384(.A1(new_n12558_), .A2(new_n12576_), .B(new_n7166_), .ZN(new_n12577_));
  NOR2_X1    g12385(.A1(new_n12561_), .A2(new_n12577_), .ZN(new_n12578_));
  AOI21_X1   g12386(.A1(new_n12578_), .A2(new_n6813_), .B(new_n12455_), .ZN(new_n12579_));
  OAI21_X1   g12387(.A1(new_n12561_), .A2(new_n12577_), .B(\asqrt[28] ), .ZN(new_n12580_));
  NAND2_X1   g12388(.A1(new_n12580_), .A2(new_n6454_), .ZN(new_n12581_));
  OAI21_X1   g12389(.A1(new_n12579_), .A2(new_n12581_), .B(new_n12451_), .ZN(new_n12582_));
  INV_X1     g12390(.I(new_n12580_), .ZN(new_n12583_));
  OAI21_X1   g12391(.A1(new_n12579_), .A2(new_n12583_), .B(\asqrt[29] ), .ZN(new_n12584_));
  NAND3_X1   g12392(.A1(new_n12582_), .A2(new_n12584_), .A3(new_n6106_), .ZN(new_n12585_));
  NAND2_X1   g12393(.A1(new_n12585_), .A2(new_n12449_), .ZN(new_n12586_));
  NAND2_X1   g12394(.A1(new_n12582_), .A2(new_n12584_), .ZN(new_n12587_));
  AOI21_X1   g12395(.A1(new_n12587_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n12588_));
  AOI21_X1   g12396(.A1(new_n12588_), .A2(new_n12586_), .B(new_n12446_), .ZN(new_n12589_));
  INV_X1     g12397(.I(new_n12451_), .ZN(new_n12590_));
  INV_X1     g12398(.I(new_n12461_), .ZN(new_n12591_));
  NOR2_X1    g12399(.A1(new_n12574_), .A2(new_n12575_), .ZN(new_n12592_));
  AOI21_X1   g12400(.A1(new_n12592_), .A2(new_n7561_), .B(new_n12591_), .ZN(new_n12593_));
  NAND2_X1   g12401(.A1(new_n12576_), .A2(new_n7166_), .ZN(new_n12594_));
  OAI21_X1   g12402(.A1(new_n12593_), .A2(new_n12594_), .B(new_n12457_), .ZN(new_n12595_));
  INV_X1     g12403(.I(new_n12576_), .ZN(new_n12596_));
  OAI21_X1   g12404(.A1(new_n12593_), .A2(new_n12596_), .B(\asqrt[27] ), .ZN(new_n12597_));
  NAND3_X1   g12405(.A1(new_n12595_), .A2(new_n12597_), .A3(new_n6813_), .ZN(new_n12598_));
  NAND2_X1   g12406(.A1(new_n12598_), .A2(new_n12454_), .ZN(new_n12599_));
  NAND2_X1   g12407(.A1(new_n12595_), .A2(new_n12597_), .ZN(new_n12600_));
  AOI21_X1   g12408(.A1(new_n12600_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n12601_));
  AOI21_X1   g12409(.A1(new_n12601_), .A2(new_n12599_), .B(new_n12590_), .ZN(new_n12602_));
  AOI21_X1   g12410(.A1(new_n12599_), .A2(new_n12580_), .B(new_n6454_), .ZN(new_n12603_));
  OAI21_X1   g12411(.A1(new_n12602_), .A2(new_n12603_), .B(\asqrt[30] ), .ZN(new_n12604_));
  AOI21_X1   g12412(.A1(new_n12586_), .A2(new_n12604_), .B(new_n5750_), .ZN(new_n12605_));
  NOR2_X1    g12413(.A1(new_n12589_), .A2(new_n12605_), .ZN(new_n12606_));
  AOI21_X1   g12414(.A1(new_n12606_), .A2(new_n5435_), .B(new_n12443_), .ZN(new_n12607_));
  OAI21_X1   g12415(.A1(new_n12589_), .A2(new_n12605_), .B(\asqrt[32] ), .ZN(new_n12608_));
  NAND2_X1   g12416(.A1(new_n12608_), .A2(new_n5110_), .ZN(new_n12609_));
  OAI21_X1   g12417(.A1(new_n12607_), .A2(new_n12609_), .B(new_n12439_), .ZN(new_n12610_));
  INV_X1     g12418(.I(new_n12608_), .ZN(new_n12611_));
  OAI21_X1   g12419(.A1(new_n12607_), .A2(new_n12611_), .B(\asqrt[33] ), .ZN(new_n12612_));
  NAND3_X1   g12420(.A1(new_n12610_), .A2(new_n12612_), .A3(new_n4810_), .ZN(new_n12613_));
  NAND2_X1   g12421(.A1(new_n12613_), .A2(new_n12437_), .ZN(new_n12614_));
  NAND2_X1   g12422(.A1(new_n12610_), .A2(new_n12612_), .ZN(new_n12615_));
  AOI21_X1   g12423(.A1(new_n12615_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n12616_));
  AOI21_X1   g12424(.A1(new_n12616_), .A2(new_n12614_), .B(new_n12434_), .ZN(new_n12617_));
  INV_X1     g12425(.I(new_n12439_), .ZN(new_n12618_));
  INV_X1     g12426(.I(new_n12449_), .ZN(new_n12619_));
  NOR2_X1    g12427(.A1(new_n12602_), .A2(new_n12603_), .ZN(new_n12620_));
  AOI21_X1   g12428(.A1(new_n12620_), .A2(new_n6106_), .B(new_n12619_), .ZN(new_n12621_));
  NAND2_X1   g12429(.A1(new_n12604_), .A2(new_n5750_), .ZN(new_n12622_));
  OAI21_X1   g12430(.A1(new_n12621_), .A2(new_n12622_), .B(new_n12445_), .ZN(new_n12623_));
  INV_X1     g12431(.I(new_n12604_), .ZN(new_n12624_));
  OAI21_X1   g12432(.A1(new_n12621_), .A2(new_n12624_), .B(\asqrt[31] ), .ZN(new_n12625_));
  NAND3_X1   g12433(.A1(new_n12623_), .A2(new_n12625_), .A3(new_n5435_), .ZN(new_n12626_));
  NAND2_X1   g12434(.A1(new_n12626_), .A2(new_n12442_), .ZN(new_n12627_));
  NAND2_X1   g12435(.A1(new_n12623_), .A2(new_n12625_), .ZN(new_n12628_));
  AOI21_X1   g12436(.A1(new_n12628_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n12629_));
  AOI21_X1   g12437(.A1(new_n12629_), .A2(new_n12627_), .B(new_n12618_), .ZN(new_n12630_));
  AOI21_X1   g12438(.A1(new_n12627_), .A2(new_n12608_), .B(new_n5110_), .ZN(new_n12631_));
  OAI21_X1   g12439(.A1(new_n12630_), .A2(new_n12631_), .B(\asqrt[34] ), .ZN(new_n12632_));
  AOI21_X1   g12440(.A1(new_n12614_), .A2(new_n12632_), .B(new_n4510_), .ZN(new_n12633_));
  NOR2_X1    g12441(.A1(new_n12617_), .A2(new_n12633_), .ZN(new_n12634_));
  AOI21_X1   g12442(.A1(new_n12634_), .A2(new_n4224_), .B(new_n12431_), .ZN(new_n12635_));
  OAI21_X1   g12443(.A1(new_n12617_), .A2(new_n12633_), .B(\asqrt[36] ), .ZN(new_n12636_));
  NAND2_X1   g12444(.A1(new_n12636_), .A2(new_n3928_), .ZN(new_n12637_));
  OAI21_X1   g12445(.A1(new_n12635_), .A2(new_n12637_), .B(new_n12427_), .ZN(new_n12638_));
  INV_X1     g12446(.I(new_n12636_), .ZN(new_n12639_));
  OAI21_X1   g12447(.A1(new_n12635_), .A2(new_n12639_), .B(\asqrt[37] ), .ZN(new_n12640_));
  NAND3_X1   g12448(.A1(new_n12638_), .A2(new_n12640_), .A3(new_n3675_), .ZN(new_n12641_));
  NAND2_X1   g12449(.A1(new_n12641_), .A2(new_n12425_), .ZN(new_n12642_));
  NAND2_X1   g12450(.A1(new_n12638_), .A2(new_n12640_), .ZN(new_n12643_));
  AOI21_X1   g12451(.A1(new_n12643_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n12644_));
  AOI21_X1   g12452(.A1(new_n12644_), .A2(new_n12642_), .B(new_n12422_), .ZN(new_n12645_));
  INV_X1     g12453(.I(new_n12427_), .ZN(new_n12646_));
  INV_X1     g12454(.I(new_n12437_), .ZN(new_n12647_));
  NOR2_X1    g12455(.A1(new_n12630_), .A2(new_n12631_), .ZN(new_n12648_));
  AOI21_X1   g12456(.A1(new_n12648_), .A2(new_n4810_), .B(new_n12647_), .ZN(new_n12649_));
  NAND2_X1   g12457(.A1(new_n12632_), .A2(new_n4510_), .ZN(new_n12650_));
  OAI21_X1   g12458(.A1(new_n12649_), .A2(new_n12650_), .B(new_n12433_), .ZN(new_n12651_));
  INV_X1     g12459(.I(new_n12632_), .ZN(new_n12652_));
  OAI21_X1   g12460(.A1(new_n12649_), .A2(new_n12652_), .B(\asqrt[35] ), .ZN(new_n12653_));
  NAND3_X1   g12461(.A1(new_n12651_), .A2(new_n12653_), .A3(new_n4224_), .ZN(new_n12654_));
  NAND2_X1   g12462(.A1(new_n12654_), .A2(new_n12430_), .ZN(new_n12655_));
  NAND2_X1   g12463(.A1(new_n12651_), .A2(new_n12653_), .ZN(new_n12656_));
  AOI21_X1   g12464(.A1(new_n12656_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n12657_));
  AOI21_X1   g12465(.A1(new_n12657_), .A2(new_n12655_), .B(new_n12646_), .ZN(new_n12658_));
  AOI21_X1   g12466(.A1(new_n12655_), .A2(new_n12636_), .B(new_n3928_), .ZN(new_n12659_));
  OAI21_X1   g12467(.A1(new_n12658_), .A2(new_n12659_), .B(\asqrt[38] ), .ZN(new_n12660_));
  AOI21_X1   g12468(.A1(new_n12642_), .A2(new_n12660_), .B(new_n3400_), .ZN(new_n12661_));
  NOR2_X1    g12469(.A1(new_n12645_), .A2(new_n12661_), .ZN(new_n12662_));
  AOI21_X1   g12470(.A1(new_n12662_), .A2(new_n3167_), .B(new_n12419_), .ZN(new_n12663_));
  OAI21_X1   g12471(.A1(new_n12645_), .A2(new_n12661_), .B(\asqrt[40] ), .ZN(new_n12664_));
  NAND2_X1   g12472(.A1(new_n12664_), .A2(new_n2912_), .ZN(new_n12665_));
  OAI21_X1   g12473(.A1(new_n12663_), .A2(new_n12665_), .B(new_n12415_), .ZN(new_n12666_));
  INV_X1     g12474(.I(new_n12664_), .ZN(new_n12667_));
  OAI21_X1   g12475(.A1(new_n12663_), .A2(new_n12667_), .B(\asqrt[41] ), .ZN(new_n12668_));
  NAND3_X1   g12476(.A1(new_n12666_), .A2(new_n12668_), .A3(new_n2699_), .ZN(new_n12669_));
  NAND2_X1   g12477(.A1(new_n12669_), .A2(new_n12413_), .ZN(new_n12670_));
  NAND2_X1   g12478(.A1(new_n12666_), .A2(new_n12668_), .ZN(new_n12671_));
  AOI21_X1   g12479(.A1(new_n12671_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n12672_));
  AOI21_X1   g12480(.A1(new_n12672_), .A2(new_n12670_), .B(new_n12410_), .ZN(new_n12673_));
  INV_X1     g12481(.I(new_n12415_), .ZN(new_n12674_));
  INV_X1     g12482(.I(new_n12425_), .ZN(new_n12675_));
  NOR2_X1    g12483(.A1(new_n12658_), .A2(new_n12659_), .ZN(new_n12676_));
  AOI21_X1   g12484(.A1(new_n12676_), .A2(new_n3675_), .B(new_n12675_), .ZN(new_n12677_));
  NAND2_X1   g12485(.A1(new_n12660_), .A2(new_n3400_), .ZN(new_n12678_));
  OAI21_X1   g12486(.A1(new_n12677_), .A2(new_n12678_), .B(new_n12421_), .ZN(new_n12679_));
  INV_X1     g12487(.I(new_n12660_), .ZN(new_n12680_));
  OAI21_X1   g12488(.A1(new_n12677_), .A2(new_n12680_), .B(\asqrt[39] ), .ZN(new_n12681_));
  NAND3_X1   g12489(.A1(new_n12679_), .A2(new_n12681_), .A3(new_n3167_), .ZN(new_n12682_));
  NAND2_X1   g12490(.A1(new_n12682_), .A2(new_n12418_), .ZN(new_n12683_));
  NAND2_X1   g12491(.A1(new_n12679_), .A2(new_n12681_), .ZN(new_n12684_));
  AOI21_X1   g12492(.A1(new_n12684_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n12685_));
  AOI21_X1   g12493(.A1(new_n12685_), .A2(new_n12683_), .B(new_n12674_), .ZN(new_n12686_));
  AOI21_X1   g12494(.A1(new_n12683_), .A2(new_n12664_), .B(new_n2912_), .ZN(new_n12687_));
  OAI21_X1   g12495(.A1(new_n12686_), .A2(new_n12687_), .B(\asqrt[42] ), .ZN(new_n12688_));
  AOI21_X1   g12496(.A1(new_n12670_), .A2(new_n12688_), .B(new_n2464_), .ZN(new_n12689_));
  NOR2_X1    g12497(.A1(new_n12673_), .A2(new_n12689_), .ZN(new_n12690_));
  AOI21_X1   g12498(.A1(new_n12690_), .A2(new_n2271_), .B(new_n12407_), .ZN(new_n12691_));
  OAI21_X1   g12499(.A1(new_n12673_), .A2(new_n12689_), .B(\asqrt[44] ), .ZN(new_n12692_));
  NAND2_X1   g12500(.A1(new_n12692_), .A2(new_n2072_), .ZN(new_n12693_));
  OAI21_X1   g12501(.A1(new_n12691_), .A2(new_n12693_), .B(new_n12403_), .ZN(new_n12694_));
  INV_X1     g12502(.I(new_n12692_), .ZN(new_n12695_));
  OAI21_X1   g12503(.A1(new_n12691_), .A2(new_n12695_), .B(\asqrt[45] ), .ZN(new_n12696_));
  NAND3_X1   g12504(.A1(new_n12694_), .A2(new_n12696_), .A3(new_n1884_), .ZN(new_n12697_));
  NAND2_X1   g12505(.A1(new_n12697_), .A2(new_n12401_), .ZN(new_n12698_));
  NAND2_X1   g12506(.A1(new_n12694_), .A2(new_n12696_), .ZN(new_n12699_));
  AOI21_X1   g12507(.A1(new_n12699_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n12700_));
  AOI21_X1   g12508(.A1(new_n12700_), .A2(new_n12698_), .B(new_n12398_), .ZN(new_n12701_));
  INV_X1     g12509(.I(new_n12403_), .ZN(new_n12702_));
  INV_X1     g12510(.I(new_n12413_), .ZN(new_n12703_));
  NOR2_X1    g12511(.A1(new_n12686_), .A2(new_n12687_), .ZN(new_n12704_));
  AOI21_X1   g12512(.A1(new_n12704_), .A2(new_n2699_), .B(new_n12703_), .ZN(new_n12705_));
  NAND2_X1   g12513(.A1(new_n12688_), .A2(new_n2464_), .ZN(new_n12706_));
  OAI21_X1   g12514(.A1(new_n12705_), .A2(new_n12706_), .B(new_n12409_), .ZN(new_n12707_));
  INV_X1     g12515(.I(new_n12688_), .ZN(new_n12708_));
  OAI21_X1   g12516(.A1(new_n12705_), .A2(new_n12708_), .B(\asqrt[43] ), .ZN(new_n12709_));
  NAND3_X1   g12517(.A1(new_n12707_), .A2(new_n12709_), .A3(new_n2271_), .ZN(new_n12710_));
  NAND2_X1   g12518(.A1(new_n12710_), .A2(new_n12406_), .ZN(new_n12711_));
  NAND2_X1   g12519(.A1(new_n12707_), .A2(new_n12709_), .ZN(new_n12712_));
  AOI21_X1   g12520(.A1(new_n12712_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n12713_));
  AOI21_X1   g12521(.A1(new_n12713_), .A2(new_n12711_), .B(new_n12702_), .ZN(new_n12714_));
  AOI21_X1   g12522(.A1(new_n12711_), .A2(new_n12692_), .B(new_n2072_), .ZN(new_n12715_));
  OAI21_X1   g12523(.A1(new_n12714_), .A2(new_n12715_), .B(\asqrt[46] ), .ZN(new_n12716_));
  AOI21_X1   g12524(.A1(new_n12698_), .A2(new_n12716_), .B(new_n1688_), .ZN(new_n12717_));
  NOR2_X1    g12525(.A1(new_n12701_), .A2(new_n12717_), .ZN(new_n12718_));
  AOI21_X1   g12526(.A1(new_n12718_), .A2(new_n1533_), .B(new_n12395_), .ZN(new_n12719_));
  OAI21_X1   g12527(.A1(new_n12701_), .A2(new_n12717_), .B(\asqrt[48] ), .ZN(new_n12720_));
  NAND2_X1   g12528(.A1(new_n12720_), .A2(new_n1368_), .ZN(new_n12721_));
  OAI21_X1   g12529(.A1(new_n12719_), .A2(new_n12721_), .B(new_n12391_), .ZN(new_n12722_));
  INV_X1     g12530(.I(new_n12720_), .ZN(new_n12723_));
  OAI21_X1   g12531(.A1(new_n12719_), .A2(new_n12723_), .B(\asqrt[49] ), .ZN(new_n12724_));
  NAND3_X1   g12532(.A1(new_n12722_), .A2(new_n12724_), .A3(new_n1228_), .ZN(new_n12725_));
  INV_X1     g12533(.I(new_n12391_), .ZN(new_n12726_));
  INV_X1     g12534(.I(new_n12401_), .ZN(new_n12727_));
  NOR2_X1    g12535(.A1(new_n12714_), .A2(new_n12715_), .ZN(new_n12728_));
  AOI21_X1   g12536(.A1(new_n12728_), .A2(new_n1884_), .B(new_n12727_), .ZN(new_n12729_));
  NAND2_X1   g12537(.A1(new_n12716_), .A2(new_n1688_), .ZN(new_n12730_));
  OAI21_X1   g12538(.A1(new_n12729_), .A2(new_n12730_), .B(new_n12397_), .ZN(new_n12731_));
  INV_X1     g12539(.I(new_n12716_), .ZN(new_n12732_));
  OAI21_X1   g12540(.A1(new_n12729_), .A2(new_n12732_), .B(\asqrt[47] ), .ZN(new_n12733_));
  NAND3_X1   g12541(.A1(new_n12731_), .A2(new_n12733_), .A3(new_n1533_), .ZN(new_n12734_));
  NAND2_X1   g12542(.A1(new_n12734_), .A2(new_n12394_), .ZN(new_n12735_));
  NAND2_X1   g12543(.A1(new_n12731_), .A2(new_n12733_), .ZN(new_n12736_));
  AOI21_X1   g12544(.A1(new_n12736_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n12737_));
  AOI21_X1   g12545(.A1(new_n12737_), .A2(new_n12735_), .B(new_n12726_), .ZN(new_n12738_));
  AOI21_X1   g12546(.A1(new_n12735_), .A2(new_n12720_), .B(new_n1368_), .ZN(new_n12739_));
  OAI21_X1   g12547(.A1(new_n12738_), .A2(new_n12739_), .B(\asqrt[50] ), .ZN(new_n12740_));
  NAND2_X1   g12548(.A1(new_n12371_), .A2(new_n11906_), .ZN(new_n12741_));
  NOR2_X1    g12549(.A1(new_n12374_), .A2(new_n11906_), .ZN(new_n12742_));
  NAND2_X1   g12550(.A1(new_n12742_), .A2(new_n12386_), .ZN(new_n12743_));
  AOI21_X1   g12551(.A1(new_n12743_), .A2(new_n12741_), .B(new_n193_), .ZN(new_n12744_));
  INV_X1     g12552(.I(new_n12744_), .ZN(new_n12745_));
  NAND3_X1   g12553(.A1(\asqrt[15] ), .A2(new_n12356_), .A3(new_n12367_), .ZN(new_n12746_));
  XOR2_X1    g12554(.A1(new_n12746_), .A2(new_n12359_), .Z(new_n12747_));
  AOI21_X1   g12555(.A1(new_n12742_), .A2(new_n12371_), .B(new_n12372_), .ZN(new_n12748_));
  OAI21_X1   g12556(.A1(new_n12326_), .A2(new_n12328_), .B(new_n12331_), .ZN(new_n12749_));
  NOR2_X1    g12557(.A1(new_n12374_), .A2(new_n12749_), .ZN(new_n12750_));
  XOR2_X1    g12558(.A1(new_n12750_), .A2(new_n11914_), .Z(new_n12751_));
  NAND3_X1   g12559(.A1(\asqrt[15] ), .A2(new_n12342_), .A3(new_n12327_), .ZN(new_n12752_));
  XOR2_X1    g12560(.A1(new_n12752_), .A2(new_n11918_), .Z(new_n12753_));
  OAI21_X1   g12561(.A1(new_n12337_), .A2(new_n12338_), .B(new_n12341_), .ZN(new_n12754_));
  NOR2_X1    g12562(.A1(new_n12374_), .A2(new_n12754_), .ZN(new_n12755_));
  XOR2_X1    g12563(.A1(new_n12755_), .A2(new_n11920_), .Z(new_n12756_));
  INV_X1     g12564(.I(new_n12756_), .ZN(new_n12757_));
  NAND3_X1   g12565(.A1(\asqrt[15] ), .A2(new_n12304_), .A3(new_n12323_), .ZN(new_n12758_));
  XOR2_X1    g12566(.A1(new_n12758_), .A2(new_n12335_), .Z(new_n12759_));
  INV_X1     g12567(.I(new_n12759_), .ZN(new_n12760_));
  OAI21_X1   g12568(.A1(new_n12298_), .A2(new_n12300_), .B(new_n12303_), .ZN(new_n12761_));
  NOR2_X1    g12569(.A1(new_n12374_), .A2(new_n12761_), .ZN(new_n12762_));
  XOR2_X1    g12570(.A1(new_n12762_), .A2(new_n11926_), .Z(new_n12763_));
  NAND3_X1   g12571(.A1(\asqrt[15] ), .A2(new_n12317_), .A3(new_n12299_), .ZN(new_n12764_));
  XOR2_X1    g12572(.A1(new_n12764_), .A2(new_n11930_), .Z(new_n12765_));
  OAI21_X1   g12573(.A1(new_n12312_), .A2(new_n12313_), .B(new_n12316_), .ZN(new_n12766_));
  NOR2_X1    g12574(.A1(new_n12374_), .A2(new_n12766_), .ZN(new_n12767_));
  XOR2_X1    g12575(.A1(new_n12767_), .A2(new_n11932_), .Z(new_n12768_));
  INV_X1     g12576(.I(new_n12768_), .ZN(new_n12769_));
  NAND3_X1   g12577(.A1(\asqrt[15] ), .A2(new_n12276_), .A3(new_n12295_), .ZN(new_n12770_));
  XOR2_X1    g12578(.A1(new_n12770_), .A2(new_n12310_), .Z(new_n12771_));
  INV_X1     g12579(.I(new_n12771_), .ZN(new_n12772_));
  OAI21_X1   g12580(.A1(new_n12270_), .A2(new_n12272_), .B(new_n12275_), .ZN(new_n12773_));
  NOR2_X1    g12581(.A1(new_n12374_), .A2(new_n12773_), .ZN(new_n12774_));
  XOR2_X1    g12582(.A1(new_n12774_), .A2(new_n11938_), .Z(new_n12775_));
  NAND3_X1   g12583(.A1(\asqrt[15] ), .A2(new_n12289_), .A3(new_n12271_), .ZN(new_n12776_));
  XOR2_X1    g12584(.A1(new_n12776_), .A2(new_n11942_), .Z(new_n12777_));
  NOR2_X1    g12585(.A1(new_n12738_), .A2(new_n12739_), .ZN(new_n12778_));
  AOI21_X1   g12586(.A1(new_n12778_), .A2(new_n1228_), .B(new_n12378_), .ZN(new_n12779_));
  NAND2_X1   g12587(.A1(new_n12740_), .A2(new_n1088_), .ZN(new_n12780_));
  OAI21_X1   g12588(.A1(new_n12779_), .A2(new_n12780_), .B(new_n12777_), .ZN(new_n12781_));
  INV_X1     g12589(.I(new_n12740_), .ZN(new_n12782_));
  OAI21_X1   g12590(.A1(new_n12779_), .A2(new_n12782_), .B(\asqrt[51] ), .ZN(new_n12783_));
  NAND3_X1   g12591(.A1(new_n12781_), .A2(new_n12783_), .A3(new_n962_), .ZN(new_n12784_));
  NAND2_X1   g12592(.A1(new_n12784_), .A2(new_n12775_), .ZN(new_n12785_));
  NAND2_X1   g12593(.A1(new_n12781_), .A2(new_n12783_), .ZN(new_n12786_));
  AOI21_X1   g12594(.A1(new_n12786_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n12787_));
  AOI21_X1   g12595(.A1(new_n12787_), .A2(new_n12785_), .B(new_n12772_), .ZN(new_n12788_));
  INV_X1     g12596(.I(new_n12777_), .ZN(new_n12789_));
  NAND2_X1   g12597(.A1(new_n12725_), .A2(new_n12377_), .ZN(new_n12790_));
  NAND2_X1   g12598(.A1(new_n12722_), .A2(new_n12724_), .ZN(new_n12791_));
  AOI21_X1   g12599(.A1(new_n12791_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n12792_));
  AOI21_X1   g12600(.A1(new_n12792_), .A2(new_n12790_), .B(new_n12789_), .ZN(new_n12793_));
  AOI21_X1   g12601(.A1(new_n12790_), .A2(new_n12740_), .B(new_n1088_), .ZN(new_n12794_));
  OAI21_X1   g12602(.A1(new_n12793_), .A2(new_n12794_), .B(\asqrt[52] ), .ZN(new_n12795_));
  AOI21_X1   g12603(.A1(new_n12785_), .A2(new_n12795_), .B(new_n842_), .ZN(new_n12796_));
  NOR2_X1    g12604(.A1(new_n12788_), .A2(new_n12796_), .ZN(new_n12797_));
  AOI21_X1   g12605(.A1(new_n12797_), .A2(new_n720_), .B(new_n12769_), .ZN(new_n12798_));
  OAI21_X1   g12606(.A1(new_n12788_), .A2(new_n12796_), .B(\asqrt[54] ), .ZN(new_n12799_));
  NAND2_X1   g12607(.A1(new_n12799_), .A2(new_n630_), .ZN(new_n12800_));
  OAI21_X1   g12608(.A1(new_n12798_), .A2(new_n12800_), .B(new_n12765_), .ZN(new_n12801_));
  INV_X1     g12609(.I(new_n12799_), .ZN(new_n12802_));
  OAI21_X1   g12610(.A1(new_n12798_), .A2(new_n12802_), .B(\asqrt[55] ), .ZN(new_n12803_));
  NAND3_X1   g12611(.A1(new_n12801_), .A2(new_n12803_), .A3(new_n545_), .ZN(new_n12804_));
  NAND2_X1   g12612(.A1(new_n12804_), .A2(new_n12763_), .ZN(new_n12805_));
  NAND2_X1   g12613(.A1(new_n12801_), .A2(new_n12803_), .ZN(new_n12806_));
  AOI21_X1   g12614(.A1(new_n12806_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n12807_));
  AOI21_X1   g12615(.A1(new_n12807_), .A2(new_n12805_), .B(new_n12760_), .ZN(new_n12808_));
  INV_X1     g12616(.I(new_n12765_), .ZN(new_n12809_));
  INV_X1     g12617(.I(new_n12775_), .ZN(new_n12810_));
  NOR2_X1    g12618(.A1(new_n12793_), .A2(new_n12794_), .ZN(new_n12811_));
  AOI21_X1   g12619(.A1(new_n12811_), .A2(new_n962_), .B(new_n12810_), .ZN(new_n12812_));
  NAND2_X1   g12620(.A1(new_n12795_), .A2(new_n842_), .ZN(new_n12813_));
  OAI21_X1   g12621(.A1(new_n12812_), .A2(new_n12813_), .B(new_n12771_), .ZN(new_n12814_));
  INV_X1     g12622(.I(new_n12795_), .ZN(new_n12815_));
  OAI21_X1   g12623(.A1(new_n12812_), .A2(new_n12815_), .B(\asqrt[53] ), .ZN(new_n12816_));
  NAND3_X1   g12624(.A1(new_n12814_), .A2(new_n12816_), .A3(new_n720_), .ZN(new_n12817_));
  NAND2_X1   g12625(.A1(new_n12817_), .A2(new_n12768_), .ZN(new_n12818_));
  NAND2_X1   g12626(.A1(new_n12814_), .A2(new_n12816_), .ZN(new_n12819_));
  AOI21_X1   g12627(.A1(new_n12819_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n12820_));
  AOI21_X1   g12628(.A1(new_n12820_), .A2(new_n12818_), .B(new_n12809_), .ZN(new_n12821_));
  AOI21_X1   g12629(.A1(new_n12818_), .A2(new_n12799_), .B(new_n630_), .ZN(new_n12822_));
  OAI21_X1   g12630(.A1(new_n12821_), .A2(new_n12822_), .B(\asqrt[56] ), .ZN(new_n12823_));
  AOI21_X1   g12631(.A1(new_n12805_), .A2(new_n12823_), .B(new_n450_), .ZN(new_n12824_));
  NOR2_X1    g12632(.A1(new_n12808_), .A2(new_n12824_), .ZN(new_n12825_));
  AOI21_X1   g12633(.A1(new_n12825_), .A2(new_n403_), .B(new_n12757_), .ZN(new_n12826_));
  OAI21_X1   g12634(.A1(new_n12808_), .A2(new_n12824_), .B(\asqrt[58] ), .ZN(new_n12827_));
  NAND2_X1   g12635(.A1(new_n12827_), .A2(new_n339_), .ZN(new_n12828_));
  OAI21_X1   g12636(.A1(new_n12826_), .A2(new_n12828_), .B(new_n12753_), .ZN(new_n12829_));
  INV_X1     g12637(.I(new_n12827_), .ZN(new_n12830_));
  OAI21_X1   g12638(.A1(new_n12826_), .A2(new_n12830_), .B(\asqrt[59] ), .ZN(new_n12831_));
  NAND3_X1   g12639(.A1(new_n12829_), .A2(new_n12831_), .A3(new_n288_), .ZN(new_n12832_));
  NAND2_X1   g12640(.A1(new_n12832_), .A2(new_n12751_), .ZN(new_n12833_));
  INV_X1     g12641(.I(new_n12753_), .ZN(new_n12834_));
  INV_X1     g12642(.I(new_n12763_), .ZN(new_n12835_));
  NOR2_X1    g12643(.A1(new_n12821_), .A2(new_n12822_), .ZN(new_n12836_));
  AOI21_X1   g12644(.A1(new_n12836_), .A2(new_n545_), .B(new_n12835_), .ZN(new_n12837_));
  NAND2_X1   g12645(.A1(new_n12823_), .A2(new_n450_), .ZN(new_n12838_));
  OAI21_X1   g12646(.A1(new_n12837_), .A2(new_n12838_), .B(new_n12759_), .ZN(new_n12839_));
  INV_X1     g12647(.I(new_n12823_), .ZN(new_n12840_));
  OAI21_X1   g12648(.A1(new_n12837_), .A2(new_n12840_), .B(\asqrt[57] ), .ZN(new_n12841_));
  NAND3_X1   g12649(.A1(new_n12839_), .A2(new_n12841_), .A3(new_n403_), .ZN(new_n12842_));
  NAND2_X1   g12650(.A1(new_n12842_), .A2(new_n12756_), .ZN(new_n12843_));
  NAND2_X1   g12651(.A1(new_n12839_), .A2(new_n12841_), .ZN(new_n12844_));
  AOI21_X1   g12652(.A1(new_n12844_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n12845_));
  AOI21_X1   g12653(.A1(new_n12845_), .A2(new_n12843_), .B(new_n12834_), .ZN(new_n12846_));
  AOI21_X1   g12654(.A1(new_n12843_), .A2(new_n12827_), .B(new_n339_), .ZN(new_n12847_));
  OAI21_X1   g12655(.A1(new_n12846_), .A2(new_n12847_), .B(\asqrt[60] ), .ZN(new_n12848_));
  AOI21_X1   g12656(.A1(new_n12833_), .A2(new_n12848_), .B(new_n242_), .ZN(new_n12849_));
  NAND3_X1   g12657(.A1(\asqrt[15] ), .A2(new_n12332_), .A3(new_n12348_), .ZN(new_n12850_));
  XOR2_X1    g12658(.A1(new_n12850_), .A2(new_n12360_), .Z(new_n12851_));
  INV_X1     g12659(.I(new_n12851_), .ZN(new_n12852_));
  NAND2_X1   g12660(.A1(new_n12829_), .A2(new_n12831_), .ZN(new_n12853_));
  AOI21_X1   g12661(.A1(new_n12853_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n12854_));
  AOI21_X1   g12662(.A1(new_n12854_), .A2(new_n12833_), .B(new_n12852_), .ZN(new_n12855_));
  OAI21_X1   g12663(.A1(new_n12855_), .A2(new_n12849_), .B(\asqrt[62] ), .ZN(new_n12856_));
  INV_X1     g12664(.I(new_n12856_), .ZN(new_n12857_));
  NOR2_X1    g12665(.A1(new_n12855_), .A2(new_n12849_), .ZN(new_n12858_));
  AOI21_X1   g12666(.A1(new_n12333_), .A2(new_n12354_), .B(new_n12349_), .ZN(new_n12859_));
  NAND2_X1   g12667(.A1(\asqrt[15] ), .A2(new_n12859_), .ZN(new_n12860_));
  XOR2_X1    g12668(.A1(new_n12860_), .A2(new_n12352_), .Z(new_n12861_));
  INV_X1     g12669(.I(new_n12861_), .ZN(new_n12862_));
  AOI21_X1   g12670(.A1(new_n12858_), .A2(new_n234_), .B(new_n12862_), .ZN(new_n12863_));
  OAI21_X1   g12671(.A1(new_n12863_), .A2(new_n12857_), .B(new_n12748_), .ZN(new_n12864_));
  OAI21_X1   g12672(.A1(new_n12864_), .A2(new_n12747_), .B(new_n193_), .ZN(new_n12865_));
  NOR2_X1    g12673(.A1(new_n12863_), .A2(new_n12857_), .ZN(new_n12866_));
  NAND2_X1   g12674(.A1(new_n12866_), .A2(new_n12747_), .ZN(new_n12867_));
  NOR2_X1    g12675(.A1(\asqrt[15] ), .A2(new_n11907_), .ZN(new_n12868_));
  INV_X1     g12676(.I(new_n12868_), .ZN(new_n12869_));
  NAND4_X1   g12677(.A1(new_n12865_), .A2(new_n12745_), .A3(new_n12867_), .A4(new_n12869_), .ZN(\asqrt[14] ));
  NAND3_X1   g12678(.A1(\asqrt[14] ), .A2(new_n12725_), .A3(new_n12740_), .ZN(new_n12871_));
  XOR2_X1    g12679(.A1(new_n12871_), .A2(new_n12378_), .Z(new_n12872_));
  INV_X1     g12680(.I(new_n12751_), .ZN(new_n12873_));
  NOR2_X1    g12681(.A1(new_n12846_), .A2(new_n12847_), .ZN(new_n12874_));
  AOI21_X1   g12682(.A1(new_n12874_), .A2(new_n288_), .B(new_n12873_), .ZN(new_n12875_));
  INV_X1     g12683(.I(new_n12848_), .ZN(new_n12876_));
  OAI21_X1   g12684(.A1(new_n12875_), .A2(new_n12876_), .B(\asqrt[61] ), .ZN(new_n12877_));
  NAND2_X1   g12685(.A1(new_n12848_), .A2(new_n242_), .ZN(new_n12878_));
  OAI21_X1   g12686(.A1(new_n12875_), .A2(new_n12878_), .B(new_n12851_), .ZN(new_n12879_));
  NAND3_X1   g12687(.A1(new_n12879_), .A2(new_n12877_), .A3(new_n234_), .ZN(new_n12880_));
  NAND2_X1   g12688(.A1(new_n12880_), .A2(new_n12861_), .ZN(new_n12881_));
  NAND2_X1   g12689(.A1(new_n12881_), .A2(new_n12856_), .ZN(new_n12882_));
  NAND2_X1   g12690(.A1(new_n12882_), .A2(new_n12747_), .ZN(new_n12883_));
  INV_X1     g12691(.I(new_n12747_), .ZN(new_n12884_));
  INV_X1     g12692(.I(new_n12748_), .ZN(new_n12885_));
  AOI21_X1   g12693(.A1(new_n12881_), .A2(new_n12856_), .B(new_n12885_), .ZN(new_n12886_));
  AOI21_X1   g12694(.A1(new_n12886_), .A2(new_n12884_), .B(\asqrt[63] ), .ZN(new_n12887_));
  NOR2_X1    g12695(.A1(new_n12882_), .A2(new_n12884_), .ZN(new_n12888_));
  NOR4_X1    g12696(.A1(new_n12887_), .A2(new_n12744_), .A3(new_n12888_), .A4(new_n12868_), .ZN(new_n12889_));
  NOR2_X1    g12697(.A1(new_n12889_), .A2(new_n12747_), .ZN(new_n12890_));
  NAND2_X1   g12698(.A1(new_n12890_), .A2(new_n12866_), .ZN(new_n12891_));
  AOI21_X1   g12699(.A1(new_n12891_), .A2(new_n12883_), .B(new_n193_), .ZN(new_n12892_));
  NAND3_X1   g12700(.A1(\asqrt[14] ), .A2(new_n12856_), .A3(new_n12880_), .ZN(new_n12893_));
  XOR2_X1    g12701(.A1(new_n12893_), .A2(new_n12861_), .Z(new_n12894_));
  INV_X1     g12702(.I(new_n12894_), .ZN(new_n12895_));
  AOI21_X1   g12703(.A1(new_n12890_), .A2(new_n12882_), .B(new_n12888_), .ZN(new_n12896_));
  INV_X1     g12704(.I(new_n12896_), .ZN(new_n12897_));
  OAI21_X1   g12705(.A1(new_n12826_), .A2(new_n12828_), .B(new_n12831_), .ZN(new_n12898_));
  NOR2_X1    g12706(.A1(new_n12889_), .A2(new_n12898_), .ZN(new_n12899_));
  XOR2_X1    g12707(.A1(new_n12899_), .A2(new_n12753_), .Z(new_n12900_));
  NAND3_X1   g12708(.A1(\asqrt[14] ), .A2(new_n12842_), .A3(new_n12827_), .ZN(new_n12901_));
  XOR2_X1    g12709(.A1(new_n12901_), .A2(new_n12757_), .Z(new_n12902_));
  OAI21_X1   g12710(.A1(new_n12837_), .A2(new_n12838_), .B(new_n12841_), .ZN(new_n12903_));
  NOR2_X1    g12711(.A1(new_n12889_), .A2(new_n12903_), .ZN(new_n12904_));
  XOR2_X1    g12712(.A1(new_n12904_), .A2(new_n12759_), .Z(new_n12905_));
  INV_X1     g12713(.I(new_n12905_), .ZN(new_n12906_));
  NAND3_X1   g12714(.A1(\asqrt[14] ), .A2(new_n12804_), .A3(new_n12823_), .ZN(new_n12907_));
  XOR2_X1    g12715(.A1(new_n12907_), .A2(new_n12835_), .Z(new_n12908_));
  INV_X1     g12716(.I(new_n12908_), .ZN(new_n12909_));
  OAI21_X1   g12717(.A1(new_n12798_), .A2(new_n12800_), .B(new_n12803_), .ZN(new_n12910_));
  NOR2_X1    g12718(.A1(new_n12889_), .A2(new_n12910_), .ZN(new_n12911_));
  XOR2_X1    g12719(.A1(new_n12911_), .A2(new_n12765_), .Z(new_n12912_));
  NAND3_X1   g12720(.A1(\asqrt[14] ), .A2(new_n12817_), .A3(new_n12799_), .ZN(new_n12913_));
  XOR2_X1    g12721(.A1(new_n12913_), .A2(new_n12769_), .Z(new_n12914_));
  OAI21_X1   g12722(.A1(new_n12812_), .A2(new_n12813_), .B(new_n12816_), .ZN(new_n12915_));
  NOR2_X1    g12723(.A1(new_n12889_), .A2(new_n12915_), .ZN(new_n12916_));
  XOR2_X1    g12724(.A1(new_n12916_), .A2(new_n12771_), .Z(new_n12917_));
  INV_X1     g12725(.I(new_n12917_), .ZN(new_n12918_));
  NAND3_X1   g12726(.A1(\asqrt[14] ), .A2(new_n12784_), .A3(new_n12795_), .ZN(new_n12919_));
  XOR2_X1    g12727(.A1(new_n12919_), .A2(new_n12810_), .Z(new_n12920_));
  INV_X1     g12728(.I(new_n12920_), .ZN(new_n12921_));
  OAI21_X1   g12729(.A1(new_n12779_), .A2(new_n12780_), .B(new_n12783_), .ZN(new_n12922_));
  NOR2_X1    g12730(.A1(new_n12889_), .A2(new_n12922_), .ZN(new_n12923_));
  XOR2_X1    g12731(.A1(new_n12923_), .A2(new_n12777_), .Z(new_n12924_));
  OAI21_X1   g12732(.A1(new_n12719_), .A2(new_n12721_), .B(new_n12724_), .ZN(new_n12925_));
  NOR2_X1    g12733(.A1(new_n12889_), .A2(new_n12925_), .ZN(new_n12926_));
  XOR2_X1    g12734(.A1(new_n12926_), .A2(new_n12391_), .Z(new_n12927_));
  INV_X1     g12735(.I(new_n12927_), .ZN(new_n12928_));
  NAND3_X1   g12736(.A1(\asqrt[14] ), .A2(new_n12734_), .A3(new_n12720_), .ZN(new_n12929_));
  XOR2_X1    g12737(.A1(new_n12929_), .A2(new_n12395_), .Z(new_n12930_));
  INV_X1     g12738(.I(new_n12930_), .ZN(new_n12931_));
  OAI21_X1   g12739(.A1(new_n12729_), .A2(new_n12730_), .B(new_n12733_), .ZN(new_n12932_));
  NOR2_X1    g12740(.A1(new_n12889_), .A2(new_n12932_), .ZN(new_n12933_));
  XOR2_X1    g12741(.A1(new_n12933_), .A2(new_n12397_), .Z(new_n12934_));
  NAND3_X1   g12742(.A1(\asqrt[14] ), .A2(new_n12697_), .A3(new_n12716_), .ZN(new_n12935_));
  XOR2_X1    g12743(.A1(new_n12935_), .A2(new_n12727_), .Z(new_n12936_));
  OAI21_X1   g12744(.A1(new_n12691_), .A2(new_n12693_), .B(new_n12696_), .ZN(new_n12937_));
  NOR2_X1    g12745(.A1(new_n12889_), .A2(new_n12937_), .ZN(new_n12938_));
  XOR2_X1    g12746(.A1(new_n12938_), .A2(new_n12403_), .Z(new_n12939_));
  INV_X1     g12747(.I(new_n12939_), .ZN(new_n12940_));
  NAND3_X1   g12748(.A1(\asqrt[14] ), .A2(new_n12710_), .A3(new_n12692_), .ZN(new_n12941_));
  XOR2_X1    g12749(.A1(new_n12941_), .A2(new_n12407_), .Z(new_n12942_));
  INV_X1     g12750(.I(new_n12942_), .ZN(new_n12943_));
  OAI21_X1   g12751(.A1(new_n12705_), .A2(new_n12706_), .B(new_n12709_), .ZN(new_n12944_));
  NOR2_X1    g12752(.A1(new_n12889_), .A2(new_n12944_), .ZN(new_n12945_));
  XOR2_X1    g12753(.A1(new_n12945_), .A2(new_n12409_), .Z(new_n12946_));
  NAND3_X1   g12754(.A1(\asqrt[14] ), .A2(new_n12669_), .A3(new_n12688_), .ZN(new_n12947_));
  XOR2_X1    g12755(.A1(new_n12947_), .A2(new_n12703_), .Z(new_n12948_));
  OAI21_X1   g12756(.A1(new_n12663_), .A2(new_n12665_), .B(new_n12668_), .ZN(new_n12949_));
  NOR2_X1    g12757(.A1(new_n12889_), .A2(new_n12949_), .ZN(new_n12950_));
  XOR2_X1    g12758(.A1(new_n12950_), .A2(new_n12415_), .Z(new_n12951_));
  INV_X1     g12759(.I(new_n12951_), .ZN(new_n12952_));
  NAND3_X1   g12760(.A1(\asqrt[14] ), .A2(new_n12682_), .A3(new_n12664_), .ZN(new_n12953_));
  XOR2_X1    g12761(.A1(new_n12953_), .A2(new_n12419_), .Z(new_n12954_));
  INV_X1     g12762(.I(new_n12954_), .ZN(new_n12955_));
  OAI21_X1   g12763(.A1(new_n12677_), .A2(new_n12678_), .B(new_n12681_), .ZN(new_n12956_));
  NOR2_X1    g12764(.A1(new_n12889_), .A2(new_n12956_), .ZN(new_n12957_));
  XOR2_X1    g12765(.A1(new_n12957_), .A2(new_n12421_), .Z(new_n12958_));
  NAND3_X1   g12766(.A1(\asqrt[14] ), .A2(new_n12641_), .A3(new_n12660_), .ZN(new_n12959_));
  XOR2_X1    g12767(.A1(new_n12959_), .A2(new_n12675_), .Z(new_n12960_));
  OAI21_X1   g12768(.A1(new_n12635_), .A2(new_n12637_), .B(new_n12640_), .ZN(new_n12961_));
  NOR2_X1    g12769(.A1(new_n12889_), .A2(new_n12961_), .ZN(new_n12962_));
  XOR2_X1    g12770(.A1(new_n12962_), .A2(new_n12427_), .Z(new_n12963_));
  INV_X1     g12771(.I(new_n12963_), .ZN(new_n12964_));
  NAND3_X1   g12772(.A1(\asqrt[14] ), .A2(new_n12654_), .A3(new_n12636_), .ZN(new_n12965_));
  XOR2_X1    g12773(.A1(new_n12965_), .A2(new_n12431_), .Z(new_n12966_));
  INV_X1     g12774(.I(new_n12966_), .ZN(new_n12967_));
  OAI21_X1   g12775(.A1(new_n12649_), .A2(new_n12650_), .B(new_n12653_), .ZN(new_n12968_));
  NOR2_X1    g12776(.A1(new_n12889_), .A2(new_n12968_), .ZN(new_n12969_));
  XOR2_X1    g12777(.A1(new_n12969_), .A2(new_n12433_), .Z(new_n12970_));
  NAND3_X1   g12778(.A1(\asqrt[14] ), .A2(new_n12613_), .A3(new_n12632_), .ZN(new_n12971_));
  XOR2_X1    g12779(.A1(new_n12971_), .A2(new_n12647_), .Z(new_n12972_));
  OAI21_X1   g12780(.A1(new_n12607_), .A2(new_n12609_), .B(new_n12612_), .ZN(new_n12973_));
  NOR2_X1    g12781(.A1(new_n12889_), .A2(new_n12973_), .ZN(new_n12974_));
  XOR2_X1    g12782(.A1(new_n12974_), .A2(new_n12439_), .Z(new_n12975_));
  INV_X1     g12783(.I(new_n12975_), .ZN(new_n12976_));
  NAND3_X1   g12784(.A1(\asqrt[14] ), .A2(new_n12626_), .A3(new_n12608_), .ZN(new_n12977_));
  XOR2_X1    g12785(.A1(new_n12977_), .A2(new_n12443_), .Z(new_n12978_));
  INV_X1     g12786(.I(new_n12978_), .ZN(new_n12979_));
  OAI21_X1   g12787(.A1(new_n12621_), .A2(new_n12622_), .B(new_n12625_), .ZN(new_n12980_));
  NOR2_X1    g12788(.A1(new_n12889_), .A2(new_n12980_), .ZN(new_n12981_));
  XOR2_X1    g12789(.A1(new_n12981_), .A2(new_n12445_), .Z(new_n12982_));
  NAND3_X1   g12790(.A1(\asqrt[14] ), .A2(new_n12585_), .A3(new_n12604_), .ZN(new_n12983_));
  XOR2_X1    g12791(.A1(new_n12983_), .A2(new_n12619_), .Z(new_n12984_));
  OAI21_X1   g12792(.A1(new_n12579_), .A2(new_n12581_), .B(new_n12584_), .ZN(new_n12985_));
  NOR2_X1    g12793(.A1(new_n12889_), .A2(new_n12985_), .ZN(new_n12986_));
  XOR2_X1    g12794(.A1(new_n12986_), .A2(new_n12451_), .Z(new_n12987_));
  INV_X1     g12795(.I(new_n12987_), .ZN(new_n12988_));
  NAND3_X1   g12796(.A1(\asqrt[14] ), .A2(new_n12598_), .A3(new_n12580_), .ZN(new_n12989_));
  XOR2_X1    g12797(.A1(new_n12989_), .A2(new_n12455_), .Z(new_n12990_));
  INV_X1     g12798(.I(new_n12990_), .ZN(new_n12991_));
  OAI21_X1   g12799(.A1(new_n12593_), .A2(new_n12594_), .B(new_n12597_), .ZN(new_n12992_));
  NOR2_X1    g12800(.A1(new_n12889_), .A2(new_n12992_), .ZN(new_n12993_));
  XOR2_X1    g12801(.A1(new_n12993_), .A2(new_n12457_), .Z(new_n12994_));
  NAND3_X1   g12802(.A1(\asqrt[14] ), .A2(new_n12557_), .A3(new_n12576_), .ZN(new_n12995_));
  XOR2_X1    g12803(.A1(new_n12995_), .A2(new_n12591_), .Z(new_n12996_));
  OAI21_X1   g12804(.A1(new_n12551_), .A2(new_n12553_), .B(new_n12556_), .ZN(new_n12997_));
  NOR2_X1    g12805(.A1(new_n12889_), .A2(new_n12997_), .ZN(new_n12998_));
  XOR2_X1    g12806(.A1(new_n12998_), .A2(new_n12463_), .Z(new_n12999_));
  INV_X1     g12807(.I(new_n12999_), .ZN(new_n13000_));
  NAND3_X1   g12808(.A1(\asqrt[14] ), .A2(new_n12570_), .A3(new_n12552_), .ZN(new_n13001_));
  XOR2_X1    g12809(.A1(new_n13001_), .A2(new_n12467_), .Z(new_n13002_));
  INV_X1     g12810(.I(new_n13002_), .ZN(new_n13003_));
  OAI21_X1   g12811(.A1(new_n12565_), .A2(new_n12566_), .B(new_n12569_), .ZN(new_n13004_));
  NOR2_X1    g12812(.A1(new_n12889_), .A2(new_n13004_), .ZN(new_n13005_));
  XOR2_X1    g12813(.A1(new_n13005_), .A2(new_n12469_), .Z(new_n13006_));
  NAND3_X1   g12814(.A1(\asqrt[14] ), .A2(new_n12529_), .A3(new_n12548_), .ZN(new_n13007_));
  XOR2_X1    g12815(.A1(new_n13007_), .A2(new_n12563_), .Z(new_n13008_));
  OAI21_X1   g12816(.A1(new_n12523_), .A2(new_n12525_), .B(new_n12528_), .ZN(new_n13009_));
  NOR2_X1    g12817(.A1(new_n12889_), .A2(new_n13009_), .ZN(new_n13010_));
  XOR2_X1    g12818(.A1(new_n13010_), .A2(new_n12476_), .Z(new_n13011_));
  INV_X1     g12819(.I(new_n13011_), .ZN(new_n13012_));
  NAND3_X1   g12820(.A1(\asqrt[14] ), .A2(new_n12542_), .A3(new_n12524_), .ZN(new_n13013_));
  XOR2_X1    g12821(.A1(new_n13013_), .A2(new_n12479_), .Z(new_n13014_));
  INV_X1     g12822(.I(new_n13014_), .ZN(new_n13015_));
  OAI21_X1   g12823(.A1(new_n12537_), .A2(new_n12538_), .B(new_n12541_), .ZN(new_n13016_));
  NOR2_X1    g12824(.A1(new_n12889_), .A2(new_n13016_), .ZN(new_n13017_));
  XOR2_X1    g12825(.A1(new_n13017_), .A2(new_n12482_), .Z(new_n13018_));
  NAND3_X1   g12826(.A1(\asqrt[14] ), .A2(new_n12502_), .A3(new_n12520_), .ZN(new_n13019_));
  XOR2_X1    g12827(.A1(new_n13019_), .A2(new_n12536_), .Z(new_n13020_));
  NOR2_X1    g12828(.A1(new_n12499_), .A2(\asqrt[17] ), .ZN(new_n13021_));
  NOR3_X1    g12829(.A1(new_n12889_), .A2(new_n13021_), .A3(new_n12519_), .ZN(new_n13022_));
  XOR2_X1    g12830(.A1(new_n13022_), .A2(new_n12490_), .Z(new_n13023_));
  INV_X1     g12831(.I(new_n13023_), .ZN(new_n13024_));
  NAND3_X1   g12832(.A1(\asqrt[14] ), .A2(new_n12491_), .A3(new_n12492_), .ZN(new_n13025_));
  NOR4_X1    g12833(.A1(new_n12887_), .A2(new_n12374_), .A3(new_n12744_), .A4(new_n12888_), .ZN(new_n13026_));
  INV_X1     g12834(.I(new_n13026_), .ZN(new_n13027_));
  AOI21_X1   g12835(.A1(new_n13025_), .A2(new_n13027_), .B(\a[30] ), .ZN(new_n13028_));
  NOR3_X1    g12836(.A1(new_n12889_), .A2(\a[28] ), .A3(\a[29] ), .ZN(new_n13029_));
  NOR3_X1    g12837(.A1(new_n13029_), .A2(new_n12038_), .A3(new_n13026_), .ZN(new_n13030_));
  NOR2_X1    g12838(.A1(new_n13030_), .A2(new_n13028_), .ZN(new_n13031_));
  INV_X1     g12839(.I(\a[26] ), .ZN(new_n13032_));
  INV_X1     g12840(.I(\a[27] ), .ZN(new_n13033_));
  NAND3_X1   g12841(.A1(new_n13032_), .A2(new_n13033_), .A3(new_n12491_), .ZN(new_n13034_));
  OAI21_X1   g12842(.A1(new_n12889_), .A2(new_n12491_), .B(new_n13034_), .ZN(new_n13035_));
  NAND2_X1   g12843(.A1(new_n13035_), .A2(\asqrt[15] ), .ZN(new_n13036_));
  OAI21_X1   g12844(.A1(new_n12889_), .A2(\a[28] ), .B(\a[29] ), .ZN(new_n13037_));
  NAND2_X1   g12845(.A1(new_n13037_), .A2(new_n13025_), .ZN(new_n13038_));
  NOR2_X1    g12846(.A1(new_n13035_), .A2(\asqrt[15] ), .ZN(new_n13039_));
  OAI21_X1   g12847(.A1(new_n13038_), .A2(new_n13039_), .B(new_n13036_), .ZN(new_n13040_));
  OAI21_X1   g12848(.A1(new_n13040_), .A2(\asqrt[16] ), .B(new_n13031_), .ZN(new_n13041_));
  NAND2_X1   g12849(.A1(new_n13040_), .A2(\asqrt[16] ), .ZN(new_n13042_));
  NAND3_X1   g12850(.A1(new_n13041_), .A2(new_n11406_), .A3(new_n13042_), .ZN(new_n13043_));
  NOR3_X1    g12851(.A1(new_n12889_), .A2(new_n12513_), .A3(new_n12498_), .ZN(new_n13044_));
  XOR2_X1    g12852(.A1(new_n13044_), .A2(new_n12515_), .Z(new_n13045_));
  AOI21_X1   g12853(.A1(new_n13041_), .A2(new_n13042_), .B(new_n11406_), .ZN(new_n13046_));
  AOI21_X1   g12854(.A1(new_n13043_), .A2(new_n13045_), .B(new_n13046_), .ZN(new_n13047_));
  AOI21_X1   g12855(.A1(new_n13047_), .A2(new_n10953_), .B(new_n13024_), .ZN(new_n13048_));
  OAI21_X1   g12856(.A1(new_n13047_), .A2(new_n10953_), .B(new_n10478_), .ZN(new_n13049_));
  OAI21_X1   g12857(.A1(new_n13048_), .A2(new_n13049_), .B(new_n13020_), .ZN(new_n13050_));
  NOR2_X1    g12858(.A1(new_n13047_), .A2(new_n10953_), .ZN(new_n13051_));
  OAI21_X1   g12859(.A1(new_n13048_), .A2(new_n13051_), .B(\asqrt[19] ), .ZN(new_n13052_));
  NAND3_X1   g12860(.A1(new_n13050_), .A2(new_n13052_), .A3(new_n10045_), .ZN(new_n13053_));
  NAND2_X1   g12861(.A1(new_n13053_), .A2(new_n13018_), .ZN(new_n13054_));
  NAND2_X1   g12862(.A1(new_n13050_), .A2(new_n13052_), .ZN(new_n13055_));
  AOI21_X1   g12863(.A1(new_n13055_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n13056_));
  AOI21_X1   g12864(.A1(new_n13056_), .A2(new_n13054_), .B(new_n13015_), .ZN(new_n13057_));
  INV_X1     g12865(.I(new_n13020_), .ZN(new_n13058_));
  OAI21_X1   g12866(.A1(new_n13029_), .A2(new_n13026_), .B(new_n12038_), .ZN(new_n13059_));
  NAND3_X1   g12867(.A1(new_n13025_), .A2(new_n13027_), .A3(\a[30] ), .ZN(new_n13060_));
  NAND2_X1   g12868(.A1(new_n13059_), .A2(new_n13060_), .ZN(new_n13061_));
  NAND2_X1   g12869(.A1(\asqrt[14] ), .A2(\a[28] ), .ZN(new_n13062_));
  AOI21_X1   g12870(.A1(new_n13062_), .A2(new_n13034_), .B(new_n12374_), .ZN(new_n13063_));
  AOI21_X1   g12871(.A1(\asqrt[14] ), .A2(new_n12491_), .B(new_n12492_), .ZN(new_n13064_));
  NOR2_X1    g12872(.A1(new_n13029_), .A2(new_n13064_), .ZN(new_n13065_));
  NAND3_X1   g12873(.A1(new_n13062_), .A2(new_n12374_), .A3(new_n13034_), .ZN(new_n13066_));
  AOI21_X1   g12874(.A1(new_n13065_), .A2(new_n13066_), .B(new_n13063_), .ZN(new_n13067_));
  AOI21_X1   g12875(.A1(new_n13067_), .A2(new_n11901_), .B(new_n13061_), .ZN(new_n13068_));
  NOR2_X1    g12876(.A1(new_n13067_), .A2(new_n11901_), .ZN(new_n13069_));
  NOR3_X1    g12877(.A1(new_n13068_), .A2(\asqrt[17] ), .A3(new_n13069_), .ZN(new_n13070_));
  INV_X1     g12878(.I(new_n13045_), .ZN(new_n13071_));
  OAI21_X1   g12879(.A1(new_n13068_), .A2(new_n13069_), .B(\asqrt[17] ), .ZN(new_n13072_));
  OAI21_X1   g12880(.A1(new_n13070_), .A2(new_n13071_), .B(new_n13072_), .ZN(new_n13073_));
  OAI21_X1   g12881(.A1(new_n13073_), .A2(\asqrt[18] ), .B(new_n13023_), .ZN(new_n13074_));
  AOI21_X1   g12882(.A1(new_n13073_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n13075_));
  AOI21_X1   g12883(.A1(new_n13075_), .A2(new_n13074_), .B(new_n13058_), .ZN(new_n13076_));
  NAND2_X1   g12884(.A1(new_n13073_), .A2(\asqrt[18] ), .ZN(new_n13077_));
  AOI21_X1   g12885(.A1(new_n13074_), .A2(new_n13077_), .B(new_n10478_), .ZN(new_n13078_));
  OAI21_X1   g12886(.A1(new_n13076_), .A2(new_n13078_), .B(\asqrt[20] ), .ZN(new_n13079_));
  AOI21_X1   g12887(.A1(new_n13054_), .A2(new_n13079_), .B(new_n9590_), .ZN(new_n13080_));
  NOR2_X1    g12888(.A1(new_n13057_), .A2(new_n13080_), .ZN(new_n13081_));
  AOI21_X1   g12889(.A1(new_n13081_), .A2(new_n9177_), .B(new_n13012_), .ZN(new_n13082_));
  OAI21_X1   g12890(.A1(new_n13057_), .A2(new_n13080_), .B(\asqrt[22] ), .ZN(new_n13083_));
  NAND2_X1   g12891(.A1(new_n13083_), .A2(new_n8742_), .ZN(new_n13084_));
  OAI21_X1   g12892(.A1(new_n13082_), .A2(new_n13084_), .B(new_n13008_), .ZN(new_n13085_));
  INV_X1     g12893(.I(new_n13083_), .ZN(new_n13086_));
  OAI21_X1   g12894(.A1(new_n13082_), .A2(new_n13086_), .B(\asqrt[23] ), .ZN(new_n13087_));
  NAND3_X1   g12895(.A1(new_n13085_), .A2(new_n13087_), .A3(new_n8349_), .ZN(new_n13088_));
  NAND2_X1   g12896(.A1(new_n13088_), .A2(new_n13006_), .ZN(new_n13089_));
  NAND2_X1   g12897(.A1(new_n13085_), .A2(new_n13087_), .ZN(new_n13090_));
  AOI21_X1   g12898(.A1(new_n13090_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n13091_));
  AOI21_X1   g12899(.A1(new_n13091_), .A2(new_n13089_), .B(new_n13003_), .ZN(new_n13092_));
  INV_X1     g12900(.I(new_n13008_), .ZN(new_n13093_));
  INV_X1     g12901(.I(new_n13018_), .ZN(new_n13094_));
  NOR2_X1    g12902(.A1(new_n13076_), .A2(new_n13078_), .ZN(new_n13095_));
  AOI21_X1   g12903(.A1(new_n13095_), .A2(new_n10045_), .B(new_n13094_), .ZN(new_n13096_));
  NAND2_X1   g12904(.A1(new_n13079_), .A2(new_n9590_), .ZN(new_n13097_));
  OAI21_X1   g12905(.A1(new_n13096_), .A2(new_n13097_), .B(new_n13014_), .ZN(new_n13098_));
  INV_X1     g12906(.I(new_n13079_), .ZN(new_n13099_));
  OAI21_X1   g12907(.A1(new_n13096_), .A2(new_n13099_), .B(\asqrt[21] ), .ZN(new_n13100_));
  NAND3_X1   g12908(.A1(new_n13098_), .A2(new_n13100_), .A3(new_n9177_), .ZN(new_n13101_));
  NAND2_X1   g12909(.A1(new_n13101_), .A2(new_n13011_), .ZN(new_n13102_));
  NAND2_X1   g12910(.A1(new_n13098_), .A2(new_n13100_), .ZN(new_n13103_));
  AOI21_X1   g12911(.A1(new_n13103_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n13104_));
  AOI21_X1   g12912(.A1(new_n13104_), .A2(new_n13102_), .B(new_n13093_), .ZN(new_n13105_));
  AOI21_X1   g12913(.A1(new_n13102_), .A2(new_n13083_), .B(new_n8742_), .ZN(new_n13106_));
  OAI21_X1   g12914(.A1(new_n13105_), .A2(new_n13106_), .B(\asqrt[24] ), .ZN(new_n13107_));
  AOI21_X1   g12915(.A1(new_n13089_), .A2(new_n13107_), .B(new_n7934_), .ZN(new_n13108_));
  NOR2_X1    g12916(.A1(new_n13092_), .A2(new_n13108_), .ZN(new_n13109_));
  AOI21_X1   g12917(.A1(new_n13109_), .A2(new_n7561_), .B(new_n13000_), .ZN(new_n13110_));
  OAI21_X1   g12918(.A1(new_n13092_), .A2(new_n13108_), .B(\asqrt[26] ), .ZN(new_n13111_));
  NAND2_X1   g12919(.A1(new_n13111_), .A2(new_n7166_), .ZN(new_n13112_));
  OAI21_X1   g12920(.A1(new_n13110_), .A2(new_n13112_), .B(new_n12996_), .ZN(new_n13113_));
  INV_X1     g12921(.I(new_n13111_), .ZN(new_n13114_));
  OAI21_X1   g12922(.A1(new_n13110_), .A2(new_n13114_), .B(\asqrt[27] ), .ZN(new_n13115_));
  NAND3_X1   g12923(.A1(new_n13113_), .A2(new_n13115_), .A3(new_n6813_), .ZN(new_n13116_));
  NAND2_X1   g12924(.A1(new_n13116_), .A2(new_n12994_), .ZN(new_n13117_));
  NAND2_X1   g12925(.A1(new_n13113_), .A2(new_n13115_), .ZN(new_n13118_));
  AOI21_X1   g12926(.A1(new_n13118_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n13119_));
  AOI21_X1   g12927(.A1(new_n13119_), .A2(new_n13117_), .B(new_n12991_), .ZN(new_n13120_));
  INV_X1     g12928(.I(new_n12996_), .ZN(new_n13121_));
  INV_X1     g12929(.I(new_n13006_), .ZN(new_n13122_));
  NOR2_X1    g12930(.A1(new_n13105_), .A2(new_n13106_), .ZN(new_n13123_));
  AOI21_X1   g12931(.A1(new_n13123_), .A2(new_n8349_), .B(new_n13122_), .ZN(new_n13124_));
  NAND2_X1   g12932(.A1(new_n13107_), .A2(new_n7934_), .ZN(new_n13125_));
  OAI21_X1   g12933(.A1(new_n13124_), .A2(new_n13125_), .B(new_n13002_), .ZN(new_n13126_));
  INV_X1     g12934(.I(new_n13107_), .ZN(new_n13127_));
  OAI21_X1   g12935(.A1(new_n13124_), .A2(new_n13127_), .B(\asqrt[25] ), .ZN(new_n13128_));
  NAND3_X1   g12936(.A1(new_n13126_), .A2(new_n13128_), .A3(new_n7561_), .ZN(new_n13129_));
  NAND2_X1   g12937(.A1(new_n13129_), .A2(new_n12999_), .ZN(new_n13130_));
  NAND2_X1   g12938(.A1(new_n13126_), .A2(new_n13128_), .ZN(new_n13131_));
  AOI21_X1   g12939(.A1(new_n13131_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n13132_));
  AOI21_X1   g12940(.A1(new_n13132_), .A2(new_n13130_), .B(new_n13121_), .ZN(new_n13133_));
  AOI21_X1   g12941(.A1(new_n13130_), .A2(new_n13111_), .B(new_n7166_), .ZN(new_n13134_));
  OAI21_X1   g12942(.A1(new_n13133_), .A2(new_n13134_), .B(\asqrt[28] ), .ZN(new_n13135_));
  AOI21_X1   g12943(.A1(new_n13117_), .A2(new_n13135_), .B(new_n6454_), .ZN(new_n13136_));
  NOR2_X1    g12944(.A1(new_n13120_), .A2(new_n13136_), .ZN(new_n13137_));
  AOI21_X1   g12945(.A1(new_n13137_), .A2(new_n6106_), .B(new_n12988_), .ZN(new_n13138_));
  OAI21_X1   g12946(.A1(new_n13120_), .A2(new_n13136_), .B(\asqrt[30] ), .ZN(new_n13139_));
  NAND2_X1   g12947(.A1(new_n13139_), .A2(new_n5750_), .ZN(new_n13140_));
  OAI21_X1   g12948(.A1(new_n13138_), .A2(new_n13140_), .B(new_n12984_), .ZN(new_n13141_));
  INV_X1     g12949(.I(new_n13139_), .ZN(new_n13142_));
  OAI21_X1   g12950(.A1(new_n13138_), .A2(new_n13142_), .B(\asqrt[31] ), .ZN(new_n13143_));
  NAND3_X1   g12951(.A1(new_n13141_), .A2(new_n13143_), .A3(new_n5435_), .ZN(new_n13144_));
  NAND2_X1   g12952(.A1(new_n13144_), .A2(new_n12982_), .ZN(new_n13145_));
  NAND2_X1   g12953(.A1(new_n13141_), .A2(new_n13143_), .ZN(new_n13146_));
  AOI21_X1   g12954(.A1(new_n13146_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n13147_));
  AOI21_X1   g12955(.A1(new_n13147_), .A2(new_n13145_), .B(new_n12979_), .ZN(new_n13148_));
  INV_X1     g12956(.I(new_n12984_), .ZN(new_n13149_));
  INV_X1     g12957(.I(new_n12994_), .ZN(new_n13150_));
  NOR2_X1    g12958(.A1(new_n13133_), .A2(new_n13134_), .ZN(new_n13151_));
  AOI21_X1   g12959(.A1(new_n13151_), .A2(new_n6813_), .B(new_n13150_), .ZN(new_n13152_));
  NAND2_X1   g12960(.A1(new_n13135_), .A2(new_n6454_), .ZN(new_n13153_));
  OAI21_X1   g12961(.A1(new_n13152_), .A2(new_n13153_), .B(new_n12990_), .ZN(new_n13154_));
  INV_X1     g12962(.I(new_n13135_), .ZN(new_n13155_));
  OAI21_X1   g12963(.A1(new_n13152_), .A2(new_n13155_), .B(\asqrt[29] ), .ZN(new_n13156_));
  NAND3_X1   g12964(.A1(new_n13154_), .A2(new_n13156_), .A3(new_n6106_), .ZN(new_n13157_));
  NAND2_X1   g12965(.A1(new_n13157_), .A2(new_n12987_), .ZN(new_n13158_));
  NAND2_X1   g12966(.A1(new_n13154_), .A2(new_n13156_), .ZN(new_n13159_));
  AOI21_X1   g12967(.A1(new_n13159_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n13160_));
  AOI21_X1   g12968(.A1(new_n13160_), .A2(new_n13158_), .B(new_n13149_), .ZN(new_n13161_));
  AOI21_X1   g12969(.A1(new_n13158_), .A2(new_n13139_), .B(new_n5750_), .ZN(new_n13162_));
  OAI21_X1   g12970(.A1(new_n13161_), .A2(new_n13162_), .B(\asqrt[32] ), .ZN(new_n13163_));
  AOI21_X1   g12971(.A1(new_n13145_), .A2(new_n13163_), .B(new_n5110_), .ZN(new_n13164_));
  NOR2_X1    g12972(.A1(new_n13148_), .A2(new_n13164_), .ZN(new_n13165_));
  AOI21_X1   g12973(.A1(new_n13165_), .A2(new_n4810_), .B(new_n12976_), .ZN(new_n13166_));
  OAI21_X1   g12974(.A1(new_n13148_), .A2(new_n13164_), .B(\asqrt[34] ), .ZN(new_n13167_));
  NAND2_X1   g12975(.A1(new_n13167_), .A2(new_n4510_), .ZN(new_n13168_));
  OAI21_X1   g12976(.A1(new_n13166_), .A2(new_n13168_), .B(new_n12972_), .ZN(new_n13169_));
  INV_X1     g12977(.I(new_n13167_), .ZN(new_n13170_));
  OAI21_X1   g12978(.A1(new_n13166_), .A2(new_n13170_), .B(\asqrt[35] ), .ZN(new_n13171_));
  NAND3_X1   g12979(.A1(new_n13169_), .A2(new_n13171_), .A3(new_n4224_), .ZN(new_n13172_));
  NAND2_X1   g12980(.A1(new_n13172_), .A2(new_n12970_), .ZN(new_n13173_));
  NAND2_X1   g12981(.A1(new_n13169_), .A2(new_n13171_), .ZN(new_n13174_));
  AOI21_X1   g12982(.A1(new_n13174_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n13175_));
  AOI21_X1   g12983(.A1(new_n13175_), .A2(new_n13173_), .B(new_n12967_), .ZN(new_n13176_));
  INV_X1     g12984(.I(new_n12972_), .ZN(new_n13177_));
  INV_X1     g12985(.I(new_n12982_), .ZN(new_n13178_));
  NOR2_X1    g12986(.A1(new_n13161_), .A2(new_n13162_), .ZN(new_n13179_));
  AOI21_X1   g12987(.A1(new_n13179_), .A2(new_n5435_), .B(new_n13178_), .ZN(new_n13180_));
  NAND2_X1   g12988(.A1(new_n13163_), .A2(new_n5110_), .ZN(new_n13181_));
  OAI21_X1   g12989(.A1(new_n13180_), .A2(new_n13181_), .B(new_n12978_), .ZN(new_n13182_));
  INV_X1     g12990(.I(new_n13163_), .ZN(new_n13183_));
  OAI21_X1   g12991(.A1(new_n13180_), .A2(new_n13183_), .B(\asqrt[33] ), .ZN(new_n13184_));
  NAND3_X1   g12992(.A1(new_n13182_), .A2(new_n13184_), .A3(new_n4810_), .ZN(new_n13185_));
  NAND2_X1   g12993(.A1(new_n13185_), .A2(new_n12975_), .ZN(new_n13186_));
  NAND2_X1   g12994(.A1(new_n13182_), .A2(new_n13184_), .ZN(new_n13187_));
  AOI21_X1   g12995(.A1(new_n13187_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n13188_));
  AOI21_X1   g12996(.A1(new_n13188_), .A2(new_n13186_), .B(new_n13177_), .ZN(new_n13189_));
  AOI21_X1   g12997(.A1(new_n13186_), .A2(new_n13167_), .B(new_n4510_), .ZN(new_n13190_));
  OAI21_X1   g12998(.A1(new_n13189_), .A2(new_n13190_), .B(\asqrt[36] ), .ZN(new_n13191_));
  AOI21_X1   g12999(.A1(new_n13173_), .A2(new_n13191_), .B(new_n3928_), .ZN(new_n13192_));
  NOR2_X1    g13000(.A1(new_n13176_), .A2(new_n13192_), .ZN(new_n13193_));
  AOI21_X1   g13001(.A1(new_n13193_), .A2(new_n3675_), .B(new_n12964_), .ZN(new_n13194_));
  OAI21_X1   g13002(.A1(new_n13176_), .A2(new_n13192_), .B(\asqrt[38] ), .ZN(new_n13195_));
  NAND2_X1   g13003(.A1(new_n13195_), .A2(new_n3400_), .ZN(new_n13196_));
  OAI21_X1   g13004(.A1(new_n13194_), .A2(new_n13196_), .B(new_n12960_), .ZN(new_n13197_));
  INV_X1     g13005(.I(new_n13195_), .ZN(new_n13198_));
  OAI21_X1   g13006(.A1(new_n13194_), .A2(new_n13198_), .B(\asqrt[39] ), .ZN(new_n13199_));
  NAND3_X1   g13007(.A1(new_n13197_), .A2(new_n13199_), .A3(new_n3167_), .ZN(new_n13200_));
  NAND2_X1   g13008(.A1(new_n13200_), .A2(new_n12958_), .ZN(new_n13201_));
  NAND2_X1   g13009(.A1(new_n13197_), .A2(new_n13199_), .ZN(new_n13202_));
  AOI21_X1   g13010(.A1(new_n13202_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n13203_));
  AOI21_X1   g13011(.A1(new_n13203_), .A2(new_n13201_), .B(new_n12955_), .ZN(new_n13204_));
  INV_X1     g13012(.I(new_n12960_), .ZN(new_n13205_));
  INV_X1     g13013(.I(new_n12970_), .ZN(new_n13206_));
  NOR2_X1    g13014(.A1(new_n13189_), .A2(new_n13190_), .ZN(new_n13207_));
  AOI21_X1   g13015(.A1(new_n13207_), .A2(new_n4224_), .B(new_n13206_), .ZN(new_n13208_));
  NAND2_X1   g13016(.A1(new_n13191_), .A2(new_n3928_), .ZN(new_n13209_));
  OAI21_X1   g13017(.A1(new_n13208_), .A2(new_n13209_), .B(new_n12966_), .ZN(new_n13210_));
  INV_X1     g13018(.I(new_n13191_), .ZN(new_n13211_));
  OAI21_X1   g13019(.A1(new_n13208_), .A2(new_n13211_), .B(\asqrt[37] ), .ZN(new_n13212_));
  NAND3_X1   g13020(.A1(new_n13210_), .A2(new_n13212_), .A3(new_n3675_), .ZN(new_n13213_));
  NAND2_X1   g13021(.A1(new_n13213_), .A2(new_n12963_), .ZN(new_n13214_));
  NAND2_X1   g13022(.A1(new_n13210_), .A2(new_n13212_), .ZN(new_n13215_));
  AOI21_X1   g13023(.A1(new_n13215_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n13216_));
  AOI21_X1   g13024(.A1(new_n13216_), .A2(new_n13214_), .B(new_n13205_), .ZN(new_n13217_));
  AOI21_X1   g13025(.A1(new_n13214_), .A2(new_n13195_), .B(new_n3400_), .ZN(new_n13218_));
  OAI21_X1   g13026(.A1(new_n13217_), .A2(new_n13218_), .B(\asqrt[40] ), .ZN(new_n13219_));
  AOI21_X1   g13027(.A1(new_n13201_), .A2(new_n13219_), .B(new_n2912_), .ZN(new_n13220_));
  NOR2_X1    g13028(.A1(new_n13204_), .A2(new_n13220_), .ZN(new_n13221_));
  AOI21_X1   g13029(.A1(new_n13221_), .A2(new_n2699_), .B(new_n12952_), .ZN(new_n13222_));
  OAI21_X1   g13030(.A1(new_n13204_), .A2(new_n13220_), .B(\asqrt[42] ), .ZN(new_n13223_));
  NAND2_X1   g13031(.A1(new_n13223_), .A2(new_n2464_), .ZN(new_n13224_));
  OAI21_X1   g13032(.A1(new_n13222_), .A2(new_n13224_), .B(new_n12948_), .ZN(new_n13225_));
  INV_X1     g13033(.I(new_n13223_), .ZN(new_n13226_));
  OAI21_X1   g13034(.A1(new_n13222_), .A2(new_n13226_), .B(\asqrt[43] ), .ZN(new_n13227_));
  NAND3_X1   g13035(.A1(new_n13225_), .A2(new_n13227_), .A3(new_n2271_), .ZN(new_n13228_));
  NAND2_X1   g13036(.A1(new_n13228_), .A2(new_n12946_), .ZN(new_n13229_));
  NAND2_X1   g13037(.A1(new_n13225_), .A2(new_n13227_), .ZN(new_n13230_));
  AOI21_X1   g13038(.A1(new_n13230_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n13231_));
  AOI21_X1   g13039(.A1(new_n13231_), .A2(new_n13229_), .B(new_n12943_), .ZN(new_n13232_));
  INV_X1     g13040(.I(new_n12948_), .ZN(new_n13233_));
  INV_X1     g13041(.I(new_n12958_), .ZN(new_n13234_));
  NOR2_X1    g13042(.A1(new_n13217_), .A2(new_n13218_), .ZN(new_n13235_));
  AOI21_X1   g13043(.A1(new_n13235_), .A2(new_n3167_), .B(new_n13234_), .ZN(new_n13236_));
  NAND2_X1   g13044(.A1(new_n13219_), .A2(new_n2912_), .ZN(new_n13237_));
  OAI21_X1   g13045(.A1(new_n13236_), .A2(new_n13237_), .B(new_n12954_), .ZN(new_n13238_));
  INV_X1     g13046(.I(new_n13219_), .ZN(new_n13239_));
  OAI21_X1   g13047(.A1(new_n13236_), .A2(new_n13239_), .B(\asqrt[41] ), .ZN(new_n13240_));
  NAND3_X1   g13048(.A1(new_n13238_), .A2(new_n13240_), .A3(new_n2699_), .ZN(new_n13241_));
  NAND2_X1   g13049(.A1(new_n13241_), .A2(new_n12951_), .ZN(new_n13242_));
  NAND2_X1   g13050(.A1(new_n13238_), .A2(new_n13240_), .ZN(new_n13243_));
  AOI21_X1   g13051(.A1(new_n13243_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n13244_));
  AOI21_X1   g13052(.A1(new_n13244_), .A2(new_n13242_), .B(new_n13233_), .ZN(new_n13245_));
  AOI21_X1   g13053(.A1(new_n13242_), .A2(new_n13223_), .B(new_n2464_), .ZN(new_n13246_));
  OAI21_X1   g13054(.A1(new_n13245_), .A2(new_n13246_), .B(\asqrt[44] ), .ZN(new_n13247_));
  AOI21_X1   g13055(.A1(new_n13229_), .A2(new_n13247_), .B(new_n2072_), .ZN(new_n13248_));
  NOR2_X1    g13056(.A1(new_n13232_), .A2(new_n13248_), .ZN(new_n13249_));
  AOI21_X1   g13057(.A1(new_n13249_), .A2(new_n1884_), .B(new_n12940_), .ZN(new_n13250_));
  OAI21_X1   g13058(.A1(new_n13232_), .A2(new_n13248_), .B(\asqrt[46] ), .ZN(new_n13251_));
  NAND2_X1   g13059(.A1(new_n13251_), .A2(new_n1688_), .ZN(new_n13252_));
  OAI21_X1   g13060(.A1(new_n13250_), .A2(new_n13252_), .B(new_n12936_), .ZN(new_n13253_));
  INV_X1     g13061(.I(new_n13251_), .ZN(new_n13254_));
  OAI21_X1   g13062(.A1(new_n13250_), .A2(new_n13254_), .B(\asqrt[47] ), .ZN(new_n13255_));
  NAND3_X1   g13063(.A1(new_n13253_), .A2(new_n13255_), .A3(new_n1533_), .ZN(new_n13256_));
  NAND2_X1   g13064(.A1(new_n13256_), .A2(new_n12934_), .ZN(new_n13257_));
  NAND2_X1   g13065(.A1(new_n13253_), .A2(new_n13255_), .ZN(new_n13258_));
  AOI21_X1   g13066(.A1(new_n13258_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n13259_));
  AOI21_X1   g13067(.A1(new_n13259_), .A2(new_n13257_), .B(new_n12931_), .ZN(new_n13260_));
  INV_X1     g13068(.I(new_n12936_), .ZN(new_n13261_));
  INV_X1     g13069(.I(new_n12946_), .ZN(new_n13262_));
  NOR2_X1    g13070(.A1(new_n13245_), .A2(new_n13246_), .ZN(new_n13263_));
  AOI21_X1   g13071(.A1(new_n13263_), .A2(new_n2271_), .B(new_n13262_), .ZN(new_n13264_));
  NAND2_X1   g13072(.A1(new_n13247_), .A2(new_n2072_), .ZN(new_n13265_));
  OAI21_X1   g13073(.A1(new_n13264_), .A2(new_n13265_), .B(new_n12942_), .ZN(new_n13266_));
  INV_X1     g13074(.I(new_n13247_), .ZN(new_n13267_));
  OAI21_X1   g13075(.A1(new_n13264_), .A2(new_n13267_), .B(\asqrt[45] ), .ZN(new_n13268_));
  NAND3_X1   g13076(.A1(new_n13266_), .A2(new_n13268_), .A3(new_n1884_), .ZN(new_n13269_));
  NAND2_X1   g13077(.A1(new_n13269_), .A2(new_n12939_), .ZN(new_n13270_));
  NAND2_X1   g13078(.A1(new_n13266_), .A2(new_n13268_), .ZN(new_n13271_));
  AOI21_X1   g13079(.A1(new_n13271_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n13272_));
  AOI21_X1   g13080(.A1(new_n13272_), .A2(new_n13270_), .B(new_n13261_), .ZN(new_n13273_));
  AOI21_X1   g13081(.A1(new_n13270_), .A2(new_n13251_), .B(new_n1688_), .ZN(new_n13274_));
  OAI21_X1   g13082(.A1(new_n13273_), .A2(new_n13274_), .B(\asqrt[48] ), .ZN(new_n13275_));
  AOI21_X1   g13083(.A1(new_n13257_), .A2(new_n13275_), .B(new_n1368_), .ZN(new_n13276_));
  NOR2_X1    g13084(.A1(new_n13260_), .A2(new_n13276_), .ZN(new_n13277_));
  AOI21_X1   g13085(.A1(new_n13277_), .A2(new_n1228_), .B(new_n12928_), .ZN(new_n13278_));
  OAI21_X1   g13086(.A1(new_n13260_), .A2(new_n13276_), .B(\asqrt[50] ), .ZN(new_n13279_));
  NAND2_X1   g13087(.A1(new_n13279_), .A2(new_n1088_), .ZN(new_n13280_));
  OAI21_X1   g13088(.A1(new_n13278_), .A2(new_n13280_), .B(new_n12872_), .ZN(new_n13281_));
  INV_X1     g13089(.I(new_n13279_), .ZN(new_n13282_));
  OAI21_X1   g13090(.A1(new_n13278_), .A2(new_n13282_), .B(\asqrt[51] ), .ZN(new_n13283_));
  NAND3_X1   g13091(.A1(new_n13281_), .A2(new_n13283_), .A3(new_n962_), .ZN(new_n13284_));
  NAND2_X1   g13092(.A1(new_n13284_), .A2(new_n12924_), .ZN(new_n13285_));
  NAND2_X1   g13093(.A1(new_n13281_), .A2(new_n13283_), .ZN(new_n13286_));
  AOI21_X1   g13094(.A1(new_n13286_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n13287_));
  AOI21_X1   g13095(.A1(new_n13287_), .A2(new_n13285_), .B(new_n12921_), .ZN(new_n13288_));
  INV_X1     g13096(.I(new_n12872_), .ZN(new_n13289_));
  INV_X1     g13097(.I(new_n12934_), .ZN(new_n13290_));
  NOR2_X1    g13098(.A1(new_n13273_), .A2(new_n13274_), .ZN(new_n13291_));
  AOI21_X1   g13099(.A1(new_n13291_), .A2(new_n1533_), .B(new_n13290_), .ZN(new_n13292_));
  NAND2_X1   g13100(.A1(new_n13275_), .A2(new_n1368_), .ZN(new_n13293_));
  OAI21_X1   g13101(.A1(new_n13292_), .A2(new_n13293_), .B(new_n12930_), .ZN(new_n13294_));
  INV_X1     g13102(.I(new_n13275_), .ZN(new_n13295_));
  OAI21_X1   g13103(.A1(new_n13292_), .A2(new_n13295_), .B(\asqrt[49] ), .ZN(new_n13296_));
  NAND3_X1   g13104(.A1(new_n13294_), .A2(new_n13296_), .A3(new_n1228_), .ZN(new_n13297_));
  NAND2_X1   g13105(.A1(new_n13297_), .A2(new_n12927_), .ZN(new_n13298_));
  NAND2_X1   g13106(.A1(new_n13294_), .A2(new_n13296_), .ZN(new_n13299_));
  AOI21_X1   g13107(.A1(new_n13299_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n13300_));
  AOI21_X1   g13108(.A1(new_n13300_), .A2(new_n13298_), .B(new_n13289_), .ZN(new_n13301_));
  AOI21_X1   g13109(.A1(new_n13298_), .A2(new_n13279_), .B(new_n1088_), .ZN(new_n13302_));
  OAI21_X1   g13110(.A1(new_n13301_), .A2(new_n13302_), .B(\asqrt[52] ), .ZN(new_n13303_));
  AOI21_X1   g13111(.A1(new_n13285_), .A2(new_n13303_), .B(new_n842_), .ZN(new_n13304_));
  NOR2_X1    g13112(.A1(new_n13288_), .A2(new_n13304_), .ZN(new_n13305_));
  AOI21_X1   g13113(.A1(new_n13305_), .A2(new_n720_), .B(new_n12918_), .ZN(new_n13306_));
  OAI21_X1   g13114(.A1(new_n13288_), .A2(new_n13304_), .B(\asqrt[54] ), .ZN(new_n13307_));
  NAND2_X1   g13115(.A1(new_n13307_), .A2(new_n630_), .ZN(new_n13308_));
  OAI21_X1   g13116(.A1(new_n13306_), .A2(new_n13308_), .B(new_n12914_), .ZN(new_n13309_));
  INV_X1     g13117(.I(new_n13307_), .ZN(new_n13310_));
  OAI21_X1   g13118(.A1(new_n13306_), .A2(new_n13310_), .B(\asqrt[55] ), .ZN(new_n13311_));
  NAND3_X1   g13119(.A1(new_n13309_), .A2(new_n13311_), .A3(new_n545_), .ZN(new_n13312_));
  NAND2_X1   g13120(.A1(new_n13312_), .A2(new_n12912_), .ZN(new_n13313_));
  NAND2_X1   g13121(.A1(new_n13309_), .A2(new_n13311_), .ZN(new_n13314_));
  AOI21_X1   g13122(.A1(new_n13314_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n13315_));
  AOI21_X1   g13123(.A1(new_n13315_), .A2(new_n13313_), .B(new_n12909_), .ZN(new_n13316_));
  INV_X1     g13124(.I(new_n12914_), .ZN(new_n13317_));
  INV_X1     g13125(.I(new_n12924_), .ZN(new_n13318_));
  NOR2_X1    g13126(.A1(new_n13301_), .A2(new_n13302_), .ZN(new_n13319_));
  AOI21_X1   g13127(.A1(new_n13319_), .A2(new_n962_), .B(new_n13318_), .ZN(new_n13320_));
  NAND2_X1   g13128(.A1(new_n13303_), .A2(new_n842_), .ZN(new_n13321_));
  OAI21_X1   g13129(.A1(new_n13320_), .A2(new_n13321_), .B(new_n12920_), .ZN(new_n13322_));
  INV_X1     g13130(.I(new_n13303_), .ZN(new_n13323_));
  OAI21_X1   g13131(.A1(new_n13320_), .A2(new_n13323_), .B(\asqrt[53] ), .ZN(new_n13324_));
  NAND3_X1   g13132(.A1(new_n13322_), .A2(new_n13324_), .A3(new_n720_), .ZN(new_n13325_));
  NAND2_X1   g13133(.A1(new_n13325_), .A2(new_n12917_), .ZN(new_n13326_));
  NAND2_X1   g13134(.A1(new_n13322_), .A2(new_n13324_), .ZN(new_n13327_));
  AOI21_X1   g13135(.A1(new_n13327_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n13328_));
  AOI21_X1   g13136(.A1(new_n13328_), .A2(new_n13326_), .B(new_n13317_), .ZN(new_n13329_));
  AOI21_X1   g13137(.A1(new_n13326_), .A2(new_n13307_), .B(new_n630_), .ZN(new_n13330_));
  OAI21_X1   g13138(.A1(new_n13329_), .A2(new_n13330_), .B(\asqrt[56] ), .ZN(new_n13331_));
  AOI21_X1   g13139(.A1(new_n13313_), .A2(new_n13331_), .B(new_n450_), .ZN(new_n13332_));
  NOR2_X1    g13140(.A1(new_n13316_), .A2(new_n13332_), .ZN(new_n13333_));
  AOI21_X1   g13141(.A1(new_n13333_), .A2(new_n403_), .B(new_n12906_), .ZN(new_n13334_));
  OAI21_X1   g13142(.A1(new_n13316_), .A2(new_n13332_), .B(\asqrt[58] ), .ZN(new_n13335_));
  NAND2_X1   g13143(.A1(new_n13335_), .A2(new_n339_), .ZN(new_n13336_));
  OAI21_X1   g13144(.A1(new_n13334_), .A2(new_n13336_), .B(new_n12902_), .ZN(new_n13337_));
  INV_X1     g13145(.I(new_n13335_), .ZN(new_n13338_));
  OAI21_X1   g13146(.A1(new_n13334_), .A2(new_n13338_), .B(\asqrt[59] ), .ZN(new_n13339_));
  NAND3_X1   g13147(.A1(new_n13337_), .A2(new_n13339_), .A3(new_n288_), .ZN(new_n13340_));
  NAND2_X1   g13148(.A1(new_n13340_), .A2(new_n12900_), .ZN(new_n13341_));
  INV_X1     g13149(.I(new_n12902_), .ZN(new_n13342_));
  INV_X1     g13150(.I(new_n12912_), .ZN(new_n13343_));
  NOR2_X1    g13151(.A1(new_n13329_), .A2(new_n13330_), .ZN(new_n13344_));
  AOI21_X1   g13152(.A1(new_n13344_), .A2(new_n545_), .B(new_n13343_), .ZN(new_n13345_));
  NAND2_X1   g13153(.A1(new_n13331_), .A2(new_n450_), .ZN(new_n13346_));
  OAI21_X1   g13154(.A1(new_n13345_), .A2(new_n13346_), .B(new_n12908_), .ZN(new_n13347_));
  INV_X1     g13155(.I(new_n13331_), .ZN(new_n13348_));
  OAI21_X1   g13156(.A1(new_n13345_), .A2(new_n13348_), .B(\asqrt[57] ), .ZN(new_n13349_));
  NAND3_X1   g13157(.A1(new_n13347_), .A2(new_n13349_), .A3(new_n403_), .ZN(new_n13350_));
  NAND2_X1   g13158(.A1(new_n13350_), .A2(new_n12905_), .ZN(new_n13351_));
  NAND2_X1   g13159(.A1(new_n13347_), .A2(new_n13349_), .ZN(new_n13352_));
  AOI21_X1   g13160(.A1(new_n13352_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n13353_));
  AOI21_X1   g13161(.A1(new_n13353_), .A2(new_n13351_), .B(new_n13342_), .ZN(new_n13354_));
  AOI21_X1   g13162(.A1(new_n13351_), .A2(new_n13335_), .B(new_n339_), .ZN(new_n13355_));
  OAI21_X1   g13163(.A1(new_n13354_), .A2(new_n13355_), .B(\asqrt[60] ), .ZN(new_n13356_));
  AOI21_X1   g13164(.A1(new_n13341_), .A2(new_n13356_), .B(new_n242_), .ZN(new_n13357_));
  NAND3_X1   g13165(.A1(\asqrt[14] ), .A2(new_n12832_), .A3(new_n12848_), .ZN(new_n13358_));
  XOR2_X1    g13166(.A1(new_n13358_), .A2(new_n12873_), .Z(new_n13359_));
  INV_X1     g13167(.I(new_n13359_), .ZN(new_n13360_));
  NAND2_X1   g13168(.A1(new_n13337_), .A2(new_n13339_), .ZN(new_n13361_));
  AOI21_X1   g13169(.A1(new_n13361_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n13362_));
  AOI21_X1   g13170(.A1(new_n13362_), .A2(new_n13341_), .B(new_n13360_), .ZN(new_n13363_));
  OAI21_X1   g13171(.A1(new_n13363_), .A2(new_n13357_), .B(\asqrt[62] ), .ZN(new_n13364_));
  AOI21_X1   g13172(.A1(new_n12833_), .A2(new_n12854_), .B(new_n12849_), .ZN(new_n13365_));
  NAND2_X1   g13173(.A1(\asqrt[14] ), .A2(new_n13365_), .ZN(new_n13366_));
  XOR2_X1    g13174(.A1(new_n13366_), .A2(new_n12852_), .Z(new_n13367_));
  INV_X1     g13175(.I(new_n12900_), .ZN(new_n13368_));
  NOR2_X1    g13176(.A1(new_n13354_), .A2(new_n13355_), .ZN(new_n13369_));
  AOI21_X1   g13177(.A1(new_n13369_), .A2(new_n288_), .B(new_n13368_), .ZN(new_n13370_));
  INV_X1     g13178(.I(new_n13356_), .ZN(new_n13371_));
  OAI21_X1   g13179(.A1(new_n13370_), .A2(new_n13371_), .B(\asqrt[61] ), .ZN(new_n13372_));
  NAND2_X1   g13180(.A1(new_n13356_), .A2(new_n242_), .ZN(new_n13373_));
  OAI21_X1   g13181(.A1(new_n13370_), .A2(new_n13373_), .B(new_n13359_), .ZN(new_n13374_));
  NAND3_X1   g13182(.A1(new_n13374_), .A2(new_n13372_), .A3(new_n234_), .ZN(new_n13375_));
  NAND2_X1   g13183(.A1(new_n13375_), .A2(new_n13367_), .ZN(new_n13376_));
  AOI21_X1   g13184(.A1(new_n13376_), .A2(new_n13364_), .B(new_n12897_), .ZN(new_n13377_));
  AOI21_X1   g13185(.A1(new_n13377_), .A2(new_n12895_), .B(\asqrt[63] ), .ZN(new_n13378_));
  NAND2_X1   g13186(.A1(new_n13376_), .A2(new_n13364_), .ZN(new_n13379_));
  NOR2_X1    g13187(.A1(new_n13379_), .A2(new_n12895_), .ZN(new_n13380_));
  NOR2_X1    g13188(.A1(\asqrt[14] ), .A2(new_n12884_), .ZN(new_n13381_));
  NOR4_X1    g13189(.A1(new_n13378_), .A2(new_n12892_), .A3(new_n13380_), .A4(new_n13381_), .ZN(new_n13382_));
  OAI21_X1   g13190(.A1(new_n13278_), .A2(new_n13280_), .B(new_n13283_), .ZN(new_n13383_));
  NOR2_X1    g13191(.A1(new_n13382_), .A2(new_n13383_), .ZN(new_n13384_));
  XOR2_X1    g13192(.A1(new_n13384_), .A2(new_n12872_), .Z(new_n13385_));
  INV_X1     g13193(.I(new_n13385_), .ZN(new_n13386_));
  INV_X1     g13194(.I(new_n12892_), .ZN(new_n13387_));
  INV_X1     g13195(.I(new_n13364_), .ZN(new_n13388_));
  NOR2_X1    g13196(.A1(new_n13363_), .A2(new_n13357_), .ZN(new_n13389_));
  INV_X1     g13197(.I(new_n13367_), .ZN(new_n13390_));
  AOI21_X1   g13198(.A1(new_n13389_), .A2(new_n234_), .B(new_n13390_), .ZN(new_n13391_));
  OAI21_X1   g13199(.A1(new_n13391_), .A2(new_n13388_), .B(new_n12896_), .ZN(new_n13392_));
  OAI21_X1   g13200(.A1(new_n13392_), .A2(new_n12894_), .B(new_n193_), .ZN(new_n13393_));
  NOR2_X1    g13201(.A1(new_n13391_), .A2(new_n13388_), .ZN(new_n13394_));
  NAND2_X1   g13202(.A1(new_n13394_), .A2(new_n12894_), .ZN(new_n13395_));
  INV_X1     g13203(.I(new_n13381_), .ZN(new_n13396_));
  NAND4_X1   g13204(.A1(new_n13393_), .A2(new_n13387_), .A3(new_n13395_), .A4(new_n13396_), .ZN(\asqrt[13] ));
  NAND3_X1   g13205(.A1(\asqrt[13] ), .A2(new_n13297_), .A3(new_n13279_), .ZN(new_n13398_));
  XOR2_X1    g13206(.A1(new_n13398_), .A2(new_n12928_), .Z(new_n13399_));
  OAI21_X1   g13207(.A1(new_n13292_), .A2(new_n13293_), .B(new_n13296_), .ZN(new_n13400_));
  NOR2_X1    g13208(.A1(new_n13382_), .A2(new_n13400_), .ZN(new_n13401_));
  XOR2_X1    g13209(.A1(new_n13401_), .A2(new_n12930_), .Z(new_n13402_));
  INV_X1     g13210(.I(new_n13402_), .ZN(new_n13403_));
  NAND3_X1   g13211(.A1(\asqrt[13] ), .A2(new_n13256_), .A3(new_n13275_), .ZN(new_n13404_));
  XOR2_X1    g13212(.A1(new_n13404_), .A2(new_n13290_), .Z(new_n13405_));
  INV_X1     g13213(.I(new_n13405_), .ZN(new_n13406_));
  OAI21_X1   g13214(.A1(new_n13250_), .A2(new_n13252_), .B(new_n13255_), .ZN(new_n13407_));
  NOR2_X1    g13215(.A1(new_n13382_), .A2(new_n13407_), .ZN(new_n13408_));
  XOR2_X1    g13216(.A1(new_n13408_), .A2(new_n12936_), .Z(new_n13409_));
  NAND3_X1   g13217(.A1(\asqrt[13] ), .A2(new_n13269_), .A3(new_n13251_), .ZN(new_n13410_));
  XOR2_X1    g13218(.A1(new_n13410_), .A2(new_n12940_), .Z(new_n13411_));
  OAI21_X1   g13219(.A1(new_n13264_), .A2(new_n13265_), .B(new_n13268_), .ZN(new_n13412_));
  NOR2_X1    g13220(.A1(new_n13382_), .A2(new_n13412_), .ZN(new_n13413_));
  XOR2_X1    g13221(.A1(new_n13413_), .A2(new_n12942_), .Z(new_n13414_));
  INV_X1     g13222(.I(new_n13414_), .ZN(new_n13415_));
  NAND3_X1   g13223(.A1(\asqrt[13] ), .A2(new_n13228_), .A3(new_n13247_), .ZN(new_n13416_));
  XOR2_X1    g13224(.A1(new_n13416_), .A2(new_n13262_), .Z(new_n13417_));
  INV_X1     g13225(.I(new_n13417_), .ZN(new_n13418_));
  OAI21_X1   g13226(.A1(new_n13222_), .A2(new_n13224_), .B(new_n13227_), .ZN(new_n13419_));
  NOR2_X1    g13227(.A1(new_n13382_), .A2(new_n13419_), .ZN(new_n13420_));
  XOR2_X1    g13228(.A1(new_n13420_), .A2(new_n12948_), .Z(new_n13421_));
  NAND3_X1   g13229(.A1(\asqrt[13] ), .A2(new_n13241_), .A3(new_n13223_), .ZN(new_n13422_));
  XOR2_X1    g13230(.A1(new_n13422_), .A2(new_n12952_), .Z(new_n13423_));
  OAI21_X1   g13231(.A1(new_n13236_), .A2(new_n13237_), .B(new_n13240_), .ZN(new_n13424_));
  NOR2_X1    g13232(.A1(new_n13382_), .A2(new_n13424_), .ZN(new_n13425_));
  XOR2_X1    g13233(.A1(new_n13425_), .A2(new_n12954_), .Z(new_n13426_));
  INV_X1     g13234(.I(new_n13426_), .ZN(new_n13427_));
  NAND3_X1   g13235(.A1(\asqrt[13] ), .A2(new_n13200_), .A3(new_n13219_), .ZN(new_n13428_));
  XOR2_X1    g13236(.A1(new_n13428_), .A2(new_n13234_), .Z(new_n13429_));
  INV_X1     g13237(.I(new_n13429_), .ZN(new_n13430_));
  OAI21_X1   g13238(.A1(new_n13194_), .A2(new_n13196_), .B(new_n13199_), .ZN(new_n13431_));
  NOR2_X1    g13239(.A1(new_n13382_), .A2(new_n13431_), .ZN(new_n13432_));
  XOR2_X1    g13240(.A1(new_n13432_), .A2(new_n12960_), .Z(new_n13433_));
  NAND3_X1   g13241(.A1(\asqrt[13] ), .A2(new_n13213_), .A3(new_n13195_), .ZN(new_n13434_));
  XOR2_X1    g13242(.A1(new_n13434_), .A2(new_n12964_), .Z(new_n13435_));
  OAI21_X1   g13243(.A1(new_n13208_), .A2(new_n13209_), .B(new_n13212_), .ZN(new_n13436_));
  NOR2_X1    g13244(.A1(new_n13382_), .A2(new_n13436_), .ZN(new_n13437_));
  XOR2_X1    g13245(.A1(new_n13437_), .A2(new_n12966_), .Z(new_n13438_));
  INV_X1     g13246(.I(new_n13438_), .ZN(new_n13439_));
  NAND3_X1   g13247(.A1(\asqrt[13] ), .A2(new_n13172_), .A3(new_n13191_), .ZN(new_n13440_));
  XOR2_X1    g13248(.A1(new_n13440_), .A2(new_n13206_), .Z(new_n13441_));
  INV_X1     g13249(.I(new_n13441_), .ZN(new_n13442_));
  OAI21_X1   g13250(.A1(new_n13166_), .A2(new_n13168_), .B(new_n13171_), .ZN(new_n13443_));
  NOR2_X1    g13251(.A1(new_n13382_), .A2(new_n13443_), .ZN(new_n13444_));
  XOR2_X1    g13252(.A1(new_n13444_), .A2(new_n12972_), .Z(new_n13445_));
  NAND3_X1   g13253(.A1(\asqrt[13] ), .A2(new_n13185_), .A3(new_n13167_), .ZN(new_n13446_));
  XOR2_X1    g13254(.A1(new_n13446_), .A2(new_n12976_), .Z(new_n13447_));
  OAI21_X1   g13255(.A1(new_n13180_), .A2(new_n13181_), .B(new_n13184_), .ZN(new_n13448_));
  NOR2_X1    g13256(.A1(new_n13382_), .A2(new_n13448_), .ZN(new_n13449_));
  XOR2_X1    g13257(.A1(new_n13449_), .A2(new_n12978_), .Z(new_n13450_));
  INV_X1     g13258(.I(new_n13450_), .ZN(new_n13451_));
  NAND3_X1   g13259(.A1(\asqrt[13] ), .A2(new_n13144_), .A3(new_n13163_), .ZN(new_n13452_));
  XOR2_X1    g13260(.A1(new_n13452_), .A2(new_n13178_), .Z(new_n13453_));
  INV_X1     g13261(.I(new_n13453_), .ZN(new_n13454_));
  OAI21_X1   g13262(.A1(new_n13138_), .A2(new_n13140_), .B(new_n13143_), .ZN(new_n13455_));
  NOR2_X1    g13263(.A1(new_n13382_), .A2(new_n13455_), .ZN(new_n13456_));
  XOR2_X1    g13264(.A1(new_n13456_), .A2(new_n12984_), .Z(new_n13457_));
  NAND3_X1   g13265(.A1(\asqrt[13] ), .A2(new_n13157_), .A3(new_n13139_), .ZN(new_n13458_));
  XOR2_X1    g13266(.A1(new_n13458_), .A2(new_n12988_), .Z(new_n13459_));
  OAI21_X1   g13267(.A1(new_n13152_), .A2(new_n13153_), .B(new_n13156_), .ZN(new_n13460_));
  NOR2_X1    g13268(.A1(new_n13382_), .A2(new_n13460_), .ZN(new_n13461_));
  XOR2_X1    g13269(.A1(new_n13461_), .A2(new_n12990_), .Z(new_n13462_));
  INV_X1     g13270(.I(new_n13462_), .ZN(new_n13463_));
  NAND3_X1   g13271(.A1(\asqrt[13] ), .A2(new_n13116_), .A3(new_n13135_), .ZN(new_n13464_));
  XOR2_X1    g13272(.A1(new_n13464_), .A2(new_n13150_), .Z(new_n13465_));
  INV_X1     g13273(.I(new_n13465_), .ZN(new_n13466_));
  OAI21_X1   g13274(.A1(new_n13110_), .A2(new_n13112_), .B(new_n13115_), .ZN(new_n13467_));
  NOR2_X1    g13275(.A1(new_n13382_), .A2(new_n13467_), .ZN(new_n13468_));
  XOR2_X1    g13276(.A1(new_n13468_), .A2(new_n12996_), .Z(new_n13469_));
  NAND3_X1   g13277(.A1(\asqrt[13] ), .A2(new_n13129_), .A3(new_n13111_), .ZN(new_n13470_));
  XOR2_X1    g13278(.A1(new_n13470_), .A2(new_n13000_), .Z(new_n13471_));
  OAI21_X1   g13279(.A1(new_n13124_), .A2(new_n13125_), .B(new_n13128_), .ZN(new_n13472_));
  NOR2_X1    g13280(.A1(new_n13382_), .A2(new_n13472_), .ZN(new_n13473_));
  XOR2_X1    g13281(.A1(new_n13473_), .A2(new_n13002_), .Z(new_n13474_));
  INV_X1     g13282(.I(new_n13474_), .ZN(new_n13475_));
  NAND3_X1   g13283(.A1(\asqrt[13] ), .A2(new_n13088_), .A3(new_n13107_), .ZN(new_n13476_));
  XOR2_X1    g13284(.A1(new_n13476_), .A2(new_n13122_), .Z(new_n13477_));
  INV_X1     g13285(.I(new_n13477_), .ZN(new_n13478_));
  OAI21_X1   g13286(.A1(new_n13082_), .A2(new_n13084_), .B(new_n13087_), .ZN(new_n13479_));
  NOR2_X1    g13287(.A1(new_n13382_), .A2(new_n13479_), .ZN(new_n13480_));
  XOR2_X1    g13288(.A1(new_n13480_), .A2(new_n13008_), .Z(new_n13481_));
  NAND3_X1   g13289(.A1(\asqrt[13] ), .A2(new_n13101_), .A3(new_n13083_), .ZN(new_n13482_));
  XOR2_X1    g13290(.A1(new_n13482_), .A2(new_n13012_), .Z(new_n13483_));
  OAI21_X1   g13291(.A1(new_n13096_), .A2(new_n13097_), .B(new_n13100_), .ZN(new_n13484_));
  NOR2_X1    g13292(.A1(new_n13382_), .A2(new_n13484_), .ZN(new_n13485_));
  XOR2_X1    g13293(.A1(new_n13485_), .A2(new_n13014_), .Z(new_n13486_));
  INV_X1     g13294(.I(new_n13486_), .ZN(new_n13487_));
  NAND3_X1   g13295(.A1(\asqrt[13] ), .A2(new_n13053_), .A3(new_n13079_), .ZN(new_n13488_));
  XOR2_X1    g13296(.A1(new_n13488_), .A2(new_n13094_), .Z(new_n13489_));
  INV_X1     g13297(.I(new_n13489_), .ZN(new_n13490_));
  AOI21_X1   g13298(.A1(new_n13074_), .A2(new_n13075_), .B(new_n13078_), .ZN(new_n13491_));
  NAND2_X1   g13299(.A1(\asqrt[13] ), .A2(new_n13491_), .ZN(new_n13492_));
  XOR2_X1    g13300(.A1(new_n13492_), .A2(new_n13058_), .Z(new_n13493_));
  NOR2_X1    g13301(.A1(new_n13073_), .A2(\asqrt[18] ), .ZN(new_n13494_));
  NOR3_X1    g13302(.A1(new_n13382_), .A2(new_n13494_), .A3(new_n13051_), .ZN(new_n13495_));
  XOR2_X1    g13303(.A1(new_n13495_), .A2(new_n13023_), .Z(new_n13496_));
  NOR3_X1    g13304(.A1(new_n13382_), .A2(new_n13070_), .A3(new_n13046_), .ZN(new_n13497_));
  XOR2_X1    g13305(.A1(new_n13497_), .A2(new_n13045_), .Z(new_n13498_));
  INV_X1     g13306(.I(new_n13498_), .ZN(new_n13499_));
  NOR2_X1    g13307(.A1(new_n13040_), .A2(\asqrt[16] ), .ZN(new_n13500_));
  NOR3_X1    g13308(.A1(new_n13382_), .A2(new_n13500_), .A3(new_n13069_), .ZN(new_n13501_));
  XOR2_X1    g13309(.A1(new_n13501_), .A2(new_n13031_), .Z(new_n13502_));
  INV_X1     g13310(.I(new_n13502_), .ZN(new_n13503_));
  NAND3_X1   g13311(.A1(\asqrt[13] ), .A2(new_n13032_), .A3(new_n13033_), .ZN(new_n13504_));
  NOR4_X1    g13312(.A1(new_n13378_), .A2(new_n12889_), .A3(new_n12892_), .A4(new_n13380_), .ZN(new_n13505_));
  INV_X1     g13313(.I(new_n13505_), .ZN(new_n13506_));
  AOI21_X1   g13314(.A1(new_n13504_), .A2(new_n13506_), .B(\a[28] ), .ZN(new_n13507_));
  NOR3_X1    g13315(.A1(new_n13382_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n13508_));
  NOR3_X1    g13316(.A1(new_n13508_), .A2(new_n12491_), .A3(new_n13505_), .ZN(new_n13509_));
  NOR2_X1    g13317(.A1(new_n13509_), .A2(new_n13507_), .ZN(new_n13510_));
  INV_X1     g13318(.I(\a[24] ), .ZN(new_n13511_));
  INV_X1     g13319(.I(\a[25] ), .ZN(new_n13512_));
  NAND3_X1   g13320(.A1(new_n13511_), .A2(new_n13512_), .A3(new_n13032_), .ZN(new_n13513_));
  OAI21_X1   g13321(.A1(new_n13382_), .A2(new_n13032_), .B(new_n13513_), .ZN(new_n13514_));
  NAND2_X1   g13322(.A1(new_n13514_), .A2(\asqrt[14] ), .ZN(new_n13515_));
  OAI21_X1   g13323(.A1(new_n13382_), .A2(\a[26] ), .B(\a[27] ), .ZN(new_n13516_));
  NAND2_X1   g13324(.A1(new_n13516_), .A2(new_n13504_), .ZN(new_n13517_));
  NOR2_X1    g13325(.A1(new_n13514_), .A2(\asqrt[14] ), .ZN(new_n13518_));
  OAI21_X1   g13326(.A1(new_n13517_), .A2(new_n13518_), .B(new_n13515_), .ZN(new_n13519_));
  OAI21_X1   g13327(.A1(\asqrt[15] ), .A2(new_n13519_), .B(new_n13510_), .ZN(new_n13520_));
  NAND2_X1   g13328(.A1(new_n13519_), .A2(\asqrt[15] ), .ZN(new_n13521_));
  NAND3_X1   g13329(.A1(new_n13520_), .A2(new_n11901_), .A3(new_n13521_), .ZN(new_n13522_));
  NOR3_X1    g13330(.A1(new_n13382_), .A2(new_n13063_), .A3(new_n13039_), .ZN(new_n13523_));
  XOR2_X1    g13331(.A1(new_n13523_), .A2(new_n13065_), .Z(new_n13524_));
  NAND2_X1   g13332(.A1(new_n13522_), .A2(new_n13524_), .ZN(new_n13525_));
  NAND2_X1   g13333(.A1(new_n13520_), .A2(new_n13521_), .ZN(new_n13526_));
  AOI21_X1   g13334(.A1(new_n13526_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n13527_));
  AOI21_X1   g13335(.A1(new_n13527_), .A2(new_n13525_), .B(new_n13503_), .ZN(new_n13528_));
  OAI21_X1   g13336(.A1(new_n13508_), .A2(new_n13505_), .B(new_n12491_), .ZN(new_n13529_));
  NAND3_X1   g13337(.A1(new_n13504_), .A2(\a[28] ), .A3(new_n13506_), .ZN(new_n13530_));
  NAND2_X1   g13338(.A1(new_n13529_), .A2(new_n13530_), .ZN(new_n13531_));
  NAND2_X1   g13339(.A1(\asqrt[13] ), .A2(\a[26] ), .ZN(new_n13532_));
  AOI21_X1   g13340(.A1(new_n13532_), .A2(new_n13513_), .B(new_n12889_), .ZN(new_n13533_));
  AOI21_X1   g13341(.A1(\asqrt[13] ), .A2(new_n13032_), .B(new_n13033_), .ZN(new_n13534_));
  NOR2_X1    g13342(.A1(new_n13534_), .A2(new_n13508_), .ZN(new_n13535_));
  NAND3_X1   g13343(.A1(new_n13532_), .A2(new_n12889_), .A3(new_n13513_), .ZN(new_n13536_));
  AOI21_X1   g13344(.A1(new_n13535_), .A2(new_n13536_), .B(new_n13533_), .ZN(new_n13537_));
  AOI21_X1   g13345(.A1(new_n13537_), .A2(new_n12374_), .B(new_n13531_), .ZN(new_n13538_));
  NOR2_X1    g13346(.A1(new_n13537_), .A2(new_n12374_), .ZN(new_n13539_));
  OAI21_X1   g13347(.A1(new_n13538_), .A2(new_n13539_), .B(\asqrt[16] ), .ZN(new_n13540_));
  AOI21_X1   g13348(.A1(new_n13525_), .A2(new_n13540_), .B(new_n11406_), .ZN(new_n13541_));
  NOR2_X1    g13349(.A1(new_n13528_), .A2(new_n13541_), .ZN(new_n13542_));
  AOI21_X1   g13350(.A1(new_n13542_), .A2(new_n10953_), .B(new_n13499_), .ZN(new_n13543_));
  OAI21_X1   g13351(.A1(new_n13528_), .A2(new_n13541_), .B(\asqrt[18] ), .ZN(new_n13544_));
  NAND2_X1   g13352(.A1(new_n13544_), .A2(new_n10478_), .ZN(new_n13545_));
  OAI21_X1   g13353(.A1(new_n13543_), .A2(new_n13545_), .B(new_n13496_), .ZN(new_n13546_));
  INV_X1     g13354(.I(new_n13544_), .ZN(new_n13547_));
  OAI21_X1   g13355(.A1(new_n13543_), .A2(new_n13547_), .B(\asqrt[19] ), .ZN(new_n13548_));
  NAND3_X1   g13356(.A1(new_n13546_), .A2(new_n13548_), .A3(new_n10045_), .ZN(new_n13549_));
  NAND2_X1   g13357(.A1(new_n13549_), .A2(new_n13493_), .ZN(new_n13550_));
  NAND2_X1   g13358(.A1(new_n13546_), .A2(new_n13548_), .ZN(new_n13551_));
  AOI21_X1   g13359(.A1(new_n13551_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n13552_));
  AOI21_X1   g13360(.A1(new_n13552_), .A2(new_n13550_), .B(new_n13490_), .ZN(new_n13553_));
  INV_X1     g13361(.I(new_n13496_), .ZN(new_n13554_));
  NOR2_X1    g13362(.A1(new_n13538_), .A2(new_n13539_), .ZN(new_n13555_));
  INV_X1     g13363(.I(new_n13524_), .ZN(new_n13556_));
  AOI21_X1   g13364(.A1(new_n13555_), .A2(new_n11901_), .B(new_n13556_), .ZN(new_n13557_));
  NAND2_X1   g13365(.A1(new_n13540_), .A2(new_n11406_), .ZN(new_n13558_));
  OAI21_X1   g13366(.A1(new_n13557_), .A2(new_n13558_), .B(new_n13502_), .ZN(new_n13559_));
  INV_X1     g13367(.I(new_n13540_), .ZN(new_n13560_));
  OAI21_X1   g13368(.A1(new_n13557_), .A2(new_n13560_), .B(\asqrt[17] ), .ZN(new_n13561_));
  NAND3_X1   g13369(.A1(new_n13559_), .A2(new_n13561_), .A3(new_n10953_), .ZN(new_n13562_));
  NAND2_X1   g13370(.A1(new_n13562_), .A2(new_n13498_), .ZN(new_n13563_));
  NAND2_X1   g13371(.A1(new_n13559_), .A2(new_n13561_), .ZN(new_n13564_));
  AOI21_X1   g13372(.A1(new_n13564_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n13565_));
  AOI21_X1   g13373(.A1(new_n13565_), .A2(new_n13563_), .B(new_n13554_), .ZN(new_n13566_));
  AOI21_X1   g13374(.A1(new_n13563_), .A2(new_n13544_), .B(new_n10478_), .ZN(new_n13567_));
  OAI21_X1   g13375(.A1(new_n13566_), .A2(new_n13567_), .B(\asqrt[20] ), .ZN(new_n13568_));
  AOI21_X1   g13376(.A1(new_n13550_), .A2(new_n13568_), .B(new_n9590_), .ZN(new_n13569_));
  NOR2_X1    g13377(.A1(new_n13553_), .A2(new_n13569_), .ZN(new_n13570_));
  AOI21_X1   g13378(.A1(new_n13570_), .A2(new_n9177_), .B(new_n13487_), .ZN(new_n13571_));
  OAI21_X1   g13379(.A1(new_n13553_), .A2(new_n13569_), .B(\asqrt[22] ), .ZN(new_n13572_));
  NAND2_X1   g13380(.A1(new_n13572_), .A2(new_n8742_), .ZN(new_n13573_));
  OAI21_X1   g13381(.A1(new_n13571_), .A2(new_n13573_), .B(new_n13483_), .ZN(new_n13574_));
  INV_X1     g13382(.I(new_n13572_), .ZN(new_n13575_));
  OAI21_X1   g13383(.A1(new_n13571_), .A2(new_n13575_), .B(\asqrt[23] ), .ZN(new_n13576_));
  NAND3_X1   g13384(.A1(new_n13574_), .A2(new_n13576_), .A3(new_n8349_), .ZN(new_n13577_));
  NAND2_X1   g13385(.A1(new_n13577_), .A2(new_n13481_), .ZN(new_n13578_));
  NAND2_X1   g13386(.A1(new_n13574_), .A2(new_n13576_), .ZN(new_n13579_));
  AOI21_X1   g13387(.A1(new_n13579_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n13580_));
  AOI21_X1   g13388(.A1(new_n13580_), .A2(new_n13578_), .B(new_n13478_), .ZN(new_n13581_));
  INV_X1     g13389(.I(new_n13483_), .ZN(new_n13582_));
  INV_X1     g13390(.I(new_n13493_), .ZN(new_n13583_));
  NOR2_X1    g13391(.A1(new_n13566_), .A2(new_n13567_), .ZN(new_n13584_));
  AOI21_X1   g13392(.A1(new_n13584_), .A2(new_n10045_), .B(new_n13583_), .ZN(new_n13585_));
  NAND2_X1   g13393(.A1(new_n13568_), .A2(new_n9590_), .ZN(new_n13586_));
  OAI21_X1   g13394(.A1(new_n13585_), .A2(new_n13586_), .B(new_n13489_), .ZN(new_n13587_));
  INV_X1     g13395(.I(new_n13568_), .ZN(new_n13588_));
  OAI21_X1   g13396(.A1(new_n13585_), .A2(new_n13588_), .B(\asqrt[21] ), .ZN(new_n13589_));
  NAND3_X1   g13397(.A1(new_n13587_), .A2(new_n13589_), .A3(new_n9177_), .ZN(new_n13590_));
  NAND2_X1   g13398(.A1(new_n13590_), .A2(new_n13486_), .ZN(new_n13591_));
  NAND2_X1   g13399(.A1(new_n13587_), .A2(new_n13589_), .ZN(new_n13592_));
  AOI21_X1   g13400(.A1(new_n13592_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n13593_));
  AOI21_X1   g13401(.A1(new_n13593_), .A2(new_n13591_), .B(new_n13582_), .ZN(new_n13594_));
  AOI21_X1   g13402(.A1(new_n13591_), .A2(new_n13572_), .B(new_n8742_), .ZN(new_n13595_));
  OAI21_X1   g13403(.A1(new_n13594_), .A2(new_n13595_), .B(\asqrt[24] ), .ZN(new_n13596_));
  AOI21_X1   g13404(.A1(new_n13578_), .A2(new_n13596_), .B(new_n7934_), .ZN(new_n13597_));
  NOR2_X1    g13405(.A1(new_n13581_), .A2(new_n13597_), .ZN(new_n13598_));
  AOI21_X1   g13406(.A1(new_n13598_), .A2(new_n7561_), .B(new_n13475_), .ZN(new_n13599_));
  OAI21_X1   g13407(.A1(new_n13581_), .A2(new_n13597_), .B(\asqrt[26] ), .ZN(new_n13600_));
  NAND2_X1   g13408(.A1(new_n13600_), .A2(new_n7166_), .ZN(new_n13601_));
  OAI21_X1   g13409(.A1(new_n13599_), .A2(new_n13601_), .B(new_n13471_), .ZN(new_n13602_));
  INV_X1     g13410(.I(new_n13600_), .ZN(new_n13603_));
  OAI21_X1   g13411(.A1(new_n13599_), .A2(new_n13603_), .B(\asqrt[27] ), .ZN(new_n13604_));
  NAND3_X1   g13412(.A1(new_n13602_), .A2(new_n13604_), .A3(new_n6813_), .ZN(new_n13605_));
  NAND2_X1   g13413(.A1(new_n13605_), .A2(new_n13469_), .ZN(new_n13606_));
  NAND2_X1   g13414(.A1(new_n13602_), .A2(new_n13604_), .ZN(new_n13607_));
  AOI21_X1   g13415(.A1(new_n13607_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n13608_));
  AOI21_X1   g13416(.A1(new_n13608_), .A2(new_n13606_), .B(new_n13466_), .ZN(new_n13609_));
  INV_X1     g13417(.I(new_n13471_), .ZN(new_n13610_));
  INV_X1     g13418(.I(new_n13481_), .ZN(new_n13611_));
  NOR2_X1    g13419(.A1(new_n13594_), .A2(new_n13595_), .ZN(new_n13612_));
  AOI21_X1   g13420(.A1(new_n13612_), .A2(new_n8349_), .B(new_n13611_), .ZN(new_n13613_));
  NAND2_X1   g13421(.A1(new_n13596_), .A2(new_n7934_), .ZN(new_n13614_));
  OAI21_X1   g13422(.A1(new_n13613_), .A2(new_n13614_), .B(new_n13477_), .ZN(new_n13615_));
  INV_X1     g13423(.I(new_n13596_), .ZN(new_n13616_));
  OAI21_X1   g13424(.A1(new_n13613_), .A2(new_n13616_), .B(\asqrt[25] ), .ZN(new_n13617_));
  NAND3_X1   g13425(.A1(new_n13615_), .A2(new_n13617_), .A3(new_n7561_), .ZN(new_n13618_));
  NAND2_X1   g13426(.A1(new_n13618_), .A2(new_n13474_), .ZN(new_n13619_));
  NAND2_X1   g13427(.A1(new_n13615_), .A2(new_n13617_), .ZN(new_n13620_));
  AOI21_X1   g13428(.A1(new_n13620_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n13621_));
  AOI21_X1   g13429(.A1(new_n13621_), .A2(new_n13619_), .B(new_n13610_), .ZN(new_n13622_));
  AOI21_X1   g13430(.A1(new_n13619_), .A2(new_n13600_), .B(new_n7166_), .ZN(new_n13623_));
  OAI21_X1   g13431(.A1(new_n13622_), .A2(new_n13623_), .B(\asqrt[28] ), .ZN(new_n13624_));
  AOI21_X1   g13432(.A1(new_n13606_), .A2(new_n13624_), .B(new_n6454_), .ZN(new_n13625_));
  NOR2_X1    g13433(.A1(new_n13609_), .A2(new_n13625_), .ZN(new_n13626_));
  AOI21_X1   g13434(.A1(new_n13626_), .A2(new_n6106_), .B(new_n13463_), .ZN(new_n13627_));
  OAI21_X1   g13435(.A1(new_n13609_), .A2(new_n13625_), .B(\asqrt[30] ), .ZN(new_n13628_));
  NAND2_X1   g13436(.A1(new_n13628_), .A2(new_n5750_), .ZN(new_n13629_));
  OAI21_X1   g13437(.A1(new_n13627_), .A2(new_n13629_), .B(new_n13459_), .ZN(new_n13630_));
  INV_X1     g13438(.I(new_n13628_), .ZN(new_n13631_));
  OAI21_X1   g13439(.A1(new_n13627_), .A2(new_n13631_), .B(\asqrt[31] ), .ZN(new_n13632_));
  NAND3_X1   g13440(.A1(new_n13630_), .A2(new_n13632_), .A3(new_n5435_), .ZN(new_n13633_));
  NAND2_X1   g13441(.A1(new_n13633_), .A2(new_n13457_), .ZN(new_n13634_));
  NAND2_X1   g13442(.A1(new_n13630_), .A2(new_n13632_), .ZN(new_n13635_));
  AOI21_X1   g13443(.A1(new_n13635_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n13636_));
  AOI21_X1   g13444(.A1(new_n13636_), .A2(new_n13634_), .B(new_n13454_), .ZN(new_n13637_));
  INV_X1     g13445(.I(new_n13459_), .ZN(new_n13638_));
  INV_X1     g13446(.I(new_n13469_), .ZN(new_n13639_));
  NOR2_X1    g13447(.A1(new_n13622_), .A2(new_n13623_), .ZN(new_n13640_));
  AOI21_X1   g13448(.A1(new_n13640_), .A2(new_n6813_), .B(new_n13639_), .ZN(new_n13641_));
  NAND2_X1   g13449(.A1(new_n13624_), .A2(new_n6454_), .ZN(new_n13642_));
  OAI21_X1   g13450(.A1(new_n13641_), .A2(new_n13642_), .B(new_n13465_), .ZN(new_n13643_));
  INV_X1     g13451(.I(new_n13624_), .ZN(new_n13644_));
  OAI21_X1   g13452(.A1(new_n13641_), .A2(new_n13644_), .B(\asqrt[29] ), .ZN(new_n13645_));
  NAND3_X1   g13453(.A1(new_n13643_), .A2(new_n13645_), .A3(new_n6106_), .ZN(new_n13646_));
  NAND2_X1   g13454(.A1(new_n13646_), .A2(new_n13462_), .ZN(new_n13647_));
  NAND2_X1   g13455(.A1(new_n13643_), .A2(new_n13645_), .ZN(new_n13648_));
  AOI21_X1   g13456(.A1(new_n13648_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n13649_));
  AOI21_X1   g13457(.A1(new_n13649_), .A2(new_n13647_), .B(new_n13638_), .ZN(new_n13650_));
  AOI21_X1   g13458(.A1(new_n13647_), .A2(new_n13628_), .B(new_n5750_), .ZN(new_n13651_));
  OAI21_X1   g13459(.A1(new_n13650_), .A2(new_n13651_), .B(\asqrt[32] ), .ZN(new_n13652_));
  AOI21_X1   g13460(.A1(new_n13634_), .A2(new_n13652_), .B(new_n5110_), .ZN(new_n13653_));
  NOR2_X1    g13461(.A1(new_n13637_), .A2(new_n13653_), .ZN(new_n13654_));
  AOI21_X1   g13462(.A1(new_n13654_), .A2(new_n4810_), .B(new_n13451_), .ZN(new_n13655_));
  OAI21_X1   g13463(.A1(new_n13637_), .A2(new_n13653_), .B(\asqrt[34] ), .ZN(new_n13656_));
  NAND2_X1   g13464(.A1(new_n13656_), .A2(new_n4510_), .ZN(new_n13657_));
  OAI21_X1   g13465(.A1(new_n13655_), .A2(new_n13657_), .B(new_n13447_), .ZN(new_n13658_));
  INV_X1     g13466(.I(new_n13656_), .ZN(new_n13659_));
  OAI21_X1   g13467(.A1(new_n13655_), .A2(new_n13659_), .B(\asqrt[35] ), .ZN(new_n13660_));
  NAND3_X1   g13468(.A1(new_n13658_), .A2(new_n13660_), .A3(new_n4224_), .ZN(new_n13661_));
  NAND2_X1   g13469(.A1(new_n13661_), .A2(new_n13445_), .ZN(new_n13662_));
  NAND2_X1   g13470(.A1(new_n13658_), .A2(new_n13660_), .ZN(new_n13663_));
  AOI21_X1   g13471(.A1(new_n13663_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n13664_));
  AOI21_X1   g13472(.A1(new_n13664_), .A2(new_n13662_), .B(new_n13442_), .ZN(new_n13665_));
  INV_X1     g13473(.I(new_n13447_), .ZN(new_n13666_));
  INV_X1     g13474(.I(new_n13457_), .ZN(new_n13667_));
  NOR2_X1    g13475(.A1(new_n13650_), .A2(new_n13651_), .ZN(new_n13668_));
  AOI21_X1   g13476(.A1(new_n13668_), .A2(new_n5435_), .B(new_n13667_), .ZN(new_n13669_));
  NAND2_X1   g13477(.A1(new_n13652_), .A2(new_n5110_), .ZN(new_n13670_));
  OAI21_X1   g13478(.A1(new_n13669_), .A2(new_n13670_), .B(new_n13453_), .ZN(new_n13671_));
  INV_X1     g13479(.I(new_n13652_), .ZN(new_n13672_));
  OAI21_X1   g13480(.A1(new_n13669_), .A2(new_n13672_), .B(\asqrt[33] ), .ZN(new_n13673_));
  NAND3_X1   g13481(.A1(new_n13671_), .A2(new_n13673_), .A3(new_n4810_), .ZN(new_n13674_));
  NAND2_X1   g13482(.A1(new_n13674_), .A2(new_n13450_), .ZN(new_n13675_));
  NAND2_X1   g13483(.A1(new_n13671_), .A2(new_n13673_), .ZN(new_n13676_));
  AOI21_X1   g13484(.A1(new_n13676_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n13677_));
  AOI21_X1   g13485(.A1(new_n13677_), .A2(new_n13675_), .B(new_n13666_), .ZN(new_n13678_));
  AOI21_X1   g13486(.A1(new_n13675_), .A2(new_n13656_), .B(new_n4510_), .ZN(new_n13679_));
  OAI21_X1   g13487(.A1(new_n13678_), .A2(new_n13679_), .B(\asqrt[36] ), .ZN(new_n13680_));
  AOI21_X1   g13488(.A1(new_n13662_), .A2(new_n13680_), .B(new_n3928_), .ZN(new_n13681_));
  NOR2_X1    g13489(.A1(new_n13665_), .A2(new_n13681_), .ZN(new_n13682_));
  AOI21_X1   g13490(.A1(new_n13682_), .A2(new_n3675_), .B(new_n13439_), .ZN(new_n13683_));
  OAI21_X1   g13491(.A1(new_n13665_), .A2(new_n13681_), .B(\asqrt[38] ), .ZN(new_n13684_));
  NAND2_X1   g13492(.A1(new_n13684_), .A2(new_n3400_), .ZN(new_n13685_));
  OAI21_X1   g13493(.A1(new_n13683_), .A2(new_n13685_), .B(new_n13435_), .ZN(new_n13686_));
  INV_X1     g13494(.I(new_n13684_), .ZN(new_n13687_));
  OAI21_X1   g13495(.A1(new_n13683_), .A2(new_n13687_), .B(\asqrt[39] ), .ZN(new_n13688_));
  NAND3_X1   g13496(.A1(new_n13686_), .A2(new_n13688_), .A3(new_n3167_), .ZN(new_n13689_));
  NAND2_X1   g13497(.A1(new_n13689_), .A2(new_n13433_), .ZN(new_n13690_));
  NAND2_X1   g13498(.A1(new_n13686_), .A2(new_n13688_), .ZN(new_n13691_));
  AOI21_X1   g13499(.A1(new_n13691_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n13692_));
  AOI21_X1   g13500(.A1(new_n13692_), .A2(new_n13690_), .B(new_n13430_), .ZN(new_n13693_));
  INV_X1     g13501(.I(new_n13435_), .ZN(new_n13694_));
  INV_X1     g13502(.I(new_n13445_), .ZN(new_n13695_));
  NOR2_X1    g13503(.A1(new_n13678_), .A2(new_n13679_), .ZN(new_n13696_));
  AOI21_X1   g13504(.A1(new_n13696_), .A2(new_n4224_), .B(new_n13695_), .ZN(new_n13697_));
  NAND2_X1   g13505(.A1(new_n13680_), .A2(new_n3928_), .ZN(new_n13698_));
  OAI21_X1   g13506(.A1(new_n13697_), .A2(new_n13698_), .B(new_n13441_), .ZN(new_n13699_));
  INV_X1     g13507(.I(new_n13680_), .ZN(new_n13700_));
  OAI21_X1   g13508(.A1(new_n13697_), .A2(new_n13700_), .B(\asqrt[37] ), .ZN(new_n13701_));
  NAND3_X1   g13509(.A1(new_n13699_), .A2(new_n13701_), .A3(new_n3675_), .ZN(new_n13702_));
  NAND2_X1   g13510(.A1(new_n13702_), .A2(new_n13438_), .ZN(new_n13703_));
  NAND2_X1   g13511(.A1(new_n13699_), .A2(new_n13701_), .ZN(new_n13704_));
  AOI21_X1   g13512(.A1(new_n13704_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n13705_));
  AOI21_X1   g13513(.A1(new_n13705_), .A2(new_n13703_), .B(new_n13694_), .ZN(new_n13706_));
  AOI21_X1   g13514(.A1(new_n13703_), .A2(new_n13684_), .B(new_n3400_), .ZN(new_n13707_));
  OAI21_X1   g13515(.A1(new_n13706_), .A2(new_n13707_), .B(\asqrt[40] ), .ZN(new_n13708_));
  AOI21_X1   g13516(.A1(new_n13690_), .A2(new_n13708_), .B(new_n2912_), .ZN(new_n13709_));
  NOR2_X1    g13517(.A1(new_n13693_), .A2(new_n13709_), .ZN(new_n13710_));
  AOI21_X1   g13518(.A1(new_n13710_), .A2(new_n2699_), .B(new_n13427_), .ZN(new_n13711_));
  OAI21_X1   g13519(.A1(new_n13693_), .A2(new_n13709_), .B(\asqrt[42] ), .ZN(new_n13712_));
  NAND2_X1   g13520(.A1(new_n13712_), .A2(new_n2464_), .ZN(new_n13713_));
  OAI21_X1   g13521(.A1(new_n13711_), .A2(new_n13713_), .B(new_n13423_), .ZN(new_n13714_));
  INV_X1     g13522(.I(new_n13712_), .ZN(new_n13715_));
  OAI21_X1   g13523(.A1(new_n13711_), .A2(new_n13715_), .B(\asqrt[43] ), .ZN(new_n13716_));
  NAND3_X1   g13524(.A1(new_n13714_), .A2(new_n13716_), .A3(new_n2271_), .ZN(new_n13717_));
  NAND2_X1   g13525(.A1(new_n13717_), .A2(new_n13421_), .ZN(new_n13718_));
  NAND2_X1   g13526(.A1(new_n13714_), .A2(new_n13716_), .ZN(new_n13719_));
  AOI21_X1   g13527(.A1(new_n13719_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n13720_));
  AOI21_X1   g13528(.A1(new_n13720_), .A2(new_n13718_), .B(new_n13418_), .ZN(new_n13721_));
  INV_X1     g13529(.I(new_n13423_), .ZN(new_n13722_));
  INV_X1     g13530(.I(new_n13433_), .ZN(new_n13723_));
  NOR2_X1    g13531(.A1(new_n13706_), .A2(new_n13707_), .ZN(new_n13724_));
  AOI21_X1   g13532(.A1(new_n13724_), .A2(new_n3167_), .B(new_n13723_), .ZN(new_n13725_));
  NAND2_X1   g13533(.A1(new_n13708_), .A2(new_n2912_), .ZN(new_n13726_));
  OAI21_X1   g13534(.A1(new_n13725_), .A2(new_n13726_), .B(new_n13429_), .ZN(new_n13727_));
  INV_X1     g13535(.I(new_n13708_), .ZN(new_n13728_));
  OAI21_X1   g13536(.A1(new_n13725_), .A2(new_n13728_), .B(\asqrt[41] ), .ZN(new_n13729_));
  NAND3_X1   g13537(.A1(new_n13727_), .A2(new_n13729_), .A3(new_n2699_), .ZN(new_n13730_));
  NAND2_X1   g13538(.A1(new_n13730_), .A2(new_n13426_), .ZN(new_n13731_));
  NAND2_X1   g13539(.A1(new_n13727_), .A2(new_n13729_), .ZN(new_n13732_));
  AOI21_X1   g13540(.A1(new_n13732_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n13733_));
  AOI21_X1   g13541(.A1(new_n13733_), .A2(new_n13731_), .B(new_n13722_), .ZN(new_n13734_));
  AOI21_X1   g13542(.A1(new_n13731_), .A2(new_n13712_), .B(new_n2464_), .ZN(new_n13735_));
  OAI21_X1   g13543(.A1(new_n13734_), .A2(new_n13735_), .B(\asqrt[44] ), .ZN(new_n13736_));
  AOI21_X1   g13544(.A1(new_n13718_), .A2(new_n13736_), .B(new_n2072_), .ZN(new_n13737_));
  NOR2_X1    g13545(.A1(new_n13721_), .A2(new_n13737_), .ZN(new_n13738_));
  AOI21_X1   g13546(.A1(new_n13738_), .A2(new_n1884_), .B(new_n13415_), .ZN(new_n13739_));
  OAI21_X1   g13547(.A1(new_n13721_), .A2(new_n13737_), .B(\asqrt[46] ), .ZN(new_n13740_));
  NAND2_X1   g13548(.A1(new_n13740_), .A2(new_n1688_), .ZN(new_n13741_));
  OAI21_X1   g13549(.A1(new_n13739_), .A2(new_n13741_), .B(new_n13411_), .ZN(new_n13742_));
  INV_X1     g13550(.I(new_n13740_), .ZN(new_n13743_));
  OAI21_X1   g13551(.A1(new_n13739_), .A2(new_n13743_), .B(\asqrt[47] ), .ZN(new_n13744_));
  NAND3_X1   g13552(.A1(new_n13742_), .A2(new_n13744_), .A3(new_n1533_), .ZN(new_n13745_));
  NAND2_X1   g13553(.A1(new_n13745_), .A2(new_n13409_), .ZN(new_n13746_));
  NAND2_X1   g13554(.A1(new_n13742_), .A2(new_n13744_), .ZN(new_n13747_));
  AOI21_X1   g13555(.A1(new_n13747_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n13748_));
  AOI21_X1   g13556(.A1(new_n13748_), .A2(new_n13746_), .B(new_n13406_), .ZN(new_n13749_));
  INV_X1     g13557(.I(new_n13411_), .ZN(new_n13750_));
  INV_X1     g13558(.I(new_n13421_), .ZN(new_n13751_));
  NOR2_X1    g13559(.A1(new_n13734_), .A2(new_n13735_), .ZN(new_n13752_));
  AOI21_X1   g13560(.A1(new_n13752_), .A2(new_n2271_), .B(new_n13751_), .ZN(new_n13753_));
  NAND2_X1   g13561(.A1(new_n13736_), .A2(new_n2072_), .ZN(new_n13754_));
  OAI21_X1   g13562(.A1(new_n13753_), .A2(new_n13754_), .B(new_n13417_), .ZN(new_n13755_));
  INV_X1     g13563(.I(new_n13736_), .ZN(new_n13756_));
  OAI21_X1   g13564(.A1(new_n13753_), .A2(new_n13756_), .B(\asqrt[45] ), .ZN(new_n13757_));
  NAND3_X1   g13565(.A1(new_n13755_), .A2(new_n13757_), .A3(new_n1884_), .ZN(new_n13758_));
  NAND2_X1   g13566(.A1(new_n13758_), .A2(new_n13414_), .ZN(new_n13759_));
  NAND2_X1   g13567(.A1(new_n13755_), .A2(new_n13757_), .ZN(new_n13760_));
  AOI21_X1   g13568(.A1(new_n13760_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n13761_));
  AOI21_X1   g13569(.A1(new_n13761_), .A2(new_n13759_), .B(new_n13750_), .ZN(new_n13762_));
  AOI21_X1   g13570(.A1(new_n13759_), .A2(new_n13740_), .B(new_n1688_), .ZN(new_n13763_));
  OAI21_X1   g13571(.A1(new_n13762_), .A2(new_n13763_), .B(\asqrt[48] ), .ZN(new_n13764_));
  AOI21_X1   g13572(.A1(new_n13746_), .A2(new_n13764_), .B(new_n1368_), .ZN(new_n13765_));
  NOR2_X1    g13573(.A1(new_n13749_), .A2(new_n13765_), .ZN(new_n13766_));
  AOI21_X1   g13574(.A1(new_n13766_), .A2(new_n1228_), .B(new_n13403_), .ZN(new_n13767_));
  OAI21_X1   g13575(.A1(new_n13749_), .A2(new_n13765_), .B(\asqrt[50] ), .ZN(new_n13768_));
  NAND2_X1   g13576(.A1(new_n13768_), .A2(new_n1088_), .ZN(new_n13769_));
  OAI21_X1   g13577(.A1(new_n13767_), .A2(new_n13769_), .B(new_n13399_), .ZN(new_n13770_));
  INV_X1     g13578(.I(new_n13768_), .ZN(new_n13771_));
  OAI21_X1   g13579(.A1(new_n13767_), .A2(new_n13771_), .B(\asqrt[51] ), .ZN(new_n13772_));
  NAND3_X1   g13580(.A1(new_n13770_), .A2(new_n13772_), .A3(new_n962_), .ZN(new_n13773_));
  INV_X1     g13581(.I(new_n13399_), .ZN(new_n13774_));
  INV_X1     g13582(.I(new_n13409_), .ZN(new_n13775_));
  NOR2_X1    g13583(.A1(new_n13762_), .A2(new_n13763_), .ZN(new_n13776_));
  AOI21_X1   g13584(.A1(new_n13776_), .A2(new_n1533_), .B(new_n13775_), .ZN(new_n13777_));
  NAND2_X1   g13585(.A1(new_n13764_), .A2(new_n1368_), .ZN(new_n13778_));
  OAI21_X1   g13586(.A1(new_n13777_), .A2(new_n13778_), .B(new_n13405_), .ZN(new_n13779_));
  INV_X1     g13587(.I(new_n13764_), .ZN(new_n13780_));
  OAI21_X1   g13588(.A1(new_n13777_), .A2(new_n13780_), .B(\asqrt[49] ), .ZN(new_n13781_));
  NAND3_X1   g13589(.A1(new_n13779_), .A2(new_n13781_), .A3(new_n1228_), .ZN(new_n13782_));
  NAND2_X1   g13590(.A1(new_n13782_), .A2(new_n13402_), .ZN(new_n13783_));
  NAND2_X1   g13591(.A1(new_n13779_), .A2(new_n13781_), .ZN(new_n13784_));
  AOI21_X1   g13592(.A1(new_n13784_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n13785_));
  AOI21_X1   g13593(.A1(new_n13785_), .A2(new_n13783_), .B(new_n13774_), .ZN(new_n13786_));
  AOI21_X1   g13594(.A1(new_n13783_), .A2(new_n13768_), .B(new_n1088_), .ZN(new_n13787_));
  OAI21_X1   g13595(.A1(new_n13786_), .A2(new_n13787_), .B(\asqrt[52] ), .ZN(new_n13788_));
  NAND2_X1   g13596(.A1(new_n13379_), .A2(new_n12894_), .ZN(new_n13789_));
  NOR2_X1    g13597(.A1(new_n13382_), .A2(new_n12894_), .ZN(new_n13790_));
  NAND2_X1   g13598(.A1(new_n13790_), .A2(new_n13394_), .ZN(new_n13791_));
  AOI21_X1   g13599(.A1(new_n13791_), .A2(new_n13789_), .B(new_n193_), .ZN(new_n13792_));
  INV_X1     g13600(.I(new_n13792_), .ZN(new_n13793_));
  NAND3_X1   g13601(.A1(\asqrt[13] ), .A2(new_n13364_), .A3(new_n13375_), .ZN(new_n13794_));
  XOR2_X1    g13602(.A1(new_n13794_), .A2(new_n13367_), .Z(new_n13795_));
  AOI21_X1   g13603(.A1(new_n13790_), .A2(new_n13379_), .B(new_n13380_), .ZN(new_n13796_));
  OAI21_X1   g13604(.A1(new_n13334_), .A2(new_n13336_), .B(new_n13339_), .ZN(new_n13797_));
  NOR2_X1    g13605(.A1(new_n13382_), .A2(new_n13797_), .ZN(new_n13798_));
  XOR2_X1    g13606(.A1(new_n13798_), .A2(new_n12902_), .Z(new_n13799_));
  NAND3_X1   g13607(.A1(\asqrt[13] ), .A2(new_n13350_), .A3(new_n13335_), .ZN(new_n13800_));
  XOR2_X1    g13608(.A1(new_n13800_), .A2(new_n12906_), .Z(new_n13801_));
  OAI21_X1   g13609(.A1(new_n13345_), .A2(new_n13346_), .B(new_n13349_), .ZN(new_n13802_));
  NOR2_X1    g13610(.A1(new_n13382_), .A2(new_n13802_), .ZN(new_n13803_));
  XOR2_X1    g13611(.A1(new_n13803_), .A2(new_n12908_), .Z(new_n13804_));
  INV_X1     g13612(.I(new_n13804_), .ZN(new_n13805_));
  NAND3_X1   g13613(.A1(\asqrt[13] ), .A2(new_n13312_), .A3(new_n13331_), .ZN(new_n13806_));
  XOR2_X1    g13614(.A1(new_n13806_), .A2(new_n13343_), .Z(new_n13807_));
  INV_X1     g13615(.I(new_n13807_), .ZN(new_n13808_));
  OAI21_X1   g13616(.A1(new_n13306_), .A2(new_n13308_), .B(new_n13311_), .ZN(new_n13809_));
  NOR2_X1    g13617(.A1(new_n13382_), .A2(new_n13809_), .ZN(new_n13810_));
  XOR2_X1    g13618(.A1(new_n13810_), .A2(new_n12914_), .Z(new_n13811_));
  NAND3_X1   g13619(.A1(\asqrt[13] ), .A2(new_n13325_), .A3(new_n13307_), .ZN(new_n13812_));
  XOR2_X1    g13620(.A1(new_n13812_), .A2(new_n12918_), .Z(new_n13813_));
  OAI21_X1   g13621(.A1(new_n13320_), .A2(new_n13321_), .B(new_n13324_), .ZN(new_n13814_));
  NOR2_X1    g13622(.A1(new_n13382_), .A2(new_n13814_), .ZN(new_n13815_));
  XOR2_X1    g13623(.A1(new_n13815_), .A2(new_n12920_), .Z(new_n13816_));
  INV_X1     g13624(.I(new_n13816_), .ZN(new_n13817_));
  NAND3_X1   g13625(.A1(\asqrt[13] ), .A2(new_n13284_), .A3(new_n13303_), .ZN(new_n13818_));
  XOR2_X1    g13626(.A1(new_n13818_), .A2(new_n13318_), .Z(new_n13819_));
  INV_X1     g13627(.I(new_n13819_), .ZN(new_n13820_));
  NAND2_X1   g13628(.A1(new_n13773_), .A2(new_n13385_), .ZN(new_n13821_));
  NAND2_X1   g13629(.A1(new_n13770_), .A2(new_n13772_), .ZN(new_n13822_));
  AOI21_X1   g13630(.A1(new_n13822_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n13823_));
  AOI21_X1   g13631(.A1(new_n13823_), .A2(new_n13821_), .B(new_n13820_), .ZN(new_n13824_));
  AOI21_X1   g13632(.A1(new_n13821_), .A2(new_n13788_), .B(new_n842_), .ZN(new_n13825_));
  NOR2_X1    g13633(.A1(new_n13824_), .A2(new_n13825_), .ZN(new_n13826_));
  AOI21_X1   g13634(.A1(new_n13826_), .A2(new_n720_), .B(new_n13817_), .ZN(new_n13827_));
  OAI21_X1   g13635(.A1(new_n13824_), .A2(new_n13825_), .B(\asqrt[54] ), .ZN(new_n13828_));
  NAND2_X1   g13636(.A1(new_n13828_), .A2(new_n630_), .ZN(new_n13829_));
  OAI21_X1   g13637(.A1(new_n13827_), .A2(new_n13829_), .B(new_n13813_), .ZN(new_n13830_));
  INV_X1     g13638(.I(new_n13828_), .ZN(new_n13831_));
  OAI21_X1   g13639(.A1(new_n13827_), .A2(new_n13831_), .B(\asqrt[55] ), .ZN(new_n13832_));
  NAND3_X1   g13640(.A1(new_n13830_), .A2(new_n13832_), .A3(new_n545_), .ZN(new_n13833_));
  NAND2_X1   g13641(.A1(new_n13833_), .A2(new_n13811_), .ZN(new_n13834_));
  NAND2_X1   g13642(.A1(new_n13830_), .A2(new_n13832_), .ZN(new_n13835_));
  AOI21_X1   g13643(.A1(new_n13835_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n13836_));
  AOI21_X1   g13644(.A1(new_n13836_), .A2(new_n13834_), .B(new_n13808_), .ZN(new_n13837_));
  INV_X1     g13645(.I(new_n13813_), .ZN(new_n13838_));
  NOR2_X1    g13646(.A1(new_n13786_), .A2(new_n13787_), .ZN(new_n13839_));
  AOI21_X1   g13647(.A1(new_n13839_), .A2(new_n962_), .B(new_n13386_), .ZN(new_n13840_));
  NAND2_X1   g13648(.A1(new_n13788_), .A2(new_n842_), .ZN(new_n13841_));
  OAI21_X1   g13649(.A1(new_n13840_), .A2(new_n13841_), .B(new_n13819_), .ZN(new_n13842_));
  INV_X1     g13650(.I(new_n13788_), .ZN(new_n13843_));
  OAI21_X1   g13651(.A1(new_n13840_), .A2(new_n13843_), .B(\asqrt[53] ), .ZN(new_n13844_));
  NAND3_X1   g13652(.A1(new_n13842_), .A2(new_n13844_), .A3(new_n720_), .ZN(new_n13845_));
  NAND2_X1   g13653(.A1(new_n13845_), .A2(new_n13816_), .ZN(new_n13846_));
  NAND2_X1   g13654(.A1(new_n13842_), .A2(new_n13844_), .ZN(new_n13847_));
  AOI21_X1   g13655(.A1(new_n13847_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n13848_));
  AOI21_X1   g13656(.A1(new_n13848_), .A2(new_n13846_), .B(new_n13838_), .ZN(new_n13849_));
  AOI21_X1   g13657(.A1(new_n13846_), .A2(new_n13828_), .B(new_n630_), .ZN(new_n13850_));
  OAI21_X1   g13658(.A1(new_n13849_), .A2(new_n13850_), .B(\asqrt[56] ), .ZN(new_n13851_));
  AOI21_X1   g13659(.A1(new_n13834_), .A2(new_n13851_), .B(new_n450_), .ZN(new_n13852_));
  NOR2_X1    g13660(.A1(new_n13837_), .A2(new_n13852_), .ZN(new_n13853_));
  AOI21_X1   g13661(.A1(new_n13853_), .A2(new_n403_), .B(new_n13805_), .ZN(new_n13854_));
  OAI21_X1   g13662(.A1(new_n13837_), .A2(new_n13852_), .B(\asqrt[58] ), .ZN(new_n13855_));
  NAND2_X1   g13663(.A1(new_n13855_), .A2(new_n339_), .ZN(new_n13856_));
  OAI21_X1   g13664(.A1(new_n13854_), .A2(new_n13856_), .B(new_n13801_), .ZN(new_n13857_));
  INV_X1     g13665(.I(new_n13855_), .ZN(new_n13858_));
  OAI21_X1   g13666(.A1(new_n13854_), .A2(new_n13858_), .B(\asqrt[59] ), .ZN(new_n13859_));
  NAND3_X1   g13667(.A1(new_n13857_), .A2(new_n13859_), .A3(new_n288_), .ZN(new_n13860_));
  NAND2_X1   g13668(.A1(new_n13860_), .A2(new_n13799_), .ZN(new_n13861_));
  INV_X1     g13669(.I(new_n13801_), .ZN(new_n13862_));
  INV_X1     g13670(.I(new_n13811_), .ZN(new_n13863_));
  NOR2_X1    g13671(.A1(new_n13849_), .A2(new_n13850_), .ZN(new_n13864_));
  AOI21_X1   g13672(.A1(new_n13864_), .A2(new_n545_), .B(new_n13863_), .ZN(new_n13865_));
  NAND2_X1   g13673(.A1(new_n13851_), .A2(new_n450_), .ZN(new_n13866_));
  OAI21_X1   g13674(.A1(new_n13865_), .A2(new_n13866_), .B(new_n13807_), .ZN(new_n13867_));
  INV_X1     g13675(.I(new_n13851_), .ZN(new_n13868_));
  OAI21_X1   g13676(.A1(new_n13865_), .A2(new_n13868_), .B(\asqrt[57] ), .ZN(new_n13869_));
  NAND3_X1   g13677(.A1(new_n13867_), .A2(new_n13869_), .A3(new_n403_), .ZN(new_n13870_));
  NAND2_X1   g13678(.A1(new_n13870_), .A2(new_n13804_), .ZN(new_n13871_));
  NAND2_X1   g13679(.A1(new_n13867_), .A2(new_n13869_), .ZN(new_n13872_));
  AOI21_X1   g13680(.A1(new_n13872_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n13873_));
  AOI21_X1   g13681(.A1(new_n13873_), .A2(new_n13871_), .B(new_n13862_), .ZN(new_n13874_));
  AOI21_X1   g13682(.A1(new_n13871_), .A2(new_n13855_), .B(new_n339_), .ZN(new_n13875_));
  OAI21_X1   g13683(.A1(new_n13874_), .A2(new_n13875_), .B(\asqrt[60] ), .ZN(new_n13876_));
  AOI21_X1   g13684(.A1(new_n13861_), .A2(new_n13876_), .B(new_n242_), .ZN(new_n13877_));
  NAND3_X1   g13685(.A1(\asqrt[13] ), .A2(new_n13340_), .A3(new_n13356_), .ZN(new_n13878_));
  XOR2_X1    g13686(.A1(new_n13878_), .A2(new_n13368_), .Z(new_n13879_));
  INV_X1     g13687(.I(new_n13879_), .ZN(new_n13880_));
  NAND2_X1   g13688(.A1(new_n13857_), .A2(new_n13859_), .ZN(new_n13881_));
  AOI21_X1   g13689(.A1(new_n13881_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n13882_));
  AOI21_X1   g13690(.A1(new_n13882_), .A2(new_n13861_), .B(new_n13880_), .ZN(new_n13883_));
  OAI21_X1   g13691(.A1(new_n13883_), .A2(new_n13877_), .B(\asqrt[62] ), .ZN(new_n13884_));
  INV_X1     g13692(.I(new_n13884_), .ZN(new_n13885_));
  NOR2_X1    g13693(.A1(new_n13883_), .A2(new_n13877_), .ZN(new_n13886_));
  AOI21_X1   g13694(.A1(new_n13341_), .A2(new_n13362_), .B(new_n13357_), .ZN(new_n13887_));
  NAND2_X1   g13695(.A1(\asqrt[13] ), .A2(new_n13887_), .ZN(new_n13888_));
  XOR2_X1    g13696(.A1(new_n13888_), .A2(new_n13360_), .Z(new_n13889_));
  INV_X1     g13697(.I(new_n13889_), .ZN(new_n13890_));
  AOI21_X1   g13698(.A1(new_n13886_), .A2(new_n234_), .B(new_n13890_), .ZN(new_n13891_));
  OAI21_X1   g13699(.A1(new_n13891_), .A2(new_n13885_), .B(new_n13796_), .ZN(new_n13892_));
  OAI21_X1   g13700(.A1(new_n13892_), .A2(new_n13795_), .B(new_n193_), .ZN(new_n13893_));
  NOR2_X1    g13701(.A1(new_n13891_), .A2(new_n13885_), .ZN(new_n13894_));
  NAND2_X1   g13702(.A1(new_n13894_), .A2(new_n13795_), .ZN(new_n13895_));
  NOR2_X1    g13703(.A1(\asqrt[13] ), .A2(new_n12895_), .ZN(new_n13896_));
  INV_X1     g13704(.I(new_n13896_), .ZN(new_n13897_));
  NAND4_X1   g13705(.A1(new_n13893_), .A2(new_n13793_), .A3(new_n13895_), .A4(new_n13897_), .ZN(\asqrt[12] ));
  NAND3_X1   g13706(.A1(\asqrt[12] ), .A2(new_n13773_), .A3(new_n13788_), .ZN(new_n13899_));
  XOR2_X1    g13707(.A1(new_n13899_), .A2(new_n13386_), .Z(new_n13900_));
  INV_X1     g13708(.I(new_n13799_), .ZN(new_n13901_));
  NOR2_X1    g13709(.A1(new_n13874_), .A2(new_n13875_), .ZN(new_n13902_));
  AOI21_X1   g13710(.A1(new_n13902_), .A2(new_n288_), .B(new_n13901_), .ZN(new_n13903_));
  INV_X1     g13711(.I(new_n13876_), .ZN(new_n13904_));
  OAI21_X1   g13712(.A1(new_n13903_), .A2(new_n13904_), .B(\asqrt[61] ), .ZN(new_n13905_));
  NAND2_X1   g13713(.A1(new_n13876_), .A2(new_n242_), .ZN(new_n13906_));
  OAI21_X1   g13714(.A1(new_n13903_), .A2(new_n13906_), .B(new_n13879_), .ZN(new_n13907_));
  NAND3_X1   g13715(.A1(new_n13907_), .A2(new_n13905_), .A3(new_n234_), .ZN(new_n13908_));
  NAND2_X1   g13716(.A1(new_n13908_), .A2(new_n13889_), .ZN(new_n13909_));
  NAND2_X1   g13717(.A1(new_n13909_), .A2(new_n13884_), .ZN(new_n13910_));
  NAND2_X1   g13718(.A1(new_n13910_), .A2(new_n13795_), .ZN(new_n13911_));
  INV_X1     g13719(.I(new_n13795_), .ZN(new_n13912_));
  INV_X1     g13720(.I(new_n13796_), .ZN(new_n13913_));
  AOI21_X1   g13721(.A1(new_n13909_), .A2(new_n13884_), .B(new_n13913_), .ZN(new_n13914_));
  AOI21_X1   g13722(.A1(new_n13914_), .A2(new_n13912_), .B(\asqrt[63] ), .ZN(new_n13915_));
  NOR2_X1    g13723(.A1(new_n13910_), .A2(new_n13912_), .ZN(new_n13916_));
  NOR4_X1    g13724(.A1(new_n13915_), .A2(new_n13792_), .A3(new_n13916_), .A4(new_n13896_), .ZN(new_n13917_));
  NOR2_X1    g13725(.A1(new_n13917_), .A2(new_n13795_), .ZN(new_n13918_));
  NAND2_X1   g13726(.A1(new_n13918_), .A2(new_n13894_), .ZN(new_n13919_));
  AOI21_X1   g13727(.A1(new_n13919_), .A2(new_n13911_), .B(new_n193_), .ZN(new_n13920_));
  NAND3_X1   g13728(.A1(\asqrt[12] ), .A2(new_n13884_), .A3(new_n13908_), .ZN(new_n13921_));
  XOR2_X1    g13729(.A1(new_n13921_), .A2(new_n13889_), .Z(new_n13922_));
  INV_X1     g13730(.I(new_n13922_), .ZN(new_n13923_));
  AOI21_X1   g13731(.A1(new_n13918_), .A2(new_n13910_), .B(new_n13916_), .ZN(new_n13924_));
  INV_X1     g13732(.I(new_n13924_), .ZN(new_n13925_));
  OAI21_X1   g13733(.A1(new_n13854_), .A2(new_n13856_), .B(new_n13859_), .ZN(new_n13926_));
  NOR2_X1    g13734(.A1(new_n13917_), .A2(new_n13926_), .ZN(new_n13927_));
  XOR2_X1    g13735(.A1(new_n13927_), .A2(new_n13801_), .Z(new_n13928_));
  NAND3_X1   g13736(.A1(\asqrt[12] ), .A2(new_n13870_), .A3(new_n13855_), .ZN(new_n13929_));
  XOR2_X1    g13737(.A1(new_n13929_), .A2(new_n13805_), .Z(new_n13930_));
  OAI21_X1   g13738(.A1(new_n13865_), .A2(new_n13866_), .B(new_n13869_), .ZN(new_n13931_));
  NOR2_X1    g13739(.A1(new_n13917_), .A2(new_n13931_), .ZN(new_n13932_));
  XOR2_X1    g13740(.A1(new_n13932_), .A2(new_n13807_), .Z(new_n13933_));
  INV_X1     g13741(.I(new_n13933_), .ZN(new_n13934_));
  NAND3_X1   g13742(.A1(\asqrt[12] ), .A2(new_n13833_), .A3(new_n13851_), .ZN(new_n13935_));
  XOR2_X1    g13743(.A1(new_n13935_), .A2(new_n13863_), .Z(new_n13936_));
  INV_X1     g13744(.I(new_n13936_), .ZN(new_n13937_));
  OAI21_X1   g13745(.A1(new_n13827_), .A2(new_n13829_), .B(new_n13832_), .ZN(new_n13938_));
  NOR2_X1    g13746(.A1(new_n13917_), .A2(new_n13938_), .ZN(new_n13939_));
  XOR2_X1    g13747(.A1(new_n13939_), .A2(new_n13813_), .Z(new_n13940_));
  NAND3_X1   g13748(.A1(\asqrt[12] ), .A2(new_n13845_), .A3(new_n13828_), .ZN(new_n13941_));
  XOR2_X1    g13749(.A1(new_n13941_), .A2(new_n13817_), .Z(new_n13942_));
  OAI21_X1   g13750(.A1(new_n13840_), .A2(new_n13841_), .B(new_n13844_), .ZN(new_n13943_));
  NOR2_X1    g13751(.A1(new_n13917_), .A2(new_n13943_), .ZN(new_n13944_));
  XOR2_X1    g13752(.A1(new_n13944_), .A2(new_n13819_), .Z(new_n13945_));
  INV_X1     g13753(.I(new_n13945_), .ZN(new_n13946_));
  INV_X1     g13754(.I(new_n13900_), .ZN(new_n13947_));
  OAI21_X1   g13755(.A1(new_n13767_), .A2(new_n13769_), .B(new_n13772_), .ZN(new_n13948_));
  NOR2_X1    g13756(.A1(new_n13917_), .A2(new_n13948_), .ZN(new_n13949_));
  XOR2_X1    g13757(.A1(new_n13949_), .A2(new_n13399_), .Z(new_n13950_));
  NAND3_X1   g13758(.A1(\asqrt[12] ), .A2(new_n13782_), .A3(new_n13768_), .ZN(new_n13951_));
  XOR2_X1    g13759(.A1(new_n13951_), .A2(new_n13403_), .Z(new_n13952_));
  OAI21_X1   g13760(.A1(new_n13777_), .A2(new_n13778_), .B(new_n13781_), .ZN(new_n13953_));
  NOR2_X1    g13761(.A1(new_n13917_), .A2(new_n13953_), .ZN(new_n13954_));
  XOR2_X1    g13762(.A1(new_n13954_), .A2(new_n13405_), .Z(new_n13955_));
  INV_X1     g13763(.I(new_n13955_), .ZN(new_n13956_));
  NAND3_X1   g13764(.A1(\asqrt[12] ), .A2(new_n13745_), .A3(new_n13764_), .ZN(new_n13957_));
  XOR2_X1    g13765(.A1(new_n13957_), .A2(new_n13775_), .Z(new_n13958_));
  INV_X1     g13766(.I(new_n13958_), .ZN(new_n13959_));
  OAI21_X1   g13767(.A1(new_n13739_), .A2(new_n13741_), .B(new_n13744_), .ZN(new_n13960_));
  NOR2_X1    g13768(.A1(new_n13917_), .A2(new_n13960_), .ZN(new_n13961_));
  XOR2_X1    g13769(.A1(new_n13961_), .A2(new_n13411_), .Z(new_n13962_));
  NAND3_X1   g13770(.A1(\asqrt[12] ), .A2(new_n13758_), .A3(new_n13740_), .ZN(new_n13963_));
  XOR2_X1    g13771(.A1(new_n13963_), .A2(new_n13415_), .Z(new_n13964_));
  OAI21_X1   g13772(.A1(new_n13753_), .A2(new_n13754_), .B(new_n13757_), .ZN(new_n13965_));
  NOR2_X1    g13773(.A1(new_n13917_), .A2(new_n13965_), .ZN(new_n13966_));
  XOR2_X1    g13774(.A1(new_n13966_), .A2(new_n13417_), .Z(new_n13967_));
  INV_X1     g13775(.I(new_n13967_), .ZN(new_n13968_));
  NAND3_X1   g13776(.A1(\asqrt[12] ), .A2(new_n13717_), .A3(new_n13736_), .ZN(new_n13969_));
  XOR2_X1    g13777(.A1(new_n13969_), .A2(new_n13751_), .Z(new_n13970_));
  INV_X1     g13778(.I(new_n13970_), .ZN(new_n13971_));
  OAI21_X1   g13779(.A1(new_n13711_), .A2(new_n13713_), .B(new_n13716_), .ZN(new_n13972_));
  NOR2_X1    g13780(.A1(new_n13917_), .A2(new_n13972_), .ZN(new_n13973_));
  XOR2_X1    g13781(.A1(new_n13973_), .A2(new_n13423_), .Z(new_n13974_));
  NAND3_X1   g13782(.A1(\asqrt[12] ), .A2(new_n13730_), .A3(new_n13712_), .ZN(new_n13975_));
  XOR2_X1    g13783(.A1(new_n13975_), .A2(new_n13427_), .Z(new_n13976_));
  OAI21_X1   g13784(.A1(new_n13725_), .A2(new_n13726_), .B(new_n13729_), .ZN(new_n13977_));
  NOR2_X1    g13785(.A1(new_n13917_), .A2(new_n13977_), .ZN(new_n13978_));
  XOR2_X1    g13786(.A1(new_n13978_), .A2(new_n13429_), .Z(new_n13979_));
  INV_X1     g13787(.I(new_n13979_), .ZN(new_n13980_));
  NAND3_X1   g13788(.A1(\asqrt[12] ), .A2(new_n13689_), .A3(new_n13708_), .ZN(new_n13981_));
  XOR2_X1    g13789(.A1(new_n13981_), .A2(new_n13723_), .Z(new_n13982_));
  INV_X1     g13790(.I(new_n13982_), .ZN(new_n13983_));
  OAI21_X1   g13791(.A1(new_n13683_), .A2(new_n13685_), .B(new_n13688_), .ZN(new_n13984_));
  NOR2_X1    g13792(.A1(new_n13917_), .A2(new_n13984_), .ZN(new_n13985_));
  XOR2_X1    g13793(.A1(new_n13985_), .A2(new_n13435_), .Z(new_n13986_));
  NAND3_X1   g13794(.A1(\asqrt[12] ), .A2(new_n13702_), .A3(new_n13684_), .ZN(new_n13987_));
  XOR2_X1    g13795(.A1(new_n13987_), .A2(new_n13439_), .Z(new_n13988_));
  OAI21_X1   g13796(.A1(new_n13697_), .A2(new_n13698_), .B(new_n13701_), .ZN(new_n13989_));
  NOR2_X1    g13797(.A1(new_n13917_), .A2(new_n13989_), .ZN(new_n13990_));
  XOR2_X1    g13798(.A1(new_n13990_), .A2(new_n13441_), .Z(new_n13991_));
  INV_X1     g13799(.I(new_n13991_), .ZN(new_n13992_));
  NAND3_X1   g13800(.A1(\asqrt[12] ), .A2(new_n13661_), .A3(new_n13680_), .ZN(new_n13993_));
  XOR2_X1    g13801(.A1(new_n13993_), .A2(new_n13695_), .Z(new_n13994_));
  INV_X1     g13802(.I(new_n13994_), .ZN(new_n13995_));
  OAI21_X1   g13803(.A1(new_n13655_), .A2(new_n13657_), .B(new_n13660_), .ZN(new_n13996_));
  NOR2_X1    g13804(.A1(new_n13917_), .A2(new_n13996_), .ZN(new_n13997_));
  XOR2_X1    g13805(.A1(new_n13997_), .A2(new_n13447_), .Z(new_n13998_));
  NAND3_X1   g13806(.A1(\asqrt[12] ), .A2(new_n13674_), .A3(new_n13656_), .ZN(new_n13999_));
  XOR2_X1    g13807(.A1(new_n13999_), .A2(new_n13451_), .Z(new_n14000_));
  OAI21_X1   g13808(.A1(new_n13669_), .A2(new_n13670_), .B(new_n13673_), .ZN(new_n14001_));
  NOR2_X1    g13809(.A1(new_n13917_), .A2(new_n14001_), .ZN(new_n14002_));
  XOR2_X1    g13810(.A1(new_n14002_), .A2(new_n13453_), .Z(new_n14003_));
  INV_X1     g13811(.I(new_n14003_), .ZN(new_n14004_));
  NAND3_X1   g13812(.A1(\asqrt[12] ), .A2(new_n13633_), .A3(new_n13652_), .ZN(new_n14005_));
  XOR2_X1    g13813(.A1(new_n14005_), .A2(new_n13667_), .Z(new_n14006_));
  INV_X1     g13814(.I(new_n14006_), .ZN(new_n14007_));
  OAI21_X1   g13815(.A1(new_n13627_), .A2(new_n13629_), .B(new_n13632_), .ZN(new_n14008_));
  NOR2_X1    g13816(.A1(new_n13917_), .A2(new_n14008_), .ZN(new_n14009_));
  XOR2_X1    g13817(.A1(new_n14009_), .A2(new_n13459_), .Z(new_n14010_));
  NAND3_X1   g13818(.A1(\asqrt[12] ), .A2(new_n13646_), .A3(new_n13628_), .ZN(new_n14011_));
  XOR2_X1    g13819(.A1(new_n14011_), .A2(new_n13463_), .Z(new_n14012_));
  OAI21_X1   g13820(.A1(new_n13641_), .A2(new_n13642_), .B(new_n13645_), .ZN(new_n14013_));
  NOR2_X1    g13821(.A1(new_n13917_), .A2(new_n14013_), .ZN(new_n14014_));
  XOR2_X1    g13822(.A1(new_n14014_), .A2(new_n13465_), .Z(new_n14015_));
  INV_X1     g13823(.I(new_n14015_), .ZN(new_n14016_));
  NAND3_X1   g13824(.A1(\asqrt[12] ), .A2(new_n13605_), .A3(new_n13624_), .ZN(new_n14017_));
  XOR2_X1    g13825(.A1(new_n14017_), .A2(new_n13639_), .Z(new_n14018_));
  INV_X1     g13826(.I(new_n14018_), .ZN(new_n14019_));
  OAI21_X1   g13827(.A1(new_n13599_), .A2(new_n13601_), .B(new_n13604_), .ZN(new_n14020_));
  NOR2_X1    g13828(.A1(new_n13917_), .A2(new_n14020_), .ZN(new_n14021_));
  XOR2_X1    g13829(.A1(new_n14021_), .A2(new_n13471_), .Z(new_n14022_));
  NAND3_X1   g13830(.A1(\asqrt[12] ), .A2(new_n13618_), .A3(new_n13600_), .ZN(new_n14023_));
  XOR2_X1    g13831(.A1(new_n14023_), .A2(new_n13475_), .Z(new_n14024_));
  OAI21_X1   g13832(.A1(new_n13613_), .A2(new_n13614_), .B(new_n13617_), .ZN(new_n14025_));
  NOR2_X1    g13833(.A1(new_n13917_), .A2(new_n14025_), .ZN(new_n14026_));
  XOR2_X1    g13834(.A1(new_n14026_), .A2(new_n13477_), .Z(new_n14027_));
  INV_X1     g13835(.I(new_n14027_), .ZN(new_n14028_));
  NAND3_X1   g13836(.A1(\asqrt[12] ), .A2(new_n13577_), .A3(new_n13596_), .ZN(new_n14029_));
  XOR2_X1    g13837(.A1(new_n14029_), .A2(new_n13611_), .Z(new_n14030_));
  INV_X1     g13838(.I(new_n14030_), .ZN(new_n14031_));
  OAI21_X1   g13839(.A1(new_n13571_), .A2(new_n13573_), .B(new_n13576_), .ZN(new_n14032_));
  NOR2_X1    g13840(.A1(new_n13917_), .A2(new_n14032_), .ZN(new_n14033_));
  XOR2_X1    g13841(.A1(new_n14033_), .A2(new_n13483_), .Z(new_n14034_));
  NAND3_X1   g13842(.A1(\asqrt[12] ), .A2(new_n13590_), .A3(new_n13572_), .ZN(new_n14035_));
  XOR2_X1    g13843(.A1(new_n14035_), .A2(new_n13487_), .Z(new_n14036_));
  OAI21_X1   g13844(.A1(new_n13585_), .A2(new_n13586_), .B(new_n13589_), .ZN(new_n14037_));
  NOR2_X1    g13845(.A1(new_n13917_), .A2(new_n14037_), .ZN(new_n14038_));
  XOR2_X1    g13846(.A1(new_n14038_), .A2(new_n13489_), .Z(new_n14039_));
  INV_X1     g13847(.I(new_n14039_), .ZN(new_n14040_));
  NAND3_X1   g13848(.A1(\asqrt[12] ), .A2(new_n13549_), .A3(new_n13568_), .ZN(new_n14041_));
  XOR2_X1    g13849(.A1(new_n14041_), .A2(new_n13583_), .Z(new_n14042_));
  INV_X1     g13850(.I(new_n14042_), .ZN(new_n14043_));
  OAI21_X1   g13851(.A1(new_n13543_), .A2(new_n13545_), .B(new_n13548_), .ZN(new_n14044_));
  NOR2_X1    g13852(.A1(new_n13917_), .A2(new_n14044_), .ZN(new_n14045_));
  XOR2_X1    g13853(.A1(new_n14045_), .A2(new_n13496_), .Z(new_n14046_));
  NAND3_X1   g13854(.A1(\asqrt[12] ), .A2(new_n13562_), .A3(new_n13544_), .ZN(new_n14047_));
  XOR2_X1    g13855(.A1(new_n14047_), .A2(new_n13499_), .Z(new_n14048_));
  OAI21_X1   g13856(.A1(new_n13557_), .A2(new_n13558_), .B(new_n13561_), .ZN(new_n14049_));
  NOR2_X1    g13857(.A1(new_n13917_), .A2(new_n14049_), .ZN(new_n14050_));
  XOR2_X1    g13858(.A1(new_n14050_), .A2(new_n13502_), .Z(new_n14051_));
  INV_X1     g13859(.I(new_n14051_), .ZN(new_n14052_));
  NAND3_X1   g13860(.A1(\asqrt[12] ), .A2(new_n13522_), .A3(new_n13540_), .ZN(new_n14053_));
  XOR2_X1    g13861(.A1(new_n14053_), .A2(new_n13556_), .Z(new_n14054_));
  INV_X1     g13862(.I(new_n14054_), .ZN(new_n14055_));
  NOR2_X1    g13863(.A1(new_n13519_), .A2(\asqrt[15] ), .ZN(new_n14056_));
  NOR3_X1    g13864(.A1(new_n13917_), .A2(new_n14056_), .A3(new_n13539_), .ZN(new_n14057_));
  XOR2_X1    g13865(.A1(new_n14057_), .A2(new_n13510_), .Z(new_n14058_));
  NOR3_X1    g13866(.A1(new_n13917_), .A2(\a[24] ), .A3(\a[25] ), .ZN(new_n14059_));
  NOR4_X1    g13867(.A1(new_n13915_), .A2(new_n13382_), .A3(new_n13792_), .A4(new_n13916_), .ZN(new_n14060_));
  OAI21_X1   g13868(.A1(new_n14059_), .A2(new_n14060_), .B(new_n13032_), .ZN(new_n14061_));
  NAND3_X1   g13869(.A1(\asqrt[12] ), .A2(new_n13511_), .A3(new_n13512_), .ZN(new_n14062_));
  INV_X1     g13870(.I(new_n14060_), .ZN(new_n14063_));
  NAND3_X1   g13871(.A1(new_n14062_), .A2(\a[26] ), .A3(new_n14063_), .ZN(new_n14064_));
  NAND2_X1   g13872(.A1(new_n14061_), .A2(new_n14064_), .ZN(new_n14065_));
  INV_X1     g13873(.I(\a[22] ), .ZN(new_n14066_));
  INV_X1     g13874(.I(\a[23] ), .ZN(new_n14067_));
  NAND3_X1   g13875(.A1(new_n14066_), .A2(new_n14067_), .A3(new_n13511_), .ZN(new_n14068_));
  NAND2_X1   g13876(.A1(\asqrt[12] ), .A2(\a[24] ), .ZN(new_n14069_));
  AOI21_X1   g13877(.A1(new_n14069_), .A2(new_n14068_), .B(new_n13382_), .ZN(new_n14070_));
  AOI21_X1   g13878(.A1(\asqrt[12] ), .A2(new_n13511_), .B(new_n13512_), .ZN(new_n14071_));
  NOR2_X1    g13879(.A1(new_n14059_), .A2(new_n14071_), .ZN(new_n14072_));
  NAND3_X1   g13880(.A1(new_n14069_), .A2(new_n13382_), .A3(new_n14068_), .ZN(new_n14073_));
  AOI21_X1   g13881(.A1(new_n14072_), .A2(new_n14073_), .B(new_n14070_), .ZN(new_n14074_));
  AOI21_X1   g13882(.A1(new_n14074_), .A2(new_n12889_), .B(new_n14065_), .ZN(new_n14075_));
  NOR2_X1    g13883(.A1(new_n14074_), .A2(new_n12889_), .ZN(new_n14076_));
  NOR3_X1    g13884(.A1(new_n14075_), .A2(\asqrt[15] ), .A3(new_n14076_), .ZN(new_n14077_));
  NOR3_X1    g13885(.A1(new_n13917_), .A2(new_n13533_), .A3(new_n13518_), .ZN(new_n14078_));
  XOR2_X1    g13886(.A1(new_n14078_), .A2(new_n13535_), .Z(new_n14079_));
  INV_X1     g13887(.I(new_n14079_), .ZN(new_n14080_));
  OAI21_X1   g13888(.A1(new_n14075_), .A2(new_n14076_), .B(\asqrt[15] ), .ZN(new_n14081_));
  OAI21_X1   g13889(.A1(new_n14077_), .A2(new_n14080_), .B(new_n14081_), .ZN(new_n14082_));
  OAI21_X1   g13890(.A1(new_n14082_), .A2(\asqrt[16] ), .B(new_n14058_), .ZN(new_n14083_));
  AOI21_X1   g13891(.A1(new_n14082_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n14084_));
  AOI21_X1   g13892(.A1(new_n14084_), .A2(new_n14083_), .B(new_n14055_), .ZN(new_n14085_));
  NAND2_X1   g13893(.A1(new_n14082_), .A2(\asqrt[16] ), .ZN(new_n14086_));
  AOI21_X1   g13894(.A1(new_n14083_), .A2(new_n14086_), .B(new_n11406_), .ZN(new_n14087_));
  NOR2_X1    g13895(.A1(new_n14085_), .A2(new_n14087_), .ZN(new_n14088_));
  AOI21_X1   g13896(.A1(new_n14088_), .A2(new_n10953_), .B(new_n14052_), .ZN(new_n14089_));
  OAI21_X1   g13897(.A1(new_n14085_), .A2(new_n14087_), .B(\asqrt[18] ), .ZN(new_n14090_));
  NAND2_X1   g13898(.A1(new_n14090_), .A2(new_n10478_), .ZN(new_n14091_));
  OAI21_X1   g13899(.A1(new_n14089_), .A2(new_n14091_), .B(new_n14048_), .ZN(new_n14092_));
  INV_X1     g13900(.I(new_n14090_), .ZN(new_n14093_));
  OAI21_X1   g13901(.A1(new_n14089_), .A2(new_n14093_), .B(\asqrt[19] ), .ZN(new_n14094_));
  NAND3_X1   g13902(.A1(new_n14092_), .A2(new_n14094_), .A3(new_n10045_), .ZN(new_n14095_));
  NAND2_X1   g13903(.A1(new_n14095_), .A2(new_n14046_), .ZN(new_n14096_));
  NAND2_X1   g13904(.A1(new_n14092_), .A2(new_n14094_), .ZN(new_n14097_));
  AOI21_X1   g13905(.A1(new_n14097_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n14098_));
  AOI21_X1   g13906(.A1(new_n14098_), .A2(new_n14096_), .B(new_n14043_), .ZN(new_n14099_));
  INV_X1     g13907(.I(new_n14048_), .ZN(new_n14100_));
  INV_X1     g13908(.I(new_n14058_), .ZN(new_n14101_));
  AOI21_X1   g13909(.A1(new_n14062_), .A2(new_n14063_), .B(\a[26] ), .ZN(new_n14102_));
  NOR3_X1    g13910(.A1(new_n14059_), .A2(new_n13032_), .A3(new_n14060_), .ZN(new_n14103_));
  NOR2_X1    g13911(.A1(new_n14103_), .A2(new_n14102_), .ZN(new_n14104_));
  OAI21_X1   g13912(.A1(new_n13917_), .A2(new_n13511_), .B(new_n14068_), .ZN(new_n14105_));
  NAND2_X1   g13913(.A1(new_n14105_), .A2(\asqrt[13] ), .ZN(new_n14106_));
  OAI21_X1   g13914(.A1(new_n13917_), .A2(\a[24] ), .B(\a[25] ), .ZN(new_n14107_));
  NAND2_X1   g13915(.A1(new_n14107_), .A2(new_n14062_), .ZN(new_n14108_));
  NOR2_X1    g13916(.A1(new_n14105_), .A2(\asqrt[13] ), .ZN(new_n14109_));
  OAI21_X1   g13917(.A1(new_n14108_), .A2(new_n14109_), .B(new_n14106_), .ZN(new_n14110_));
  OAI21_X1   g13918(.A1(\asqrt[14] ), .A2(new_n14110_), .B(new_n14104_), .ZN(new_n14111_));
  NAND2_X1   g13919(.A1(new_n14110_), .A2(\asqrt[14] ), .ZN(new_n14112_));
  NAND3_X1   g13920(.A1(new_n14111_), .A2(new_n12374_), .A3(new_n14112_), .ZN(new_n14113_));
  AOI21_X1   g13921(.A1(new_n14111_), .A2(new_n14112_), .B(new_n12374_), .ZN(new_n14114_));
  AOI21_X1   g13922(.A1(new_n14113_), .A2(new_n14079_), .B(new_n14114_), .ZN(new_n14115_));
  AOI21_X1   g13923(.A1(new_n14115_), .A2(new_n11901_), .B(new_n14101_), .ZN(new_n14116_));
  OAI21_X1   g13924(.A1(new_n14115_), .A2(new_n11901_), .B(new_n11406_), .ZN(new_n14117_));
  OAI21_X1   g13925(.A1(new_n14116_), .A2(new_n14117_), .B(new_n14054_), .ZN(new_n14118_));
  NOR2_X1    g13926(.A1(new_n14115_), .A2(new_n11901_), .ZN(new_n14119_));
  OAI21_X1   g13927(.A1(new_n14116_), .A2(new_n14119_), .B(\asqrt[17] ), .ZN(new_n14120_));
  NAND3_X1   g13928(.A1(new_n14118_), .A2(new_n14120_), .A3(new_n10953_), .ZN(new_n14121_));
  NAND2_X1   g13929(.A1(new_n14121_), .A2(new_n14051_), .ZN(new_n14122_));
  NAND2_X1   g13930(.A1(new_n14118_), .A2(new_n14120_), .ZN(new_n14123_));
  AOI21_X1   g13931(.A1(new_n14123_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n14124_));
  AOI21_X1   g13932(.A1(new_n14124_), .A2(new_n14122_), .B(new_n14100_), .ZN(new_n14125_));
  AOI21_X1   g13933(.A1(new_n14122_), .A2(new_n14090_), .B(new_n10478_), .ZN(new_n14126_));
  OAI21_X1   g13934(.A1(new_n14125_), .A2(new_n14126_), .B(\asqrt[20] ), .ZN(new_n14127_));
  AOI21_X1   g13935(.A1(new_n14096_), .A2(new_n14127_), .B(new_n9590_), .ZN(new_n14128_));
  NOR2_X1    g13936(.A1(new_n14099_), .A2(new_n14128_), .ZN(new_n14129_));
  AOI21_X1   g13937(.A1(new_n14129_), .A2(new_n9177_), .B(new_n14040_), .ZN(new_n14130_));
  OAI21_X1   g13938(.A1(new_n14099_), .A2(new_n14128_), .B(\asqrt[22] ), .ZN(new_n14131_));
  NAND2_X1   g13939(.A1(new_n14131_), .A2(new_n8742_), .ZN(new_n14132_));
  OAI21_X1   g13940(.A1(new_n14130_), .A2(new_n14132_), .B(new_n14036_), .ZN(new_n14133_));
  INV_X1     g13941(.I(new_n14131_), .ZN(new_n14134_));
  OAI21_X1   g13942(.A1(new_n14130_), .A2(new_n14134_), .B(\asqrt[23] ), .ZN(new_n14135_));
  NAND3_X1   g13943(.A1(new_n14133_), .A2(new_n14135_), .A3(new_n8349_), .ZN(new_n14136_));
  NAND2_X1   g13944(.A1(new_n14136_), .A2(new_n14034_), .ZN(new_n14137_));
  NAND2_X1   g13945(.A1(new_n14133_), .A2(new_n14135_), .ZN(new_n14138_));
  AOI21_X1   g13946(.A1(new_n14138_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n14139_));
  AOI21_X1   g13947(.A1(new_n14139_), .A2(new_n14137_), .B(new_n14031_), .ZN(new_n14140_));
  INV_X1     g13948(.I(new_n14036_), .ZN(new_n14141_));
  INV_X1     g13949(.I(new_n14046_), .ZN(new_n14142_));
  NOR2_X1    g13950(.A1(new_n14125_), .A2(new_n14126_), .ZN(new_n14143_));
  AOI21_X1   g13951(.A1(new_n14143_), .A2(new_n10045_), .B(new_n14142_), .ZN(new_n14144_));
  NAND2_X1   g13952(.A1(new_n14127_), .A2(new_n9590_), .ZN(new_n14145_));
  OAI21_X1   g13953(.A1(new_n14144_), .A2(new_n14145_), .B(new_n14042_), .ZN(new_n14146_));
  INV_X1     g13954(.I(new_n14127_), .ZN(new_n14147_));
  OAI21_X1   g13955(.A1(new_n14144_), .A2(new_n14147_), .B(\asqrt[21] ), .ZN(new_n14148_));
  NAND3_X1   g13956(.A1(new_n14146_), .A2(new_n14148_), .A3(new_n9177_), .ZN(new_n14149_));
  NAND2_X1   g13957(.A1(new_n14149_), .A2(new_n14039_), .ZN(new_n14150_));
  NAND2_X1   g13958(.A1(new_n14146_), .A2(new_n14148_), .ZN(new_n14151_));
  AOI21_X1   g13959(.A1(new_n14151_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n14152_));
  AOI21_X1   g13960(.A1(new_n14152_), .A2(new_n14150_), .B(new_n14141_), .ZN(new_n14153_));
  AOI21_X1   g13961(.A1(new_n14150_), .A2(new_n14131_), .B(new_n8742_), .ZN(new_n14154_));
  OAI21_X1   g13962(.A1(new_n14153_), .A2(new_n14154_), .B(\asqrt[24] ), .ZN(new_n14155_));
  AOI21_X1   g13963(.A1(new_n14137_), .A2(new_n14155_), .B(new_n7934_), .ZN(new_n14156_));
  NOR2_X1    g13964(.A1(new_n14140_), .A2(new_n14156_), .ZN(new_n14157_));
  AOI21_X1   g13965(.A1(new_n14157_), .A2(new_n7561_), .B(new_n14028_), .ZN(new_n14158_));
  OAI21_X1   g13966(.A1(new_n14140_), .A2(new_n14156_), .B(\asqrt[26] ), .ZN(new_n14159_));
  NAND2_X1   g13967(.A1(new_n14159_), .A2(new_n7166_), .ZN(new_n14160_));
  OAI21_X1   g13968(.A1(new_n14158_), .A2(new_n14160_), .B(new_n14024_), .ZN(new_n14161_));
  INV_X1     g13969(.I(new_n14159_), .ZN(new_n14162_));
  OAI21_X1   g13970(.A1(new_n14158_), .A2(new_n14162_), .B(\asqrt[27] ), .ZN(new_n14163_));
  NAND3_X1   g13971(.A1(new_n14161_), .A2(new_n14163_), .A3(new_n6813_), .ZN(new_n14164_));
  NAND2_X1   g13972(.A1(new_n14164_), .A2(new_n14022_), .ZN(new_n14165_));
  NAND2_X1   g13973(.A1(new_n14161_), .A2(new_n14163_), .ZN(new_n14166_));
  AOI21_X1   g13974(.A1(new_n14166_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n14167_));
  AOI21_X1   g13975(.A1(new_n14167_), .A2(new_n14165_), .B(new_n14019_), .ZN(new_n14168_));
  INV_X1     g13976(.I(new_n14024_), .ZN(new_n14169_));
  INV_X1     g13977(.I(new_n14034_), .ZN(new_n14170_));
  NOR2_X1    g13978(.A1(new_n14153_), .A2(new_n14154_), .ZN(new_n14171_));
  AOI21_X1   g13979(.A1(new_n14171_), .A2(new_n8349_), .B(new_n14170_), .ZN(new_n14172_));
  NAND2_X1   g13980(.A1(new_n14155_), .A2(new_n7934_), .ZN(new_n14173_));
  OAI21_X1   g13981(.A1(new_n14172_), .A2(new_n14173_), .B(new_n14030_), .ZN(new_n14174_));
  INV_X1     g13982(.I(new_n14155_), .ZN(new_n14175_));
  OAI21_X1   g13983(.A1(new_n14172_), .A2(new_n14175_), .B(\asqrt[25] ), .ZN(new_n14176_));
  NAND3_X1   g13984(.A1(new_n14174_), .A2(new_n14176_), .A3(new_n7561_), .ZN(new_n14177_));
  NAND2_X1   g13985(.A1(new_n14177_), .A2(new_n14027_), .ZN(new_n14178_));
  NAND2_X1   g13986(.A1(new_n14174_), .A2(new_n14176_), .ZN(new_n14179_));
  AOI21_X1   g13987(.A1(new_n14179_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n14180_));
  AOI21_X1   g13988(.A1(new_n14180_), .A2(new_n14178_), .B(new_n14169_), .ZN(new_n14181_));
  AOI21_X1   g13989(.A1(new_n14178_), .A2(new_n14159_), .B(new_n7166_), .ZN(new_n14182_));
  OAI21_X1   g13990(.A1(new_n14181_), .A2(new_n14182_), .B(\asqrt[28] ), .ZN(new_n14183_));
  AOI21_X1   g13991(.A1(new_n14165_), .A2(new_n14183_), .B(new_n6454_), .ZN(new_n14184_));
  NOR2_X1    g13992(.A1(new_n14168_), .A2(new_n14184_), .ZN(new_n14185_));
  AOI21_X1   g13993(.A1(new_n14185_), .A2(new_n6106_), .B(new_n14016_), .ZN(new_n14186_));
  OAI21_X1   g13994(.A1(new_n14168_), .A2(new_n14184_), .B(\asqrt[30] ), .ZN(new_n14187_));
  NAND2_X1   g13995(.A1(new_n14187_), .A2(new_n5750_), .ZN(new_n14188_));
  OAI21_X1   g13996(.A1(new_n14186_), .A2(new_n14188_), .B(new_n14012_), .ZN(new_n14189_));
  INV_X1     g13997(.I(new_n14187_), .ZN(new_n14190_));
  OAI21_X1   g13998(.A1(new_n14186_), .A2(new_n14190_), .B(\asqrt[31] ), .ZN(new_n14191_));
  NAND3_X1   g13999(.A1(new_n14189_), .A2(new_n14191_), .A3(new_n5435_), .ZN(new_n14192_));
  NAND2_X1   g14000(.A1(new_n14192_), .A2(new_n14010_), .ZN(new_n14193_));
  NAND2_X1   g14001(.A1(new_n14189_), .A2(new_n14191_), .ZN(new_n14194_));
  AOI21_X1   g14002(.A1(new_n14194_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n14195_));
  AOI21_X1   g14003(.A1(new_n14195_), .A2(new_n14193_), .B(new_n14007_), .ZN(new_n14196_));
  INV_X1     g14004(.I(new_n14012_), .ZN(new_n14197_));
  INV_X1     g14005(.I(new_n14022_), .ZN(new_n14198_));
  NOR2_X1    g14006(.A1(new_n14181_), .A2(new_n14182_), .ZN(new_n14199_));
  AOI21_X1   g14007(.A1(new_n14199_), .A2(new_n6813_), .B(new_n14198_), .ZN(new_n14200_));
  NAND2_X1   g14008(.A1(new_n14183_), .A2(new_n6454_), .ZN(new_n14201_));
  OAI21_X1   g14009(.A1(new_n14200_), .A2(new_n14201_), .B(new_n14018_), .ZN(new_n14202_));
  INV_X1     g14010(.I(new_n14183_), .ZN(new_n14203_));
  OAI21_X1   g14011(.A1(new_n14200_), .A2(new_n14203_), .B(\asqrt[29] ), .ZN(new_n14204_));
  NAND3_X1   g14012(.A1(new_n14202_), .A2(new_n14204_), .A3(new_n6106_), .ZN(new_n14205_));
  NAND2_X1   g14013(.A1(new_n14205_), .A2(new_n14015_), .ZN(new_n14206_));
  NAND2_X1   g14014(.A1(new_n14202_), .A2(new_n14204_), .ZN(new_n14207_));
  AOI21_X1   g14015(.A1(new_n14207_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n14208_));
  AOI21_X1   g14016(.A1(new_n14208_), .A2(new_n14206_), .B(new_n14197_), .ZN(new_n14209_));
  AOI21_X1   g14017(.A1(new_n14206_), .A2(new_n14187_), .B(new_n5750_), .ZN(new_n14210_));
  OAI21_X1   g14018(.A1(new_n14209_), .A2(new_n14210_), .B(\asqrt[32] ), .ZN(new_n14211_));
  AOI21_X1   g14019(.A1(new_n14193_), .A2(new_n14211_), .B(new_n5110_), .ZN(new_n14212_));
  NOR2_X1    g14020(.A1(new_n14196_), .A2(new_n14212_), .ZN(new_n14213_));
  AOI21_X1   g14021(.A1(new_n14213_), .A2(new_n4810_), .B(new_n14004_), .ZN(new_n14214_));
  OAI21_X1   g14022(.A1(new_n14196_), .A2(new_n14212_), .B(\asqrt[34] ), .ZN(new_n14215_));
  NAND2_X1   g14023(.A1(new_n14215_), .A2(new_n4510_), .ZN(new_n14216_));
  OAI21_X1   g14024(.A1(new_n14214_), .A2(new_n14216_), .B(new_n14000_), .ZN(new_n14217_));
  INV_X1     g14025(.I(new_n14215_), .ZN(new_n14218_));
  OAI21_X1   g14026(.A1(new_n14214_), .A2(new_n14218_), .B(\asqrt[35] ), .ZN(new_n14219_));
  NAND3_X1   g14027(.A1(new_n14217_), .A2(new_n14219_), .A3(new_n4224_), .ZN(new_n14220_));
  NAND2_X1   g14028(.A1(new_n14220_), .A2(new_n13998_), .ZN(new_n14221_));
  NAND2_X1   g14029(.A1(new_n14217_), .A2(new_n14219_), .ZN(new_n14222_));
  AOI21_X1   g14030(.A1(new_n14222_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n14223_));
  AOI21_X1   g14031(.A1(new_n14223_), .A2(new_n14221_), .B(new_n13995_), .ZN(new_n14224_));
  INV_X1     g14032(.I(new_n14000_), .ZN(new_n14225_));
  INV_X1     g14033(.I(new_n14010_), .ZN(new_n14226_));
  NOR2_X1    g14034(.A1(new_n14209_), .A2(new_n14210_), .ZN(new_n14227_));
  AOI21_X1   g14035(.A1(new_n14227_), .A2(new_n5435_), .B(new_n14226_), .ZN(new_n14228_));
  NAND2_X1   g14036(.A1(new_n14211_), .A2(new_n5110_), .ZN(new_n14229_));
  OAI21_X1   g14037(.A1(new_n14228_), .A2(new_n14229_), .B(new_n14006_), .ZN(new_n14230_));
  INV_X1     g14038(.I(new_n14211_), .ZN(new_n14231_));
  OAI21_X1   g14039(.A1(new_n14228_), .A2(new_n14231_), .B(\asqrt[33] ), .ZN(new_n14232_));
  NAND3_X1   g14040(.A1(new_n14230_), .A2(new_n14232_), .A3(new_n4810_), .ZN(new_n14233_));
  NAND2_X1   g14041(.A1(new_n14233_), .A2(new_n14003_), .ZN(new_n14234_));
  NAND2_X1   g14042(.A1(new_n14230_), .A2(new_n14232_), .ZN(new_n14235_));
  AOI21_X1   g14043(.A1(new_n14235_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n14236_));
  AOI21_X1   g14044(.A1(new_n14236_), .A2(new_n14234_), .B(new_n14225_), .ZN(new_n14237_));
  AOI21_X1   g14045(.A1(new_n14234_), .A2(new_n14215_), .B(new_n4510_), .ZN(new_n14238_));
  OAI21_X1   g14046(.A1(new_n14237_), .A2(new_n14238_), .B(\asqrt[36] ), .ZN(new_n14239_));
  AOI21_X1   g14047(.A1(new_n14221_), .A2(new_n14239_), .B(new_n3928_), .ZN(new_n14240_));
  NOR2_X1    g14048(.A1(new_n14224_), .A2(new_n14240_), .ZN(new_n14241_));
  AOI21_X1   g14049(.A1(new_n14241_), .A2(new_n3675_), .B(new_n13992_), .ZN(new_n14242_));
  OAI21_X1   g14050(.A1(new_n14224_), .A2(new_n14240_), .B(\asqrt[38] ), .ZN(new_n14243_));
  NAND2_X1   g14051(.A1(new_n14243_), .A2(new_n3400_), .ZN(new_n14244_));
  OAI21_X1   g14052(.A1(new_n14242_), .A2(new_n14244_), .B(new_n13988_), .ZN(new_n14245_));
  INV_X1     g14053(.I(new_n14243_), .ZN(new_n14246_));
  OAI21_X1   g14054(.A1(new_n14242_), .A2(new_n14246_), .B(\asqrt[39] ), .ZN(new_n14247_));
  NAND3_X1   g14055(.A1(new_n14245_), .A2(new_n14247_), .A3(new_n3167_), .ZN(new_n14248_));
  NAND2_X1   g14056(.A1(new_n14248_), .A2(new_n13986_), .ZN(new_n14249_));
  NAND2_X1   g14057(.A1(new_n14245_), .A2(new_n14247_), .ZN(new_n14250_));
  AOI21_X1   g14058(.A1(new_n14250_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n14251_));
  AOI21_X1   g14059(.A1(new_n14251_), .A2(new_n14249_), .B(new_n13983_), .ZN(new_n14252_));
  INV_X1     g14060(.I(new_n13988_), .ZN(new_n14253_));
  INV_X1     g14061(.I(new_n13998_), .ZN(new_n14254_));
  NOR2_X1    g14062(.A1(new_n14237_), .A2(new_n14238_), .ZN(new_n14255_));
  AOI21_X1   g14063(.A1(new_n14255_), .A2(new_n4224_), .B(new_n14254_), .ZN(new_n14256_));
  NAND2_X1   g14064(.A1(new_n14239_), .A2(new_n3928_), .ZN(new_n14257_));
  OAI21_X1   g14065(.A1(new_n14256_), .A2(new_n14257_), .B(new_n13994_), .ZN(new_n14258_));
  INV_X1     g14066(.I(new_n14239_), .ZN(new_n14259_));
  OAI21_X1   g14067(.A1(new_n14256_), .A2(new_n14259_), .B(\asqrt[37] ), .ZN(new_n14260_));
  NAND3_X1   g14068(.A1(new_n14258_), .A2(new_n14260_), .A3(new_n3675_), .ZN(new_n14261_));
  NAND2_X1   g14069(.A1(new_n14261_), .A2(new_n13991_), .ZN(new_n14262_));
  NAND2_X1   g14070(.A1(new_n14258_), .A2(new_n14260_), .ZN(new_n14263_));
  AOI21_X1   g14071(.A1(new_n14263_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n14264_));
  AOI21_X1   g14072(.A1(new_n14264_), .A2(new_n14262_), .B(new_n14253_), .ZN(new_n14265_));
  AOI21_X1   g14073(.A1(new_n14262_), .A2(new_n14243_), .B(new_n3400_), .ZN(new_n14266_));
  OAI21_X1   g14074(.A1(new_n14265_), .A2(new_n14266_), .B(\asqrt[40] ), .ZN(new_n14267_));
  AOI21_X1   g14075(.A1(new_n14249_), .A2(new_n14267_), .B(new_n2912_), .ZN(new_n14268_));
  NOR2_X1    g14076(.A1(new_n14252_), .A2(new_n14268_), .ZN(new_n14269_));
  AOI21_X1   g14077(.A1(new_n14269_), .A2(new_n2699_), .B(new_n13980_), .ZN(new_n14270_));
  OAI21_X1   g14078(.A1(new_n14252_), .A2(new_n14268_), .B(\asqrt[42] ), .ZN(new_n14271_));
  NAND2_X1   g14079(.A1(new_n14271_), .A2(new_n2464_), .ZN(new_n14272_));
  OAI21_X1   g14080(.A1(new_n14270_), .A2(new_n14272_), .B(new_n13976_), .ZN(new_n14273_));
  INV_X1     g14081(.I(new_n14271_), .ZN(new_n14274_));
  OAI21_X1   g14082(.A1(new_n14270_), .A2(new_n14274_), .B(\asqrt[43] ), .ZN(new_n14275_));
  NAND3_X1   g14083(.A1(new_n14273_), .A2(new_n14275_), .A3(new_n2271_), .ZN(new_n14276_));
  NAND2_X1   g14084(.A1(new_n14276_), .A2(new_n13974_), .ZN(new_n14277_));
  NAND2_X1   g14085(.A1(new_n14273_), .A2(new_n14275_), .ZN(new_n14278_));
  AOI21_X1   g14086(.A1(new_n14278_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n14279_));
  AOI21_X1   g14087(.A1(new_n14279_), .A2(new_n14277_), .B(new_n13971_), .ZN(new_n14280_));
  INV_X1     g14088(.I(new_n13976_), .ZN(new_n14281_));
  INV_X1     g14089(.I(new_n13986_), .ZN(new_n14282_));
  NOR2_X1    g14090(.A1(new_n14265_), .A2(new_n14266_), .ZN(new_n14283_));
  AOI21_X1   g14091(.A1(new_n14283_), .A2(new_n3167_), .B(new_n14282_), .ZN(new_n14284_));
  NAND2_X1   g14092(.A1(new_n14267_), .A2(new_n2912_), .ZN(new_n14285_));
  OAI21_X1   g14093(.A1(new_n14284_), .A2(new_n14285_), .B(new_n13982_), .ZN(new_n14286_));
  INV_X1     g14094(.I(new_n14267_), .ZN(new_n14287_));
  OAI21_X1   g14095(.A1(new_n14284_), .A2(new_n14287_), .B(\asqrt[41] ), .ZN(new_n14288_));
  NAND3_X1   g14096(.A1(new_n14286_), .A2(new_n14288_), .A3(new_n2699_), .ZN(new_n14289_));
  NAND2_X1   g14097(.A1(new_n14289_), .A2(new_n13979_), .ZN(new_n14290_));
  NAND2_X1   g14098(.A1(new_n14286_), .A2(new_n14288_), .ZN(new_n14291_));
  AOI21_X1   g14099(.A1(new_n14291_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n14292_));
  AOI21_X1   g14100(.A1(new_n14292_), .A2(new_n14290_), .B(new_n14281_), .ZN(new_n14293_));
  AOI21_X1   g14101(.A1(new_n14290_), .A2(new_n14271_), .B(new_n2464_), .ZN(new_n14294_));
  OAI21_X1   g14102(.A1(new_n14293_), .A2(new_n14294_), .B(\asqrt[44] ), .ZN(new_n14295_));
  AOI21_X1   g14103(.A1(new_n14277_), .A2(new_n14295_), .B(new_n2072_), .ZN(new_n14296_));
  NOR2_X1    g14104(.A1(new_n14280_), .A2(new_n14296_), .ZN(new_n14297_));
  AOI21_X1   g14105(.A1(new_n14297_), .A2(new_n1884_), .B(new_n13968_), .ZN(new_n14298_));
  OAI21_X1   g14106(.A1(new_n14280_), .A2(new_n14296_), .B(\asqrt[46] ), .ZN(new_n14299_));
  NAND2_X1   g14107(.A1(new_n14299_), .A2(new_n1688_), .ZN(new_n14300_));
  OAI21_X1   g14108(.A1(new_n14298_), .A2(new_n14300_), .B(new_n13964_), .ZN(new_n14301_));
  INV_X1     g14109(.I(new_n14299_), .ZN(new_n14302_));
  OAI21_X1   g14110(.A1(new_n14298_), .A2(new_n14302_), .B(\asqrt[47] ), .ZN(new_n14303_));
  NAND3_X1   g14111(.A1(new_n14301_), .A2(new_n14303_), .A3(new_n1533_), .ZN(new_n14304_));
  NAND2_X1   g14112(.A1(new_n14304_), .A2(new_n13962_), .ZN(new_n14305_));
  NAND2_X1   g14113(.A1(new_n14301_), .A2(new_n14303_), .ZN(new_n14306_));
  AOI21_X1   g14114(.A1(new_n14306_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n14307_));
  AOI21_X1   g14115(.A1(new_n14307_), .A2(new_n14305_), .B(new_n13959_), .ZN(new_n14308_));
  INV_X1     g14116(.I(new_n13964_), .ZN(new_n14309_));
  INV_X1     g14117(.I(new_n13974_), .ZN(new_n14310_));
  NOR2_X1    g14118(.A1(new_n14293_), .A2(new_n14294_), .ZN(new_n14311_));
  AOI21_X1   g14119(.A1(new_n14311_), .A2(new_n2271_), .B(new_n14310_), .ZN(new_n14312_));
  NAND2_X1   g14120(.A1(new_n14295_), .A2(new_n2072_), .ZN(new_n14313_));
  OAI21_X1   g14121(.A1(new_n14312_), .A2(new_n14313_), .B(new_n13970_), .ZN(new_n14314_));
  INV_X1     g14122(.I(new_n14295_), .ZN(new_n14315_));
  OAI21_X1   g14123(.A1(new_n14312_), .A2(new_n14315_), .B(\asqrt[45] ), .ZN(new_n14316_));
  NAND3_X1   g14124(.A1(new_n14314_), .A2(new_n14316_), .A3(new_n1884_), .ZN(new_n14317_));
  NAND2_X1   g14125(.A1(new_n14317_), .A2(new_n13967_), .ZN(new_n14318_));
  NAND2_X1   g14126(.A1(new_n14314_), .A2(new_n14316_), .ZN(new_n14319_));
  AOI21_X1   g14127(.A1(new_n14319_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n14320_));
  AOI21_X1   g14128(.A1(new_n14320_), .A2(new_n14318_), .B(new_n14309_), .ZN(new_n14321_));
  AOI21_X1   g14129(.A1(new_n14318_), .A2(new_n14299_), .B(new_n1688_), .ZN(new_n14322_));
  OAI21_X1   g14130(.A1(new_n14321_), .A2(new_n14322_), .B(\asqrt[48] ), .ZN(new_n14323_));
  AOI21_X1   g14131(.A1(new_n14305_), .A2(new_n14323_), .B(new_n1368_), .ZN(new_n14324_));
  NOR2_X1    g14132(.A1(new_n14308_), .A2(new_n14324_), .ZN(new_n14325_));
  AOI21_X1   g14133(.A1(new_n14325_), .A2(new_n1228_), .B(new_n13956_), .ZN(new_n14326_));
  OAI21_X1   g14134(.A1(new_n14308_), .A2(new_n14324_), .B(\asqrt[50] ), .ZN(new_n14327_));
  NAND2_X1   g14135(.A1(new_n14327_), .A2(new_n1088_), .ZN(new_n14328_));
  OAI21_X1   g14136(.A1(new_n14326_), .A2(new_n14328_), .B(new_n13952_), .ZN(new_n14329_));
  INV_X1     g14137(.I(new_n14327_), .ZN(new_n14330_));
  OAI21_X1   g14138(.A1(new_n14326_), .A2(new_n14330_), .B(\asqrt[51] ), .ZN(new_n14331_));
  NAND3_X1   g14139(.A1(new_n14329_), .A2(new_n14331_), .A3(new_n962_), .ZN(new_n14332_));
  NAND2_X1   g14140(.A1(new_n14332_), .A2(new_n13950_), .ZN(new_n14333_));
  NAND2_X1   g14141(.A1(new_n14329_), .A2(new_n14331_), .ZN(new_n14334_));
  AOI21_X1   g14142(.A1(new_n14334_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n14335_));
  AOI21_X1   g14143(.A1(new_n14335_), .A2(new_n14333_), .B(new_n13947_), .ZN(new_n14336_));
  INV_X1     g14144(.I(new_n13952_), .ZN(new_n14337_));
  INV_X1     g14145(.I(new_n13962_), .ZN(new_n14338_));
  NOR2_X1    g14146(.A1(new_n14321_), .A2(new_n14322_), .ZN(new_n14339_));
  AOI21_X1   g14147(.A1(new_n14339_), .A2(new_n1533_), .B(new_n14338_), .ZN(new_n14340_));
  NAND2_X1   g14148(.A1(new_n14323_), .A2(new_n1368_), .ZN(new_n14341_));
  OAI21_X1   g14149(.A1(new_n14340_), .A2(new_n14341_), .B(new_n13958_), .ZN(new_n14342_));
  INV_X1     g14150(.I(new_n14323_), .ZN(new_n14343_));
  OAI21_X1   g14151(.A1(new_n14340_), .A2(new_n14343_), .B(\asqrt[49] ), .ZN(new_n14344_));
  NAND3_X1   g14152(.A1(new_n14342_), .A2(new_n14344_), .A3(new_n1228_), .ZN(new_n14345_));
  NAND2_X1   g14153(.A1(new_n14345_), .A2(new_n13955_), .ZN(new_n14346_));
  NAND2_X1   g14154(.A1(new_n14342_), .A2(new_n14344_), .ZN(new_n14347_));
  AOI21_X1   g14155(.A1(new_n14347_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n14348_));
  AOI21_X1   g14156(.A1(new_n14348_), .A2(new_n14346_), .B(new_n14337_), .ZN(new_n14349_));
  AOI21_X1   g14157(.A1(new_n14346_), .A2(new_n14327_), .B(new_n1088_), .ZN(new_n14350_));
  OAI21_X1   g14158(.A1(new_n14349_), .A2(new_n14350_), .B(\asqrt[52] ), .ZN(new_n14351_));
  AOI21_X1   g14159(.A1(new_n14333_), .A2(new_n14351_), .B(new_n842_), .ZN(new_n14352_));
  NOR2_X1    g14160(.A1(new_n14336_), .A2(new_n14352_), .ZN(new_n14353_));
  AOI21_X1   g14161(.A1(new_n14353_), .A2(new_n720_), .B(new_n13946_), .ZN(new_n14354_));
  OAI21_X1   g14162(.A1(new_n14336_), .A2(new_n14352_), .B(\asqrt[54] ), .ZN(new_n14355_));
  NAND2_X1   g14163(.A1(new_n14355_), .A2(new_n630_), .ZN(new_n14356_));
  OAI21_X1   g14164(.A1(new_n14354_), .A2(new_n14356_), .B(new_n13942_), .ZN(new_n14357_));
  INV_X1     g14165(.I(new_n14355_), .ZN(new_n14358_));
  OAI21_X1   g14166(.A1(new_n14354_), .A2(new_n14358_), .B(\asqrt[55] ), .ZN(new_n14359_));
  NAND3_X1   g14167(.A1(new_n14357_), .A2(new_n14359_), .A3(new_n545_), .ZN(new_n14360_));
  NAND2_X1   g14168(.A1(new_n14360_), .A2(new_n13940_), .ZN(new_n14361_));
  NAND2_X1   g14169(.A1(new_n14357_), .A2(new_n14359_), .ZN(new_n14362_));
  AOI21_X1   g14170(.A1(new_n14362_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n14363_));
  AOI21_X1   g14171(.A1(new_n14363_), .A2(new_n14361_), .B(new_n13937_), .ZN(new_n14364_));
  INV_X1     g14172(.I(new_n13942_), .ZN(new_n14365_));
  INV_X1     g14173(.I(new_n13950_), .ZN(new_n14366_));
  NOR2_X1    g14174(.A1(new_n14349_), .A2(new_n14350_), .ZN(new_n14367_));
  AOI21_X1   g14175(.A1(new_n14367_), .A2(new_n962_), .B(new_n14366_), .ZN(new_n14368_));
  NAND2_X1   g14176(.A1(new_n14351_), .A2(new_n842_), .ZN(new_n14369_));
  OAI21_X1   g14177(.A1(new_n14368_), .A2(new_n14369_), .B(new_n13900_), .ZN(new_n14370_));
  INV_X1     g14178(.I(new_n14351_), .ZN(new_n14371_));
  OAI21_X1   g14179(.A1(new_n14368_), .A2(new_n14371_), .B(\asqrt[53] ), .ZN(new_n14372_));
  NAND3_X1   g14180(.A1(new_n14370_), .A2(new_n14372_), .A3(new_n720_), .ZN(new_n14373_));
  NAND2_X1   g14181(.A1(new_n14373_), .A2(new_n13945_), .ZN(new_n14374_));
  NAND2_X1   g14182(.A1(new_n14370_), .A2(new_n14372_), .ZN(new_n14375_));
  AOI21_X1   g14183(.A1(new_n14375_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n14376_));
  AOI21_X1   g14184(.A1(new_n14376_), .A2(new_n14374_), .B(new_n14365_), .ZN(new_n14377_));
  AOI21_X1   g14185(.A1(new_n14374_), .A2(new_n14355_), .B(new_n630_), .ZN(new_n14378_));
  OAI21_X1   g14186(.A1(new_n14377_), .A2(new_n14378_), .B(\asqrt[56] ), .ZN(new_n14379_));
  AOI21_X1   g14187(.A1(new_n14361_), .A2(new_n14379_), .B(new_n450_), .ZN(new_n14380_));
  NOR2_X1    g14188(.A1(new_n14364_), .A2(new_n14380_), .ZN(new_n14381_));
  AOI21_X1   g14189(.A1(new_n14381_), .A2(new_n403_), .B(new_n13934_), .ZN(new_n14382_));
  OAI21_X1   g14190(.A1(new_n14364_), .A2(new_n14380_), .B(\asqrt[58] ), .ZN(new_n14383_));
  NAND2_X1   g14191(.A1(new_n14383_), .A2(new_n339_), .ZN(new_n14384_));
  OAI21_X1   g14192(.A1(new_n14382_), .A2(new_n14384_), .B(new_n13930_), .ZN(new_n14385_));
  INV_X1     g14193(.I(new_n14383_), .ZN(new_n14386_));
  OAI21_X1   g14194(.A1(new_n14382_), .A2(new_n14386_), .B(\asqrt[59] ), .ZN(new_n14387_));
  NAND3_X1   g14195(.A1(new_n14385_), .A2(new_n14387_), .A3(new_n288_), .ZN(new_n14388_));
  NAND2_X1   g14196(.A1(new_n14388_), .A2(new_n13928_), .ZN(new_n14389_));
  INV_X1     g14197(.I(new_n13930_), .ZN(new_n14390_));
  INV_X1     g14198(.I(new_n13940_), .ZN(new_n14391_));
  NOR2_X1    g14199(.A1(new_n14377_), .A2(new_n14378_), .ZN(new_n14392_));
  AOI21_X1   g14200(.A1(new_n14392_), .A2(new_n545_), .B(new_n14391_), .ZN(new_n14393_));
  NAND2_X1   g14201(.A1(new_n14379_), .A2(new_n450_), .ZN(new_n14394_));
  OAI21_X1   g14202(.A1(new_n14393_), .A2(new_n14394_), .B(new_n13936_), .ZN(new_n14395_));
  INV_X1     g14203(.I(new_n14379_), .ZN(new_n14396_));
  OAI21_X1   g14204(.A1(new_n14393_), .A2(new_n14396_), .B(\asqrt[57] ), .ZN(new_n14397_));
  NAND3_X1   g14205(.A1(new_n14395_), .A2(new_n14397_), .A3(new_n403_), .ZN(new_n14398_));
  NAND2_X1   g14206(.A1(new_n14398_), .A2(new_n13933_), .ZN(new_n14399_));
  NAND2_X1   g14207(.A1(new_n14395_), .A2(new_n14397_), .ZN(new_n14400_));
  AOI21_X1   g14208(.A1(new_n14400_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n14401_));
  AOI21_X1   g14209(.A1(new_n14401_), .A2(new_n14399_), .B(new_n14390_), .ZN(new_n14402_));
  AOI21_X1   g14210(.A1(new_n14399_), .A2(new_n14383_), .B(new_n339_), .ZN(new_n14403_));
  OAI21_X1   g14211(.A1(new_n14402_), .A2(new_n14403_), .B(\asqrt[60] ), .ZN(new_n14404_));
  AOI21_X1   g14212(.A1(new_n14389_), .A2(new_n14404_), .B(new_n242_), .ZN(new_n14405_));
  NAND3_X1   g14213(.A1(\asqrt[12] ), .A2(new_n13860_), .A3(new_n13876_), .ZN(new_n14406_));
  XOR2_X1    g14214(.A1(new_n14406_), .A2(new_n13901_), .Z(new_n14407_));
  INV_X1     g14215(.I(new_n14407_), .ZN(new_n14408_));
  NAND2_X1   g14216(.A1(new_n14385_), .A2(new_n14387_), .ZN(new_n14409_));
  AOI21_X1   g14217(.A1(new_n14409_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n14410_));
  AOI21_X1   g14218(.A1(new_n14410_), .A2(new_n14389_), .B(new_n14408_), .ZN(new_n14411_));
  OAI21_X1   g14219(.A1(new_n14411_), .A2(new_n14405_), .B(\asqrt[62] ), .ZN(new_n14412_));
  AOI21_X1   g14220(.A1(new_n13861_), .A2(new_n13882_), .B(new_n13877_), .ZN(new_n14413_));
  NAND2_X1   g14221(.A1(\asqrt[12] ), .A2(new_n14413_), .ZN(new_n14414_));
  XOR2_X1    g14222(.A1(new_n14414_), .A2(new_n13880_), .Z(new_n14415_));
  INV_X1     g14223(.I(new_n13928_), .ZN(new_n14416_));
  NOR2_X1    g14224(.A1(new_n14402_), .A2(new_n14403_), .ZN(new_n14417_));
  AOI21_X1   g14225(.A1(new_n14417_), .A2(new_n288_), .B(new_n14416_), .ZN(new_n14418_));
  INV_X1     g14226(.I(new_n14404_), .ZN(new_n14419_));
  OAI21_X1   g14227(.A1(new_n14418_), .A2(new_n14419_), .B(\asqrt[61] ), .ZN(new_n14420_));
  NAND2_X1   g14228(.A1(new_n14404_), .A2(new_n242_), .ZN(new_n14421_));
  OAI21_X1   g14229(.A1(new_n14418_), .A2(new_n14421_), .B(new_n14407_), .ZN(new_n14422_));
  NAND3_X1   g14230(.A1(new_n14422_), .A2(new_n14420_), .A3(new_n234_), .ZN(new_n14423_));
  NAND2_X1   g14231(.A1(new_n14423_), .A2(new_n14415_), .ZN(new_n14424_));
  AOI21_X1   g14232(.A1(new_n14424_), .A2(new_n14412_), .B(new_n13925_), .ZN(new_n14425_));
  AOI21_X1   g14233(.A1(new_n14425_), .A2(new_n13923_), .B(\asqrt[63] ), .ZN(new_n14426_));
  NAND2_X1   g14234(.A1(new_n14424_), .A2(new_n14412_), .ZN(new_n14427_));
  NOR2_X1    g14235(.A1(new_n14427_), .A2(new_n13923_), .ZN(new_n14428_));
  NOR2_X1    g14236(.A1(\asqrt[12] ), .A2(new_n13912_), .ZN(new_n14429_));
  NOR4_X1    g14237(.A1(new_n14426_), .A2(new_n13920_), .A3(new_n14428_), .A4(new_n14429_), .ZN(new_n14430_));
  OAI21_X1   g14238(.A1(new_n14368_), .A2(new_n14369_), .B(new_n14372_), .ZN(new_n14431_));
  NOR2_X1    g14239(.A1(new_n14430_), .A2(new_n14431_), .ZN(new_n14432_));
  XOR2_X1    g14240(.A1(new_n14432_), .A2(new_n13900_), .Z(new_n14433_));
  INV_X1     g14241(.I(new_n14433_), .ZN(new_n14434_));
  INV_X1     g14242(.I(new_n13920_), .ZN(new_n14435_));
  INV_X1     g14243(.I(new_n14412_), .ZN(new_n14436_));
  NOR2_X1    g14244(.A1(new_n14411_), .A2(new_n14405_), .ZN(new_n14437_));
  INV_X1     g14245(.I(new_n14415_), .ZN(new_n14438_));
  AOI21_X1   g14246(.A1(new_n14437_), .A2(new_n234_), .B(new_n14438_), .ZN(new_n14439_));
  OAI21_X1   g14247(.A1(new_n14439_), .A2(new_n14436_), .B(new_n13924_), .ZN(new_n14440_));
  OAI21_X1   g14248(.A1(new_n14440_), .A2(new_n13922_), .B(new_n193_), .ZN(new_n14441_));
  NOR2_X1    g14249(.A1(new_n14439_), .A2(new_n14436_), .ZN(new_n14442_));
  NAND2_X1   g14250(.A1(new_n14442_), .A2(new_n13922_), .ZN(new_n14443_));
  INV_X1     g14251(.I(new_n14429_), .ZN(new_n14444_));
  NAND4_X1   g14252(.A1(new_n14441_), .A2(new_n14435_), .A3(new_n14443_), .A4(new_n14444_), .ZN(\asqrt[11] ));
  NAND3_X1   g14253(.A1(\asqrt[11] ), .A2(new_n14332_), .A3(new_n14351_), .ZN(new_n14446_));
  XOR2_X1    g14254(.A1(new_n14446_), .A2(new_n14366_), .Z(new_n14447_));
  OAI21_X1   g14255(.A1(new_n14326_), .A2(new_n14328_), .B(new_n14331_), .ZN(new_n14448_));
  NOR2_X1    g14256(.A1(new_n14430_), .A2(new_n14448_), .ZN(new_n14449_));
  XOR2_X1    g14257(.A1(new_n14449_), .A2(new_n13952_), .Z(new_n14450_));
  INV_X1     g14258(.I(new_n14450_), .ZN(new_n14451_));
  NAND3_X1   g14259(.A1(\asqrt[11] ), .A2(new_n14345_), .A3(new_n14327_), .ZN(new_n14452_));
  XOR2_X1    g14260(.A1(new_n14452_), .A2(new_n13956_), .Z(new_n14453_));
  INV_X1     g14261(.I(new_n14453_), .ZN(new_n14454_));
  OAI21_X1   g14262(.A1(new_n14340_), .A2(new_n14341_), .B(new_n14344_), .ZN(new_n14455_));
  NOR2_X1    g14263(.A1(new_n14430_), .A2(new_n14455_), .ZN(new_n14456_));
  XOR2_X1    g14264(.A1(new_n14456_), .A2(new_n13958_), .Z(new_n14457_));
  NAND3_X1   g14265(.A1(\asqrt[11] ), .A2(new_n14304_), .A3(new_n14323_), .ZN(new_n14458_));
  XOR2_X1    g14266(.A1(new_n14458_), .A2(new_n14338_), .Z(new_n14459_));
  OAI21_X1   g14267(.A1(new_n14298_), .A2(new_n14300_), .B(new_n14303_), .ZN(new_n14460_));
  NOR2_X1    g14268(.A1(new_n14430_), .A2(new_n14460_), .ZN(new_n14461_));
  XOR2_X1    g14269(.A1(new_n14461_), .A2(new_n13964_), .Z(new_n14462_));
  INV_X1     g14270(.I(new_n14462_), .ZN(new_n14463_));
  NAND3_X1   g14271(.A1(\asqrt[11] ), .A2(new_n14317_), .A3(new_n14299_), .ZN(new_n14464_));
  XOR2_X1    g14272(.A1(new_n14464_), .A2(new_n13968_), .Z(new_n14465_));
  INV_X1     g14273(.I(new_n14465_), .ZN(new_n14466_));
  OAI21_X1   g14274(.A1(new_n14312_), .A2(new_n14313_), .B(new_n14316_), .ZN(new_n14467_));
  NOR2_X1    g14275(.A1(new_n14430_), .A2(new_n14467_), .ZN(new_n14468_));
  XOR2_X1    g14276(.A1(new_n14468_), .A2(new_n13970_), .Z(new_n14469_));
  NAND3_X1   g14277(.A1(\asqrt[11] ), .A2(new_n14276_), .A3(new_n14295_), .ZN(new_n14470_));
  XOR2_X1    g14278(.A1(new_n14470_), .A2(new_n14310_), .Z(new_n14471_));
  OAI21_X1   g14279(.A1(new_n14270_), .A2(new_n14272_), .B(new_n14275_), .ZN(new_n14472_));
  NOR2_X1    g14280(.A1(new_n14430_), .A2(new_n14472_), .ZN(new_n14473_));
  XOR2_X1    g14281(.A1(new_n14473_), .A2(new_n13976_), .Z(new_n14474_));
  INV_X1     g14282(.I(new_n14474_), .ZN(new_n14475_));
  NAND3_X1   g14283(.A1(\asqrt[11] ), .A2(new_n14289_), .A3(new_n14271_), .ZN(new_n14476_));
  XOR2_X1    g14284(.A1(new_n14476_), .A2(new_n13980_), .Z(new_n14477_));
  INV_X1     g14285(.I(new_n14477_), .ZN(new_n14478_));
  OAI21_X1   g14286(.A1(new_n14284_), .A2(new_n14285_), .B(new_n14288_), .ZN(new_n14479_));
  NOR2_X1    g14287(.A1(new_n14430_), .A2(new_n14479_), .ZN(new_n14480_));
  XOR2_X1    g14288(.A1(new_n14480_), .A2(new_n13982_), .Z(new_n14481_));
  NAND3_X1   g14289(.A1(\asqrt[11] ), .A2(new_n14248_), .A3(new_n14267_), .ZN(new_n14482_));
  XOR2_X1    g14290(.A1(new_n14482_), .A2(new_n14282_), .Z(new_n14483_));
  OAI21_X1   g14291(.A1(new_n14242_), .A2(new_n14244_), .B(new_n14247_), .ZN(new_n14484_));
  NOR2_X1    g14292(.A1(new_n14430_), .A2(new_n14484_), .ZN(new_n14485_));
  XOR2_X1    g14293(.A1(new_n14485_), .A2(new_n13988_), .Z(new_n14486_));
  INV_X1     g14294(.I(new_n14486_), .ZN(new_n14487_));
  NAND3_X1   g14295(.A1(\asqrt[11] ), .A2(new_n14261_), .A3(new_n14243_), .ZN(new_n14488_));
  XOR2_X1    g14296(.A1(new_n14488_), .A2(new_n13992_), .Z(new_n14489_));
  INV_X1     g14297(.I(new_n14489_), .ZN(new_n14490_));
  OAI21_X1   g14298(.A1(new_n14256_), .A2(new_n14257_), .B(new_n14260_), .ZN(new_n14491_));
  NOR2_X1    g14299(.A1(new_n14430_), .A2(new_n14491_), .ZN(new_n14492_));
  XOR2_X1    g14300(.A1(new_n14492_), .A2(new_n13994_), .Z(new_n14493_));
  NAND3_X1   g14301(.A1(\asqrt[11] ), .A2(new_n14220_), .A3(new_n14239_), .ZN(new_n14494_));
  XOR2_X1    g14302(.A1(new_n14494_), .A2(new_n14254_), .Z(new_n14495_));
  OAI21_X1   g14303(.A1(new_n14214_), .A2(new_n14216_), .B(new_n14219_), .ZN(new_n14496_));
  NOR2_X1    g14304(.A1(new_n14430_), .A2(new_n14496_), .ZN(new_n14497_));
  XOR2_X1    g14305(.A1(new_n14497_), .A2(new_n14000_), .Z(new_n14498_));
  INV_X1     g14306(.I(new_n14498_), .ZN(new_n14499_));
  NAND3_X1   g14307(.A1(\asqrt[11] ), .A2(new_n14233_), .A3(new_n14215_), .ZN(new_n14500_));
  XOR2_X1    g14308(.A1(new_n14500_), .A2(new_n14004_), .Z(new_n14501_));
  INV_X1     g14309(.I(new_n14501_), .ZN(new_n14502_));
  OAI21_X1   g14310(.A1(new_n14228_), .A2(new_n14229_), .B(new_n14232_), .ZN(new_n14503_));
  NOR2_X1    g14311(.A1(new_n14430_), .A2(new_n14503_), .ZN(new_n14504_));
  XOR2_X1    g14312(.A1(new_n14504_), .A2(new_n14006_), .Z(new_n14505_));
  NAND3_X1   g14313(.A1(\asqrt[11] ), .A2(new_n14192_), .A3(new_n14211_), .ZN(new_n14506_));
  XOR2_X1    g14314(.A1(new_n14506_), .A2(new_n14226_), .Z(new_n14507_));
  OAI21_X1   g14315(.A1(new_n14186_), .A2(new_n14188_), .B(new_n14191_), .ZN(new_n14508_));
  NOR2_X1    g14316(.A1(new_n14430_), .A2(new_n14508_), .ZN(new_n14509_));
  XOR2_X1    g14317(.A1(new_n14509_), .A2(new_n14012_), .Z(new_n14510_));
  INV_X1     g14318(.I(new_n14510_), .ZN(new_n14511_));
  NAND3_X1   g14319(.A1(\asqrt[11] ), .A2(new_n14205_), .A3(new_n14187_), .ZN(new_n14512_));
  XOR2_X1    g14320(.A1(new_n14512_), .A2(new_n14016_), .Z(new_n14513_));
  INV_X1     g14321(.I(new_n14513_), .ZN(new_n14514_));
  OAI21_X1   g14322(.A1(new_n14200_), .A2(new_n14201_), .B(new_n14204_), .ZN(new_n14515_));
  NOR2_X1    g14323(.A1(new_n14430_), .A2(new_n14515_), .ZN(new_n14516_));
  XOR2_X1    g14324(.A1(new_n14516_), .A2(new_n14018_), .Z(new_n14517_));
  NAND3_X1   g14325(.A1(\asqrt[11] ), .A2(new_n14164_), .A3(new_n14183_), .ZN(new_n14518_));
  XOR2_X1    g14326(.A1(new_n14518_), .A2(new_n14198_), .Z(new_n14519_));
  OAI21_X1   g14327(.A1(new_n14158_), .A2(new_n14160_), .B(new_n14163_), .ZN(new_n14520_));
  NOR2_X1    g14328(.A1(new_n14430_), .A2(new_n14520_), .ZN(new_n14521_));
  XOR2_X1    g14329(.A1(new_n14521_), .A2(new_n14024_), .Z(new_n14522_));
  INV_X1     g14330(.I(new_n14522_), .ZN(new_n14523_));
  NAND3_X1   g14331(.A1(\asqrt[11] ), .A2(new_n14177_), .A3(new_n14159_), .ZN(new_n14524_));
  XOR2_X1    g14332(.A1(new_n14524_), .A2(new_n14028_), .Z(new_n14525_));
  INV_X1     g14333(.I(new_n14525_), .ZN(new_n14526_));
  OAI21_X1   g14334(.A1(new_n14172_), .A2(new_n14173_), .B(new_n14176_), .ZN(new_n14527_));
  NOR2_X1    g14335(.A1(new_n14430_), .A2(new_n14527_), .ZN(new_n14528_));
  XOR2_X1    g14336(.A1(new_n14528_), .A2(new_n14030_), .Z(new_n14529_));
  NAND3_X1   g14337(.A1(\asqrt[11] ), .A2(new_n14136_), .A3(new_n14155_), .ZN(new_n14530_));
  XOR2_X1    g14338(.A1(new_n14530_), .A2(new_n14170_), .Z(new_n14531_));
  OAI21_X1   g14339(.A1(new_n14130_), .A2(new_n14132_), .B(new_n14135_), .ZN(new_n14532_));
  NOR2_X1    g14340(.A1(new_n14430_), .A2(new_n14532_), .ZN(new_n14533_));
  XOR2_X1    g14341(.A1(new_n14533_), .A2(new_n14036_), .Z(new_n14534_));
  INV_X1     g14342(.I(new_n14534_), .ZN(new_n14535_));
  NAND3_X1   g14343(.A1(\asqrt[11] ), .A2(new_n14149_), .A3(new_n14131_), .ZN(new_n14536_));
  XOR2_X1    g14344(.A1(new_n14536_), .A2(new_n14040_), .Z(new_n14537_));
  INV_X1     g14345(.I(new_n14537_), .ZN(new_n14538_));
  OAI21_X1   g14346(.A1(new_n14144_), .A2(new_n14145_), .B(new_n14148_), .ZN(new_n14539_));
  NOR2_X1    g14347(.A1(new_n14430_), .A2(new_n14539_), .ZN(new_n14540_));
  XOR2_X1    g14348(.A1(new_n14540_), .A2(new_n14042_), .Z(new_n14541_));
  NAND3_X1   g14349(.A1(\asqrt[11] ), .A2(new_n14095_), .A3(new_n14127_), .ZN(new_n14542_));
  XOR2_X1    g14350(.A1(new_n14542_), .A2(new_n14142_), .Z(new_n14543_));
  OAI21_X1   g14351(.A1(new_n14089_), .A2(new_n14091_), .B(new_n14094_), .ZN(new_n14544_));
  NOR2_X1    g14352(.A1(new_n14430_), .A2(new_n14544_), .ZN(new_n14545_));
  XOR2_X1    g14353(.A1(new_n14545_), .A2(new_n14048_), .Z(new_n14546_));
  INV_X1     g14354(.I(new_n14546_), .ZN(new_n14547_));
  NAND3_X1   g14355(.A1(\asqrt[11] ), .A2(new_n14121_), .A3(new_n14090_), .ZN(new_n14548_));
  XOR2_X1    g14356(.A1(new_n14548_), .A2(new_n14052_), .Z(new_n14549_));
  INV_X1     g14357(.I(new_n14549_), .ZN(new_n14550_));
  AOI21_X1   g14358(.A1(new_n14083_), .A2(new_n14084_), .B(new_n14087_), .ZN(new_n14551_));
  NAND2_X1   g14359(.A1(\asqrt[11] ), .A2(new_n14551_), .ZN(new_n14552_));
  XOR2_X1    g14360(.A1(new_n14552_), .A2(new_n14055_), .Z(new_n14553_));
  NOR2_X1    g14361(.A1(new_n14082_), .A2(\asqrt[16] ), .ZN(new_n14554_));
  NOR3_X1    g14362(.A1(new_n14430_), .A2(new_n14554_), .A3(new_n14119_), .ZN(new_n14555_));
  XOR2_X1    g14363(.A1(new_n14555_), .A2(new_n14058_), .Z(new_n14556_));
  NOR3_X1    g14364(.A1(new_n14430_), .A2(new_n14077_), .A3(new_n14114_), .ZN(new_n14557_));
  XOR2_X1    g14365(.A1(new_n14557_), .A2(new_n14079_), .Z(new_n14558_));
  INV_X1     g14366(.I(new_n14558_), .ZN(new_n14559_));
  NOR2_X1    g14367(.A1(new_n14110_), .A2(\asqrt[14] ), .ZN(new_n14560_));
  NOR3_X1    g14368(.A1(new_n14430_), .A2(new_n14560_), .A3(new_n14076_), .ZN(new_n14561_));
  XOR2_X1    g14369(.A1(new_n14561_), .A2(new_n14104_), .Z(new_n14562_));
  INV_X1     g14370(.I(new_n14562_), .ZN(new_n14563_));
  NAND3_X1   g14371(.A1(\asqrt[11] ), .A2(new_n14066_), .A3(new_n14067_), .ZN(new_n14564_));
  NAND4_X1   g14372(.A1(new_n14441_), .A2(\asqrt[12] ), .A3(new_n14443_), .A4(new_n14435_), .ZN(new_n14565_));
  AOI21_X1   g14373(.A1(new_n14564_), .A2(new_n14565_), .B(\a[24] ), .ZN(new_n14566_));
  NOR3_X1    g14374(.A1(new_n14430_), .A2(\a[22] ), .A3(\a[23] ), .ZN(new_n14567_));
  INV_X1     g14375(.I(new_n14565_), .ZN(new_n14568_));
  NOR3_X1    g14376(.A1(new_n14567_), .A2(new_n13511_), .A3(new_n14568_), .ZN(new_n14569_));
  NOR2_X1    g14377(.A1(new_n14569_), .A2(new_n14566_), .ZN(new_n14570_));
  INV_X1     g14378(.I(\a[20] ), .ZN(new_n14571_));
  INV_X1     g14379(.I(\a[21] ), .ZN(new_n14572_));
  NAND3_X1   g14380(.A1(new_n14571_), .A2(new_n14572_), .A3(new_n14066_), .ZN(new_n14573_));
  OAI21_X1   g14381(.A1(new_n14430_), .A2(new_n14066_), .B(new_n14573_), .ZN(new_n14574_));
  NAND2_X1   g14382(.A1(new_n14574_), .A2(\asqrt[12] ), .ZN(new_n14575_));
  OAI21_X1   g14383(.A1(new_n14430_), .A2(\a[22] ), .B(\a[23] ), .ZN(new_n14576_));
  NAND2_X1   g14384(.A1(new_n14576_), .A2(new_n14564_), .ZN(new_n14577_));
  NOR2_X1    g14385(.A1(new_n14574_), .A2(\asqrt[12] ), .ZN(new_n14578_));
  OAI21_X1   g14386(.A1(new_n14577_), .A2(new_n14578_), .B(new_n14575_), .ZN(new_n14579_));
  OAI21_X1   g14387(.A1(new_n14579_), .A2(\asqrt[13] ), .B(new_n14570_), .ZN(new_n14580_));
  NAND2_X1   g14388(.A1(new_n14579_), .A2(\asqrt[13] ), .ZN(new_n14581_));
  NAND3_X1   g14389(.A1(new_n14580_), .A2(new_n12889_), .A3(new_n14581_), .ZN(new_n14582_));
  NOR3_X1    g14390(.A1(new_n14430_), .A2(new_n14070_), .A3(new_n14109_), .ZN(new_n14583_));
  XOR2_X1    g14391(.A1(new_n14583_), .A2(new_n14072_), .Z(new_n14584_));
  NAND2_X1   g14392(.A1(new_n14582_), .A2(new_n14584_), .ZN(new_n14585_));
  NAND2_X1   g14393(.A1(new_n14580_), .A2(new_n14581_), .ZN(new_n14586_));
  AOI21_X1   g14394(.A1(new_n14586_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n14587_));
  AOI21_X1   g14395(.A1(new_n14587_), .A2(new_n14585_), .B(new_n14563_), .ZN(new_n14588_));
  OAI21_X1   g14396(.A1(new_n14567_), .A2(new_n14568_), .B(new_n13511_), .ZN(new_n14589_));
  NAND3_X1   g14397(.A1(new_n14564_), .A2(\a[24] ), .A3(new_n14565_), .ZN(new_n14590_));
  NAND2_X1   g14398(.A1(new_n14589_), .A2(new_n14590_), .ZN(new_n14591_));
  NAND2_X1   g14399(.A1(\asqrt[11] ), .A2(\a[22] ), .ZN(new_n14592_));
  AOI21_X1   g14400(.A1(new_n14592_), .A2(new_n14573_), .B(new_n13917_), .ZN(new_n14593_));
  AOI21_X1   g14401(.A1(\asqrt[11] ), .A2(new_n14066_), .B(new_n14067_), .ZN(new_n14594_));
  NOR2_X1    g14402(.A1(new_n14567_), .A2(new_n14594_), .ZN(new_n14595_));
  NAND3_X1   g14403(.A1(new_n14592_), .A2(new_n13917_), .A3(new_n14573_), .ZN(new_n14596_));
  AOI21_X1   g14404(.A1(new_n14595_), .A2(new_n14596_), .B(new_n14593_), .ZN(new_n14597_));
  AOI21_X1   g14405(.A1(new_n14597_), .A2(new_n13382_), .B(new_n14591_), .ZN(new_n14598_));
  NOR2_X1    g14406(.A1(new_n14597_), .A2(new_n13382_), .ZN(new_n14599_));
  OAI21_X1   g14407(.A1(new_n14598_), .A2(new_n14599_), .B(\asqrt[14] ), .ZN(new_n14600_));
  AOI21_X1   g14408(.A1(new_n14585_), .A2(new_n14600_), .B(new_n12374_), .ZN(new_n14601_));
  NOR2_X1    g14409(.A1(new_n14588_), .A2(new_n14601_), .ZN(new_n14602_));
  AOI21_X1   g14410(.A1(new_n14602_), .A2(new_n11901_), .B(new_n14559_), .ZN(new_n14603_));
  OAI21_X1   g14411(.A1(new_n14588_), .A2(new_n14601_), .B(\asqrt[16] ), .ZN(new_n14604_));
  NAND2_X1   g14412(.A1(new_n14604_), .A2(new_n11406_), .ZN(new_n14605_));
  OAI21_X1   g14413(.A1(new_n14603_), .A2(new_n14605_), .B(new_n14556_), .ZN(new_n14606_));
  INV_X1     g14414(.I(new_n14604_), .ZN(new_n14607_));
  OAI21_X1   g14415(.A1(new_n14603_), .A2(new_n14607_), .B(\asqrt[17] ), .ZN(new_n14608_));
  NAND3_X1   g14416(.A1(new_n14606_), .A2(new_n14608_), .A3(new_n10953_), .ZN(new_n14609_));
  NAND2_X1   g14417(.A1(new_n14609_), .A2(new_n14553_), .ZN(new_n14610_));
  NAND2_X1   g14418(.A1(new_n14606_), .A2(new_n14608_), .ZN(new_n14611_));
  AOI21_X1   g14419(.A1(new_n14611_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n14612_));
  AOI21_X1   g14420(.A1(new_n14612_), .A2(new_n14610_), .B(new_n14550_), .ZN(new_n14613_));
  INV_X1     g14421(.I(new_n14556_), .ZN(new_n14614_));
  NOR2_X1    g14422(.A1(new_n14598_), .A2(new_n14599_), .ZN(new_n14615_));
  INV_X1     g14423(.I(new_n14584_), .ZN(new_n14616_));
  AOI21_X1   g14424(.A1(new_n14615_), .A2(new_n12889_), .B(new_n14616_), .ZN(new_n14617_));
  NAND2_X1   g14425(.A1(new_n14600_), .A2(new_n12374_), .ZN(new_n14618_));
  OAI21_X1   g14426(.A1(new_n14617_), .A2(new_n14618_), .B(new_n14562_), .ZN(new_n14619_));
  INV_X1     g14427(.I(new_n14600_), .ZN(new_n14620_));
  OAI21_X1   g14428(.A1(new_n14617_), .A2(new_n14620_), .B(\asqrt[15] ), .ZN(new_n14621_));
  NAND3_X1   g14429(.A1(new_n14619_), .A2(new_n14621_), .A3(new_n11901_), .ZN(new_n14622_));
  NAND2_X1   g14430(.A1(new_n14622_), .A2(new_n14558_), .ZN(new_n14623_));
  NAND2_X1   g14431(.A1(new_n14619_), .A2(new_n14621_), .ZN(new_n14624_));
  AOI21_X1   g14432(.A1(new_n14624_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n14625_));
  AOI21_X1   g14433(.A1(new_n14625_), .A2(new_n14623_), .B(new_n14614_), .ZN(new_n14626_));
  AOI21_X1   g14434(.A1(new_n14623_), .A2(new_n14604_), .B(new_n11406_), .ZN(new_n14627_));
  OAI21_X1   g14435(.A1(new_n14626_), .A2(new_n14627_), .B(\asqrt[18] ), .ZN(new_n14628_));
  AOI21_X1   g14436(.A1(new_n14610_), .A2(new_n14628_), .B(new_n10478_), .ZN(new_n14629_));
  NOR2_X1    g14437(.A1(new_n14613_), .A2(new_n14629_), .ZN(new_n14630_));
  AOI21_X1   g14438(.A1(new_n14630_), .A2(new_n10045_), .B(new_n14547_), .ZN(new_n14631_));
  OAI21_X1   g14439(.A1(new_n14613_), .A2(new_n14629_), .B(\asqrt[20] ), .ZN(new_n14632_));
  NAND2_X1   g14440(.A1(new_n14632_), .A2(new_n9590_), .ZN(new_n14633_));
  OAI21_X1   g14441(.A1(new_n14631_), .A2(new_n14633_), .B(new_n14543_), .ZN(new_n14634_));
  INV_X1     g14442(.I(new_n14632_), .ZN(new_n14635_));
  OAI21_X1   g14443(.A1(new_n14631_), .A2(new_n14635_), .B(\asqrt[21] ), .ZN(new_n14636_));
  NAND3_X1   g14444(.A1(new_n14634_), .A2(new_n14636_), .A3(new_n9177_), .ZN(new_n14637_));
  NAND2_X1   g14445(.A1(new_n14637_), .A2(new_n14541_), .ZN(new_n14638_));
  NAND2_X1   g14446(.A1(new_n14634_), .A2(new_n14636_), .ZN(new_n14639_));
  AOI21_X1   g14447(.A1(new_n14639_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n14640_));
  AOI21_X1   g14448(.A1(new_n14640_), .A2(new_n14638_), .B(new_n14538_), .ZN(new_n14641_));
  INV_X1     g14449(.I(new_n14543_), .ZN(new_n14642_));
  INV_X1     g14450(.I(new_n14553_), .ZN(new_n14643_));
  NOR2_X1    g14451(.A1(new_n14626_), .A2(new_n14627_), .ZN(new_n14644_));
  AOI21_X1   g14452(.A1(new_n14644_), .A2(new_n10953_), .B(new_n14643_), .ZN(new_n14645_));
  NAND2_X1   g14453(.A1(new_n14628_), .A2(new_n10478_), .ZN(new_n14646_));
  OAI21_X1   g14454(.A1(new_n14645_), .A2(new_n14646_), .B(new_n14549_), .ZN(new_n14647_));
  INV_X1     g14455(.I(new_n14628_), .ZN(new_n14648_));
  OAI21_X1   g14456(.A1(new_n14645_), .A2(new_n14648_), .B(\asqrt[19] ), .ZN(new_n14649_));
  NAND3_X1   g14457(.A1(new_n14647_), .A2(new_n14649_), .A3(new_n10045_), .ZN(new_n14650_));
  NAND2_X1   g14458(.A1(new_n14650_), .A2(new_n14546_), .ZN(new_n14651_));
  NAND2_X1   g14459(.A1(new_n14647_), .A2(new_n14649_), .ZN(new_n14652_));
  AOI21_X1   g14460(.A1(new_n14652_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n14653_));
  AOI21_X1   g14461(.A1(new_n14653_), .A2(new_n14651_), .B(new_n14642_), .ZN(new_n14654_));
  AOI21_X1   g14462(.A1(new_n14651_), .A2(new_n14632_), .B(new_n9590_), .ZN(new_n14655_));
  OAI21_X1   g14463(.A1(new_n14654_), .A2(new_n14655_), .B(\asqrt[22] ), .ZN(new_n14656_));
  AOI21_X1   g14464(.A1(new_n14638_), .A2(new_n14656_), .B(new_n8742_), .ZN(new_n14657_));
  NOR2_X1    g14465(.A1(new_n14641_), .A2(new_n14657_), .ZN(new_n14658_));
  AOI21_X1   g14466(.A1(new_n14658_), .A2(new_n8349_), .B(new_n14535_), .ZN(new_n14659_));
  OAI21_X1   g14467(.A1(new_n14641_), .A2(new_n14657_), .B(\asqrt[24] ), .ZN(new_n14660_));
  NAND2_X1   g14468(.A1(new_n14660_), .A2(new_n7934_), .ZN(new_n14661_));
  OAI21_X1   g14469(.A1(new_n14659_), .A2(new_n14661_), .B(new_n14531_), .ZN(new_n14662_));
  INV_X1     g14470(.I(new_n14660_), .ZN(new_n14663_));
  OAI21_X1   g14471(.A1(new_n14659_), .A2(new_n14663_), .B(\asqrt[25] ), .ZN(new_n14664_));
  NAND3_X1   g14472(.A1(new_n14662_), .A2(new_n14664_), .A3(new_n7561_), .ZN(new_n14665_));
  NAND2_X1   g14473(.A1(new_n14665_), .A2(new_n14529_), .ZN(new_n14666_));
  NAND2_X1   g14474(.A1(new_n14662_), .A2(new_n14664_), .ZN(new_n14667_));
  AOI21_X1   g14475(.A1(new_n14667_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n14668_));
  AOI21_X1   g14476(.A1(new_n14668_), .A2(new_n14666_), .B(new_n14526_), .ZN(new_n14669_));
  INV_X1     g14477(.I(new_n14531_), .ZN(new_n14670_));
  INV_X1     g14478(.I(new_n14541_), .ZN(new_n14671_));
  NOR2_X1    g14479(.A1(new_n14654_), .A2(new_n14655_), .ZN(new_n14672_));
  AOI21_X1   g14480(.A1(new_n14672_), .A2(new_n9177_), .B(new_n14671_), .ZN(new_n14673_));
  NAND2_X1   g14481(.A1(new_n14656_), .A2(new_n8742_), .ZN(new_n14674_));
  OAI21_X1   g14482(.A1(new_n14673_), .A2(new_n14674_), .B(new_n14537_), .ZN(new_n14675_));
  INV_X1     g14483(.I(new_n14656_), .ZN(new_n14676_));
  OAI21_X1   g14484(.A1(new_n14673_), .A2(new_n14676_), .B(\asqrt[23] ), .ZN(new_n14677_));
  NAND3_X1   g14485(.A1(new_n14675_), .A2(new_n14677_), .A3(new_n8349_), .ZN(new_n14678_));
  NAND2_X1   g14486(.A1(new_n14678_), .A2(new_n14534_), .ZN(new_n14679_));
  NAND2_X1   g14487(.A1(new_n14675_), .A2(new_n14677_), .ZN(new_n14680_));
  AOI21_X1   g14488(.A1(new_n14680_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n14681_));
  AOI21_X1   g14489(.A1(new_n14681_), .A2(new_n14679_), .B(new_n14670_), .ZN(new_n14682_));
  AOI21_X1   g14490(.A1(new_n14679_), .A2(new_n14660_), .B(new_n7934_), .ZN(new_n14683_));
  OAI21_X1   g14491(.A1(new_n14682_), .A2(new_n14683_), .B(\asqrt[26] ), .ZN(new_n14684_));
  AOI21_X1   g14492(.A1(new_n14666_), .A2(new_n14684_), .B(new_n7166_), .ZN(new_n14685_));
  NOR2_X1    g14493(.A1(new_n14669_), .A2(new_n14685_), .ZN(new_n14686_));
  AOI21_X1   g14494(.A1(new_n14686_), .A2(new_n6813_), .B(new_n14523_), .ZN(new_n14687_));
  OAI21_X1   g14495(.A1(new_n14669_), .A2(new_n14685_), .B(\asqrt[28] ), .ZN(new_n14688_));
  NAND2_X1   g14496(.A1(new_n14688_), .A2(new_n6454_), .ZN(new_n14689_));
  OAI21_X1   g14497(.A1(new_n14687_), .A2(new_n14689_), .B(new_n14519_), .ZN(new_n14690_));
  INV_X1     g14498(.I(new_n14688_), .ZN(new_n14691_));
  OAI21_X1   g14499(.A1(new_n14687_), .A2(new_n14691_), .B(\asqrt[29] ), .ZN(new_n14692_));
  NAND3_X1   g14500(.A1(new_n14690_), .A2(new_n14692_), .A3(new_n6106_), .ZN(new_n14693_));
  NAND2_X1   g14501(.A1(new_n14693_), .A2(new_n14517_), .ZN(new_n14694_));
  NAND2_X1   g14502(.A1(new_n14690_), .A2(new_n14692_), .ZN(new_n14695_));
  AOI21_X1   g14503(.A1(new_n14695_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n14696_));
  AOI21_X1   g14504(.A1(new_n14696_), .A2(new_n14694_), .B(new_n14514_), .ZN(new_n14697_));
  INV_X1     g14505(.I(new_n14519_), .ZN(new_n14698_));
  INV_X1     g14506(.I(new_n14529_), .ZN(new_n14699_));
  NOR2_X1    g14507(.A1(new_n14682_), .A2(new_n14683_), .ZN(new_n14700_));
  AOI21_X1   g14508(.A1(new_n14700_), .A2(new_n7561_), .B(new_n14699_), .ZN(new_n14701_));
  NAND2_X1   g14509(.A1(new_n14684_), .A2(new_n7166_), .ZN(new_n14702_));
  OAI21_X1   g14510(.A1(new_n14701_), .A2(new_n14702_), .B(new_n14525_), .ZN(new_n14703_));
  INV_X1     g14511(.I(new_n14684_), .ZN(new_n14704_));
  OAI21_X1   g14512(.A1(new_n14701_), .A2(new_n14704_), .B(\asqrt[27] ), .ZN(new_n14705_));
  NAND3_X1   g14513(.A1(new_n14703_), .A2(new_n14705_), .A3(new_n6813_), .ZN(new_n14706_));
  NAND2_X1   g14514(.A1(new_n14706_), .A2(new_n14522_), .ZN(new_n14707_));
  NAND2_X1   g14515(.A1(new_n14703_), .A2(new_n14705_), .ZN(new_n14708_));
  AOI21_X1   g14516(.A1(new_n14708_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n14709_));
  AOI21_X1   g14517(.A1(new_n14709_), .A2(new_n14707_), .B(new_n14698_), .ZN(new_n14710_));
  AOI21_X1   g14518(.A1(new_n14707_), .A2(new_n14688_), .B(new_n6454_), .ZN(new_n14711_));
  OAI21_X1   g14519(.A1(new_n14710_), .A2(new_n14711_), .B(\asqrt[30] ), .ZN(new_n14712_));
  AOI21_X1   g14520(.A1(new_n14694_), .A2(new_n14712_), .B(new_n5750_), .ZN(new_n14713_));
  NOR2_X1    g14521(.A1(new_n14697_), .A2(new_n14713_), .ZN(new_n14714_));
  AOI21_X1   g14522(.A1(new_n14714_), .A2(new_n5435_), .B(new_n14511_), .ZN(new_n14715_));
  OAI21_X1   g14523(.A1(new_n14697_), .A2(new_n14713_), .B(\asqrt[32] ), .ZN(new_n14716_));
  NAND2_X1   g14524(.A1(new_n14716_), .A2(new_n5110_), .ZN(new_n14717_));
  OAI21_X1   g14525(.A1(new_n14715_), .A2(new_n14717_), .B(new_n14507_), .ZN(new_n14718_));
  INV_X1     g14526(.I(new_n14716_), .ZN(new_n14719_));
  OAI21_X1   g14527(.A1(new_n14715_), .A2(new_n14719_), .B(\asqrt[33] ), .ZN(new_n14720_));
  NAND3_X1   g14528(.A1(new_n14718_), .A2(new_n14720_), .A3(new_n4810_), .ZN(new_n14721_));
  NAND2_X1   g14529(.A1(new_n14721_), .A2(new_n14505_), .ZN(new_n14722_));
  NAND2_X1   g14530(.A1(new_n14718_), .A2(new_n14720_), .ZN(new_n14723_));
  AOI21_X1   g14531(.A1(new_n14723_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n14724_));
  AOI21_X1   g14532(.A1(new_n14724_), .A2(new_n14722_), .B(new_n14502_), .ZN(new_n14725_));
  INV_X1     g14533(.I(new_n14507_), .ZN(new_n14726_));
  INV_X1     g14534(.I(new_n14517_), .ZN(new_n14727_));
  NOR2_X1    g14535(.A1(new_n14710_), .A2(new_n14711_), .ZN(new_n14728_));
  AOI21_X1   g14536(.A1(new_n14728_), .A2(new_n6106_), .B(new_n14727_), .ZN(new_n14729_));
  NAND2_X1   g14537(.A1(new_n14712_), .A2(new_n5750_), .ZN(new_n14730_));
  OAI21_X1   g14538(.A1(new_n14729_), .A2(new_n14730_), .B(new_n14513_), .ZN(new_n14731_));
  INV_X1     g14539(.I(new_n14712_), .ZN(new_n14732_));
  OAI21_X1   g14540(.A1(new_n14729_), .A2(new_n14732_), .B(\asqrt[31] ), .ZN(new_n14733_));
  NAND3_X1   g14541(.A1(new_n14731_), .A2(new_n14733_), .A3(new_n5435_), .ZN(new_n14734_));
  NAND2_X1   g14542(.A1(new_n14734_), .A2(new_n14510_), .ZN(new_n14735_));
  NAND2_X1   g14543(.A1(new_n14731_), .A2(new_n14733_), .ZN(new_n14736_));
  AOI21_X1   g14544(.A1(new_n14736_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n14737_));
  AOI21_X1   g14545(.A1(new_n14737_), .A2(new_n14735_), .B(new_n14726_), .ZN(new_n14738_));
  AOI21_X1   g14546(.A1(new_n14735_), .A2(new_n14716_), .B(new_n5110_), .ZN(new_n14739_));
  OAI21_X1   g14547(.A1(new_n14738_), .A2(new_n14739_), .B(\asqrt[34] ), .ZN(new_n14740_));
  AOI21_X1   g14548(.A1(new_n14722_), .A2(new_n14740_), .B(new_n4510_), .ZN(new_n14741_));
  NOR2_X1    g14549(.A1(new_n14725_), .A2(new_n14741_), .ZN(new_n14742_));
  AOI21_X1   g14550(.A1(new_n14742_), .A2(new_n4224_), .B(new_n14499_), .ZN(new_n14743_));
  OAI21_X1   g14551(.A1(new_n14725_), .A2(new_n14741_), .B(\asqrt[36] ), .ZN(new_n14744_));
  NAND2_X1   g14552(.A1(new_n14744_), .A2(new_n3928_), .ZN(new_n14745_));
  OAI21_X1   g14553(.A1(new_n14743_), .A2(new_n14745_), .B(new_n14495_), .ZN(new_n14746_));
  INV_X1     g14554(.I(new_n14744_), .ZN(new_n14747_));
  OAI21_X1   g14555(.A1(new_n14743_), .A2(new_n14747_), .B(\asqrt[37] ), .ZN(new_n14748_));
  NAND3_X1   g14556(.A1(new_n14746_), .A2(new_n14748_), .A3(new_n3675_), .ZN(new_n14749_));
  NAND2_X1   g14557(.A1(new_n14749_), .A2(new_n14493_), .ZN(new_n14750_));
  NAND2_X1   g14558(.A1(new_n14746_), .A2(new_n14748_), .ZN(new_n14751_));
  AOI21_X1   g14559(.A1(new_n14751_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n14752_));
  AOI21_X1   g14560(.A1(new_n14752_), .A2(new_n14750_), .B(new_n14490_), .ZN(new_n14753_));
  INV_X1     g14561(.I(new_n14495_), .ZN(new_n14754_));
  INV_X1     g14562(.I(new_n14505_), .ZN(new_n14755_));
  NOR2_X1    g14563(.A1(new_n14738_), .A2(new_n14739_), .ZN(new_n14756_));
  AOI21_X1   g14564(.A1(new_n14756_), .A2(new_n4810_), .B(new_n14755_), .ZN(new_n14757_));
  NAND2_X1   g14565(.A1(new_n14740_), .A2(new_n4510_), .ZN(new_n14758_));
  OAI21_X1   g14566(.A1(new_n14757_), .A2(new_n14758_), .B(new_n14501_), .ZN(new_n14759_));
  INV_X1     g14567(.I(new_n14740_), .ZN(new_n14760_));
  OAI21_X1   g14568(.A1(new_n14757_), .A2(new_n14760_), .B(\asqrt[35] ), .ZN(new_n14761_));
  NAND3_X1   g14569(.A1(new_n14759_), .A2(new_n14761_), .A3(new_n4224_), .ZN(new_n14762_));
  NAND2_X1   g14570(.A1(new_n14762_), .A2(new_n14498_), .ZN(new_n14763_));
  NAND2_X1   g14571(.A1(new_n14759_), .A2(new_n14761_), .ZN(new_n14764_));
  AOI21_X1   g14572(.A1(new_n14764_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n14765_));
  AOI21_X1   g14573(.A1(new_n14765_), .A2(new_n14763_), .B(new_n14754_), .ZN(new_n14766_));
  AOI21_X1   g14574(.A1(new_n14763_), .A2(new_n14744_), .B(new_n3928_), .ZN(new_n14767_));
  OAI21_X1   g14575(.A1(new_n14766_), .A2(new_n14767_), .B(\asqrt[38] ), .ZN(new_n14768_));
  AOI21_X1   g14576(.A1(new_n14750_), .A2(new_n14768_), .B(new_n3400_), .ZN(new_n14769_));
  NOR2_X1    g14577(.A1(new_n14753_), .A2(new_n14769_), .ZN(new_n14770_));
  AOI21_X1   g14578(.A1(new_n14770_), .A2(new_n3167_), .B(new_n14487_), .ZN(new_n14771_));
  OAI21_X1   g14579(.A1(new_n14753_), .A2(new_n14769_), .B(\asqrt[40] ), .ZN(new_n14772_));
  NAND2_X1   g14580(.A1(new_n14772_), .A2(new_n2912_), .ZN(new_n14773_));
  OAI21_X1   g14581(.A1(new_n14771_), .A2(new_n14773_), .B(new_n14483_), .ZN(new_n14774_));
  INV_X1     g14582(.I(new_n14772_), .ZN(new_n14775_));
  OAI21_X1   g14583(.A1(new_n14771_), .A2(new_n14775_), .B(\asqrt[41] ), .ZN(new_n14776_));
  NAND3_X1   g14584(.A1(new_n14774_), .A2(new_n14776_), .A3(new_n2699_), .ZN(new_n14777_));
  NAND2_X1   g14585(.A1(new_n14777_), .A2(new_n14481_), .ZN(new_n14778_));
  NAND2_X1   g14586(.A1(new_n14774_), .A2(new_n14776_), .ZN(new_n14779_));
  AOI21_X1   g14587(.A1(new_n14779_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n14780_));
  AOI21_X1   g14588(.A1(new_n14780_), .A2(new_n14778_), .B(new_n14478_), .ZN(new_n14781_));
  INV_X1     g14589(.I(new_n14483_), .ZN(new_n14782_));
  INV_X1     g14590(.I(new_n14493_), .ZN(new_n14783_));
  NOR2_X1    g14591(.A1(new_n14766_), .A2(new_n14767_), .ZN(new_n14784_));
  AOI21_X1   g14592(.A1(new_n14784_), .A2(new_n3675_), .B(new_n14783_), .ZN(new_n14785_));
  NAND2_X1   g14593(.A1(new_n14768_), .A2(new_n3400_), .ZN(new_n14786_));
  OAI21_X1   g14594(.A1(new_n14785_), .A2(new_n14786_), .B(new_n14489_), .ZN(new_n14787_));
  INV_X1     g14595(.I(new_n14768_), .ZN(new_n14788_));
  OAI21_X1   g14596(.A1(new_n14785_), .A2(new_n14788_), .B(\asqrt[39] ), .ZN(new_n14789_));
  NAND3_X1   g14597(.A1(new_n14787_), .A2(new_n14789_), .A3(new_n3167_), .ZN(new_n14790_));
  NAND2_X1   g14598(.A1(new_n14790_), .A2(new_n14486_), .ZN(new_n14791_));
  NAND2_X1   g14599(.A1(new_n14787_), .A2(new_n14789_), .ZN(new_n14792_));
  AOI21_X1   g14600(.A1(new_n14792_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n14793_));
  AOI21_X1   g14601(.A1(new_n14793_), .A2(new_n14791_), .B(new_n14782_), .ZN(new_n14794_));
  AOI21_X1   g14602(.A1(new_n14791_), .A2(new_n14772_), .B(new_n2912_), .ZN(new_n14795_));
  OAI21_X1   g14603(.A1(new_n14794_), .A2(new_n14795_), .B(\asqrt[42] ), .ZN(new_n14796_));
  AOI21_X1   g14604(.A1(new_n14778_), .A2(new_n14796_), .B(new_n2464_), .ZN(new_n14797_));
  NOR2_X1    g14605(.A1(new_n14781_), .A2(new_n14797_), .ZN(new_n14798_));
  AOI21_X1   g14606(.A1(new_n14798_), .A2(new_n2271_), .B(new_n14475_), .ZN(new_n14799_));
  OAI21_X1   g14607(.A1(new_n14781_), .A2(new_n14797_), .B(\asqrt[44] ), .ZN(new_n14800_));
  NAND2_X1   g14608(.A1(new_n14800_), .A2(new_n2072_), .ZN(new_n14801_));
  OAI21_X1   g14609(.A1(new_n14799_), .A2(new_n14801_), .B(new_n14471_), .ZN(new_n14802_));
  INV_X1     g14610(.I(new_n14800_), .ZN(new_n14803_));
  OAI21_X1   g14611(.A1(new_n14799_), .A2(new_n14803_), .B(\asqrt[45] ), .ZN(new_n14804_));
  NAND3_X1   g14612(.A1(new_n14802_), .A2(new_n14804_), .A3(new_n1884_), .ZN(new_n14805_));
  NAND2_X1   g14613(.A1(new_n14805_), .A2(new_n14469_), .ZN(new_n14806_));
  NAND2_X1   g14614(.A1(new_n14802_), .A2(new_n14804_), .ZN(new_n14807_));
  AOI21_X1   g14615(.A1(new_n14807_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n14808_));
  AOI21_X1   g14616(.A1(new_n14808_), .A2(new_n14806_), .B(new_n14466_), .ZN(new_n14809_));
  INV_X1     g14617(.I(new_n14471_), .ZN(new_n14810_));
  INV_X1     g14618(.I(new_n14481_), .ZN(new_n14811_));
  NOR2_X1    g14619(.A1(new_n14794_), .A2(new_n14795_), .ZN(new_n14812_));
  AOI21_X1   g14620(.A1(new_n14812_), .A2(new_n2699_), .B(new_n14811_), .ZN(new_n14813_));
  NAND2_X1   g14621(.A1(new_n14796_), .A2(new_n2464_), .ZN(new_n14814_));
  OAI21_X1   g14622(.A1(new_n14813_), .A2(new_n14814_), .B(new_n14477_), .ZN(new_n14815_));
  INV_X1     g14623(.I(new_n14796_), .ZN(new_n14816_));
  OAI21_X1   g14624(.A1(new_n14813_), .A2(new_n14816_), .B(\asqrt[43] ), .ZN(new_n14817_));
  NAND3_X1   g14625(.A1(new_n14815_), .A2(new_n14817_), .A3(new_n2271_), .ZN(new_n14818_));
  NAND2_X1   g14626(.A1(new_n14818_), .A2(new_n14474_), .ZN(new_n14819_));
  NAND2_X1   g14627(.A1(new_n14815_), .A2(new_n14817_), .ZN(new_n14820_));
  AOI21_X1   g14628(.A1(new_n14820_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n14821_));
  AOI21_X1   g14629(.A1(new_n14821_), .A2(new_n14819_), .B(new_n14810_), .ZN(new_n14822_));
  AOI21_X1   g14630(.A1(new_n14819_), .A2(new_n14800_), .B(new_n2072_), .ZN(new_n14823_));
  OAI21_X1   g14631(.A1(new_n14822_), .A2(new_n14823_), .B(\asqrt[46] ), .ZN(new_n14824_));
  AOI21_X1   g14632(.A1(new_n14806_), .A2(new_n14824_), .B(new_n1688_), .ZN(new_n14825_));
  NOR2_X1    g14633(.A1(new_n14809_), .A2(new_n14825_), .ZN(new_n14826_));
  AOI21_X1   g14634(.A1(new_n14826_), .A2(new_n1533_), .B(new_n14463_), .ZN(new_n14827_));
  OAI21_X1   g14635(.A1(new_n14809_), .A2(new_n14825_), .B(\asqrt[48] ), .ZN(new_n14828_));
  NAND2_X1   g14636(.A1(new_n14828_), .A2(new_n1368_), .ZN(new_n14829_));
  OAI21_X1   g14637(.A1(new_n14827_), .A2(new_n14829_), .B(new_n14459_), .ZN(new_n14830_));
  INV_X1     g14638(.I(new_n14828_), .ZN(new_n14831_));
  OAI21_X1   g14639(.A1(new_n14827_), .A2(new_n14831_), .B(\asqrt[49] ), .ZN(new_n14832_));
  NAND3_X1   g14640(.A1(new_n14830_), .A2(new_n14832_), .A3(new_n1228_), .ZN(new_n14833_));
  NAND2_X1   g14641(.A1(new_n14833_), .A2(new_n14457_), .ZN(new_n14834_));
  NAND2_X1   g14642(.A1(new_n14830_), .A2(new_n14832_), .ZN(new_n14835_));
  AOI21_X1   g14643(.A1(new_n14835_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n14836_));
  AOI21_X1   g14644(.A1(new_n14836_), .A2(new_n14834_), .B(new_n14454_), .ZN(new_n14837_));
  INV_X1     g14645(.I(new_n14459_), .ZN(new_n14838_));
  INV_X1     g14646(.I(new_n14469_), .ZN(new_n14839_));
  NOR2_X1    g14647(.A1(new_n14822_), .A2(new_n14823_), .ZN(new_n14840_));
  AOI21_X1   g14648(.A1(new_n14840_), .A2(new_n1884_), .B(new_n14839_), .ZN(new_n14841_));
  NAND2_X1   g14649(.A1(new_n14824_), .A2(new_n1688_), .ZN(new_n14842_));
  OAI21_X1   g14650(.A1(new_n14841_), .A2(new_n14842_), .B(new_n14465_), .ZN(new_n14843_));
  INV_X1     g14651(.I(new_n14824_), .ZN(new_n14844_));
  OAI21_X1   g14652(.A1(new_n14841_), .A2(new_n14844_), .B(\asqrt[47] ), .ZN(new_n14845_));
  NAND3_X1   g14653(.A1(new_n14843_), .A2(new_n14845_), .A3(new_n1533_), .ZN(new_n14846_));
  NAND2_X1   g14654(.A1(new_n14846_), .A2(new_n14462_), .ZN(new_n14847_));
  NAND2_X1   g14655(.A1(new_n14843_), .A2(new_n14845_), .ZN(new_n14848_));
  AOI21_X1   g14656(.A1(new_n14848_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n14849_));
  AOI21_X1   g14657(.A1(new_n14849_), .A2(new_n14847_), .B(new_n14838_), .ZN(new_n14850_));
  AOI21_X1   g14658(.A1(new_n14847_), .A2(new_n14828_), .B(new_n1368_), .ZN(new_n14851_));
  OAI21_X1   g14659(.A1(new_n14850_), .A2(new_n14851_), .B(\asqrt[50] ), .ZN(new_n14852_));
  AOI21_X1   g14660(.A1(new_n14834_), .A2(new_n14852_), .B(new_n1088_), .ZN(new_n14853_));
  NOR2_X1    g14661(.A1(new_n14837_), .A2(new_n14853_), .ZN(new_n14854_));
  AOI21_X1   g14662(.A1(new_n14854_), .A2(new_n962_), .B(new_n14451_), .ZN(new_n14855_));
  OAI21_X1   g14663(.A1(new_n14837_), .A2(new_n14853_), .B(\asqrt[52] ), .ZN(new_n14856_));
  NAND2_X1   g14664(.A1(new_n14856_), .A2(new_n842_), .ZN(new_n14857_));
  OAI21_X1   g14665(.A1(new_n14855_), .A2(new_n14857_), .B(new_n14447_), .ZN(new_n14858_));
  INV_X1     g14666(.I(new_n14856_), .ZN(new_n14859_));
  OAI21_X1   g14667(.A1(new_n14855_), .A2(new_n14859_), .B(\asqrt[53] ), .ZN(new_n14860_));
  NAND3_X1   g14668(.A1(new_n14858_), .A2(new_n14860_), .A3(new_n720_), .ZN(new_n14861_));
  INV_X1     g14669(.I(new_n14447_), .ZN(new_n14862_));
  INV_X1     g14670(.I(new_n14457_), .ZN(new_n14863_));
  NOR2_X1    g14671(.A1(new_n14850_), .A2(new_n14851_), .ZN(new_n14864_));
  AOI21_X1   g14672(.A1(new_n14864_), .A2(new_n1228_), .B(new_n14863_), .ZN(new_n14865_));
  NAND2_X1   g14673(.A1(new_n14852_), .A2(new_n1088_), .ZN(new_n14866_));
  OAI21_X1   g14674(.A1(new_n14865_), .A2(new_n14866_), .B(new_n14453_), .ZN(new_n14867_));
  INV_X1     g14675(.I(new_n14852_), .ZN(new_n14868_));
  OAI21_X1   g14676(.A1(new_n14865_), .A2(new_n14868_), .B(\asqrt[51] ), .ZN(new_n14869_));
  NAND3_X1   g14677(.A1(new_n14867_), .A2(new_n14869_), .A3(new_n962_), .ZN(new_n14870_));
  NAND2_X1   g14678(.A1(new_n14870_), .A2(new_n14450_), .ZN(new_n14871_));
  NAND2_X1   g14679(.A1(new_n14867_), .A2(new_n14869_), .ZN(new_n14872_));
  AOI21_X1   g14680(.A1(new_n14872_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n14873_));
  AOI21_X1   g14681(.A1(new_n14873_), .A2(new_n14871_), .B(new_n14862_), .ZN(new_n14874_));
  AOI21_X1   g14682(.A1(new_n14871_), .A2(new_n14856_), .B(new_n842_), .ZN(new_n14875_));
  OAI21_X1   g14683(.A1(new_n14874_), .A2(new_n14875_), .B(\asqrt[54] ), .ZN(new_n14876_));
  NAND2_X1   g14684(.A1(new_n14427_), .A2(new_n13922_), .ZN(new_n14877_));
  NOR2_X1    g14685(.A1(new_n14430_), .A2(new_n13922_), .ZN(new_n14878_));
  NAND2_X1   g14686(.A1(new_n14878_), .A2(new_n14442_), .ZN(new_n14879_));
  AOI21_X1   g14687(.A1(new_n14879_), .A2(new_n14877_), .B(new_n193_), .ZN(new_n14880_));
  INV_X1     g14688(.I(new_n14880_), .ZN(new_n14881_));
  NAND3_X1   g14689(.A1(\asqrt[11] ), .A2(new_n14412_), .A3(new_n14423_), .ZN(new_n14882_));
  XOR2_X1    g14690(.A1(new_n14882_), .A2(new_n14415_), .Z(new_n14883_));
  AOI21_X1   g14691(.A1(new_n14878_), .A2(new_n14427_), .B(new_n14428_), .ZN(new_n14884_));
  OAI21_X1   g14692(.A1(new_n14382_), .A2(new_n14384_), .B(new_n14387_), .ZN(new_n14885_));
  NOR2_X1    g14693(.A1(new_n14430_), .A2(new_n14885_), .ZN(new_n14886_));
  XOR2_X1    g14694(.A1(new_n14886_), .A2(new_n13930_), .Z(new_n14887_));
  NAND3_X1   g14695(.A1(\asqrt[11] ), .A2(new_n14398_), .A3(new_n14383_), .ZN(new_n14888_));
  XOR2_X1    g14696(.A1(new_n14888_), .A2(new_n13934_), .Z(new_n14889_));
  OAI21_X1   g14697(.A1(new_n14393_), .A2(new_n14394_), .B(new_n14397_), .ZN(new_n14890_));
  NOR2_X1    g14698(.A1(new_n14430_), .A2(new_n14890_), .ZN(new_n14891_));
  XOR2_X1    g14699(.A1(new_n14891_), .A2(new_n13936_), .Z(new_n14892_));
  INV_X1     g14700(.I(new_n14892_), .ZN(new_n14893_));
  NAND3_X1   g14701(.A1(\asqrt[11] ), .A2(new_n14360_), .A3(new_n14379_), .ZN(new_n14894_));
  XOR2_X1    g14702(.A1(new_n14894_), .A2(new_n14391_), .Z(new_n14895_));
  INV_X1     g14703(.I(new_n14895_), .ZN(new_n14896_));
  OAI21_X1   g14704(.A1(new_n14354_), .A2(new_n14356_), .B(new_n14359_), .ZN(new_n14897_));
  NOR2_X1    g14705(.A1(new_n14430_), .A2(new_n14897_), .ZN(new_n14898_));
  XOR2_X1    g14706(.A1(new_n14898_), .A2(new_n13942_), .Z(new_n14899_));
  NAND3_X1   g14707(.A1(\asqrt[11] ), .A2(new_n14373_), .A3(new_n14355_), .ZN(new_n14900_));
  XOR2_X1    g14708(.A1(new_n14900_), .A2(new_n13946_), .Z(new_n14901_));
  NOR2_X1    g14709(.A1(new_n14874_), .A2(new_n14875_), .ZN(new_n14902_));
  AOI21_X1   g14710(.A1(new_n14902_), .A2(new_n720_), .B(new_n14434_), .ZN(new_n14903_));
  NAND2_X1   g14711(.A1(new_n14876_), .A2(new_n630_), .ZN(new_n14904_));
  OAI21_X1   g14712(.A1(new_n14903_), .A2(new_n14904_), .B(new_n14901_), .ZN(new_n14905_));
  INV_X1     g14713(.I(new_n14876_), .ZN(new_n14906_));
  OAI21_X1   g14714(.A1(new_n14903_), .A2(new_n14906_), .B(\asqrt[55] ), .ZN(new_n14907_));
  NAND3_X1   g14715(.A1(new_n14905_), .A2(new_n14907_), .A3(new_n545_), .ZN(new_n14908_));
  NAND2_X1   g14716(.A1(new_n14908_), .A2(new_n14899_), .ZN(new_n14909_));
  NAND2_X1   g14717(.A1(new_n14905_), .A2(new_n14907_), .ZN(new_n14910_));
  AOI21_X1   g14718(.A1(new_n14910_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n14911_));
  AOI21_X1   g14719(.A1(new_n14911_), .A2(new_n14909_), .B(new_n14896_), .ZN(new_n14912_));
  INV_X1     g14720(.I(new_n14901_), .ZN(new_n14913_));
  NAND2_X1   g14721(.A1(new_n14861_), .A2(new_n14433_), .ZN(new_n14914_));
  NAND2_X1   g14722(.A1(new_n14858_), .A2(new_n14860_), .ZN(new_n14915_));
  AOI21_X1   g14723(.A1(new_n14915_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n14916_));
  AOI21_X1   g14724(.A1(new_n14916_), .A2(new_n14914_), .B(new_n14913_), .ZN(new_n14917_));
  AOI21_X1   g14725(.A1(new_n14914_), .A2(new_n14876_), .B(new_n630_), .ZN(new_n14918_));
  OAI21_X1   g14726(.A1(new_n14917_), .A2(new_n14918_), .B(\asqrt[56] ), .ZN(new_n14919_));
  AOI21_X1   g14727(.A1(new_n14909_), .A2(new_n14919_), .B(new_n450_), .ZN(new_n14920_));
  NOR2_X1    g14728(.A1(new_n14912_), .A2(new_n14920_), .ZN(new_n14921_));
  AOI21_X1   g14729(.A1(new_n14921_), .A2(new_n403_), .B(new_n14893_), .ZN(new_n14922_));
  OAI21_X1   g14730(.A1(new_n14912_), .A2(new_n14920_), .B(\asqrt[58] ), .ZN(new_n14923_));
  NAND2_X1   g14731(.A1(new_n14923_), .A2(new_n339_), .ZN(new_n14924_));
  OAI21_X1   g14732(.A1(new_n14922_), .A2(new_n14924_), .B(new_n14889_), .ZN(new_n14925_));
  INV_X1     g14733(.I(new_n14923_), .ZN(new_n14926_));
  OAI21_X1   g14734(.A1(new_n14922_), .A2(new_n14926_), .B(\asqrt[59] ), .ZN(new_n14927_));
  NAND3_X1   g14735(.A1(new_n14925_), .A2(new_n14927_), .A3(new_n288_), .ZN(new_n14928_));
  NAND2_X1   g14736(.A1(new_n14928_), .A2(new_n14887_), .ZN(new_n14929_));
  INV_X1     g14737(.I(new_n14889_), .ZN(new_n14930_));
  INV_X1     g14738(.I(new_n14899_), .ZN(new_n14931_));
  NOR2_X1    g14739(.A1(new_n14917_), .A2(new_n14918_), .ZN(new_n14932_));
  AOI21_X1   g14740(.A1(new_n14932_), .A2(new_n545_), .B(new_n14931_), .ZN(new_n14933_));
  NAND2_X1   g14741(.A1(new_n14919_), .A2(new_n450_), .ZN(new_n14934_));
  OAI21_X1   g14742(.A1(new_n14933_), .A2(new_n14934_), .B(new_n14895_), .ZN(new_n14935_));
  INV_X1     g14743(.I(new_n14919_), .ZN(new_n14936_));
  OAI21_X1   g14744(.A1(new_n14933_), .A2(new_n14936_), .B(\asqrt[57] ), .ZN(new_n14937_));
  NAND3_X1   g14745(.A1(new_n14935_), .A2(new_n14937_), .A3(new_n403_), .ZN(new_n14938_));
  NAND2_X1   g14746(.A1(new_n14938_), .A2(new_n14892_), .ZN(new_n14939_));
  NAND2_X1   g14747(.A1(new_n14935_), .A2(new_n14937_), .ZN(new_n14940_));
  AOI21_X1   g14748(.A1(new_n14940_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n14941_));
  AOI21_X1   g14749(.A1(new_n14941_), .A2(new_n14939_), .B(new_n14930_), .ZN(new_n14942_));
  AOI21_X1   g14750(.A1(new_n14939_), .A2(new_n14923_), .B(new_n339_), .ZN(new_n14943_));
  OAI21_X1   g14751(.A1(new_n14942_), .A2(new_n14943_), .B(\asqrt[60] ), .ZN(new_n14944_));
  AOI21_X1   g14752(.A1(new_n14929_), .A2(new_n14944_), .B(new_n242_), .ZN(new_n14945_));
  NAND3_X1   g14753(.A1(\asqrt[11] ), .A2(new_n14388_), .A3(new_n14404_), .ZN(new_n14946_));
  XOR2_X1    g14754(.A1(new_n14946_), .A2(new_n14416_), .Z(new_n14947_));
  INV_X1     g14755(.I(new_n14947_), .ZN(new_n14948_));
  NAND2_X1   g14756(.A1(new_n14925_), .A2(new_n14927_), .ZN(new_n14949_));
  AOI21_X1   g14757(.A1(new_n14949_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n14950_));
  AOI21_X1   g14758(.A1(new_n14950_), .A2(new_n14929_), .B(new_n14948_), .ZN(new_n14951_));
  OAI21_X1   g14759(.A1(new_n14951_), .A2(new_n14945_), .B(\asqrt[62] ), .ZN(new_n14952_));
  INV_X1     g14760(.I(new_n14952_), .ZN(new_n14953_));
  NOR2_X1    g14761(.A1(new_n14951_), .A2(new_n14945_), .ZN(new_n14954_));
  AOI21_X1   g14762(.A1(new_n14389_), .A2(new_n14410_), .B(new_n14405_), .ZN(new_n14955_));
  NAND2_X1   g14763(.A1(\asqrt[11] ), .A2(new_n14955_), .ZN(new_n14956_));
  XOR2_X1    g14764(.A1(new_n14956_), .A2(new_n14408_), .Z(new_n14957_));
  INV_X1     g14765(.I(new_n14957_), .ZN(new_n14958_));
  AOI21_X1   g14766(.A1(new_n14954_), .A2(new_n234_), .B(new_n14958_), .ZN(new_n14959_));
  OAI21_X1   g14767(.A1(new_n14959_), .A2(new_n14953_), .B(new_n14884_), .ZN(new_n14960_));
  OAI21_X1   g14768(.A1(new_n14960_), .A2(new_n14883_), .B(new_n193_), .ZN(new_n14961_));
  NOR2_X1    g14769(.A1(new_n14959_), .A2(new_n14953_), .ZN(new_n14962_));
  NAND2_X1   g14770(.A1(new_n14962_), .A2(new_n14883_), .ZN(new_n14963_));
  NOR2_X1    g14771(.A1(\asqrt[11] ), .A2(new_n13923_), .ZN(new_n14964_));
  INV_X1     g14772(.I(new_n14964_), .ZN(new_n14965_));
  NAND4_X1   g14773(.A1(new_n14961_), .A2(new_n14881_), .A3(new_n14963_), .A4(new_n14965_), .ZN(\asqrt[10] ));
  NAND3_X1   g14774(.A1(\asqrt[10] ), .A2(new_n14861_), .A3(new_n14876_), .ZN(new_n14967_));
  XOR2_X1    g14775(.A1(new_n14967_), .A2(new_n14434_), .Z(new_n14968_));
  INV_X1     g14776(.I(new_n14887_), .ZN(new_n14969_));
  NOR2_X1    g14777(.A1(new_n14942_), .A2(new_n14943_), .ZN(new_n14970_));
  AOI21_X1   g14778(.A1(new_n14970_), .A2(new_n288_), .B(new_n14969_), .ZN(new_n14971_));
  INV_X1     g14779(.I(new_n14944_), .ZN(new_n14972_));
  OAI21_X1   g14780(.A1(new_n14971_), .A2(new_n14972_), .B(\asqrt[61] ), .ZN(new_n14973_));
  NAND2_X1   g14781(.A1(new_n14944_), .A2(new_n242_), .ZN(new_n14974_));
  OAI21_X1   g14782(.A1(new_n14971_), .A2(new_n14974_), .B(new_n14947_), .ZN(new_n14975_));
  NAND3_X1   g14783(.A1(new_n14975_), .A2(new_n14973_), .A3(new_n234_), .ZN(new_n14976_));
  NAND2_X1   g14784(.A1(new_n14976_), .A2(new_n14957_), .ZN(new_n14977_));
  NAND2_X1   g14785(.A1(new_n14977_), .A2(new_n14952_), .ZN(new_n14978_));
  NAND2_X1   g14786(.A1(new_n14978_), .A2(new_n14883_), .ZN(new_n14979_));
  INV_X1     g14787(.I(new_n14883_), .ZN(new_n14980_));
  INV_X1     g14788(.I(new_n14884_), .ZN(new_n14981_));
  AOI21_X1   g14789(.A1(new_n14977_), .A2(new_n14952_), .B(new_n14981_), .ZN(new_n14982_));
  AOI21_X1   g14790(.A1(new_n14982_), .A2(new_n14980_), .B(\asqrt[63] ), .ZN(new_n14983_));
  NOR2_X1    g14791(.A1(new_n14978_), .A2(new_n14980_), .ZN(new_n14984_));
  NOR4_X1    g14792(.A1(new_n14983_), .A2(new_n14880_), .A3(new_n14984_), .A4(new_n14964_), .ZN(new_n14985_));
  NOR2_X1    g14793(.A1(new_n14985_), .A2(new_n14883_), .ZN(new_n14986_));
  NAND2_X1   g14794(.A1(new_n14986_), .A2(new_n14962_), .ZN(new_n14987_));
  AOI21_X1   g14795(.A1(new_n14987_), .A2(new_n14979_), .B(new_n193_), .ZN(new_n14988_));
  NAND3_X1   g14796(.A1(\asqrt[10] ), .A2(new_n14952_), .A3(new_n14976_), .ZN(new_n14989_));
  XOR2_X1    g14797(.A1(new_n14989_), .A2(new_n14957_), .Z(new_n14990_));
  INV_X1     g14798(.I(new_n14990_), .ZN(new_n14991_));
  AOI21_X1   g14799(.A1(new_n14986_), .A2(new_n14978_), .B(new_n14984_), .ZN(new_n14992_));
  INV_X1     g14800(.I(new_n14992_), .ZN(new_n14993_));
  OAI21_X1   g14801(.A1(new_n14922_), .A2(new_n14924_), .B(new_n14927_), .ZN(new_n14994_));
  NOR2_X1    g14802(.A1(new_n14985_), .A2(new_n14994_), .ZN(new_n14995_));
  XOR2_X1    g14803(.A1(new_n14995_), .A2(new_n14889_), .Z(new_n14996_));
  NAND3_X1   g14804(.A1(\asqrt[10] ), .A2(new_n14938_), .A3(new_n14923_), .ZN(new_n14997_));
  XOR2_X1    g14805(.A1(new_n14997_), .A2(new_n14893_), .Z(new_n14998_));
  OAI21_X1   g14806(.A1(new_n14933_), .A2(new_n14934_), .B(new_n14937_), .ZN(new_n14999_));
  NOR2_X1    g14807(.A1(new_n14985_), .A2(new_n14999_), .ZN(new_n15000_));
  XOR2_X1    g14808(.A1(new_n15000_), .A2(new_n14895_), .Z(new_n15001_));
  INV_X1     g14809(.I(new_n15001_), .ZN(new_n15002_));
  NAND3_X1   g14810(.A1(\asqrt[10] ), .A2(new_n14908_), .A3(new_n14919_), .ZN(new_n15003_));
  XOR2_X1    g14811(.A1(new_n15003_), .A2(new_n14931_), .Z(new_n15004_));
  INV_X1     g14812(.I(new_n15004_), .ZN(new_n15005_));
  OAI21_X1   g14813(.A1(new_n14903_), .A2(new_n14904_), .B(new_n14907_), .ZN(new_n15006_));
  NOR2_X1    g14814(.A1(new_n14985_), .A2(new_n15006_), .ZN(new_n15007_));
  XOR2_X1    g14815(.A1(new_n15007_), .A2(new_n14901_), .Z(new_n15008_));
  OAI21_X1   g14816(.A1(new_n14855_), .A2(new_n14857_), .B(new_n14860_), .ZN(new_n15009_));
  NOR2_X1    g14817(.A1(new_n14985_), .A2(new_n15009_), .ZN(new_n15010_));
  XOR2_X1    g14818(.A1(new_n15010_), .A2(new_n14447_), .Z(new_n15011_));
  INV_X1     g14819(.I(new_n15011_), .ZN(new_n15012_));
  NAND3_X1   g14820(.A1(\asqrt[10] ), .A2(new_n14870_), .A3(new_n14856_), .ZN(new_n15013_));
  XOR2_X1    g14821(.A1(new_n15013_), .A2(new_n14451_), .Z(new_n15014_));
  INV_X1     g14822(.I(new_n15014_), .ZN(new_n15015_));
  OAI21_X1   g14823(.A1(new_n14865_), .A2(new_n14866_), .B(new_n14869_), .ZN(new_n15016_));
  NOR2_X1    g14824(.A1(new_n14985_), .A2(new_n15016_), .ZN(new_n15017_));
  XOR2_X1    g14825(.A1(new_n15017_), .A2(new_n14453_), .Z(new_n15018_));
  NAND3_X1   g14826(.A1(\asqrt[10] ), .A2(new_n14833_), .A3(new_n14852_), .ZN(new_n15019_));
  XOR2_X1    g14827(.A1(new_n15019_), .A2(new_n14863_), .Z(new_n15020_));
  OAI21_X1   g14828(.A1(new_n14827_), .A2(new_n14829_), .B(new_n14832_), .ZN(new_n15021_));
  NOR2_X1    g14829(.A1(new_n14985_), .A2(new_n15021_), .ZN(new_n15022_));
  XOR2_X1    g14830(.A1(new_n15022_), .A2(new_n14459_), .Z(new_n15023_));
  INV_X1     g14831(.I(new_n15023_), .ZN(new_n15024_));
  NAND3_X1   g14832(.A1(\asqrt[10] ), .A2(new_n14846_), .A3(new_n14828_), .ZN(new_n15025_));
  XOR2_X1    g14833(.A1(new_n15025_), .A2(new_n14463_), .Z(new_n15026_));
  INV_X1     g14834(.I(new_n15026_), .ZN(new_n15027_));
  OAI21_X1   g14835(.A1(new_n14841_), .A2(new_n14842_), .B(new_n14845_), .ZN(new_n15028_));
  NOR2_X1    g14836(.A1(new_n14985_), .A2(new_n15028_), .ZN(new_n15029_));
  XOR2_X1    g14837(.A1(new_n15029_), .A2(new_n14465_), .Z(new_n15030_));
  NAND3_X1   g14838(.A1(\asqrt[10] ), .A2(new_n14805_), .A3(new_n14824_), .ZN(new_n15031_));
  XOR2_X1    g14839(.A1(new_n15031_), .A2(new_n14839_), .Z(new_n15032_));
  OAI21_X1   g14840(.A1(new_n14799_), .A2(new_n14801_), .B(new_n14804_), .ZN(new_n15033_));
  NOR2_X1    g14841(.A1(new_n14985_), .A2(new_n15033_), .ZN(new_n15034_));
  XOR2_X1    g14842(.A1(new_n15034_), .A2(new_n14471_), .Z(new_n15035_));
  INV_X1     g14843(.I(new_n15035_), .ZN(new_n15036_));
  NAND3_X1   g14844(.A1(\asqrt[10] ), .A2(new_n14818_), .A3(new_n14800_), .ZN(new_n15037_));
  XOR2_X1    g14845(.A1(new_n15037_), .A2(new_n14475_), .Z(new_n15038_));
  INV_X1     g14846(.I(new_n15038_), .ZN(new_n15039_));
  OAI21_X1   g14847(.A1(new_n14813_), .A2(new_n14814_), .B(new_n14817_), .ZN(new_n15040_));
  NOR2_X1    g14848(.A1(new_n14985_), .A2(new_n15040_), .ZN(new_n15041_));
  XOR2_X1    g14849(.A1(new_n15041_), .A2(new_n14477_), .Z(new_n15042_));
  NAND3_X1   g14850(.A1(\asqrt[10] ), .A2(new_n14777_), .A3(new_n14796_), .ZN(new_n15043_));
  XOR2_X1    g14851(.A1(new_n15043_), .A2(new_n14811_), .Z(new_n15044_));
  OAI21_X1   g14852(.A1(new_n14771_), .A2(new_n14773_), .B(new_n14776_), .ZN(new_n15045_));
  NOR2_X1    g14853(.A1(new_n14985_), .A2(new_n15045_), .ZN(new_n15046_));
  XOR2_X1    g14854(.A1(new_n15046_), .A2(new_n14483_), .Z(new_n15047_));
  INV_X1     g14855(.I(new_n15047_), .ZN(new_n15048_));
  NAND3_X1   g14856(.A1(\asqrt[10] ), .A2(new_n14790_), .A3(new_n14772_), .ZN(new_n15049_));
  XOR2_X1    g14857(.A1(new_n15049_), .A2(new_n14487_), .Z(new_n15050_));
  INV_X1     g14858(.I(new_n15050_), .ZN(new_n15051_));
  OAI21_X1   g14859(.A1(new_n14785_), .A2(new_n14786_), .B(new_n14789_), .ZN(new_n15052_));
  NOR2_X1    g14860(.A1(new_n14985_), .A2(new_n15052_), .ZN(new_n15053_));
  XOR2_X1    g14861(.A1(new_n15053_), .A2(new_n14489_), .Z(new_n15054_));
  NAND3_X1   g14862(.A1(\asqrt[10] ), .A2(new_n14749_), .A3(new_n14768_), .ZN(new_n15055_));
  XOR2_X1    g14863(.A1(new_n15055_), .A2(new_n14783_), .Z(new_n15056_));
  OAI21_X1   g14864(.A1(new_n14743_), .A2(new_n14745_), .B(new_n14748_), .ZN(new_n15057_));
  NOR2_X1    g14865(.A1(new_n14985_), .A2(new_n15057_), .ZN(new_n15058_));
  XOR2_X1    g14866(.A1(new_n15058_), .A2(new_n14495_), .Z(new_n15059_));
  INV_X1     g14867(.I(new_n15059_), .ZN(new_n15060_));
  NAND3_X1   g14868(.A1(\asqrt[10] ), .A2(new_n14762_), .A3(new_n14744_), .ZN(new_n15061_));
  XOR2_X1    g14869(.A1(new_n15061_), .A2(new_n14499_), .Z(new_n15062_));
  INV_X1     g14870(.I(new_n15062_), .ZN(new_n15063_));
  OAI21_X1   g14871(.A1(new_n14757_), .A2(new_n14758_), .B(new_n14761_), .ZN(new_n15064_));
  NOR2_X1    g14872(.A1(new_n14985_), .A2(new_n15064_), .ZN(new_n15065_));
  XOR2_X1    g14873(.A1(new_n15065_), .A2(new_n14501_), .Z(new_n15066_));
  NAND3_X1   g14874(.A1(\asqrt[10] ), .A2(new_n14721_), .A3(new_n14740_), .ZN(new_n15067_));
  XOR2_X1    g14875(.A1(new_n15067_), .A2(new_n14755_), .Z(new_n15068_));
  OAI21_X1   g14876(.A1(new_n14715_), .A2(new_n14717_), .B(new_n14720_), .ZN(new_n15069_));
  NOR2_X1    g14877(.A1(new_n14985_), .A2(new_n15069_), .ZN(new_n15070_));
  XOR2_X1    g14878(.A1(new_n15070_), .A2(new_n14507_), .Z(new_n15071_));
  INV_X1     g14879(.I(new_n15071_), .ZN(new_n15072_));
  NAND3_X1   g14880(.A1(\asqrt[10] ), .A2(new_n14734_), .A3(new_n14716_), .ZN(new_n15073_));
  XOR2_X1    g14881(.A1(new_n15073_), .A2(new_n14511_), .Z(new_n15074_));
  INV_X1     g14882(.I(new_n15074_), .ZN(new_n15075_));
  OAI21_X1   g14883(.A1(new_n14729_), .A2(new_n14730_), .B(new_n14733_), .ZN(new_n15076_));
  NOR2_X1    g14884(.A1(new_n14985_), .A2(new_n15076_), .ZN(new_n15077_));
  XOR2_X1    g14885(.A1(new_n15077_), .A2(new_n14513_), .Z(new_n15078_));
  NAND3_X1   g14886(.A1(\asqrt[10] ), .A2(new_n14693_), .A3(new_n14712_), .ZN(new_n15079_));
  XOR2_X1    g14887(.A1(new_n15079_), .A2(new_n14727_), .Z(new_n15080_));
  OAI21_X1   g14888(.A1(new_n14687_), .A2(new_n14689_), .B(new_n14692_), .ZN(new_n15081_));
  NOR2_X1    g14889(.A1(new_n14985_), .A2(new_n15081_), .ZN(new_n15082_));
  XOR2_X1    g14890(.A1(new_n15082_), .A2(new_n14519_), .Z(new_n15083_));
  INV_X1     g14891(.I(new_n15083_), .ZN(new_n15084_));
  NAND3_X1   g14892(.A1(\asqrt[10] ), .A2(new_n14706_), .A3(new_n14688_), .ZN(new_n15085_));
  XOR2_X1    g14893(.A1(new_n15085_), .A2(new_n14523_), .Z(new_n15086_));
  INV_X1     g14894(.I(new_n15086_), .ZN(new_n15087_));
  OAI21_X1   g14895(.A1(new_n14701_), .A2(new_n14702_), .B(new_n14705_), .ZN(new_n15088_));
  NOR2_X1    g14896(.A1(new_n14985_), .A2(new_n15088_), .ZN(new_n15089_));
  XOR2_X1    g14897(.A1(new_n15089_), .A2(new_n14525_), .Z(new_n15090_));
  NAND3_X1   g14898(.A1(\asqrt[10] ), .A2(new_n14665_), .A3(new_n14684_), .ZN(new_n15091_));
  XOR2_X1    g14899(.A1(new_n15091_), .A2(new_n14699_), .Z(new_n15092_));
  OAI21_X1   g14900(.A1(new_n14659_), .A2(new_n14661_), .B(new_n14664_), .ZN(new_n15093_));
  NOR2_X1    g14901(.A1(new_n14985_), .A2(new_n15093_), .ZN(new_n15094_));
  XOR2_X1    g14902(.A1(new_n15094_), .A2(new_n14531_), .Z(new_n15095_));
  INV_X1     g14903(.I(new_n15095_), .ZN(new_n15096_));
  NAND3_X1   g14904(.A1(\asqrt[10] ), .A2(new_n14678_), .A3(new_n14660_), .ZN(new_n15097_));
  XOR2_X1    g14905(.A1(new_n15097_), .A2(new_n14535_), .Z(new_n15098_));
  INV_X1     g14906(.I(new_n15098_), .ZN(new_n15099_));
  OAI21_X1   g14907(.A1(new_n14673_), .A2(new_n14674_), .B(new_n14677_), .ZN(new_n15100_));
  NOR2_X1    g14908(.A1(new_n14985_), .A2(new_n15100_), .ZN(new_n15101_));
  XOR2_X1    g14909(.A1(new_n15101_), .A2(new_n14537_), .Z(new_n15102_));
  NAND3_X1   g14910(.A1(\asqrt[10] ), .A2(new_n14637_), .A3(new_n14656_), .ZN(new_n15103_));
  XOR2_X1    g14911(.A1(new_n15103_), .A2(new_n14671_), .Z(new_n15104_));
  OAI21_X1   g14912(.A1(new_n14631_), .A2(new_n14633_), .B(new_n14636_), .ZN(new_n15105_));
  NOR2_X1    g14913(.A1(new_n14985_), .A2(new_n15105_), .ZN(new_n15106_));
  XOR2_X1    g14914(.A1(new_n15106_), .A2(new_n14543_), .Z(new_n15107_));
  INV_X1     g14915(.I(new_n15107_), .ZN(new_n15108_));
  NAND3_X1   g14916(.A1(\asqrt[10] ), .A2(new_n14650_), .A3(new_n14632_), .ZN(new_n15109_));
  XOR2_X1    g14917(.A1(new_n15109_), .A2(new_n14547_), .Z(new_n15110_));
  INV_X1     g14918(.I(new_n15110_), .ZN(new_n15111_));
  OAI21_X1   g14919(.A1(new_n14645_), .A2(new_n14646_), .B(new_n14649_), .ZN(new_n15112_));
  NOR2_X1    g14920(.A1(new_n14985_), .A2(new_n15112_), .ZN(new_n15113_));
  XOR2_X1    g14921(.A1(new_n15113_), .A2(new_n14549_), .Z(new_n15114_));
  NAND3_X1   g14922(.A1(\asqrt[10] ), .A2(new_n14609_), .A3(new_n14628_), .ZN(new_n15115_));
  XOR2_X1    g14923(.A1(new_n15115_), .A2(new_n14643_), .Z(new_n15116_));
  OAI21_X1   g14924(.A1(new_n14603_), .A2(new_n14605_), .B(new_n14608_), .ZN(new_n15117_));
  NOR2_X1    g14925(.A1(new_n14985_), .A2(new_n15117_), .ZN(new_n15118_));
  XOR2_X1    g14926(.A1(new_n15118_), .A2(new_n14556_), .Z(new_n15119_));
  INV_X1     g14927(.I(new_n15119_), .ZN(new_n15120_));
  NAND3_X1   g14928(.A1(\asqrt[10] ), .A2(new_n14622_), .A3(new_n14604_), .ZN(new_n15121_));
  XOR2_X1    g14929(.A1(new_n15121_), .A2(new_n14559_), .Z(new_n15122_));
  INV_X1     g14930(.I(new_n15122_), .ZN(new_n15123_));
  OAI21_X1   g14931(.A1(new_n14617_), .A2(new_n14618_), .B(new_n14621_), .ZN(new_n15124_));
  NOR2_X1    g14932(.A1(new_n14985_), .A2(new_n15124_), .ZN(new_n15125_));
  XOR2_X1    g14933(.A1(new_n15125_), .A2(new_n14562_), .Z(new_n15126_));
  NAND3_X1   g14934(.A1(\asqrt[10] ), .A2(new_n14582_), .A3(new_n14600_), .ZN(new_n15127_));
  XOR2_X1    g14935(.A1(new_n15127_), .A2(new_n14616_), .Z(new_n15128_));
  NOR2_X1    g14936(.A1(new_n14579_), .A2(\asqrt[13] ), .ZN(new_n15129_));
  NOR3_X1    g14937(.A1(new_n14985_), .A2(new_n15129_), .A3(new_n14599_), .ZN(new_n15130_));
  XOR2_X1    g14938(.A1(new_n15130_), .A2(new_n14570_), .Z(new_n15131_));
  INV_X1     g14939(.I(new_n15131_), .ZN(new_n15132_));
  NAND3_X1   g14940(.A1(\asqrt[10] ), .A2(new_n14571_), .A3(new_n14572_), .ZN(new_n15133_));
  NOR4_X1    g14941(.A1(new_n14983_), .A2(new_n14430_), .A3(new_n14880_), .A4(new_n14984_), .ZN(new_n15134_));
  INV_X1     g14942(.I(new_n15134_), .ZN(new_n15135_));
  AOI21_X1   g14943(.A1(new_n15133_), .A2(new_n15135_), .B(\a[22] ), .ZN(new_n15136_));
  NOR3_X1    g14944(.A1(new_n14985_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n15137_));
  NOR3_X1    g14945(.A1(new_n15137_), .A2(new_n14066_), .A3(new_n15134_), .ZN(new_n15138_));
  NOR2_X1    g14946(.A1(new_n15138_), .A2(new_n15136_), .ZN(new_n15139_));
  INV_X1     g14947(.I(\a[18] ), .ZN(new_n15140_));
  INV_X1     g14948(.I(\a[19] ), .ZN(new_n15141_));
  NAND3_X1   g14949(.A1(new_n15140_), .A2(new_n15141_), .A3(new_n14571_), .ZN(new_n15142_));
  OAI21_X1   g14950(.A1(new_n14985_), .A2(new_n14571_), .B(new_n15142_), .ZN(new_n15143_));
  NAND2_X1   g14951(.A1(new_n15143_), .A2(\asqrt[11] ), .ZN(new_n15144_));
  OAI21_X1   g14952(.A1(new_n14985_), .A2(\a[20] ), .B(\a[21] ), .ZN(new_n15145_));
  NAND2_X1   g14953(.A1(new_n15145_), .A2(new_n15133_), .ZN(new_n15146_));
  NOR2_X1    g14954(.A1(new_n15143_), .A2(\asqrt[11] ), .ZN(new_n15147_));
  OAI21_X1   g14955(.A1(new_n15146_), .A2(new_n15147_), .B(new_n15144_), .ZN(new_n15148_));
  OAI21_X1   g14956(.A1(new_n15148_), .A2(\asqrt[12] ), .B(new_n15139_), .ZN(new_n15149_));
  NAND2_X1   g14957(.A1(new_n15148_), .A2(\asqrt[12] ), .ZN(new_n15150_));
  NAND3_X1   g14958(.A1(new_n15149_), .A2(new_n13382_), .A3(new_n15150_), .ZN(new_n15151_));
  NOR3_X1    g14959(.A1(new_n14985_), .A2(new_n14593_), .A3(new_n14578_), .ZN(new_n15152_));
  XOR2_X1    g14960(.A1(new_n15152_), .A2(new_n14595_), .Z(new_n15153_));
  AOI21_X1   g14961(.A1(new_n15149_), .A2(new_n15150_), .B(new_n13382_), .ZN(new_n15154_));
  AOI21_X1   g14962(.A1(new_n15151_), .A2(new_n15153_), .B(new_n15154_), .ZN(new_n15155_));
  AOI21_X1   g14963(.A1(new_n15155_), .A2(new_n12889_), .B(new_n15132_), .ZN(new_n15156_));
  OAI21_X1   g14964(.A1(new_n15155_), .A2(new_n12889_), .B(new_n12374_), .ZN(new_n15157_));
  OAI21_X1   g14965(.A1(new_n15156_), .A2(new_n15157_), .B(new_n15128_), .ZN(new_n15158_));
  NOR2_X1    g14966(.A1(new_n15155_), .A2(new_n12889_), .ZN(new_n15159_));
  OAI21_X1   g14967(.A1(new_n15156_), .A2(new_n15159_), .B(\asqrt[15] ), .ZN(new_n15160_));
  NAND3_X1   g14968(.A1(new_n15158_), .A2(new_n15160_), .A3(new_n11901_), .ZN(new_n15161_));
  NAND2_X1   g14969(.A1(new_n15161_), .A2(new_n15126_), .ZN(new_n15162_));
  NAND2_X1   g14970(.A1(new_n15158_), .A2(new_n15160_), .ZN(new_n15163_));
  AOI21_X1   g14971(.A1(new_n15163_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n15164_));
  AOI21_X1   g14972(.A1(new_n15164_), .A2(new_n15162_), .B(new_n15123_), .ZN(new_n15165_));
  INV_X1     g14973(.I(new_n15128_), .ZN(new_n15166_));
  OAI21_X1   g14974(.A1(new_n15137_), .A2(new_n15134_), .B(new_n14066_), .ZN(new_n15167_));
  NAND3_X1   g14975(.A1(new_n15133_), .A2(new_n15135_), .A3(\a[22] ), .ZN(new_n15168_));
  NAND2_X1   g14976(.A1(new_n15167_), .A2(new_n15168_), .ZN(new_n15169_));
  NAND2_X1   g14977(.A1(\asqrt[10] ), .A2(\a[20] ), .ZN(new_n15170_));
  AOI21_X1   g14978(.A1(new_n15170_), .A2(new_n15142_), .B(new_n14430_), .ZN(new_n15171_));
  AOI21_X1   g14979(.A1(\asqrt[10] ), .A2(new_n14571_), .B(new_n14572_), .ZN(new_n15172_));
  NOR2_X1    g14980(.A1(new_n15137_), .A2(new_n15172_), .ZN(new_n15173_));
  NAND3_X1   g14981(.A1(new_n15170_), .A2(new_n14430_), .A3(new_n15142_), .ZN(new_n15174_));
  AOI21_X1   g14982(.A1(new_n15173_), .A2(new_n15174_), .B(new_n15171_), .ZN(new_n15175_));
  AOI21_X1   g14983(.A1(new_n15175_), .A2(new_n13917_), .B(new_n15169_), .ZN(new_n15176_));
  NOR2_X1    g14984(.A1(new_n15175_), .A2(new_n13917_), .ZN(new_n15177_));
  NOR3_X1    g14985(.A1(new_n15176_), .A2(\asqrt[13] ), .A3(new_n15177_), .ZN(new_n15178_));
  INV_X1     g14986(.I(new_n15153_), .ZN(new_n15179_));
  OAI21_X1   g14987(.A1(new_n15176_), .A2(new_n15177_), .B(\asqrt[13] ), .ZN(new_n15180_));
  OAI21_X1   g14988(.A1(new_n15178_), .A2(new_n15179_), .B(new_n15180_), .ZN(new_n15181_));
  OAI21_X1   g14989(.A1(new_n15181_), .A2(\asqrt[14] ), .B(new_n15131_), .ZN(new_n15182_));
  AOI21_X1   g14990(.A1(new_n15181_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n15183_));
  AOI21_X1   g14991(.A1(new_n15183_), .A2(new_n15182_), .B(new_n15166_), .ZN(new_n15184_));
  NAND2_X1   g14992(.A1(new_n15181_), .A2(\asqrt[14] ), .ZN(new_n15185_));
  AOI21_X1   g14993(.A1(new_n15182_), .A2(new_n15185_), .B(new_n12374_), .ZN(new_n15186_));
  OAI21_X1   g14994(.A1(new_n15184_), .A2(new_n15186_), .B(\asqrt[16] ), .ZN(new_n15187_));
  AOI21_X1   g14995(.A1(new_n15162_), .A2(new_n15187_), .B(new_n11406_), .ZN(new_n15188_));
  NOR2_X1    g14996(.A1(new_n15165_), .A2(new_n15188_), .ZN(new_n15189_));
  AOI21_X1   g14997(.A1(new_n15189_), .A2(new_n10953_), .B(new_n15120_), .ZN(new_n15190_));
  OAI21_X1   g14998(.A1(new_n15165_), .A2(new_n15188_), .B(\asqrt[18] ), .ZN(new_n15191_));
  NAND2_X1   g14999(.A1(new_n15191_), .A2(new_n10478_), .ZN(new_n15192_));
  OAI21_X1   g15000(.A1(new_n15190_), .A2(new_n15192_), .B(new_n15116_), .ZN(new_n15193_));
  INV_X1     g15001(.I(new_n15191_), .ZN(new_n15194_));
  OAI21_X1   g15002(.A1(new_n15190_), .A2(new_n15194_), .B(\asqrt[19] ), .ZN(new_n15195_));
  NAND3_X1   g15003(.A1(new_n15193_), .A2(new_n15195_), .A3(new_n10045_), .ZN(new_n15196_));
  NAND2_X1   g15004(.A1(new_n15196_), .A2(new_n15114_), .ZN(new_n15197_));
  NAND2_X1   g15005(.A1(new_n15193_), .A2(new_n15195_), .ZN(new_n15198_));
  AOI21_X1   g15006(.A1(new_n15198_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n15199_));
  AOI21_X1   g15007(.A1(new_n15199_), .A2(new_n15197_), .B(new_n15111_), .ZN(new_n15200_));
  INV_X1     g15008(.I(new_n15116_), .ZN(new_n15201_));
  INV_X1     g15009(.I(new_n15126_), .ZN(new_n15202_));
  NOR2_X1    g15010(.A1(new_n15184_), .A2(new_n15186_), .ZN(new_n15203_));
  AOI21_X1   g15011(.A1(new_n15203_), .A2(new_n11901_), .B(new_n15202_), .ZN(new_n15204_));
  NAND2_X1   g15012(.A1(new_n15187_), .A2(new_n11406_), .ZN(new_n15205_));
  OAI21_X1   g15013(.A1(new_n15204_), .A2(new_n15205_), .B(new_n15122_), .ZN(new_n15206_));
  INV_X1     g15014(.I(new_n15187_), .ZN(new_n15207_));
  OAI21_X1   g15015(.A1(new_n15204_), .A2(new_n15207_), .B(\asqrt[17] ), .ZN(new_n15208_));
  NAND3_X1   g15016(.A1(new_n15206_), .A2(new_n15208_), .A3(new_n10953_), .ZN(new_n15209_));
  NAND2_X1   g15017(.A1(new_n15209_), .A2(new_n15119_), .ZN(new_n15210_));
  NAND2_X1   g15018(.A1(new_n15206_), .A2(new_n15208_), .ZN(new_n15211_));
  AOI21_X1   g15019(.A1(new_n15211_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n15212_));
  AOI21_X1   g15020(.A1(new_n15212_), .A2(new_n15210_), .B(new_n15201_), .ZN(new_n15213_));
  AOI21_X1   g15021(.A1(new_n15210_), .A2(new_n15191_), .B(new_n10478_), .ZN(new_n15214_));
  OAI21_X1   g15022(.A1(new_n15213_), .A2(new_n15214_), .B(\asqrt[20] ), .ZN(new_n15215_));
  AOI21_X1   g15023(.A1(new_n15197_), .A2(new_n15215_), .B(new_n9590_), .ZN(new_n15216_));
  NOR2_X1    g15024(.A1(new_n15200_), .A2(new_n15216_), .ZN(new_n15217_));
  AOI21_X1   g15025(.A1(new_n15217_), .A2(new_n9177_), .B(new_n15108_), .ZN(new_n15218_));
  OAI21_X1   g15026(.A1(new_n15200_), .A2(new_n15216_), .B(\asqrt[22] ), .ZN(new_n15219_));
  NAND2_X1   g15027(.A1(new_n15219_), .A2(new_n8742_), .ZN(new_n15220_));
  OAI21_X1   g15028(.A1(new_n15218_), .A2(new_n15220_), .B(new_n15104_), .ZN(new_n15221_));
  INV_X1     g15029(.I(new_n15219_), .ZN(new_n15222_));
  OAI21_X1   g15030(.A1(new_n15218_), .A2(new_n15222_), .B(\asqrt[23] ), .ZN(new_n15223_));
  NAND3_X1   g15031(.A1(new_n15221_), .A2(new_n15223_), .A3(new_n8349_), .ZN(new_n15224_));
  NAND2_X1   g15032(.A1(new_n15224_), .A2(new_n15102_), .ZN(new_n15225_));
  NAND2_X1   g15033(.A1(new_n15221_), .A2(new_n15223_), .ZN(new_n15226_));
  AOI21_X1   g15034(.A1(new_n15226_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n15227_));
  AOI21_X1   g15035(.A1(new_n15227_), .A2(new_n15225_), .B(new_n15099_), .ZN(new_n15228_));
  INV_X1     g15036(.I(new_n15104_), .ZN(new_n15229_));
  INV_X1     g15037(.I(new_n15114_), .ZN(new_n15230_));
  NOR2_X1    g15038(.A1(new_n15213_), .A2(new_n15214_), .ZN(new_n15231_));
  AOI21_X1   g15039(.A1(new_n15231_), .A2(new_n10045_), .B(new_n15230_), .ZN(new_n15232_));
  NAND2_X1   g15040(.A1(new_n15215_), .A2(new_n9590_), .ZN(new_n15233_));
  OAI21_X1   g15041(.A1(new_n15232_), .A2(new_n15233_), .B(new_n15110_), .ZN(new_n15234_));
  INV_X1     g15042(.I(new_n15215_), .ZN(new_n15235_));
  OAI21_X1   g15043(.A1(new_n15232_), .A2(new_n15235_), .B(\asqrt[21] ), .ZN(new_n15236_));
  NAND3_X1   g15044(.A1(new_n15234_), .A2(new_n15236_), .A3(new_n9177_), .ZN(new_n15237_));
  NAND2_X1   g15045(.A1(new_n15237_), .A2(new_n15107_), .ZN(new_n15238_));
  NAND2_X1   g15046(.A1(new_n15234_), .A2(new_n15236_), .ZN(new_n15239_));
  AOI21_X1   g15047(.A1(new_n15239_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n15240_));
  AOI21_X1   g15048(.A1(new_n15240_), .A2(new_n15238_), .B(new_n15229_), .ZN(new_n15241_));
  AOI21_X1   g15049(.A1(new_n15238_), .A2(new_n15219_), .B(new_n8742_), .ZN(new_n15242_));
  OAI21_X1   g15050(.A1(new_n15241_), .A2(new_n15242_), .B(\asqrt[24] ), .ZN(new_n15243_));
  AOI21_X1   g15051(.A1(new_n15225_), .A2(new_n15243_), .B(new_n7934_), .ZN(new_n15244_));
  NOR2_X1    g15052(.A1(new_n15228_), .A2(new_n15244_), .ZN(new_n15245_));
  AOI21_X1   g15053(.A1(new_n15245_), .A2(new_n7561_), .B(new_n15096_), .ZN(new_n15246_));
  OAI21_X1   g15054(.A1(new_n15228_), .A2(new_n15244_), .B(\asqrt[26] ), .ZN(new_n15247_));
  NAND2_X1   g15055(.A1(new_n15247_), .A2(new_n7166_), .ZN(new_n15248_));
  OAI21_X1   g15056(.A1(new_n15246_), .A2(new_n15248_), .B(new_n15092_), .ZN(new_n15249_));
  INV_X1     g15057(.I(new_n15247_), .ZN(new_n15250_));
  OAI21_X1   g15058(.A1(new_n15246_), .A2(new_n15250_), .B(\asqrt[27] ), .ZN(new_n15251_));
  NAND3_X1   g15059(.A1(new_n15249_), .A2(new_n15251_), .A3(new_n6813_), .ZN(new_n15252_));
  NAND2_X1   g15060(.A1(new_n15252_), .A2(new_n15090_), .ZN(new_n15253_));
  NAND2_X1   g15061(.A1(new_n15249_), .A2(new_n15251_), .ZN(new_n15254_));
  AOI21_X1   g15062(.A1(new_n15254_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n15255_));
  AOI21_X1   g15063(.A1(new_n15255_), .A2(new_n15253_), .B(new_n15087_), .ZN(new_n15256_));
  INV_X1     g15064(.I(new_n15092_), .ZN(new_n15257_));
  INV_X1     g15065(.I(new_n15102_), .ZN(new_n15258_));
  NOR2_X1    g15066(.A1(new_n15241_), .A2(new_n15242_), .ZN(new_n15259_));
  AOI21_X1   g15067(.A1(new_n15259_), .A2(new_n8349_), .B(new_n15258_), .ZN(new_n15260_));
  NAND2_X1   g15068(.A1(new_n15243_), .A2(new_n7934_), .ZN(new_n15261_));
  OAI21_X1   g15069(.A1(new_n15260_), .A2(new_n15261_), .B(new_n15098_), .ZN(new_n15262_));
  INV_X1     g15070(.I(new_n15243_), .ZN(new_n15263_));
  OAI21_X1   g15071(.A1(new_n15260_), .A2(new_n15263_), .B(\asqrt[25] ), .ZN(new_n15264_));
  NAND3_X1   g15072(.A1(new_n15262_), .A2(new_n15264_), .A3(new_n7561_), .ZN(new_n15265_));
  NAND2_X1   g15073(.A1(new_n15265_), .A2(new_n15095_), .ZN(new_n15266_));
  NAND2_X1   g15074(.A1(new_n15262_), .A2(new_n15264_), .ZN(new_n15267_));
  AOI21_X1   g15075(.A1(new_n15267_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n15268_));
  AOI21_X1   g15076(.A1(new_n15268_), .A2(new_n15266_), .B(new_n15257_), .ZN(new_n15269_));
  AOI21_X1   g15077(.A1(new_n15266_), .A2(new_n15247_), .B(new_n7166_), .ZN(new_n15270_));
  OAI21_X1   g15078(.A1(new_n15269_), .A2(new_n15270_), .B(\asqrt[28] ), .ZN(new_n15271_));
  AOI21_X1   g15079(.A1(new_n15253_), .A2(new_n15271_), .B(new_n6454_), .ZN(new_n15272_));
  NOR2_X1    g15080(.A1(new_n15256_), .A2(new_n15272_), .ZN(new_n15273_));
  AOI21_X1   g15081(.A1(new_n15273_), .A2(new_n6106_), .B(new_n15084_), .ZN(new_n15274_));
  OAI21_X1   g15082(.A1(new_n15256_), .A2(new_n15272_), .B(\asqrt[30] ), .ZN(new_n15275_));
  NAND2_X1   g15083(.A1(new_n15275_), .A2(new_n5750_), .ZN(new_n15276_));
  OAI21_X1   g15084(.A1(new_n15274_), .A2(new_n15276_), .B(new_n15080_), .ZN(new_n15277_));
  INV_X1     g15085(.I(new_n15275_), .ZN(new_n15278_));
  OAI21_X1   g15086(.A1(new_n15274_), .A2(new_n15278_), .B(\asqrt[31] ), .ZN(new_n15279_));
  NAND3_X1   g15087(.A1(new_n15277_), .A2(new_n15279_), .A3(new_n5435_), .ZN(new_n15280_));
  NAND2_X1   g15088(.A1(new_n15280_), .A2(new_n15078_), .ZN(new_n15281_));
  NAND2_X1   g15089(.A1(new_n15277_), .A2(new_n15279_), .ZN(new_n15282_));
  AOI21_X1   g15090(.A1(new_n15282_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n15283_));
  AOI21_X1   g15091(.A1(new_n15283_), .A2(new_n15281_), .B(new_n15075_), .ZN(new_n15284_));
  INV_X1     g15092(.I(new_n15080_), .ZN(new_n15285_));
  INV_X1     g15093(.I(new_n15090_), .ZN(new_n15286_));
  NOR2_X1    g15094(.A1(new_n15269_), .A2(new_n15270_), .ZN(new_n15287_));
  AOI21_X1   g15095(.A1(new_n15287_), .A2(new_n6813_), .B(new_n15286_), .ZN(new_n15288_));
  NAND2_X1   g15096(.A1(new_n15271_), .A2(new_n6454_), .ZN(new_n15289_));
  OAI21_X1   g15097(.A1(new_n15288_), .A2(new_n15289_), .B(new_n15086_), .ZN(new_n15290_));
  INV_X1     g15098(.I(new_n15271_), .ZN(new_n15291_));
  OAI21_X1   g15099(.A1(new_n15288_), .A2(new_n15291_), .B(\asqrt[29] ), .ZN(new_n15292_));
  NAND3_X1   g15100(.A1(new_n15290_), .A2(new_n15292_), .A3(new_n6106_), .ZN(new_n15293_));
  NAND2_X1   g15101(.A1(new_n15293_), .A2(new_n15083_), .ZN(new_n15294_));
  NAND2_X1   g15102(.A1(new_n15290_), .A2(new_n15292_), .ZN(new_n15295_));
  AOI21_X1   g15103(.A1(new_n15295_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n15296_));
  AOI21_X1   g15104(.A1(new_n15296_), .A2(new_n15294_), .B(new_n15285_), .ZN(new_n15297_));
  AOI21_X1   g15105(.A1(new_n15294_), .A2(new_n15275_), .B(new_n5750_), .ZN(new_n15298_));
  OAI21_X1   g15106(.A1(new_n15297_), .A2(new_n15298_), .B(\asqrt[32] ), .ZN(new_n15299_));
  AOI21_X1   g15107(.A1(new_n15281_), .A2(new_n15299_), .B(new_n5110_), .ZN(new_n15300_));
  NOR2_X1    g15108(.A1(new_n15284_), .A2(new_n15300_), .ZN(new_n15301_));
  AOI21_X1   g15109(.A1(new_n15301_), .A2(new_n4810_), .B(new_n15072_), .ZN(new_n15302_));
  OAI21_X1   g15110(.A1(new_n15284_), .A2(new_n15300_), .B(\asqrt[34] ), .ZN(new_n15303_));
  NAND2_X1   g15111(.A1(new_n15303_), .A2(new_n4510_), .ZN(new_n15304_));
  OAI21_X1   g15112(.A1(new_n15302_), .A2(new_n15304_), .B(new_n15068_), .ZN(new_n15305_));
  INV_X1     g15113(.I(new_n15303_), .ZN(new_n15306_));
  OAI21_X1   g15114(.A1(new_n15302_), .A2(new_n15306_), .B(\asqrt[35] ), .ZN(new_n15307_));
  NAND3_X1   g15115(.A1(new_n15305_), .A2(new_n15307_), .A3(new_n4224_), .ZN(new_n15308_));
  NAND2_X1   g15116(.A1(new_n15308_), .A2(new_n15066_), .ZN(new_n15309_));
  NAND2_X1   g15117(.A1(new_n15305_), .A2(new_n15307_), .ZN(new_n15310_));
  AOI21_X1   g15118(.A1(new_n15310_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n15311_));
  AOI21_X1   g15119(.A1(new_n15311_), .A2(new_n15309_), .B(new_n15063_), .ZN(new_n15312_));
  INV_X1     g15120(.I(new_n15068_), .ZN(new_n15313_));
  INV_X1     g15121(.I(new_n15078_), .ZN(new_n15314_));
  NOR2_X1    g15122(.A1(new_n15297_), .A2(new_n15298_), .ZN(new_n15315_));
  AOI21_X1   g15123(.A1(new_n15315_), .A2(new_n5435_), .B(new_n15314_), .ZN(new_n15316_));
  NAND2_X1   g15124(.A1(new_n15299_), .A2(new_n5110_), .ZN(new_n15317_));
  OAI21_X1   g15125(.A1(new_n15316_), .A2(new_n15317_), .B(new_n15074_), .ZN(new_n15318_));
  INV_X1     g15126(.I(new_n15299_), .ZN(new_n15319_));
  OAI21_X1   g15127(.A1(new_n15316_), .A2(new_n15319_), .B(\asqrt[33] ), .ZN(new_n15320_));
  NAND3_X1   g15128(.A1(new_n15318_), .A2(new_n15320_), .A3(new_n4810_), .ZN(new_n15321_));
  NAND2_X1   g15129(.A1(new_n15321_), .A2(new_n15071_), .ZN(new_n15322_));
  NAND2_X1   g15130(.A1(new_n15318_), .A2(new_n15320_), .ZN(new_n15323_));
  AOI21_X1   g15131(.A1(new_n15323_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n15324_));
  AOI21_X1   g15132(.A1(new_n15324_), .A2(new_n15322_), .B(new_n15313_), .ZN(new_n15325_));
  AOI21_X1   g15133(.A1(new_n15322_), .A2(new_n15303_), .B(new_n4510_), .ZN(new_n15326_));
  OAI21_X1   g15134(.A1(new_n15325_), .A2(new_n15326_), .B(\asqrt[36] ), .ZN(new_n15327_));
  AOI21_X1   g15135(.A1(new_n15309_), .A2(new_n15327_), .B(new_n3928_), .ZN(new_n15328_));
  NOR2_X1    g15136(.A1(new_n15312_), .A2(new_n15328_), .ZN(new_n15329_));
  AOI21_X1   g15137(.A1(new_n15329_), .A2(new_n3675_), .B(new_n15060_), .ZN(new_n15330_));
  OAI21_X1   g15138(.A1(new_n15312_), .A2(new_n15328_), .B(\asqrt[38] ), .ZN(new_n15331_));
  NAND2_X1   g15139(.A1(new_n15331_), .A2(new_n3400_), .ZN(new_n15332_));
  OAI21_X1   g15140(.A1(new_n15330_), .A2(new_n15332_), .B(new_n15056_), .ZN(new_n15333_));
  INV_X1     g15141(.I(new_n15331_), .ZN(new_n15334_));
  OAI21_X1   g15142(.A1(new_n15330_), .A2(new_n15334_), .B(\asqrt[39] ), .ZN(new_n15335_));
  NAND3_X1   g15143(.A1(new_n15333_), .A2(new_n15335_), .A3(new_n3167_), .ZN(new_n15336_));
  NAND2_X1   g15144(.A1(new_n15336_), .A2(new_n15054_), .ZN(new_n15337_));
  NAND2_X1   g15145(.A1(new_n15333_), .A2(new_n15335_), .ZN(new_n15338_));
  AOI21_X1   g15146(.A1(new_n15338_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n15339_));
  AOI21_X1   g15147(.A1(new_n15339_), .A2(new_n15337_), .B(new_n15051_), .ZN(new_n15340_));
  INV_X1     g15148(.I(new_n15056_), .ZN(new_n15341_));
  INV_X1     g15149(.I(new_n15066_), .ZN(new_n15342_));
  NOR2_X1    g15150(.A1(new_n15325_), .A2(new_n15326_), .ZN(new_n15343_));
  AOI21_X1   g15151(.A1(new_n15343_), .A2(new_n4224_), .B(new_n15342_), .ZN(new_n15344_));
  NAND2_X1   g15152(.A1(new_n15327_), .A2(new_n3928_), .ZN(new_n15345_));
  OAI21_X1   g15153(.A1(new_n15344_), .A2(new_n15345_), .B(new_n15062_), .ZN(new_n15346_));
  INV_X1     g15154(.I(new_n15327_), .ZN(new_n15347_));
  OAI21_X1   g15155(.A1(new_n15344_), .A2(new_n15347_), .B(\asqrt[37] ), .ZN(new_n15348_));
  NAND3_X1   g15156(.A1(new_n15346_), .A2(new_n15348_), .A3(new_n3675_), .ZN(new_n15349_));
  NAND2_X1   g15157(.A1(new_n15349_), .A2(new_n15059_), .ZN(new_n15350_));
  NAND2_X1   g15158(.A1(new_n15346_), .A2(new_n15348_), .ZN(new_n15351_));
  AOI21_X1   g15159(.A1(new_n15351_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n15352_));
  AOI21_X1   g15160(.A1(new_n15352_), .A2(new_n15350_), .B(new_n15341_), .ZN(new_n15353_));
  AOI21_X1   g15161(.A1(new_n15350_), .A2(new_n15331_), .B(new_n3400_), .ZN(new_n15354_));
  OAI21_X1   g15162(.A1(new_n15353_), .A2(new_n15354_), .B(\asqrt[40] ), .ZN(new_n15355_));
  AOI21_X1   g15163(.A1(new_n15337_), .A2(new_n15355_), .B(new_n2912_), .ZN(new_n15356_));
  NOR2_X1    g15164(.A1(new_n15340_), .A2(new_n15356_), .ZN(new_n15357_));
  AOI21_X1   g15165(.A1(new_n15357_), .A2(new_n2699_), .B(new_n15048_), .ZN(new_n15358_));
  OAI21_X1   g15166(.A1(new_n15340_), .A2(new_n15356_), .B(\asqrt[42] ), .ZN(new_n15359_));
  NAND2_X1   g15167(.A1(new_n15359_), .A2(new_n2464_), .ZN(new_n15360_));
  OAI21_X1   g15168(.A1(new_n15358_), .A2(new_n15360_), .B(new_n15044_), .ZN(new_n15361_));
  INV_X1     g15169(.I(new_n15359_), .ZN(new_n15362_));
  OAI21_X1   g15170(.A1(new_n15358_), .A2(new_n15362_), .B(\asqrt[43] ), .ZN(new_n15363_));
  NAND3_X1   g15171(.A1(new_n15361_), .A2(new_n15363_), .A3(new_n2271_), .ZN(new_n15364_));
  NAND2_X1   g15172(.A1(new_n15364_), .A2(new_n15042_), .ZN(new_n15365_));
  NAND2_X1   g15173(.A1(new_n15361_), .A2(new_n15363_), .ZN(new_n15366_));
  AOI21_X1   g15174(.A1(new_n15366_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n15367_));
  AOI21_X1   g15175(.A1(new_n15367_), .A2(new_n15365_), .B(new_n15039_), .ZN(new_n15368_));
  INV_X1     g15176(.I(new_n15044_), .ZN(new_n15369_));
  INV_X1     g15177(.I(new_n15054_), .ZN(new_n15370_));
  NOR2_X1    g15178(.A1(new_n15353_), .A2(new_n15354_), .ZN(new_n15371_));
  AOI21_X1   g15179(.A1(new_n15371_), .A2(new_n3167_), .B(new_n15370_), .ZN(new_n15372_));
  NAND2_X1   g15180(.A1(new_n15355_), .A2(new_n2912_), .ZN(new_n15373_));
  OAI21_X1   g15181(.A1(new_n15372_), .A2(new_n15373_), .B(new_n15050_), .ZN(new_n15374_));
  INV_X1     g15182(.I(new_n15355_), .ZN(new_n15375_));
  OAI21_X1   g15183(.A1(new_n15372_), .A2(new_n15375_), .B(\asqrt[41] ), .ZN(new_n15376_));
  NAND3_X1   g15184(.A1(new_n15374_), .A2(new_n15376_), .A3(new_n2699_), .ZN(new_n15377_));
  NAND2_X1   g15185(.A1(new_n15377_), .A2(new_n15047_), .ZN(new_n15378_));
  NAND2_X1   g15186(.A1(new_n15374_), .A2(new_n15376_), .ZN(new_n15379_));
  AOI21_X1   g15187(.A1(new_n15379_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n15380_));
  AOI21_X1   g15188(.A1(new_n15380_), .A2(new_n15378_), .B(new_n15369_), .ZN(new_n15381_));
  AOI21_X1   g15189(.A1(new_n15378_), .A2(new_n15359_), .B(new_n2464_), .ZN(new_n15382_));
  OAI21_X1   g15190(.A1(new_n15381_), .A2(new_n15382_), .B(\asqrt[44] ), .ZN(new_n15383_));
  AOI21_X1   g15191(.A1(new_n15365_), .A2(new_n15383_), .B(new_n2072_), .ZN(new_n15384_));
  NOR2_X1    g15192(.A1(new_n15368_), .A2(new_n15384_), .ZN(new_n15385_));
  AOI21_X1   g15193(.A1(new_n15385_), .A2(new_n1884_), .B(new_n15036_), .ZN(new_n15386_));
  OAI21_X1   g15194(.A1(new_n15368_), .A2(new_n15384_), .B(\asqrt[46] ), .ZN(new_n15387_));
  NAND2_X1   g15195(.A1(new_n15387_), .A2(new_n1688_), .ZN(new_n15388_));
  OAI21_X1   g15196(.A1(new_n15386_), .A2(new_n15388_), .B(new_n15032_), .ZN(new_n15389_));
  INV_X1     g15197(.I(new_n15387_), .ZN(new_n15390_));
  OAI21_X1   g15198(.A1(new_n15386_), .A2(new_n15390_), .B(\asqrt[47] ), .ZN(new_n15391_));
  NAND3_X1   g15199(.A1(new_n15389_), .A2(new_n15391_), .A3(new_n1533_), .ZN(new_n15392_));
  NAND2_X1   g15200(.A1(new_n15392_), .A2(new_n15030_), .ZN(new_n15393_));
  NAND2_X1   g15201(.A1(new_n15389_), .A2(new_n15391_), .ZN(new_n15394_));
  AOI21_X1   g15202(.A1(new_n15394_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n15395_));
  AOI21_X1   g15203(.A1(new_n15395_), .A2(new_n15393_), .B(new_n15027_), .ZN(new_n15396_));
  INV_X1     g15204(.I(new_n15032_), .ZN(new_n15397_));
  INV_X1     g15205(.I(new_n15042_), .ZN(new_n15398_));
  NOR2_X1    g15206(.A1(new_n15381_), .A2(new_n15382_), .ZN(new_n15399_));
  AOI21_X1   g15207(.A1(new_n15399_), .A2(new_n2271_), .B(new_n15398_), .ZN(new_n15400_));
  NAND2_X1   g15208(.A1(new_n15383_), .A2(new_n2072_), .ZN(new_n15401_));
  OAI21_X1   g15209(.A1(new_n15400_), .A2(new_n15401_), .B(new_n15038_), .ZN(new_n15402_));
  INV_X1     g15210(.I(new_n15383_), .ZN(new_n15403_));
  OAI21_X1   g15211(.A1(new_n15400_), .A2(new_n15403_), .B(\asqrt[45] ), .ZN(new_n15404_));
  NAND3_X1   g15212(.A1(new_n15402_), .A2(new_n15404_), .A3(new_n1884_), .ZN(new_n15405_));
  NAND2_X1   g15213(.A1(new_n15405_), .A2(new_n15035_), .ZN(new_n15406_));
  NAND2_X1   g15214(.A1(new_n15402_), .A2(new_n15404_), .ZN(new_n15407_));
  AOI21_X1   g15215(.A1(new_n15407_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n15408_));
  AOI21_X1   g15216(.A1(new_n15408_), .A2(new_n15406_), .B(new_n15397_), .ZN(new_n15409_));
  AOI21_X1   g15217(.A1(new_n15406_), .A2(new_n15387_), .B(new_n1688_), .ZN(new_n15410_));
  OAI21_X1   g15218(.A1(new_n15409_), .A2(new_n15410_), .B(\asqrt[48] ), .ZN(new_n15411_));
  AOI21_X1   g15219(.A1(new_n15393_), .A2(new_n15411_), .B(new_n1368_), .ZN(new_n15412_));
  NOR2_X1    g15220(.A1(new_n15396_), .A2(new_n15412_), .ZN(new_n15413_));
  AOI21_X1   g15221(.A1(new_n15413_), .A2(new_n1228_), .B(new_n15024_), .ZN(new_n15414_));
  OAI21_X1   g15222(.A1(new_n15396_), .A2(new_n15412_), .B(\asqrt[50] ), .ZN(new_n15415_));
  NAND2_X1   g15223(.A1(new_n15415_), .A2(new_n1088_), .ZN(new_n15416_));
  OAI21_X1   g15224(.A1(new_n15414_), .A2(new_n15416_), .B(new_n15020_), .ZN(new_n15417_));
  INV_X1     g15225(.I(new_n15415_), .ZN(new_n15418_));
  OAI21_X1   g15226(.A1(new_n15414_), .A2(new_n15418_), .B(\asqrt[51] ), .ZN(new_n15419_));
  NAND3_X1   g15227(.A1(new_n15417_), .A2(new_n15419_), .A3(new_n962_), .ZN(new_n15420_));
  NAND2_X1   g15228(.A1(new_n15420_), .A2(new_n15018_), .ZN(new_n15421_));
  NAND2_X1   g15229(.A1(new_n15417_), .A2(new_n15419_), .ZN(new_n15422_));
  AOI21_X1   g15230(.A1(new_n15422_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n15423_));
  AOI21_X1   g15231(.A1(new_n15423_), .A2(new_n15421_), .B(new_n15015_), .ZN(new_n15424_));
  INV_X1     g15232(.I(new_n15020_), .ZN(new_n15425_));
  INV_X1     g15233(.I(new_n15030_), .ZN(new_n15426_));
  NOR2_X1    g15234(.A1(new_n15409_), .A2(new_n15410_), .ZN(new_n15427_));
  AOI21_X1   g15235(.A1(new_n15427_), .A2(new_n1533_), .B(new_n15426_), .ZN(new_n15428_));
  NAND2_X1   g15236(.A1(new_n15411_), .A2(new_n1368_), .ZN(new_n15429_));
  OAI21_X1   g15237(.A1(new_n15428_), .A2(new_n15429_), .B(new_n15026_), .ZN(new_n15430_));
  INV_X1     g15238(.I(new_n15411_), .ZN(new_n15431_));
  OAI21_X1   g15239(.A1(new_n15428_), .A2(new_n15431_), .B(\asqrt[49] ), .ZN(new_n15432_));
  NAND3_X1   g15240(.A1(new_n15430_), .A2(new_n15432_), .A3(new_n1228_), .ZN(new_n15433_));
  NAND2_X1   g15241(.A1(new_n15433_), .A2(new_n15023_), .ZN(new_n15434_));
  NAND2_X1   g15242(.A1(new_n15430_), .A2(new_n15432_), .ZN(new_n15435_));
  AOI21_X1   g15243(.A1(new_n15435_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n15436_));
  AOI21_X1   g15244(.A1(new_n15436_), .A2(new_n15434_), .B(new_n15425_), .ZN(new_n15437_));
  AOI21_X1   g15245(.A1(new_n15434_), .A2(new_n15415_), .B(new_n1088_), .ZN(new_n15438_));
  OAI21_X1   g15246(.A1(new_n15437_), .A2(new_n15438_), .B(\asqrt[52] ), .ZN(new_n15439_));
  AOI21_X1   g15247(.A1(new_n15421_), .A2(new_n15439_), .B(new_n842_), .ZN(new_n15440_));
  NOR2_X1    g15248(.A1(new_n15424_), .A2(new_n15440_), .ZN(new_n15441_));
  AOI21_X1   g15249(.A1(new_n15441_), .A2(new_n720_), .B(new_n15012_), .ZN(new_n15442_));
  OAI21_X1   g15250(.A1(new_n15424_), .A2(new_n15440_), .B(\asqrt[54] ), .ZN(new_n15443_));
  NAND2_X1   g15251(.A1(new_n15443_), .A2(new_n630_), .ZN(new_n15444_));
  OAI21_X1   g15252(.A1(new_n15442_), .A2(new_n15444_), .B(new_n14968_), .ZN(new_n15445_));
  INV_X1     g15253(.I(new_n15443_), .ZN(new_n15446_));
  OAI21_X1   g15254(.A1(new_n15442_), .A2(new_n15446_), .B(\asqrt[55] ), .ZN(new_n15447_));
  NAND3_X1   g15255(.A1(new_n15445_), .A2(new_n15447_), .A3(new_n545_), .ZN(new_n15448_));
  NAND2_X1   g15256(.A1(new_n15448_), .A2(new_n15008_), .ZN(new_n15449_));
  NAND2_X1   g15257(.A1(new_n15445_), .A2(new_n15447_), .ZN(new_n15450_));
  AOI21_X1   g15258(.A1(new_n15450_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n15451_));
  AOI21_X1   g15259(.A1(new_n15451_), .A2(new_n15449_), .B(new_n15005_), .ZN(new_n15452_));
  INV_X1     g15260(.I(new_n14968_), .ZN(new_n15453_));
  INV_X1     g15261(.I(new_n15018_), .ZN(new_n15454_));
  NOR2_X1    g15262(.A1(new_n15437_), .A2(new_n15438_), .ZN(new_n15455_));
  AOI21_X1   g15263(.A1(new_n15455_), .A2(new_n962_), .B(new_n15454_), .ZN(new_n15456_));
  NAND2_X1   g15264(.A1(new_n15439_), .A2(new_n842_), .ZN(new_n15457_));
  OAI21_X1   g15265(.A1(new_n15456_), .A2(new_n15457_), .B(new_n15014_), .ZN(new_n15458_));
  INV_X1     g15266(.I(new_n15439_), .ZN(new_n15459_));
  OAI21_X1   g15267(.A1(new_n15456_), .A2(new_n15459_), .B(\asqrt[53] ), .ZN(new_n15460_));
  NAND3_X1   g15268(.A1(new_n15458_), .A2(new_n15460_), .A3(new_n720_), .ZN(new_n15461_));
  NAND2_X1   g15269(.A1(new_n15461_), .A2(new_n15011_), .ZN(new_n15462_));
  NAND2_X1   g15270(.A1(new_n15458_), .A2(new_n15460_), .ZN(new_n15463_));
  AOI21_X1   g15271(.A1(new_n15463_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n15464_));
  AOI21_X1   g15272(.A1(new_n15464_), .A2(new_n15462_), .B(new_n15453_), .ZN(new_n15465_));
  AOI21_X1   g15273(.A1(new_n15462_), .A2(new_n15443_), .B(new_n630_), .ZN(new_n15466_));
  OAI21_X1   g15274(.A1(new_n15465_), .A2(new_n15466_), .B(\asqrt[56] ), .ZN(new_n15467_));
  AOI21_X1   g15275(.A1(new_n15449_), .A2(new_n15467_), .B(new_n450_), .ZN(new_n15468_));
  NOR2_X1    g15276(.A1(new_n15452_), .A2(new_n15468_), .ZN(new_n15469_));
  AOI21_X1   g15277(.A1(new_n15469_), .A2(new_n403_), .B(new_n15002_), .ZN(new_n15470_));
  OAI21_X1   g15278(.A1(new_n15452_), .A2(new_n15468_), .B(\asqrt[58] ), .ZN(new_n15471_));
  NAND2_X1   g15279(.A1(new_n15471_), .A2(new_n339_), .ZN(new_n15472_));
  OAI21_X1   g15280(.A1(new_n15470_), .A2(new_n15472_), .B(new_n14998_), .ZN(new_n15473_));
  INV_X1     g15281(.I(new_n15471_), .ZN(new_n15474_));
  OAI21_X1   g15282(.A1(new_n15470_), .A2(new_n15474_), .B(\asqrt[59] ), .ZN(new_n15475_));
  NAND3_X1   g15283(.A1(new_n15473_), .A2(new_n15475_), .A3(new_n288_), .ZN(new_n15476_));
  NAND2_X1   g15284(.A1(new_n15476_), .A2(new_n14996_), .ZN(new_n15477_));
  INV_X1     g15285(.I(new_n14998_), .ZN(new_n15478_));
  INV_X1     g15286(.I(new_n15008_), .ZN(new_n15479_));
  NOR2_X1    g15287(.A1(new_n15465_), .A2(new_n15466_), .ZN(new_n15480_));
  AOI21_X1   g15288(.A1(new_n15480_), .A2(new_n545_), .B(new_n15479_), .ZN(new_n15481_));
  NAND2_X1   g15289(.A1(new_n15467_), .A2(new_n450_), .ZN(new_n15482_));
  OAI21_X1   g15290(.A1(new_n15481_), .A2(new_n15482_), .B(new_n15004_), .ZN(new_n15483_));
  INV_X1     g15291(.I(new_n15467_), .ZN(new_n15484_));
  OAI21_X1   g15292(.A1(new_n15481_), .A2(new_n15484_), .B(\asqrt[57] ), .ZN(new_n15485_));
  NAND3_X1   g15293(.A1(new_n15483_), .A2(new_n15485_), .A3(new_n403_), .ZN(new_n15486_));
  NAND2_X1   g15294(.A1(new_n15486_), .A2(new_n15001_), .ZN(new_n15487_));
  NAND2_X1   g15295(.A1(new_n15483_), .A2(new_n15485_), .ZN(new_n15488_));
  AOI21_X1   g15296(.A1(new_n15488_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n15489_));
  AOI21_X1   g15297(.A1(new_n15489_), .A2(new_n15487_), .B(new_n15478_), .ZN(new_n15490_));
  AOI21_X1   g15298(.A1(new_n15487_), .A2(new_n15471_), .B(new_n339_), .ZN(new_n15491_));
  OAI21_X1   g15299(.A1(new_n15490_), .A2(new_n15491_), .B(\asqrt[60] ), .ZN(new_n15492_));
  AOI21_X1   g15300(.A1(new_n15477_), .A2(new_n15492_), .B(new_n242_), .ZN(new_n15493_));
  NAND3_X1   g15301(.A1(\asqrt[10] ), .A2(new_n14928_), .A3(new_n14944_), .ZN(new_n15494_));
  XOR2_X1    g15302(.A1(new_n15494_), .A2(new_n14969_), .Z(new_n15495_));
  INV_X1     g15303(.I(new_n15495_), .ZN(new_n15496_));
  NAND2_X1   g15304(.A1(new_n15473_), .A2(new_n15475_), .ZN(new_n15497_));
  AOI21_X1   g15305(.A1(new_n15497_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n15498_));
  AOI21_X1   g15306(.A1(new_n15498_), .A2(new_n15477_), .B(new_n15496_), .ZN(new_n15499_));
  OAI21_X1   g15307(.A1(new_n15499_), .A2(new_n15493_), .B(\asqrt[62] ), .ZN(new_n15500_));
  AOI21_X1   g15308(.A1(new_n14929_), .A2(new_n14950_), .B(new_n14945_), .ZN(new_n15501_));
  NAND2_X1   g15309(.A1(\asqrt[10] ), .A2(new_n15501_), .ZN(new_n15502_));
  XOR2_X1    g15310(.A1(new_n15502_), .A2(new_n14948_), .Z(new_n15503_));
  INV_X1     g15311(.I(new_n14996_), .ZN(new_n15504_));
  NOR2_X1    g15312(.A1(new_n15490_), .A2(new_n15491_), .ZN(new_n15505_));
  AOI21_X1   g15313(.A1(new_n15505_), .A2(new_n288_), .B(new_n15504_), .ZN(new_n15506_));
  INV_X1     g15314(.I(new_n15492_), .ZN(new_n15507_));
  OAI21_X1   g15315(.A1(new_n15506_), .A2(new_n15507_), .B(\asqrt[61] ), .ZN(new_n15508_));
  NAND2_X1   g15316(.A1(new_n15492_), .A2(new_n242_), .ZN(new_n15509_));
  OAI21_X1   g15317(.A1(new_n15506_), .A2(new_n15509_), .B(new_n15495_), .ZN(new_n15510_));
  NAND3_X1   g15318(.A1(new_n15510_), .A2(new_n15508_), .A3(new_n234_), .ZN(new_n15511_));
  NAND2_X1   g15319(.A1(new_n15511_), .A2(new_n15503_), .ZN(new_n15512_));
  AOI21_X1   g15320(.A1(new_n15512_), .A2(new_n15500_), .B(new_n14993_), .ZN(new_n15513_));
  AOI21_X1   g15321(.A1(new_n15513_), .A2(new_n14991_), .B(\asqrt[63] ), .ZN(new_n15514_));
  NAND2_X1   g15322(.A1(new_n15512_), .A2(new_n15500_), .ZN(new_n15515_));
  NOR2_X1    g15323(.A1(new_n15515_), .A2(new_n14991_), .ZN(new_n15516_));
  NOR2_X1    g15324(.A1(\asqrt[10] ), .A2(new_n14980_), .ZN(new_n15517_));
  NOR4_X1    g15325(.A1(new_n15514_), .A2(new_n14988_), .A3(new_n15516_), .A4(new_n15517_), .ZN(new_n15518_));
  OAI21_X1   g15326(.A1(new_n15442_), .A2(new_n15444_), .B(new_n15447_), .ZN(new_n15519_));
  NOR2_X1    g15327(.A1(new_n15518_), .A2(new_n15519_), .ZN(new_n15520_));
  XOR2_X1    g15328(.A1(new_n15520_), .A2(new_n14968_), .Z(new_n15521_));
  INV_X1     g15329(.I(new_n15521_), .ZN(new_n15522_));
  INV_X1     g15330(.I(new_n14988_), .ZN(new_n15523_));
  INV_X1     g15331(.I(new_n15500_), .ZN(new_n15524_));
  NOR2_X1    g15332(.A1(new_n15499_), .A2(new_n15493_), .ZN(new_n15525_));
  INV_X1     g15333(.I(new_n15503_), .ZN(new_n15526_));
  AOI21_X1   g15334(.A1(new_n15525_), .A2(new_n234_), .B(new_n15526_), .ZN(new_n15527_));
  OAI21_X1   g15335(.A1(new_n15527_), .A2(new_n15524_), .B(new_n14992_), .ZN(new_n15528_));
  OAI21_X1   g15336(.A1(new_n15528_), .A2(new_n14990_), .B(new_n193_), .ZN(new_n15529_));
  NOR2_X1    g15337(.A1(new_n15527_), .A2(new_n15524_), .ZN(new_n15530_));
  NAND2_X1   g15338(.A1(new_n15530_), .A2(new_n14990_), .ZN(new_n15531_));
  INV_X1     g15339(.I(new_n15517_), .ZN(new_n15532_));
  NAND4_X1   g15340(.A1(new_n15529_), .A2(new_n15523_), .A3(new_n15531_), .A4(new_n15532_), .ZN(\asqrt[9] ));
  NAND3_X1   g15341(.A1(\asqrt[9] ), .A2(new_n15461_), .A3(new_n15443_), .ZN(new_n15534_));
  XOR2_X1    g15342(.A1(new_n15534_), .A2(new_n15012_), .Z(new_n15535_));
  OAI21_X1   g15343(.A1(new_n15456_), .A2(new_n15457_), .B(new_n15460_), .ZN(new_n15536_));
  NOR2_X1    g15344(.A1(new_n15518_), .A2(new_n15536_), .ZN(new_n15537_));
  XOR2_X1    g15345(.A1(new_n15537_), .A2(new_n15014_), .Z(new_n15538_));
  INV_X1     g15346(.I(new_n15538_), .ZN(new_n15539_));
  NAND3_X1   g15347(.A1(\asqrt[9] ), .A2(new_n15420_), .A3(new_n15439_), .ZN(new_n15540_));
  XOR2_X1    g15348(.A1(new_n15540_), .A2(new_n15454_), .Z(new_n15541_));
  INV_X1     g15349(.I(new_n15541_), .ZN(new_n15542_));
  OAI21_X1   g15350(.A1(new_n15414_), .A2(new_n15416_), .B(new_n15419_), .ZN(new_n15543_));
  NOR2_X1    g15351(.A1(new_n15518_), .A2(new_n15543_), .ZN(new_n15544_));
  XOR2_X1    g15352(.A1(new_n15544_), .A2(new_n15020_), .Z(new_n15545_));
  NAND3_X1   g15353(.A1(\asqrt[9] ), .A2(new_n15433_), .A3(new_n15415_), .ZN(new_n15546_));
  XOR2_X1    g15354(.A1(new_n15546_), .A2(new_n15024_), .Z(new_n15547_));
  OAI21_X1   g15355(.A1(new_n15428_), .A2(new_n15429_), .B(new_n15432_), .ZN(new_n15548_));
  NOR2_X1    g15356(.A1(new_n15518_), .A2(new_n15548_), .ZN(new_n15549_));
  XOR2_X1    g15357(.A1(new_n15549_), .A2(new_n15026_), .Z(new_n15550_));
  INV_X1     g15358(.I(new_n15550_), .ZN(new_n15551_));
  NAND3_X1   g15359(.A1(\asqrt[9] ), .A2(new_n15392_), .A3(new_n15411_), .ZN(new_n15552_));
  XOR2_X1    g15360(.A1(new_n15552_), .A2(new_n15426_), .Z(new_n15553_));
  INV_X1     g15361(.I(new_n15553_), .ZN(new_n15554_));
  OAI21_X1   g15362(.A1(new_n15386_), .A2(new_n15388_), .B(new_n15391_), .ZN(new_n15555_));
  NOR2_X1    g15363(.A1(new_n15518_), .A2(new_n15555_), .ZN(new_n15556_));
  XOR2_X1    g15364(.A1(new_n15556_), .A2(new_n15032_), .Z(new_n15557_));
  NAND3_X1   g15365(.A1(\asqrt[9] ), .A2(new_n15405_), .A3(new_n15387_), .ZN(new_n15558_));
  XOR2_X1    g15366(.A1(new_n15558_), .A2(new_n15036_), .Z(new_n15559_));
  OAI21_X1   g15367(.A1(new_n15400_), .A2(new_n15401_), .B(new_n15404_), .ZN(new_n15560_));
  NOR2_X1    g15368(.A1(new_n15518_), .A2(new_n15560_), .ZN(new_n15561_));
  XOR2_X1    g15369(.A1(new_n15561_), .A2(new_n15038_), .Z(new_n15562_));
  INV_X1     g15370(.I(new_n15562_), .ZN(new_n15563_));
  NAND3_X1   g15371(.A1(\asqrt[9] ), .A2(new_n15364_), .A3(new_n15383_), .ZN(new_n15564_));
  XOR2_X1    g15372(.A1(new_n15564_), .A2(new_n15398_), .Z(new_n15565_));
  INV_X1     g15373(.I(new_n15565_), .ZN(new_n15566_));
  OAI21_X1   g15374(.A1(new_n15358_), .A2(new_n15360_), .B(new_n15363_), .ZN(new_n15567_));
  NOR2_X1    g15375(.A1(new_n15518_), .A2(new_n15567_), .ZN(new_n15568_));
  XOR2_X1    g15376(.A1(new_n15568_), .A2(new_n15044_), .Z(new_n15569_));
  NAND3_X1   g15377(.A1(\asqrt[9] ), .A2(new_n15377_), .A3(new_n15359_), .ZN(new_n15570_));
  XOR2_X1    g15378(.A1(new_n15570_), .A2(new_n15048_), .Z(new_n15571_));
  OAI21_X1   g15379(.A1(new_n15372_), .A2(new_n15373_), .B(new_n15376_), .ZN(new_n15572_));
  NOR2_X1    g15380(.A1(new_n15518_), .A2(new_n15572_), .ZN(new_n15573_));
  XOR2_X1    g15381(.A1(new_n15573_), .A2(new_n15050_), .Z(new_n15574_));
  INV_X1     g15382(.I(new_n15574_), .ZN(new_n15575_));
  NAND3_X1   g15383(.A1(\asqrt[9] ), .A2(new_n15336_), .A3(new_n15355_), .ZN(new_n15576_));
  XOR2_X1    g15384(.A1(new_n15576_), .A2(new_n15370_), .Z(new_n15577_));
  INV_X1     g15385(.I(new_n15577_), .ZN(new_n15578_));
  OAI21_X1   g15386(.A1(new_n15330_), .A2(new_n15332_), .B(new_n15335_), .ZN(new_n15579_));
  NOR2_X1    g15387(.A1(new_n15518_), .A2(new_n15579_), .ZN(new_n15580_));
  XOR2_X1    g15388(.A1(new_n15580_), .A2(new_n15056_), .Z(new_n15581_));
  NAND3_X1   g15389(.A1(\asqrt[9] ), .A2(new_n15349_), .A3(new_n15331_), .ZN(new_n15582_));
  XOR2_X1    g15390(.A1(new_n15582_), .A2(new_n15060_), .Z(new_n15583_));
  OAI21_X1   g15391(.A1(new_n15344_), .A2(new_n15345_), .B(new_n15348_), .ZN(new_n15584_));
  NOR2_X1    g15392(.A1(new_n15518_), .A2(new_n15584_), .ZN(new_n15585_));
  XOR2_X1    g15393(.A1(new_n15585_), .A2(new_n15062_), .Z(new_n15586_));
  INV_X1     g15394(.I(new_n15586_), .ZN(new_n15587_));
  NAND3_X1   g15395(.A1(\asqrt[9] ), .A2(new_n15308_), .A3(new_n15327_), .ZN(new_n15588_));
  XOR2_X1    g15396(.A1(new_n15588_), .A2(new_n15342_), .Z(new_n15589_));
  INV_X1     g15397(.I(new_n15589_), .ZN(new_n15590_));
  OAI21_X1   g15398(.A1(new_n15302_), .A2(new_n15304_), .B(new_n15307_), .ZN(new_n15591_));
  NOR2_X1    g15399(.A1(new_n15518_), .A2(new_n15591_), .ZN(new_n15592_));
  XOR2_X1    g15400(.A1(new_n15592_), .A2(new_n15068_), .Z(new_n15593_));
  NAND3_X1   g15401(.A1(\asqrt[9] ), .A2(new_n15321_), .A3(new_n15303_), .ZN(new_n15594_));
  XOR2_X1    g15402(.A1(new_n15594_), .A2(new_n15072_), .Z(new_n15595_));
  OAI21_X1   g15403(.A1(new_n15316_), .A2(new_n15317_), .B(new_n15320_), .ZN(new_n15596_));
  NOR2_X1    g15404(.A1(new_n15518_), .A2(new_n15596_), .ZN(new_n15597_));
  XOR2_X1    g15405(.A1(new_n15597_), .A2(new_n15074_), .Z(new_n15598_));
  INV_X1     g15406(.I(new_n15598_), .ZN(new_n15599_));
  NAND3_X1   g15407(.A1(\asqrt[9] ), .A2(new_n15280_), .A3(new_n15299_), .ZN(new_n15600_));
  XOR2_X1    g15408(.A1(new_n15600_), .A2(new_n15314_), .Z(new_n15601_));
  INV_X1     g15409(.I(new_n15601_), .ZN(new_n15602_));
  OAI21_X1   g15410(.A1(new_n15274_), .A2(new_n15276_), .B(new_n15279_), .ZN(new_n15603_));
  NOR2_X1    g15411(.A1(new_n15518_), .A2(new_n15603_), .ZN(new_n15604_));
  XOR2_X1    g15412(.A1(new_n15604_), .A2(new_n15080_), .Z(new_n15605_));
  NAND3_X1   g15413(.A1(\asqrt[9] ), .A2(new_n15293_), .A3(new_n15275_), .ZN(new_n15606_));
  XOR2_X1    g15414(.A1(new_n15606_), .A2(new_n15084_), .Z(new_n15607_));
  OAI21_X1   g15415(.A1(new_n15288_), .A2(new_n15289_), .B(new_n15292_), .ZN(new_n15608_));
  NOR2_X1    g15416(.A1(new_n15518_), .A2(new_n15608_), .ZN(new_n15609_));
  XOR2_X1    g15417(.A1(new_n15609_), .A2(new_n15086_), .Z(new_n15610_));
  INV_X1     g15418(.I(new_n15610_), .ZN(new_n15611_));
  NAND3_X1   g15419(.A1(\asqrt[9] ), .A2(new_n15252_), .A3(new_n15271_), .ZN(new_n15612_));
  XOR2_X1    g15420(.A1(new_n15612_), .A2(new_n15286_), .Z(new_n15613_));
  INV_X1     g15421(.I(new_n15613_), .ZN(new_n15614_));
  OAI21_X1   g15422(.A1(new_n15246_), .A2(new_n15248_), .B(new_n15251_), .ZN(new_n15615_));
  NOR2_X1    g15423(.A1(new_n15518_), .A2(new_n15615_), .ZN(new_n15616_));
  XOR2_X1    g15424(.A1(new_n15616_), .A2(new_n15092_), .Z(new_n15617_));
  NAND3_X1   g15425(.A1(\asqrt[9] ), .A2(new_n15265_), .A3(new_n15247_), .ZN(new_n15618_));
  XOR2_X1    g15426(.A1(new_n15618_), .A2(new_n15096_), .Z(new_n15619_));
  OAI21_X1   g15427(.A1(new_n15260_), .A2(new_n15261_), .B(new_n15264_), .ZN(new_n15620_));
  NOR2_X1    g15428(.A1(new_n15518_), .A2(new_n15620_), .ZN(new_n15621_));
  XOR2_X1    g15429(.A1(new_n15621_), .A2(new_n15098_), .Z(new_n15622_));
  INV_X1     g15430(.I(new_n15622_), .ZN(new_n15623_));
  NAND3_X1   g15431(.A1(\asqrt[9] ), .A2(new_n15224_), .A3(new_n15243_), .ZN(new_n15624_));
  XOR2_X1    g15432(.A1(new_n15624_), .A2(new_n15258_), .Z(new_n15625_));
  INV_X1     g15433(.I(new_n15625_), .ZN(new_n15626_));
  OAI21_X1   g15434(.A1(new_n15218_), .A2(new_n15220_), .B(new_n15223_), .ZN(new_n15627_));
  NOR2_X1    g15435(.A1(new_n15518_), .A2(new_n15627_), .ZN(new_n15628_));
  XOR2_X1    g15436(.A1(new_n15628_), .A2(new_n15104_), .Z(new_n15629_));
  NAND3_X1   g15437(.A1(\asqrt[9] ), .A2(new_n15237_), .A3(new_n15219_), .ZN(new_n15630_));
  XOR2_X1    g15438(.A1(new_n15630_), .A2(new_n15108_), .Z(new_n15631_));
  OAI21_X1   g15439(.A1(new_n15232_), .A2(new_n15233_), .B(new_n15236_), .ZN(new_n15632_));
  NOR2_X1    g15440(.A1(new_n15518_), .A2(new_n15632_), .ZN(new_n15633_));
  XOR2_X1    g15441(.A1(new_n15633_), .A2(new_n15110_), .Z(new_n15634_));
  INV_X1     g15442(.I(new_n15634_), .ZN(new_n15635_));
  NAND3_X1   g15443(.A1(\asqrt[9] ), .A2(new_n15196_), .A3(new_n15215_), .ZN(new_n15636_));
  XOR2_X1    g15444(.A1(new_n15636_), .A2(new_n15230_), .Z(new_n15637_));
  INV_X1     g15445(.I(new_n15637_), .ZN(new_n15638_));
  OAI21_X1   g15446(.A1(new_n15190_), .A2(new_n15192_), .B(new_n15195_), .ZN(new_n15639_));
  NOR2_X1    g15447(.A1(new_n15518_), .A2(new_n15639_), .ZN(new_n15640_));
  XOR2_X1    g15448(.A1(new_n15640_), .A2(new_n15116_), .Z(new_n15641_));
  NAND3_X1   g15449(.A1(\asqrt[9] ), .A2(new_n15209_), .A3(new_n15191_), .ZN(new_n15642_));
  XOR2_X1    g15450(.A1(new_n15642_), .A2(new_n15120_), .Z(new_n15643_));
  OAI21_X1   g15451(.A1(new_n15204_), .A2(new_n15205_), .B(new_n15208_), .ZN(new_n15644_));
  NOR2_X1    g15452(.A1(new_n15518_), .A2(new_n15644_), .ZN(new_n15645_));
  XOR2_X1    g15453(.A1(new_n15645_), .A2(new_n15122_), .Z(new_n15646_));
  INV_X1     g15454(.I(new_n15646_), .ZN(new_n15647_));
  NAND3_X1   g15455(.A1(\asqrt[9] ), .A2(new_n15161_), .A3(new_n15187_), .ZN(new_n15648_));
  XOR2_X1    g15456(.A1(new_n15648_), .A2(new_n15202_), .Z(new_n15649_));
  INV_X1     g15457(.I(new_n15649_), .ZN(new_n15650_));
  AOI21_X1   g15458(.A1(new_n15182_), .A2(new_n15183_), .B(new_n15186_), .ZN(new_n15651_));
  NAND2_X1   g15459(.A1(\asqrt[9] ), .A2(new_n15651_), .ZN(new_n15652_));
  XOR2_X1    g15460(.A1(new_n15652_), .A2(new_n15166_), .Z(new_n15653_));
  NOR2_X1    g15461(.A1(new_n15181_), .A2(\asqrt[14] ), .ZN(new_n15654_));
  NOR3_X1    g15462(.A1(new_n15518_), .A2(new_n15654_), .A3(new_n15159_), .ZN(new_n15655_));
  XOR2_X1    g15463(.A1(new_n15655_), .A2(new_n15131_), .Z(new_n15656_));
  NOR3_X1    g15464(.A1(new_n15518_), .A2(new_n15178_), .A3(new_n15154_), .ZN(new_n15657_));
  XOR2_X1    g15465(.A1(new_n15657_), .A2(new_n15153_), .Z(new_n15658_));
  INV_X1     g15466(.I(new_n15658_), .ZN(new_n15659_));
  NOR2_X1    g15467(.A1(new_n15148_), .A2(\asqrt[12] ), .ZN(new_n15660_));
  NOR3_X1    g15468(.A1(new_n15518_), .A2(new_n15660_), .A3(new_n15177_), .ZN(new_n15661_));
  XOR2_X1    g15469(.A1(new_n15661_), .A2(new_n15139_), .Z(new_n15662_));
  INV_X1     g15470(.I(new_n15662_), .ZN(new_n15663_));
  NAND3_X1   g15471(.A1(\asqrt[9] ), .A2(new_n15140_), .A3(new_n15141_), .ZN(new_n15664_));
  NOR4_X1    g15472(.A1(new_n15514_), .A2(new_n14985_), .A3(new_n14988_), .A4(new_n15516_), .ZN(new_n15665_));
  INV_X1     g15473(.I(new_n15665_), .ZN(new_n15666_));
  AOI21_X1   g15474(.A1(new_n15664_), .A2(new_n15666_), .B(\a[20] ), .ZN(new_n15667_));
  NOR3_X1    g15475(.A1(new_n15518_), .A2(\a[18] ), .A3(\a[19] ), .ZN(new_n15668_));
  NOR3_X1    g15476(.A1(new_n15668_), .A2(new_n14571_), .A3(new_n15665_), .ZN(new_n15669_));
  NOR2_X1    g15477(.A1(new_n15669_), .A2(new_n15667_), .ZN(new_n15670_));
  INV_X1     g15478(.I(\a[16] ), .ZN(new_n15671_));
  INV_X1     g15479(.I(\a[17] ), .ZN(new_n15672_));
  NAND3_X1   g15480(.A1(new_n15671_), .A2(new_n15672_), .A3(new_n15140_), .ZN(new_n15673_));
  OAI21_X1   g15481(.A1(new_n15518_), .A2(new_n15140_), .B(new_n15673_), .ZN(new_n15674_));
  NAND2_X1   g15482(.A1(new_n15674_), .A2(\asqrt[10] ), .ZN(new_n15675_));
  OAI21_X1   g15483(.A1(new_n15518_), .A2(\a[18] ), .B(\a[19] ), .ZN(new_n15676_));
  NAND2_X1   g15484(.A1(new_n15676_), .A2(new_n15664_), .ZN(new_n15677_));
  NOR2_X1    g15485(.A1(new_n15674_), .A2(\asqrt[10] ), .ZN(new_n15678_));
  OAI21_X1   g15486(.A1(new_n15677_), .A2(new_n15678_), .B(new_n15675_), .ZN(new_n15679_));
  OAI21_X1   g15487(.A1(\asqrt[11] ), .A2(new_n15679_), .B(new_n15670_), .ZN(new_n15680_));
  NAND2_X1   g15488(.A1(new_n15679_), .A2(\asqrt[11] ), .ZN(new_n15681_));
  NAND3_X1   g15489(.A1(new_n15680_), .A2(new_n13917_), .A3(new_n15681_), .ZN(new_n15682_));
  NOR3_X1    g15490(.A1(new_n15518_), .A2(new_n15171_), .A3(new_n15147_), .ZN(new_n15683_));
  XOR2_X1    g15491(.A1(new_n15683_), .A2(new_n15173_), .Z(new_n15684_));
  NAND2_X1   g15492(.A1(new_n15682_), .A2(new_n15684_), .ZN(new_n15685_));
  NAND2_X1   g15493(.A1(new_n15680_), .A2(new_n15681_), .ZN(new_n15686_));
  AOI21_X1   g15494(.A1(new_n15686_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n15687_));
  AOI21_X1   g15495(.A1(new_n15687_), .A2(new_n15685_), .B(new_n15663_), .ZN(new_n15688_));
  OAI21_X1   g15496(.A1(new_n15668_), .A2(new_n15665_), .B(new_n14571_), .ZN(new_n15689_));
  NAND3_X1   g15497(.A1(new_n15664_), .A2(\a[20] ), .A3(new_n15666_), .ZN(new_n15690_));
  NAND2_X1   g15498(.A1(new_n15689_), .A2(new_n15690_), .ZN(new_n15691_));
  NAND2_X1   g15499(.A1(\asqrt[9] ), .A2(\a[18] ), .ZN(new_n15692_));
  AOI21_X1   g15500(.A1(new_n15692_), .A2(new_n15673_), .B(new_n14985_), .ZN(new_n15693_));
  AOI21_X1   g15501(.A1(\asqrt[9] ), .A2(new_n15140_), .B(new_n15141_), .ZN(new_n15694_));
  NOR2_X1    g15502(.A1(new_n15694_), .A2(new_n15668_), .ZN(new_n15695_));
  NAND3_X1   g15503(.A1(new_n15692_), .A2(new_n14985_), .A3(new_n15673_), .ZN(new_n15696_));
  AOI21_X1   g15504(.A1(new_n15695_), .A2(new_n15696_), .B(new_n15693_), .ZN(new_n15697_));
  AOI21_X1   g15505(.A1(new_n15697_), .A2(new_n14430_), .B(new_n15691_), .ZN(new_n15698_));
  NOR2_X1    g15506(.A1(new_n15697_), .A2(new_n14430_), .ZN(new_n15699_));
  OAI21_X1   g15507(.A1(new_n15698_), .A2(new_n15699_), .B(\asqrt[12] ), .ZN(new_n15700_));
  AOI21_X1   g15508(.A1(new_n15685_), .A2(new_n15700_), .B(new_n13382_), .ZN(new_n15701_));
  NOR2_X1    g15509(.A1(new_n15688_), .A2(new_n15701_), .ZN(new_n15702_));
  AOI21_X1   g15510(.A1(new_n15702_), .A2(new_n12889_), .B(new_n15659_), .ZN(new_n15703_));
  OAI21_X1   g15511(.A1(new_n15688_), .A2(new_n15701_), .B(\asqrt[14] ), .ZN(new_n15704_));
  NAND2_X1   g15512(.A1(new_n15704_), .A2(new_n12374_), .ZN(new_n15705_));
  OAI21_X1   g15513(.A1(new_n15703_), .A2(new_n15705_), .B(new_n15656_), .ZN(new_n15706_));
  INV_X1     g15514(.I(new_n15704_), .ZN(new_n15707_));
  OAI21_X1   g15515(.A1(new_n15703_), .A2(new_n15707_), .B(\asqrt[15] ), .ZN(new_n15708_));
  NAND3_X1   g15516(.A1(new_n15706_), .A2(new_n15708_), .A3(new_n11901_), .ZN(new_n15709_));
  NAND2_X1   g15517(.A1(new_n15709_), .A2(new_n15653_), .ZN(new_n15710_));
  NAND2_X1   g15518(.A1(new_n15706_), .A2(new_n15708_), .ZN(new_n15711_));
  AOI21_X1   g15519(.A1(new_n15711_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n15712_));
  AOI21_X1   g15520(.A1(new_n15712_), .A2(new_n15710_), .B(new_n15650_), .ZN(new_n15713_));
  INV_X1     g15521(.I(new_n15656_), .ZN(new_n15714_));
  NOR2_X1    g15522(.A1(new_n15698_), .A2(new_n15699_), .ZN(new_n15715_));
  INV_X1     g15523(.I(new_n15684_), .ZN(new_n15716_));
  AOI21_X1   g15524(.A1(new_n15715_), .A2(new_n13917_), .B(new_n15716_), .ZN(new_n15717_));
  NAND2_X1   g15525(.A1(new_n15700_), .A2(new_n13382_), .ZN(new_n15718_));
  OAI21_X1   g15526(.A1(new_n15717_), .A2(new_n15718_), .B(new_n15662_), .ZN(new_n15719_));
  INV_X1     g15527(.I(new_n15700_), .ZN(new_n15720_));
  OAI21_X1   g15528(.A1(new_n15717_), .A2(new_n15720_), .B(\asqrt[13] ), .ZN(new_n15721_));
  NAND3_X1   g15529(.A1(new_n15719_), .A2(new_n15721_), .A3(new_n12889_), .ZN(new_n15722_));
  NAND2_X1   g15530(.A1(new_n15722_), .A2(new_n15658_), .ZN(new_n15723_));
  NAND2_X1   g15531(.A1(new_n15719_), .A2(new_n15721_), .ZN(new_n15724_));
  AOI21_X1   g15532(.A1(new_n15724_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n15725_));
  AOI21_X1   g15533(.A1(new_n15725_), .A2(new_n15723_), .B(new_n15714_), .ZN(new_n15726_));
  AOI21_X1   g15534(.A1(new_n15723_), .A2(new_n15704_), .B(new_n12374_), .ZN(new_n15727_));
  OAI21_X1   g15535(.A1(new_n15726_), .A2(new_n15727_), .B(\asqrt[16] ), .ZN(new_n15728_));
  AOI21_X1   g15536(.A1(new_n15710_), .A2(new_n15728_), .B(new_n11406_), .ZN(new_n15729_));
  NOR2_X1    g15537(.A1(new_n15713_), .A2(new_n15729_), .ZN(new_n15730_));
  AOI21_X1   g15538(.A1(new_n15730_), .A2(new_n10953_), .B(new_n15647_), .ZN(new_n15731_));
  OAI21_X1   g15539(.A1(new_n15713_), .A2(new_n15729_), .B(\asqrt[18] ), .ZN(new_n15732_));
  NAND2_X1   g15540(.A1(new_n15732_), .A2(new_n10478_), .ZN(new_n15733_));
  OAI21_X1   g15541(.A1(new_n15731_), .A2(new_n15733_), .B(new_n15643_), .ZN(new_n15734_));
  INV_X1     g15542(.I(new_n15732_), .ZN(new_n15735_));
  OAI21_X1   g15543(.A1(new_n15731_), .A2(new_n15735_), .B(\asqrt[19] ), .ZN(new_n15736_));
  NAND3_X1   g15544(.A1(new_n15734_), .A2(new_n15736_), .A3(new_n10045_), .ZN(new_n15737_));
  NAND2_X1   g15545(.A1(new_n15737_), .A2(new_n15641_), .ZN(new_n15738_));
  NAND2_X1   g15546(.A1(new_n15734_), .A2(new_n15736_), .ZN(new_n15739_));
  AOI21_X1   g15547(.A1(new_n15739_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n15740_));
  AOI21_X1   g15548(.A1(new_n15740_), .A2(new_n15738_), .B(new_n15638_), .ZN(new_n15741_));
  INV_X1     g15549(.I(new_n15643_), .ZN(new_n15742_));
  INV_X1     g15550(.I(new_n15653_), .ZN(new_n15743_));
  NOR2_X1    g15551(.A1(new_n15726_), .A2(new_n15727_), .ZN(new_n15744_));
  AOI21_X1   g15552(.A1(new_n15744_), .A2(new_n11901_), .B(new_n15743_), .ZN(new_n15745_));
  NAND2_X1   g15553(.A1(new_n15728_), .A2(new_n11406_), .ZN(new_n15746_));
  OAI21_X1   g15554(.A1(new_n15745_), .A2(new_n15746_), .B(new_n15649_), .ZN(new_n15747_));
  INV_X1     g15555(.I(new_n15728_), .ZN(new_n15748_));
  OAI21_X1   g15556(.A1(new_n15745_), .A2(new_n15748_), .B(\asqrt[17] ), .ZN(new_n15749_));
  NAND3_X1   g15557(.A1(new_n15747_), .A2(new_n15749_), .A3(new_n10953_), .ZN(new_n15750_));
  NAND2_X1   g15558(.A1(new_n15750_), .A2(new_n15646_), .ZN(new_n15751_));
  NAND2_X1   g15559(.A1(new_n15747_), .A2(new_n15749_), .ZN(new_n15752_));
  AOI21_X1   g15560(.A1(new_n15752_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n15753_));
  AOI21_X1   g15561(.A1(new_n15753_), .A2(new_n15751_), .B(new_n15742_), .ZN(new_n15754_));
  AOI21_X1   g15562(.A1(new_n15751_), .A2(new_n15732_), .B(new_n10478_), .ZN(new_n15755_));
  OAI21_X1   g15563(.A1(new_n15754_), .A2(new_n15755_), .B(\asqrt[20] ), .ZN(new_n15756_));
  AOI21_X1   g15564(.A1(new_n15738_), .A2(new_n15756_), .B(new_n9590_), .ZN(new_n15757_));
  NOR2_X1    g15565(.A1(new_n15741_), .A2(new_n15757_), .ZN(new_n15758_));
  AOI21_X1   g15566(.A1(new_n15758_), .A2(new_n9177_), .B(new_n15635_), .ZN(new_n15759_));
  OAI21_X1   g15567(.A1(new_n15741_), .A2(new_n15757_), .B(\asqrt[22] ), .ZN(new_n15760_));
  NAND2_X1   g15568(.A1(new_n15760_), .A2(new_n8742_), .ZN(new_n15761_));
  OAI21_X1   g15569(.A1(new_n15759_), .A2(new_n15761_), .B(new_n15631_), .ZN(new_n15762_));
  INV_X1     g15570(.I(new_n15760_), .ZN(new_n15763_));
  OAI21_X1   g15571(.A1(new_n15759_), .A2(new_n15763_), .B(\asqrt[23] ), .ZN(new_n15764_));
  NAND3_X1   g15572(.A1(new_n15762_), .A2(new_n15764_), .A3(new_n8349_), .ZN(new_n15765_));
  NAND2_X1   g15573(.A1(new_n15765_), .A2(new_n15629_), .ZN(new_n15766_));
  NAND2_X1   g15574(.A1(new_n15762_), .A2(new_n15764_), .ZN(new_n15767_));
  AOI21_X1   g15575(.A1(new_n15767_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n15768_));
  AOI21_X1   g15576(.A1(new_n15768_), .A2(new_n15766_), .B(new_n15626_), .ZN(new_n15769_));
  INV_X1     g15577(.I(new_n15631_), .ZN(new_n15770_));
  INV_X1     g15578(.I(new_n15641_), .ZN(new_n15771_));
  NOR2_X1    g15579(.A1(new_n15754_), .A2(new_n15755_), .ZN(new_n15772_));
  AOI21_X1   g15580(.A1(new_n15772_), .A2(new_n10045_), .B(new_n15771_), .ZN(new_n15773_));
  NAND2_X1   g15581(.A1(new_n15756_), .A2(new_n9590_), .ZN(new_n15774_));
  OAI21_X1   g15582(.A1(new_n15773_), .A2(new_n15774_), .B(new_n15637_), .ZN(new_n15775_));
  INV_X1     g15583(.I(new_n15756_), .ZN(new_n15776_));
  OAI21_X1   g15584(.A1(new_n15773_), .A2(new_n15776_), .B(\asqrt[21] ), .ZN(new_n15777_));
  NAND3_X1   g15585(.A1(new_n15775_), .A2(new_n15777_), .A3(new_n9177_), .ZN(new_n15778_));
  NAND2_X1   g15586(.A1(new_n15778_), .A2(new_n15634_), .ZN(new_n15779_));
  NAND2_X1   g15587(.A1(new_n15775_), .A2(new_n15777_), .ZN(new_n15780_));
  AOI21_X1   g15588(.A1(new_n15780_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n15781_));
  AOI21_X1   g15589(.A1(new_n15781_), .A2(new_n15779_), .B(new_n15770_), .ZN(new_n15782_));
  AOI21_X1   g15590(.A1(new_n15779_), .A2(new_n15760_), .B(new_n8742_), .ZN(new_n15783_));
  OAI21_X1   g15591(.A1(new_n15782_), .A2(new_n15783_), .B(\asqrt[24] ), .ZN(new_n15784_));
  AOI21_X1   g15592(.A1(new_n15766_), .A2(new_n15784_), .B(new_n7934_), .ZN(new_n15785_));
  NOR2_X1    g15593(.A1(new_n15769_), .A2(new_n15785_), .ZN(new_n15786_));
  AOI21_X1   g15594(.A1(new_n15786_), .A2(new_n7561_), .B(new_n15623_), .ZN(new_n15787_));
  OAI21_X1   g15595(.A1(new_n15769_), .A2(new_n15785_), .B(\asqrt[26] ), .ZN(new_n15788_));
  NAND2_X1   g15596(.A1(new_n15788_), .A2(new_n7166_), .ZN(new_n15789_));
  OAI21_X1   g15597(.A1(new_n15787_), .A2(new_n15789_), .B(new_n15619_), .ZN(new_n15790_));
  INV_X1     g15598(.I(new_n15788_), .ZN(new_n15791_));
  OAI21_X1   g15599(.A1(new_n15787_), .A2(new_n15791_), .B(\asqrt[27] ), .ZN(new_n15792_));
  NAND3_X1   g15600(.A1(new_n15790_), .A2(new_n15792_), .A3(new_n6813_), .ZN(new_n15793_));
  NAND2_X1   g15601(.A1(new_n15793_), .A2(new_n15617_), .ZN(new_n15794_));
  NAND2_X1   g15602(.A1(new_n15790_), .A2(new_n15792_), .ZN(new_n15795_));
  AOI21_X1   g15603(.A1(new_n15795_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n15796_));
  AOI21_X1   g15604(.A1(new_n15796_), .A2(new_n15794_), .B(new_n15614_), .ZN(new_n15797_));
  INV_X1     g15605(.I(new_n15619_), .ZN(new_n15798_));
  INV_X1     g15606(.I(new_n15629_), .ZN(new_n15799_));
  NOR2_X1    g15607(.A1(new_n15782_), .A2(new_n15783_), .ZN(new_n15800_));
  AOI21_X1   g15608(.A1(new_n15800_), .A2(new_n8349_), .B(new_n15799_), .ZN(new_n15801_));
  NAND2_X1   g15609(.A1(new_n15784_), .A2(new_n7934_), .ZN(new_n15802_));
  OAI21_X1   g15610(.A1(new_n15801_), .A2(new_n15802_), .B(new_n15625_), .ZN(new_n15803_));
  INV_X1     g15611(.I(new_n15784_), .ZN(new_n15804_));
  OAI21_X1   g15612(.A1(new_n15801_), .A2(new_n15804_), .B(\asqrt[25] ), .ZN(new_n15805_));
  NAND3_X1   g15613(.A1(new_n15803_), .A2(new_n15805_), .A3(new_n7561_), .ZN(new_n15806_));
  NAND2_X1   g15614(.A1(new_n15806_), .A2(new_n15622_), .ZN(new_n15807_));
  NAND2_X1   g15615(.A1(new_n15803_), .A2(new_n15805_), .ZN(new_n15808_));
  AOI21_X1   g15616(.A1(new_n15808_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n15809_));
  AOI21_X1   g15617(.A1(new_n15809_), .A2(new_n15807_), .B(new_n15798_), .ZN(new_n15810_));
  AOI21_X1   g15618(.A1(new_n15807_), .A2(new_n15788_), .B(new_n7166_), .ZN(new_n15811_));
  OAI21_X1   g15619(.A1(new_n15810_), .A2(new_n15811_), .B(\asqrt[28] ), .ZN(new_n15812_));
  AOI21_X1   g15620(.A1(new_n15794_), .A2(new_n15812_), .B(new_n6454_), .ZN(new_n15813_));
  NOR2_X1    g15621(.A1(new_n15797_), .A2(new_n15813_), .ZN(new_n15814_));
  AOI21_X1   g15622(.A1(new_n15814_), .A2(new_n6106_), .B(new_n15611_), .ZN(new_n15815_));
  OAI21_X1   g15623(.A1(new_n15797_), .A2(new_n15813_), .B(\asqrt[30] ), .ZN(new_n15816_));
  NAND2_X1   g15624(.A1(new_n15816_), .A2(new_n5750_), .ZN(new_n15817_));
  OAI21_X1   g15625(.A1(new_n15815_), .A2(new_n15817_), .B(new_n15607_), .ZN(new_n15818_));
  INV_X1     g15626(.I(new_n15816_), .ZN(new_n15819_));
  OAI21_X1   g15627(.A1(new_n15815_), .A2(new_n15819_), .B(\asqrt[31] ), .ZN(new_n15820_));
  NAND3_X1   g15628(.A1(new_n15818_), .A2(new_n15820_), .A3(new_n5435_), .ZN(new_n15821_));
  NAND2_X1   g15629(.A1(new_n15821_), .A2(new_n15605_), .ZN(new_n15822_));
  NAND2_X1   g15630(.A1(new_n15818_), .A2(new_n15820_), .ZN(new_n15823_));
  AOI21_X1   g15631(.A1(new_n15823_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n15824_));
  AOI21_X1   g15632(.A1(new_n15824_), .A2(new_n15822_), .B(new_n15602_), .ZN(new_n15825_));
  INV_X1     g15633(.I(new_n15607_), .ZN(new_n15826_));
  INV_X1     g15634(.I(new_n15617_), .ZN(new_n15827_));
  NOR2_X1    g15635(.A1(new_n15810_), .A2(new_n15811_), .ZN(new_n15828_));
  AOI21_X1   g15636(.A1(new_n15828_), .A2(new_n6813_), .B(new_n15827_), .ZN(new_n15829_));
  NAND2_X1   g15637(.A1(new_n15812_), .A2(new_n6454_), .ZN(new_n15830_));
  OAI21_X1   g15638(.A1(new_n15829_), .A2(new_n15830_), .B(new_n15613_), .ZN(new_n15831_));
  INV_X1     g15639(.I(new_n15812_), .ZN(new_n15832_));
  OAI21_X1   g15640(.A1(new_n15829_), .A2(new_n15832_), .B(\asqrt[29] ), .ZN(new_n15833_));
  NAND3_X1   g15641(.A1(new_n15831_), .A2(new_n15833_), .A3(new_n6106_), .ZN(new_n15834_));
  NAND2_X1   g15642(.A1(new_n15834_), .A2(new_n15610_), .ZN(new_n15835_));
  NAND2_X1   g15643(.A1(new_n15831_), .A2(new_n15833_), .ZN(new_n15836_));
  AOI21_X1   g15644(.A1(new_n15836_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n15837_));
  AOI21_X1   g15645(.A1(new_n15837_), .A2(new_n15835_), .B(new_n15826_), .ZN(new_n15838_));
  AOI21_X1   g15646(.A1(new_n15835_), .A2(new_n15816_), .B(new_n5750_), .ZN(new_n15839_));
  OAI21_X1   g15647(.A1(new_n15838_), .A2(new_n15839_), .B(\asqrt[32] ), .ZN(new_n15840_));
  AOI21_X1   g15648(.A1(new_n15822_), .A2(new_n15840_), .B(new_n5110_), .ZN(new_n15841_));
  NOR2_X1    g15649(.A1(new_n15825_), .A2(new_n15841_), .ZN(new_n15842_));
  AOI21_X1   g15650(.A1(new_n15842_), .A2(new_n4810_), .B(new_n15599_), .ZN(new_n15843_));
  OAI21_X1   g15651(.A1(new_n15825_), .A2(new_n15841_), .B(\asqrt[34] ), .ZN(new_n15844_));
  NAND2_X1   g15652(.A1(new_n15844_), .A2(new_n4510_), .ZN(new_n15845_));
  OAI21_X1   g15653(.A1(new_n15843_), .A2(new_n15845_), .B(new_n15595_), .ZN(new_n15846_));
  INV_X1     g15654(.I(new_n15844_), .ZN(new_n15847_));
  OAI21_X1   g15655(.A1(new_n15843_), .A2(new_n15847_), .B(\asqrt[35] ), .ZN(new_n15848_));
  NAND3_X1   g15656(.A1(new_n15846_), .A2(new_n15848_), .A3(new_n4224_), .ZN(new_n15849_));
  NAND2_X1   g15657(.A1(new_n15849_), .A2(new_n15593_), .ZN(new_n15850_));
  NAND2_X1   g15658(.A1(new_n15846_), .A2(new_n15848_), .ZN(new_n15851_));
  AOI21_X1   g15659(.A1(new_n15851_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n15852_));
  AOI21_X1   g15660(.A1(new_n15852_), .A2(new_n15850_), .B(new_n15590_), .ZN(new_n15853_));
  INV_X1     g15661(.I(new_n15595_), .ZN(new_n15854_));
  INV_X1     g15662(.I(new_n15605_), .ZN(new_n15855_));
  NOR2_X1    g15663(.A1(new_n15838_), .A2(new_n15839_), .ZN(new_n15856_));
  AOI21_X1   g15664(.A1(new_n15856_), .A2(new_n5435_), .B(new_n15855_), .ZN(new_n15857_));
  NAND2_X1   g15665(.A1(new_n15840_), .A2(new_n5110_), .ZN(new_n15858_));
  OAI21_X1   g15666(.A1(new_n15857_), .A2(new_n15858_), .B(new_n15601_), .ZN(new_n15859_));
  INV_X1     g15667(.I(new_n15840_), .ZN(new_n15860_));
  OAI21_X1   g15668(.A1(new_n15857_), .A2(new_n15860_), .B(\asqrt[33] ), .ZN(new_n15861_));
  NAND3_X1   g15669(.A1(new_n15859_), .A2(new_n15861_), .A3(new_n4810_), .ZN(new_n15862_));
  NAND2_X1   g15670(.A1(new_n15862_), .A2(new_n15598_), .ZN(new_n15863_));
  NAND2_X1   g15671(.A1(new_n15859_), .A2(new_n15861_), .ZN(new_n15864_));
  AOI21_X1   g15672(.A1(new_n15864_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n15865_));
  AOI21_X1   g15673(.A1(new_n15865_), .A2(new_n15863_), .B(new_n15854_), .ZN(new_n15866_));
  AOI21_X1   g15674(.A1(new_n15863_), .A2(new_n15844_), .B(new_n4510_), .ZN(new_n15867_));
  OAI21_X1   g15675(.A1(new_n15866_), .A2(new_n15867_), .B(\asqrt[36] ), .ZN(new_n15868_));
  AOI21_X1   g15676(.A1(new_n15850_), .A2(new_n15868_), .B(new_n3928_), .ZN(new_n15869_));
  NOR2_X1    g15677(.A1(new_n15853_), .A2(new_n15869_), .ZN(new_n15870_));
  AOI21_X1   g15678(.A1(new_n15870_), .A2(new_n3675_), .B(new_n15587_), .ZN(new_n15871_));
  OAI21_X1   g15679(.A1(new_n15853_), .A2(new_n15869_), .B(\asqrt[38] ), .ZN(new_n15872_));
  NAND2_X1   g15680(.A1(new_n15872_), .A2(new_n3400_), .ZN(new_n15873_));
  OAI21_X1   g15681(.A1(new_n15871_), .A2(new_n15873_), .B(new_n15583_), .ZN(new_n15874_));
  INV_X1     g15682(.I(new_n15872_), .ZN(new_n15875_));
  OAI21_X1   g15683(.A1(new_n15871_), .A2(new_n15875_), .B(\asqrt[39] ), .ZN(new_n15876_));
  NAND3_X1   g15684(.A1(new_n15874_), .A2(new_n15876_), .A3(new_n3167_), .ZN(new_n15877_));
  NAND2_X1   g15685(.A1(new_n15877_), .A2(new_n15581_), .ZN(new_n15878_));
  NAND2_X1   g15686(.A1(new_n15874_), .A2(new_n15876_), .ZN(new_n15879_));
  AOI21_X1   g15687(.A1(new_n15879_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n15880_));
  AOI21_X1   g15688(.A1(new_n15880_), .A2(new_n15878_), .B(new_n15578_), .ZN(new_n15881_));
  INV_X1     g15689(.I(new_n15583_), .ZN(new_n15882_));
  INV_X1     g15690(.I(new_n15593_), .ZN(new_n15883_));
  NOR2_X1    g15691(.A1(new_n15866_), .A2(new_n15867_), .ZN(new_n15884_));
  AOI21_X1   g15692(.A1(new_n15884_), .A2(new_n4224_), .B(new_n15883_), .ZN(new_n15885_));
  NAND2_X1   g15693(.A1(new_n15868_), .A2(new_n3928_), .ZN(new_n15886_));
  OAI21_X1   g15694(.A1(new_n15885_), .A2(new_n15886_), .B(new_n15589_), .ZN(new_n15887_));
  INV_X1     g15695(.I(new_n15868_), .ZN(new_n15888_));
  OAI21_X1   g15696(.A1(new_n15885_), .A2(new_n15888_), .B(\asqrt[37] ), .ZN(new_n15889_));
  NAND3_X1   g15697(.A1(new_n15887_), .A2(new_n15889_), .A3(new_n3675_), .ZN(new_n15890_));
  NAND2_X1   g15698(.A1(new_n15890_), .A2(new_n15586_), .ZN(new_n15891_));
  NAND2_X1   g15699(.A1(new_n15887_), .A2(new_n15889_), .ZN(new_n15892_));
  AOI21_X1   g15700(.A1(new_n15892_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n15893_));
  AOI21_X1   g15701(.A1(new_n15893_), .A2(new_n15891_), .B(new_n15882_), .ZN(new_n15894_));
  AOI21_X1   g15702(.A1(new_n15891_), .A2(new_n15872_), .B(new_n3400_), .ZN(new_n15895_));
  OAI21_X1   g15703(.A1(new_n15894_), .A2(new_n15895_), .B(\asqrt[40] ), .ZN(new_n15896_));
  AOI21_X1   g15704(.A1(new_n15878_), .A2(new_n15896_), .B(new_n2912_), .ZN(new_n15897_));
  NOR2_X1    g15705(.A1(new_n15881_), .A2(new_n15897_), .ZN(new_n15898_));
  AOI21_X1   g15706(.A1(new_n15898_), .A2(new_n2699_), .B(new_n15575_), .ZN(new_n15899_));
  OAI21_X1   g15707(.A1(new_n15881_), .A2(new_n15897_), .B(\asqrt[42] ), .ZN(new_n15900_));
  NAND2_X1   g15708(.A1(new_n15900_), .A2(new_n2464_), .ZN(new_n15901_));
  OAI21_X1   g15709(.A1(new_n15899_), .A2(new_n15901_), .B(new_n15571_), .ZN(new_n15902_));
  INV_X1     g15710(.I(new_n15900_), .ZN(new_n15903_));
  OAI21_X1   g15711(.A1(new_n15899_), .A2(new_n15903_), .B(\asqrt[43] ), .ZN(new_n15904_));
  NAND3_X1   g15712(.A1(new_n15902_), .A2(new_n15904_), .A3(new_n2271_), .ZN(new_n15905_));
  NAND2_X1   g15713(.A1(new_n15905_), .A2(new_n15569_), .ZN(new_n15906_));
  NAND2_X1   g15714(.A1(new_n15902_), .A2(new_n15904_), .ZN(new_n15907_));
  AOI21_X1   g15715(.A1(new_n15907_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n15908_));
  AOI21_X1   g15716(.A1(new_n15908_), .A2(new_n15906_), .B(new_n15566_), .ZN(new_n15909_));
  INV_X1     g15717(.I(new_n15571_), .ZN(new_n15910_));
  INV_X1     g15718(.I(new_n15581_), .ZN(new_n15911_));
  NOR2_X1    g15719(.A1(new_n15894_), .A2(new_n15895_), .ZN(new_n15912_));
  AOI21_X1   g15720(.A1(new_n15912_), .A2(new_n3167_), .B(new_n15911_), .ZN(new_n15913_));
  NAND2_X1   g15721(.A1(new_n15896_), .A2(new_n2912_), .ZN(new_n15914_));
  OAI21_X1   g15722(.A1(new_n15913_), .A2(new_n15914_), .B(new_n15577_), .ZN(new_n15915_));
  INV_X1     g15723(.I(new_n15896_), .ZN(new_n15916_));
  OAI21_X1   g15724(.A1(new_n15913_), .A2(new_n15916_), .B(\asqrt[41] ), .ZN(new_n15917_));
  NAND3_X1   g15725(.A1(new_n15915_), .A2(new_n15917_), .A3(new_n2699_), .ZN(new_n15918_));
  NAND2_X1   g15726(.A1(new_n15918_), .A2(new_n15574_), .ZN(new_n15919_));
  NAND2_X1   g15727(.A1(new_n15915_), .A2(new_n15917_), .ZN(new_n15920_));
  AOI21_X1   g15728(.A1(new_n15920_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n15921_));
  AOI21_X1   g15729(.A1(new_n15921_), .A2(new_n15919_), .B(new_n15910_), .ZN(new_n15922_));
  AOI21_X1   g15730(.A1(new_n15919_), .A2(new_n15900_), .B(new_n2464_), .ZN(new_n15923_));
  OAI21_X1   g15731(.A1(new_n15922_), .A2(new_n15923_), .B(\asqrt[44] ), .ZN(new_n15924_));
  AOI21_X1   g15732(.A1(new_n15906_), .A2(new_n15924_), .B(new_n2072_), .ZN(new_n15925_));
  NOR2_X1    g15733(.A1(new_n15909_), .A2(new_n15925_), .ZN(new_n15926_));
  AOI21_X1   g15734(.A1(new_n15926_), .A2(new_n1884_), .B(new_n15563_), .ZN(new_n15927_));
  OAI21_X1   g15735(.A1(new_n15909_), .A2(new_n15925_), .B(\asqrt[46] ), .ZN(new_n15928_));
  NAND2_X1   g15736(.A1(new_n15928_), .A2(new_n1688_), .ZN(new_n15929_));
  OAI21_X1   g15737(.A1(new_n15927_), .A2(new_n15929_), .B(new_n15559_), .ZN(new_n15930_));
  INV_X1     g15738(.I(new_n15928_), .ZN(new_n15931_));
  OAI21_X1   g15739(.A1(new_n15927_), .A2(new_n15931_), .B(\asqrt[47] ), .ZN(new_n15932_));
  NAND3_X1   g15740(.A1(new_n15930_), .A2(new_n15932_), .A3(new_n1533_), .ZN(new_n15933_));
  NAND2_X1   g15741(.A1(new_n15933_), .A2(new_n15557_), .ZN(new_n15934_));
  NAND2_X1   g15742(.A1(new_n15930_), .A2(new_n15932_), .ZN(new_n15935_));
  AOI21_X1   g15743(.A1(new_n15935_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n15936_));
  AOI21_X1   g15744(.A1(new_n15936_), .A2(new_n15934_), .B(new_n15554_), .ZN(new_n15937_));
  INV_X1     g15745(.I(new_n15559_), .ZN(new_n15938_));
  INV_X1     g15746(.I(new_n15569_), .ZN(new_n15939_));
  NOR2_X1    g15747(.A1(new_n15922_), .A2(new_n15923_), .ZN(new_n15940_));
  AOI21_X1   g15748(.A1(new_n15940_), .A2(new_n2271_), .B(new_n15939_), .ZN(new_n15941_));
  NAND2_X1   g15749(.A1(new_n15924_), .A2(new_n2072_), .ZN(new_n15942_));
  OAI21_X1   g15750(.A1(new_n15941_), .A2(new_n15942_), .B(new_n15565_), .ZN(new_n15943_));
  INV_X1     g15751(.I(new_n15924_), .ZN(new_n15944_));
  OAI21_X1   g15752(.A1(new_n15941_), .A2(new_n15944_), .B(\asqrt[45] ), .ZN(new_n15945_));
  NAND3_X1   g15753(.A1(new_n15943_), .A2(new_n15945_), .A3(new_n1884_), .ZN(new_n15946_));
  NAND2_X1   g15754(.A1(new_n15946_), .A2(new_n15562_), .ZN(new_n15947_));
  NAND2_X1   g15755(.A1(new_n15943_), .A2(new_n15945_), .ZN(new_n15948_));
  AOI21_X1   g15756(.A1(new_n15948_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n15949_));
  AOI21_X1   g15757(.A1(new_n15949_), .A2(new_n15947_), .B(new_n15938_), .ZN(new_n15950_));
  AOI21_X1   g15758(.A1(new_n15947_), .A2(new_n15928_), .B(new_n1688_), .ZN(new_n15951_));
  OAI21_X1   g15759(.A1(new_n15950_), .A2(new_n15951_), .B(\asqrt[48] ), .ZN(new_n15952_));
  AOI21_X1   g15760(.A1(new_n15934_), .A2(new_n15952_), .B(new_n1368_), .ZN(new_n15953_));
  NOR2_X1    g15761(.A1(new_n15937_), .A2(new_n15953_), .ZN(new_n15954_));
  AOI21_X1   g15762(.A1(new_n15954_), .A2(new_n1228_), .B(new_n15551_), .ZN(new_n15955_));
  OAI21_X1   g15763(.A1(new_n15937_), .A2(new_n15953_), .B(\asqrt[50] ), .ZN(new_n15956_));
  NAND2_X1   g15764(.A1(new_n15956_), .A2(new_n1088_), .ZN(new_n15957_));
  OAI21_X1   g15765(.A1(new_n15955_), .A2(new_n15957_), .B(new_n15547_), .ZN(new_n15958_));
  INV_X1     g15766(.I(new_n15956_), .ZN(new_n15959_));
  OAI21_X1   g15767(.A1(new_n15955_), .A2(new_n15959_), .B(\asqrt[51] ), .ZN(new_n15960_));
  NAND3_X1   g15768(.A1(new_n15958_), .A2(new_n15960_), .A3(new_n962_), .ZN(new_n15961_));
  NAND2_X1   g15769(.A1(new_n15961_), .A2(new_n15545_), .ZN(new_n15962_));
  NAND2_X1   g15770(.A1(new_n15958_), .A2(new_n15960_), .ZN(new_n15963_));
  AOI21_X1   g15771(.A1(new_n15963_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n15964_));
  AOI21_X1   g15772(.A1(new_n15964_), .A2(new_n15962_), .B(new_n15542_), .ZN(new_n15965_));
  INV_X1     g15773(.I(new_n15547_), .ZN(new_n15966_));
  INV_X1     g15774(.I(new_n15557_), .ZN(new_n15967_));
  NOR2_X1    g15775(.A1(new_n15950_), .A2(new_n15951_), .ZN(new_n15968_));
  AOI21_X1   g15776(.A1(new_n15968_), .A2(new_n1533_), .B(new_n15967_), .ZN(new_n15969_));
  NAND2_X1   g15777(.A1(new_n15952_), .A2(new_n1368_), .ZN(new_n15970_));
  OAI21_X1   g15778(.A1(new_n15969_), .A2(new_n15970_), .B(new_n15553_), .ZN(new_n15971_));
  INV_X1     g15779(.I(new_n15952_), .ZN(new_n15972_));
  OAI21_X1   g15780(.A1(new_n15969_), .A2(new_n15972_), .B(\asqrt[49] ), .ZN(new_n15973_));
  NAND3_X1   g15781(.A1(new_n15971_), .A2(new_n15973_), .A3(new_n1228_), .ZN(new_n15974_));
  NAND2_X1   g15782(.A1(new_n15974_), .A2(new_n15550_), .ZN(new_n15975_));
  NAND2_X1   g15783(.A1(new_n15971_), .A2(new_n15973_), .ZN(new_n15976_));
  AOI21_X1   g15784(.A1(new_n15976_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n15977_));
  AOI21_X1   g15785(.A1(new_n15977_), .A2(new_n15975_), .B(new_n15966_), .ZN(new_n15978_));
  AOI21_X1   g15786(.A1(new_n15975_), .A2(new_n15956_), .B(new_n1088_), .ZN(new_n15979_));
  OAI21_X1   g15787(.A1(new_n15978_), .A2(new_n15979_), .B(\asqrt[52] ), .ZN(new_n15980_));
  AOI21_X1   g15788(.A1(new_n15962_), .A2(new_n15980_), .B(new_n842_), .ZN(new_n15981_));
  NOR2_X1    g15789(.A1(new_n15965_), .A2(new_n15981_), .ZN(new_n15982_));
  AOI21_X1   g15790(.A1(new_n15982_), .A2(new_n720_), .B(new_n15539_), .ZN(new_n15983_));
  OAI21_X1   g15791(.A1(new_n15965_), .A2(new_n15981_), .B(\asqrt[54] ), .ZN(new_n15984_));
  NAND2_X1   g15792(.A1(new_n15984_), .A2(new_n630_), .ZN(new_n15985_));
  OAI21_X1   g15793(.A1(new_n15983_), .A2(new_n15985_), .B(new_n15535_), .ZN(new_n15986_));
  INV_X1     g15794(.I(new_n15984_), .ZN(new_n15987_));
  OAI21_X1   g15795(.A1(new_n15983_), .A2(new_n15987_), .B(\asqrt[55] ), .ZN(new_n15988_));
  NAND3_X1   g15796(.A1(new_n15986_), .A2(new_n15988_), .A3(new_n545_), .ZN(new_n15989_));
  INV_X1     g15797(.I(new_n15535_), .ZN(new_n15990_));
  INV_X1     g15798(.I(new_n15545_), .ZN(new_n15991_));
  NOR2_X1    g15799(.A1(new_n15978_), .A2(new_n15979_), .ZN(new_n15992_));
  AOI21_X1   g15800(.A1(new_n15992_), .A2(new_n962_), .B(new_n15991_), .ZN(new_n15993_));
  NAND2_X1   g15801(.A1(new_n15980_), .A2(new_n842_), .ZN(new_n15994_));
  OAI21_X1   g15802(.A1(new_n15993_), .A2(new_n15994_), .B(new_n15541_), .ZN(new_n15995_));
  INV_X1     g15803(.I(new_n15980_), .ZN(new_n15996_));
  OAI21_X1   g15804(.A1(new_n15993_), .A2(new_n15996_), .B(\asqrt[53] ), .ZN(new_n15997_));
  NAND3_X1   g15805(.A1(new_n15995_), .A2(new_n15997_), .A3(new_n720_), .ZN(new_n15998_));
  NAND2_X1   g15806(.A1(new_n15998_), .A2(new_n15538_), .ZN(new_n15999_));
  NAND2_X1   g15807(.A1(new_n15995_), .A2(new_n15997_), .ZN(new_n16000_));
  AOI21_X1   g15808(.A1(new_n16000_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n16001_));
  AOI21_X1   g15809(.A1(new_n16001_), .A2(new_n15999_), .B(new_n15990_), .ZN(new_n16002_));
  AOI21_X1   g15810(.A1(new_n15999_), .A2(new_n15984_), .B(new_n630_), .ZN(new_n16003_));
  OAI21_X1   g15811(.A1(new_n16002_), .A2(new_n16003_), .B(\asqrt[56] ), .ZN(new_n16004_));
  NAND2_X1   g15812(.A1(new_n15515_), .A2(new_n14990_), .ZN(new_n16005_));
  NOR2_X1    g15813(.A1(new_n15518_), .A2(new_n14990_), .ZN(new_n16006_));
  NAND2_X1   g15814(.A1(new_n16006_), .A2(new_n15530_), .ZN(new_n16007_));
  AOI21_X1   g15815(.A1(new_n16007_), .A2(new_n16005_), .B(new_n193_), .ZN(new_n16008_));
  INV_X1     g15816(.I(new_n16008_), .ZN(new_n16009_));
  NAND3_X1   g15817(.A1(\asqrt[9] ), .A2(new_n15500_), .A3(new_n15511_), .ZN(new_n16010_));
  XOR2_X1    g15818(.A1(new_n16010_), .A2(new_n15503_), .Z(new_n16011_));
  AOI21_X1   g15819(.A1(new_n16006_), .A2(new_n15515_), .B(new_n15516_), .ZN(new_n16012_));
  OAI21_X1   g15820(.A1(new_n15470_), .A2(new_n15472_), .B(new_n15475_), .ZN(new_n16013_));
  NOR2_X1    g15821(.A1(new_n15518_), .A2(new_n16013_), .ZN(new_n16014_));
  XOR2_X1    g15822(.A1(new_n16014_), .A2(new_n14998_), .Z(new_n16015_));
  NAND3_X1   g15823(.A1(\asqrt[9] ), .A2(new_n15486_), .A3(new_n15471_), .ZN(new_n16016_));
  XOR2_X1    g15824(.A1(new_n16016_), .A2(new_n15002_), .Z(new_n16017_));
  OAI21_X1   g15825(.A1(new_n15481_), .A2(new_n15482_), .B(new_n15485_), .ZN(new_n16018_));
  NOR2_X1    g15826(.A1(new_n15518_), .A2(new_n16018_), .ZN(new_n16019_));
  XOR2_X1    g15827(.A1(new_n16019_), .A2(new_n15004_), .Z(new_n16020_));
  INV_X1     g15828(.I(new_n16020_), .ZN(new_n16021_));
  NAND3_X1   g15829(.A1(\asqrt[9] ), .A2(new_n15448_), .A3(new_n15467_), .ZN(new_n16022_));
  XOR2_X1    g15830(.A1(new_n16022_), .A2(new_n15479_), .Z(new_n16023_));
  INV_X1     g15831(.I(new_n16023_), .ZN(new_n16024_));
  NAND2_X1   g15832(.A1(new_n15989_), .A2(new_n15521_), .ZN(new_n16025_));
  NAND2_X1   g15833(.A1(new_n15986_), .A2(new_n15988_), .ZN(new_n16026_));
  AOI21_X1   g15834(.A1(new_n16026_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n16027_));
  AOI21_X1   g15835(.A1(new_n16027_), .A2(new_n16025_), .B(new_n16024_), .ZN(new_n16028_));
  AOI21_X1   g15836(.A1(new_n16025_), .A2(new_n16004_), .B(new_n450_), .ZN(new_n16029_));
  NOR2_X1    g15837(.A1(new_n16028_), .A2(new_n16029_), .ZN(new_n16030_));
  AOI21_X1   g15838(.A1(new_n16030_), .A2(new_n403_), .B(new_n16021_), .ZN(new_n16031_));
  OAI21_X1   g15839(.A1(new_n16028_), .A2(new_n16029_), .B(\asqrt[58] ), .ZN(new_n16032_));
  NAND2_X1   g15840(.A1(new_n16032_), .A2(new_n339_), .ZN(new_n16033_));
  OAI21_X1   g15841(.A1(new_n16031_), .A2(new_n16033_), .B(new_n16017_), .ZN(new_n16034_));
  INV_X1     g15842(.I(new_n16032_), .ZN(new_n16035_));
  OAI21_X1   g15843(.A1(new_n16031_), .A2(new_n16035_), .B(\asqrt[59] ), .ZN(new_n16036_));
  NAND3_X1   g15844(.A1(new_n16034_), .A2(new_n16036_), .A3(new_n288_), .ZN(new_n16037_));
  NAND2_X1   g15845(.A1(new_n16037_), .A2(new_n16015_), .ZN(new_n16038_));
  INV_X1     g15846(.I(new_n16017_), .ZN(new_n16039_));
  NOR2_X1    g15847(.A1(new_n16002_), .A2(new_n16003_), .ZN(new_n16040_));
  AOI21_X1   g15848(.A1(new_n16040_), .A2(new_n545_), .B(new_n15522_), .ZN(new_n16041_));
  NAND2_X1   g15849(.A1(new_n16004_), .A2(new_n450_), .ZN(new_n16042_));
  OAI21_X1   g15850(.A1(new_n16041_), .A2(new_n16042_), .B(new_n16023_), .ZN(new_n16043_));
  INV_X1     g15851(.I(new_n16004_), .ZN(new_n16044_));
  OAI21_X1   g15852(.A1(new_n16041_), .A2(new_n16044_), .B(\asqrt[57] ), .ZN(new_n16045_));
  NAND3_X1   g15853(.A1(new_n16043_), .A2(new_n16045_), .A3(new_n403_), .ZN(new_n16046_));
  NAND2_X1   g15854(.A1(new_n16046_), .A2(new_n16020_), .ZN(new_n16047_));
  NAND2_X1   g15855(.A1(new_n16043_), .A2(new_n16045_), .ZN(new_n16048_));
  AOI21_X1   g15856(.A1(new_n16048_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n16049_));
  AOI21_X1   g15857(.A1(new_n16049_), .A2(new_n16047_), .B(new_n16039_), .ZN(new_n16050_));
  AOI21_X1   g15858(.A1(new_n16047_), .A2(new_n16032_), .B(new_n339_), .ZN(new_n16051_));
  OAI21_X1   g15859(.A1(new_n16050_), .A2(new_n16051_), .B(\asqrt[60] ), .ZN(new_n16052_));
  AOI21_X1   g15860(.A1(new_n16038_), .A2(new_n16052_), .B(new_n242_), .ZN(new_n16053_));
  NAND3_X1   g15861(.A1(\asqrt[9] ), .A2(new_n15476_), .A3(new_n15492_), .ZN(new_n16054_));
  XOR2_X1    g15862(.A1(new_n16054_), .A2(new_n15504_), .Z(new_n16055_));
  INV_X1     g15863(.I(new_n16055_), .ZN(new_n16056_));
  NAND2_X1   g15864(.A1(new_n16034_), .A2(new_n16036_), .ZN(new_n16057_));
  AOI21_X1   g15865(.A1(new_n16057_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n16058_));
  AOI21_X1   g15866(.A1(new_n16058_), .A2(new_n16038_), .B(new_n16056_), .ZN(new_n16059_));
  OAI21_X1   g15867(.A1(new_n16059_), .A2(new_n16053_), .B(\asqrt[62] ), .ZN(new_n16060_));
  INV_X1     g15868(.I(new_n16060_), .ZN(new_n16061_));
  NOR2_X1    g15869(.A1(new_n16059_), .A2(new_n16053_), .ZN(new_n16062_));
  AOI21_X1   g15870(.A1(new_n15477_), .A2(new_n15498_), .B(new_n15493_), .ZN(new_n16063_));
  NAND2_X1   g15871(.A1(\asqrt[9] ), .A2(new_n16063_), .ZN(new_n16064_));
  XOR2_X1    g15872(.A1(new_n16064_), .A2(new_n15496_), .Z(new_n16065_));
  INV_X1     g15873(.I(new_n16065_), .ZN(new_n16066_));
  AOI21_X1   g15874(.A1(new_n16062_), .A2(new_n234_), .B(new_n16066_), .ZN(new_n16067_));
  OAI21_X1   g15875(.A1(new_n16067_), .A2(new_n16061_), .B(new_n16012_), .ZN(new_n16068_));
  OAI21_X1   g15876(.A1(new_n16068_), .A2(new_n16011_), .B(new_n193_), .ZN(new_n16069_));
  NOR2_X1    g15877(.A1(new_n16067_), .A2(new_n16061_), .ZN(new_n16070_));
  NAND2_X1   g15878(.A1(new_n16070_), .A2(new_n16011_), .ZN(new_n16071_));
  NOR2_X1    g15879(.A1(\asqrt[9] ), .A2(new_n14991_), .ZN(new_n16072_));
  INV_X1     g15880(.I(new_n16072_), .ZN(new_n16073_));
  NAND4_X1   g15881(.A1(new_n16069_), .A2(new_n16009_), .A3(new_n16071_), .A4(new_n16073_), .ZN(\asqrt[8] ));
  NAND3_X1   g15882(.A1(\asqrt[8] ), .A2(new_n15989_), .A3(new_n16004_), .ZN(new_n16075_));
  XOR2_X1    g15883(.A1(new_n16075_), .A2(new_n15522_), .Z(new_n16076_));
  INV_X1     g15884(.I(new_n16015_), .ZN(new_n16077_));
  NOR2_X1    g15885(.A1(new_n16050_), .A2(new_n16051_), .ZN(new_n16078_));
  AOI21_X1   g15886(.A1(new_n16078_), .A2(new_n288_), .B(new_n16077_), .ZN(new_n16079_));
  INV_X1     g15887(.I(new_n16052_), .ZN(new_n16080_));
  OAI21_X1   g15888(.A1(new_n16079_), .A2(new_n16080_), .B(\asqrt[61] ), .ZN(new_n16081_));
  NAND2_X1   g15889(.A1(new_n16052_), .A2(new_n242_), .ZN(new_n16082_));
  OAI21_X1   g15890(.A1(new_n16079_), .A2(new_n16082_), .B(new_n16055_), .ZN(new_n16083_));
  NAND3_X1   g15891(.A1(new_n16083_), .A2(new_n16081_), .A3(new_n234_), .ZN(new_n16084_));
  NAND2_X1   g15892(.A1(new_n16084_), .A2(new_n16065_), .ZN(new_n16085_));
  NAND2_X1   g15893(.A1(new_n16085_), .A2(new_n16060_), .ZN(new_n16086_));
  NAND2_X1   g15894(.A1(new_n16086_), .A2(new_n16011_), .ZN(new_n16087_));
  INV_X1     g15895(.I(new_n16011_), .ZN(new_n16088_));
  INV_X1     g15896(.I(new_n16012_), .ZN(new_n16089_));
  AOI21_X1   g15897(.A1(new_n16085_), .A2(new_n16060_), .B(new_n16089_), .ZN(new_n16090_));
  AOI21_X1   g15898(.A1(new_n16090_), .A2(new_n16088_), .B(\asqrt[63] ), .ZN(new_n16091_));
  NOR2_X1    g15899(.A1(new_n16086_), .A2(new_n16088_), .ZN(new_n16092_));
  NOR4_X1    g15900(.A1(new_n16091_), .A2(new_n16008_), .A3(new_n16092_), .A4(new_n16072_), .ZN(new_n16093_));
  NOR2_X1    g15901(.A1(new_n16093_), .A2(new_n16011_), .ZN(new_n16094_));
  NAND2_X1   g15902(.A1(new_n16094_), .A2(new_n16070_), .ZN(new_n16095_));
  AOI21_X1   g15903(.A1(new_n16095_), .A2(new_n16087_), .B(new_n193_), .ZN(new_n16096_));
  NAND3_X1   g15904(.A1(\asqrt[8] ), .A2(new_n16060_), .A3(new_n16084_), .ZN(new_n16097_));
  XOR2_X1    g15905(.A1(new_n16097_), .A2(new_n16065_), .Z(new_n16098_));
  INV_X1     g15906(.I(new_n16098_), .ZN(new_n16099_));
  AOI21_X1   g15907(.A1(new_n16094_), .A2(new_n16086_), .B(new_n16092_), .ZN(new_n16100_));
  INV_X1     g15908(.I(new_n16100_), .ZN(new_n16101_));
  OAI21_X1   g15909(.A1(new_n16031_), .A2(new_n16033_), .B(new_n16036_), .ZN(new_n16102_));
  NOR2_X1    g15910(.A1(new_n16093_), .A2(new_n16102_), .ZN(new_n16103_));
  XOR2_X1    g15911(.A1(new_n16103_), .A2(new_n16017_), .Z(new_n16104_));
  NAND3_X1   g15912(.A1(\asqrt[8] ), .A2(new_n16046_), .A3(new_n16032_), .ZN(new_n16105_));
  XOR2_X1    g15913(.A1(new_n16105_), .A2(new_n16021_), .Z(new_n16106_));
  OAI21_X1   g15914(.A1(new_n16041_), .A2(new_n16042_), .B(new_n16045_), .ZN(new_n16107_));
  NOR2_X1    g15915(.A1(new_n16093_), .A2(new_n16107_), .ZN(new_n16108_));
  XOR2_X1    g15916(.A1(new_n16108_), .A2(new_n16023_), .Z(new_n16109_));
  INV_X1     g15917(.I(new_n16109_), .ZN(new_n16110_));
  INV_X1     g15918(.I(new_n16076_), .ZN(new_n16111_));
  OAI21_X1   g15919(.A1(new_n15983_), .A2(new_n15985_), .B(new_n15988_), .ZN(new_n16112_));
  NOR2_X1    g15920(.A1(new_n16093_), .A2(new_n16112_), .ZN(new_n16113_));
  XOR2_X1    g15921(.A1(new_n16113_), .A2(new_n15535_), .Z(new_n16114_));
  NAND3_X1   g15922(.A1(\asqrt[8] ), .A2(new_n15998_), .A3(new_n15984_), .ZN(new_n16115_));
  XOR2_X1    g15923(.A1(new_n16115_), .A2(new_n15539_), .Z(new_n16116_));
  OAI21_X1   g15924(.A1(new_n15993_), .A2(new_n15994_), .B(new_n15997_), .ZN(new_n16117_));
  NOR2_X1    g15925(.A1(new_n16093_), .A2(new_n16117_), .ZN(new_n16118_));
  XOR2_X1    g15926(.A1(new_n16118_), .A2(new_n15541_), .Z(new_n16119_));
  INV_X1     g15927(.I(new_n16119_), .ZN(new_n16120_));
  NAND3_X1   g15928(.A1(\asqrt[8] ), .A2(new_n15961_), .A3(new_n15980_), .ZN(new_n16121_));
  XOR2_X1    g15929(.A1(new_n16121_), .A2(new_n15991_), .Z(new_n16122_));
  INV_X1     g15930(.I(new_n16122_), .ZN(new_n16123_));
  OAI21_X1   g15931(.A1(new_n15955_), .A2(new_n15957_), .B(new_n15960_), .ZN(new_n16124_));
  NOR2_X1    g15932(.A1(new_n16093_), .A2(new_n16124_), .ZN(new_n16125_));
  XOR2_X1    g15933(.A1(new_n16125_), .A2(new_n15547_), .Z(new_n16126_));
  NAND3_X1   g15934(.A1(\asqrt[8] ), .A2(new_n15974_), .A3(new_n15956_), .ZN(new_n16127_));
  XOR2_X1    g15935(.A1(new_n16127_), .A2(new_n15551_), .Z(new_n16128_));
  OAI21_X1   g15936(.A1(new_n15969_), .A2(new_n15970_), .B(new_n15973_), .ZN(new_n16129_));
  NOR2_X1    g15937(.A1(new_n16093_), .A2(new_n16129_), .ZN(new_n16130_));
  XOR2_X1    g15938(.A1(new_n16130_), .A2(new_n15553_), .Z(new_n16131_));
  INV_X1     g15939(.I(new_n16131_), .ZN(new_n16132_));
  NAND3_X1   g15940(.A1(\asqrt[8] ), .A2(new_n15933_), .A3(new_n15952_), .ZN(new_n16133_));
  XOR2_X1    g15941(.A1(new_n16133_), .A2(new_n15967_), .Z(new_n16134_));
  INV_X1     g15942(.I(new_n16134_), .ZN(new_n16135_));
  OAI21_X1   g15943(.A1(new_n15927_), .A2(new_n15929_), .B(new_n15932_), .ZN(new_n16136_));
  NOR2_X1    g15944(.A1(new_n16093_), .A2(new_n16136_), .ZN(new_n16137_));
  XOR2_X1    g15945(.A1(new_n16137_), .A2(new_n15559_), .Z(new_n16138_));
  NAND3_X1   g15946(.A1(\asqrt[8] ), .A2(new_n15946_), .A3(new_n15928_), .ZN(new_n16139_));
  XOR2_X1    g15947(.A1(new_n16139_), .A2(new_n15563_), .Z(new_n16140_));
  OAI21_X1   g15948(.A1(new_n15941_), .A2(new_n15942_), .B(new_n15945_), .ZN(new_n16141_));
  NOR2_X1    g15949(.A1(new_n16093_), .A2(new_n16141_), .ZN(new_n16142_));
  XOR2_X1    g15950(.A1(new_n16142_), .A2(new_n15565_), .Z(new_n16143_));
  INV_X1     g15951(.I(new_n16143_), .ZN(new_n16144_));
  NAND3_X1   g15952(.A1(\asqrt[8] ), .A2(new_n15905_), .A3(new_n15924_), .ZN(new_n16145_));
  XOR2_X1    g15953(.A1(new_n16145_), .A2(new_n15939_), .Z(new_n16146_));
  INV_X1     g15954(.I(new_n16146_), .ZN(new_n16147_));
  OAI21_X1   g15955(.A1(new_n15899_), .A2(new_n15901_), .B(new_n15904_), .ZN(new_n16148_));
  NOR2_X1    g15956(.A1(new_n16093_), .A2(new_n16148_), .ZN(new_n16149_));
  XOR2_X1    g15957(.A1(new_n16149_), .A2(new_n15571_), .Z(new_n16150_));
  NAND3_X1   g15958(.A1(\asqrt[8] ), .A2(new_n15918_), .A3(new_n15900_), .ZN(new_n16151_));
  XOR2_X1    g15959(.A1(new_n16151_), .A2(new_n15575_), .Z(new_n16152_));
  OAI21_X1   g15960(.A1(new_n15913_), .A2(new_n15914_), .B(new_n15917_), .ZN(new_n16153_));
  NOR2_X1    g15961(.A1(new_n16093_), .A2(new_n16153_), .ZN(new_n16154_));
  XOR2_X1    g15962(.A1(new_n16154_), .A2(new_n15577_), .Z(new_n16155_));
  INV_X1     g15963(.I(new_n16155_), .ZN(new_n16156_));
  NAND3_X1   g15964(.A1(\asqrt[8] ), .A2(new_n15877_), .A3(new_n15896_), .ZN(new_n16157_));
  XOR2_X1    g15965(.A1(new_n16157_), .A2(new_n15911_), .Z(new_n16158_));
  INV_X1     g15966(.I(new_n16158_), .ZN(new_n16159_));
  OAI21_X1   g15967(.A1(new_n15871_), .A2(new_n15873_), .B(new_n15876_), .ZN(new_n16160_));
  NOR2_X1    g15968(.A1(new_n16093_), .A2(new_n16160_), .ZN(new_n16161_));
  XOR2_X1    g15969(.A1(new_n16161_), .A2(new_n15583_), .Z(new_n16162_));
  NAND3_X1   g15970(.A1(\asqrt[8] ), .A2(new_n15890_), .A3(new_n15872_), .ZN(new_n16163_));
  XOR2_X1    g15971(.A1(new_n16163_), .A2(new_n15587_), .Z(new_n16164_));
  OAI21_X1   g15972(.A1(new_n15885_), .A2(new_n15886_), .B(new_n15889_), .ZN(new_n16165_));
  NOR2_X1    g15973(.A1(new_n16093_), .A2(new_n16165_), .ZN(new_n16166_));
  XOR2_X1    g15974(.A1(new_n16166_), .A2(new_n15589_), .Z(new_n16167_));
  INV_X1     g15975(.I(new_n16167_), .ZN(new_n16168_));
  NAND3_X1   g15976(.A1(\asqrt[8] ), .A2(new_n15849_), .A3(new_n15868_), .ZN(new_n16169_));
  XOR2_X1    g15977(.A1(new_n16169_), .A2(new_n15883_), .Z(new_n16170_));
  INV_X1     g15978(.I(new_n16170_), .ZN(new_n16171_));
  OAI21_X1   g15979(.A1(new_n15843_), .A2(new_n15845_), .B(new_n15848_), .ZN(new_n16172_));
  NOR2_X1    g15980(.A1(new_n16093_), .A2(new_n16172_), .ZN(new_n16173_));
  XOR2_X1    g15981(.A1(new_n16173_), .A2(new_n15595_), .Z(new_n16174_));
  NAND3_X1   g15982(.A1(\asqrt[8] ), .A2(new_n15862_), .A3(new_n15844_), .ZN(new_n16175_));
  XOR2_X1    g15983(.A1(new_n16175_), .A2(new_n15599_), .Z(new_n16176_));
  OAI21_X1   g15984(.A1(new_n15857_), .A2(new_n15858_), .B(new_n15861_), .ZN(new_n16177_));
  NOR2_X1    g15985(.A1(new_n16093_), .A2(new_n16177_), .ZN(new_n16178_));
  XOR2_X1    g15986(.A1(new_n16178_), .A2(new_n15601_), .Z(new_n16179_));
  INV_X1     g15987(.I(new_n16179_), .ZN(new_n16180_));
  NAND3_X1   g15988(.A1(\asqrt[8] ), .A2(new_n15821_), .A3(new_n15840_), .ZN(new_n16181_));
  XOR2_X1    g15989(.A1(new_n16181_), .A2(new_n15855_), .Z(new_n16182_));
  INV_X1     g15990(.I(new_n16182_), .ZN(new_n16183_));
  OAI21_X1   g15991(.A1(new_n15815_), .A2(new_n15817_), .B(new_n15820_), .ZN(new_n16184_));
  NOR2_X1    g15992(.A1(new_n16093_), .A2(new_n16184_), .ZN(new_n16185_));
  XOR2_X1    g15993(.A1(new_n16185_), .A2(new_n15607_), .Z(new_n16186_));
  NAND3_X1   g15994(.A1(\asqrt[8] ), .A2(new_n15834_), .A3(new_n15816_), .ZN(new_n16187_));
  XOR2_X1    g15995(.A1(new_n16187_), .A2(new_n15611_), .Z(new_n16188_));
  OAI21_X1   g15996(.A1(new_n15829_), .A2(new_n15830_), .B(new_n15833_), .ZN(new_n16189_));
  NOR2_X1    g15997(.A1(new_n16093_), .A2(new_n16189_), .ZN(new_n16190_));
  XOR2_X1    g15998(.A1(new_n16190_), .A2(new_n15613_), .Z(new_n16191_));
  INV_X1     g15999(.I(new_n16191_), .ZN(new_n16192_));
  NAND3_X1   g16000(.A1(\asqrt[8] ), .A2(new_n15793_), .A3(new_n15812_), .ZN(new_n16193_));
  XOR2_X1    g16001(.A1(new_n16193_), .A2(new_n15827_), .Z(new_n16194_));
  INV_X1     g16002(.I(new_n16194_), .ZN(new_n16195_));
  OAI21_X1   g16003(.A1(new_n15787_), .A2(new_n15789_), .B(new_n15792_), .ZN(new_n16196_));
  NOR2_X1    g16004(.A1(new_n16093_), .A2(new_n16196_), .ZN(new_n16197_));
  XOR2_X1    g16005(.A1(new_n16197_), .A2(new_n15619_), .Z(new_n16198_));
  NAND3_X1   g16006(.A1(\asqrt[8] ), .A2(new_n15806_), .A3(new_n15788_), .ZN(new_n16199_));
  XOR2_X1    g16007(.A1(new_n16199_), .A2(new_n15623_), .Z(new_n16200_));
  OAI21_X1   g16008(.A1(new_n15801_), .A2(new_n15802_), .B(new_n15805_), .ZN(new_n16201_));
  NOR2_X1    g16009(.A1(new_n16093_), .A2(new_n16201_), .ZN(new_n16202_));
  XOR2_X1    g16010(.A1(new_n16202_), .A2(new_n15625_), .Z(new_n16203_));
  INV_X1     g16011(.I(new_n16203_), .ZN(new_n16204_));
  NAND3_X1   g16012(.A1(\asqrt[8] ), .A2(new_n15765_), .A3(new_n15784_), .ZN(new_n16205_));
  XOR2_X1    g16013(.A1(new_n16205_), .A2(new_n15799_), .Z(new_n16206_));
  INV_X1     g16014(.I(new_n16206_), .ZN(new_n16207_));
  OAI21_X1   g16015(.A1(new_n15759_), .A2(new_n15761_), .B(new_n15764_), .ZN(new_n16208_));
  NOR2_X1    g16016(.A1(new_n16093_), .A2(new_n16208_), .ZN(new_n16209_));
  XOR2_X1    g16017(.A1(new_n16209_), .A2(new_n15631_), .Z(new_n16210_));
  NAND3_X1   g16018(.A1(\asqrt[8] ), .A2(new_n15778_), .A3(new_n15760_), .ZN(new_n16211_));
  XOR2_X1    g16019(.A1(new_n16211_), .A2(new_n15635_), .Z(new_n16212_));
  OAI21_X1   g16020(.A1(new_n15773_), .A2(new_n15774_), .B(new_n15777_), .ZN(new_n16213_));
  NOR2_X1    g16021(.A1(new_n16093_), .A2(new_n16213_), .ZN(new_n16214_));
  XOR2_X1    g16022(.A1(new_n16214_), .A2(new_n15637_), .Z(new_n16215_));
  INV_X1     g16023(.I(new_n16215_), .ZN(new_n16216_));
  NAND3_X1   g16024(.A1(\asqrt[8] ), .A2(new_n15737_), .A3(new_n15756_), .ZN(new_n16217_));
  XOR2_X1    g16025(.A1(new_n16217_), .A2(new_n15771_), .Z(new_n16218_));
  INV_X1     g16026(.I(new_n16218_), .ZN(new_n16219_));
  OAI21_X1   g16027(.A1(new_n15731_), .A2(new_n15733_), .B(new_n15736_), .ZN(new_n16220_));
  NOR2_X1    g16028(.A1(new_n16093_), .A2(new_n16220_), .ZN(new_n16221_));
  XOR2_X1    g16029(.A1(new_n16221_), .A2(new_n15643_), .Z(new_n16222_));
  NAND3_X1   g16030(.A1(\asqrt[8] ), .A2(new_n15750_), .A3(new_n15732_), .ZN(new_n16223_));
  XOR2_X1    g16031(.A1(new_n16223_), .A2(new_n15647_), .Z(new_n16224_));
  OAI21_X1   g16032(.A1(new_n15745_), .A2(new_n15746_), .B(new_n15749_), .ZN(new_n16225_));
  NOR2_X1    g16033(.A1(new_n16093_), .A2(new_n16225_), .ZN(new_n16226_));
  XOR2_X1    g16034(.A1(new_n16226_), .A2(new_n15649_), .Z(new_n16227_));
  INV_X1     g16035(.I(new_n16227_), .ZN(new_n16228_));
  NAND3_X1   g16036(.A1(\asqrt[8] ), .A2(new_n15709_), .A3(new_n15728_), .ZN(new_n16229_));
  XOR2_X1    g16037(.A1(new_n16229_), .A2(new_n15743_), .Z(new_n16230_));
  INV_X1     g16038(.I(new_n16230_), .ZN(new_n16231_));
  OAI21_X1   g16039(.A1(new_n15703_), .A2(new_n15705_), .B(new_n15708_), .ZN(new_n16232_));
  NOR2_X1    g16040(.A1(new_n16093_), .A2(new_n16232_), .ZN(new_n16233_));
  XOR2_X1    g16041(.A1(new_n16233_), .A2(new_n15656_), .Z(new_n16234_));
  NAND3_X1   g16042(.A1(\asqrt[8] ), .A2(new_n15722_), .A3(new_n15704_), .ZN(new_n16235_));
  XOR2_X1    g16043(.A1(new_n16235_), .A2(new_n15659_), .Z(new_n16236_));
  OAI21_X1   g16044(.A1(new_n15717_), .A2(new_n15718_), .B(new_n15721_), .ZN(new_n16237_));
  NOR2_X1    g16045(.A1(new_n16093_), .A2(new_n16237_), .ZN(new_n16238_));
  XOR2_X1    g16046(.A1(new_n16238_), .A2(new_n15662_), .Z(new_n16239_));
  INV_X1     g16047(.I(new_n16239_), .ZN(new_n16240_));
  NAND3_X1   g16048(.A1(\asqrt[8] ), .A2(new_n15682_), .A3(new_n15700_), .ZN(new_n16241_));
  XOR2_X1    g16049(.A1(new_n16241_), .A2(new_n15716_), .Z(new_n16242_));
  INV_X1     g16050(.I(new_n16242_), .ZN(new_n16243_));
  NOR2_X1    g16051(.A1(new_n15679_), .A2(\asqrt[11] ), .ZN(new_n16244_));
  NOR3_X1    g16052(.A1(new_n16093_), .A2(new_n16244_), .A3(new_n15699_), .ZN(new_n16245_));
  XOR2_X1    g16053(.A1(new_n16245_), .A2(new_n15670_), .Z(new_n16246_));
  NOR3_X1    g16054(.A1(new_n16093_), .A2(\a[16] ), .A3(\a[17] ), .ZN(new_n16247_));
  NOR4_X1    g16055(.A1(new_n16091_), .A2(new_n15518_), .A3(new_n16008_), .A4(new_n16092_), .ZN(new_n16248_));
  OAI21_X1   g16056(.A1(new_n16247_), .A2(new_n16248_), .B(new_n15140_), .ZN(new_n16249_));
  NAND3_X1   g16057(.A1(\asqrt[8] ), .A2(new_n15671_), .A3(new_n15672_), .ZN(new_n16250_));
  INV_X1     g16058(.I(new_n16248_), .ZN(new_n16251_));
  NAND3_X1   g16059(.A1(new_n16250_), .A2(\a[18] ), .A3(new_n16251_), .ZN(new_n16252_));
  NAND2_X1   g16060(.A1(new_n16249_), .A2(new_n16252_), .ZN(new_n16253_));
  INV_X1     g16061(.I(\a[14] ), .ZN(new_n16254_));
  INV_X1     g16062(.I(\a[15] ), .ZN(new_n16255_));
  NAND3_X1   g16063(.A1(new_n16254_), .A2(new_n16255_), .A3(new_n15671_), .ZN(new_n16256_));
  NAND2_X1   g16064(.A1(\asqrt[8] ), .A2(\a[16] ), .ZN(new_n16257_));
  AOI21_X1   g16065(.A1(new_n16257_), .A2(new_n16256_), .B(new_n15518_), .ZN(new_n16258_));
  AOI21_X1   g16066(.A1(\asqrt[8] ), .A2(new_n15671_), .B(new_n15672_), .ZN(new_n16259_));
  NOR2_X1    g16067(.A1(new_n16247_), .A2(new_n16259_), .ZN(new_n16260_));
  NAND3_X1   g16068(.A1(new_n16257_), .A2(new_n15518_), .A3(new_n16256_), .ZN(new_n16261_));
  AOI21_X1   g16069(.A1(new_n16260_), .A2(new_n16261_), .B(new_n16258_), .ZN(new_n16262_));
  AOI21_X1   g16070(.A1(new_n16262_), .A2(new_n14985_), .B(new_n16253_), .ZN(new_n16263_));
  NOR2_X1    g16071(.A1(new_n16262_), .A2(new_n14985_), .ZN(new_n16264_));
  NOR3_X1    g16072(.A1(new_n16263_), .A2(\asqrt[11] ), .A3(new_n16264_), .ZN(new_n16265_));
  NOR3_X1    g16073(.A1(new_n16093_), .A2(new_n15693_), .A3(new_n15678_), .ZN(new_n16266_));
  XOR2_X1    g16074(.A1(new_n16266_), .A2(new_n15695_), .Z(new_n16267_));
  INV_X1     g16075(.I(new_n16267_), .ZN(new_n16268_));
  OAI21_X1   g16076(.A1(new_n16263_), .A2(new_n16264_), .B(\asqrt[11] ), .ZN(new_n16269_));
  OAI21_X1   g16077(.A1(new_n16265_), .A2(new_n16268_), .B(new_n16269_), .ZN(new_n16270_));
  OAI21_X1   g16078(.A1(new_n16270_), .A2(\asqrt[12] ), .B(new_n16246_), .ZN(new_n16271_));
  AOI21_X1   g16079(.A1(new_n16270_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n16272_));
  AOI21_X1   g16080(.A1(new_n16272_), .A2(new_n16271_), .B(new_n16243_), .ZN(new_n16273_));
  NAND2_X1   g16081(.A1(new_n16270_), .A2(\asqrt[12] ), .ZN(new_n16274_));
  AOI21_X1   g16082(.A1(new_n16271_), .A2(new_n16274_), .B(new_n13382_), .ZN(new_n16275_));
  NOR2_X1    g16083(.A1(new_n16273_), .A2(new_n16275_), .ZN(new_n16276_));
  AOI21_X1   g16084(.A1(new_n16276_), .A2(new_n12889_), .B(new_n16240_), .ZN(new_n16277_));
  OAI21_X1   g16085(.A1(new_n16273_), .A2(new_n16275_), .B(\asqrt[14] ), .ZN(new_n16278_));
  NAND2_X1   g16086(.A1(new_n16278_), .A2(new_n12374_), .ZN(new_n16279_));
  OAI21_X1   g16087(.A1(new_n16277_), .A2(new_n16279_), .B(new_n16236_), .ZN(new_n16280_));
  INV_X1     g16088(.I(new_n16278_), .ZN(new_n16281_));
  OAI21_X1   g16089(.A1(new_n16277_), .A2(new_n16281_), .B(\asqrt[15] ), .ZN(new_n16282_));
  NAND3_X1   g16090(.A1(new_n16280_), .A2(new_n16282_), .A3(new_n11901_), .ZN(new_n16283_));
  NAND2_X1   g16091(.A1(new_n16283_), .A2(new_n16234_), .ZN(new_n16284_));
  NAND2_X1   g16092(.A1(new_n16280_), .A2(new_n16282_), .ZN(new_n16285_));
  AOI21_X1   g16093(.A1(new_n16285_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n16286_));
  AOI21_X1   g16094(.A1(new_n16286_), .A2(new_n16284_), .B(new_n16231_), .ZN(new_n16287_));
  INV_X1     g16095(.I(new_n16236_), .ZN(new_n16288_));
  INV_X1     g16096(.I(new_n16246_), .ZN(new_n16289_));
  AOI21_X1   g16097(.A1(new_n16250_), .A2(new_n16251_), .B(\a[18] ), .ZN(new_n16290_));
  NOR3_X1    g16098(.A1(new_n16247_), .A2(new_n15140_), .A3(new_n16248_), .ZN(new_n16291_));
  NOR2_X1    g16099(.A1(new_n16291_), .A2(new_n16290_), .ZN(new_n16292_));
  OAI21_X1   g16100(.A1(new_n16093_), .A2(new_n15671_), .B(new_n16256_), .ZN(new_n16293_));
  NAND2_X1   g16101(.A1(new_n16293_), .A2(\asqrt[9] ), .ZN(new_n16294_));
  OAI21_X1   g16102(.A1(new_n16093_), .A2(\a[16] ), .B(\a[17] ), .ZN(new_n16295_));
  NAND2_X1   g16103(.A1(new_n16295_), .A2(new_n16250_), .ZN(new_n16296_));
  NOR2_X1    g16104(.A1(new_n16293_), .A2(\asqrt[9] ), .ZN(new_n16297_));
  OAI21_X1   g16105(.A1(new_n16296_), .A2(new_n16297_), .B(new_n16294_), .ZN(new_n16298_));
  OAI21_X1   g16106(.A1(\asqrt[10] ), .A2(new_n16298_), .B(new_n16292_), .ZN(new_n16299_));
  NAND2_X1   g16107(.A1(new_n16298_), .A2(\asqrt[10] ), .ZN(new_n16300_));
  NAND3_X1   g16108(.A1(new_n16299_), .A2(new_n14430_), .A3(new_n16300_), .ZN(new_n16301_));
  AOI21_X1   g16109(.A1(new_n16299_), .A2(new_n16300_), .B(new_n14430_), .ZN(new_n16302_));
  AOI21_X1   g16110(.A1(new_n16301_), .A2(new_n16267_), .B(new_n16302_), .ZN(new_n16303_));
  AOI21_X1   g16111(.A1(new_n16303_), .A2(new_n13917_), .B(new_n16289_), .ZN(new_n16304_));
  OAI21_X1   g16112(.A1(new_n16303_), .A2(new_n13917_), .B(new_n13382_), .ZN(new_n16305_));
  OAI21_X1   g16113(.A1(new_n16304_), .A2(new_n16305_), .B(new_n16242_), .ZN(new_n16306_));
  NOR2_X1    g16114(.A1(new_n16303_), .A2(new_n13917_), .ZN(new_n16307_));
  OAI21_X1   g16115(.A1(new_n16304_), .A2(new_n16307_), .B(\asqrt[13] ), .ZN(new_n16308_));
  NAND3_X1   g16116(.A1(new_n16306_), .A2(new_n16308_), .A3(new_n12889_), .ZN(new_n16309_));
  NAND2_X1   g16117(.A1(new_n16309_), .A2(new_n16239_), .ZN(new_n16310_));
  NAND2_X1   g16118(.A1(new_n16306_), .A2(new_n16308_), .ZN(new_n16311_));
  AOI21_X1   g16119(.A1(new_n16311_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n16312_));
  AOI21_X1   g16120(.A1(new_n16312_), .A2(new_n16310_), .B(new_n16288_), .ZN(new_n16313_));
  AOI21_X1   g16121(.A1(new_n16310_), .A2(new_n16278_), .B(new_n12374_), .ZN(new_n16314_));
  OAI21_X1   g16122(.A1(new_n16313_), .A2(new_n16314_), .B(\asqrt[16] ), .ZN(new_n16315_));
  AOI21_X1   g16123(.A1(new_n16284_), .A2(new_n16315_), .B(new_n11406_), .ZN(new_n16316_));
  NOR2_X1    g16124(.A1(new_n16287_), .A2(new_n16316_), .ZN(new_n16317_));
  AOI21_X1   g16125(.A1(new_n16317_), .A2(new_n10953_), .B(new_n16228_), .ZN(new_n16318_));
  OAI21_X1   g16126(.A1(new_n16287_), .A2(new_n16316_), .B(\asqrt[18] ), .ZN(new_n16319_));
  NAND2_X1   g16127(.A1(new_n16319_), .A2(new_n10478_), .ZN(new_n16320_));
  OAI21_X1   g16128(.A1(new_n16318_), .A2(new_n16320_), .B(new_n16224_), .ZN(new_n16321_));
  INV_X1     g16129(.I(new_n16319_), .ZN(new_n16322_));
  OAI21_X1   g16130(.A1(new_n16318_), .A2(new_n16322_), .B(\asqrt[19] ), .ZN(new_n16323_));
  NAND3_X1   g16131(.A1(new_n16321_), .A2(new_n16323_), .A3(new_n10045_), .ZN(new_n16324_));
  NAND2_X1   g16132(.A1(new_n16324_), .A2(new_n16222_), .ZN(new_n16325_));
  NAND2_X1   g16133(.A1(new_n16321_), .A2(new_n16323_), .ZN(new_n16326_));
  AOI21_X1   g16134(.A1(new_n16326_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n16327_));
  AOI21_X1   g16135(.A1(new_n16327_), .A2(new_n16325_), .B(new_n16219_), .ZN(new_n16328_));
  INV_X1     g16136(.I(new_n16224_), .ZN(new_n16329_));
  INV_X1     g16137(.I(new_n16234_), .ZN(new_n16330_));
  NOR2_X1    g16138(.A1(new_n16313_), .A2(new_n16314_), .ZN(new_n16331_));
  AOI21_X1   g16139(.A1(new_n16331_), .A2(new_n11901_), .B(new_n16330_), .ZN(new_n16332_));
  NAND2_X1   g16140(.A1(new_n16315_), .A2(new_n11406_), .ZN(new_n16333_));
  OAI21_X1   g16141(.A1(new_n16332_), .A2(new_n16333_), .B(new_n16230_), .ZN(new_n16334_));
  INV_X1     g16142(.I(new_n16315_), .ZN(new_n16335_));
  OAI21_X1   g16143(.A1(new_n16332_), .A2(new_n16335_), .B(\asqrt[17] ), .ZN(new_n16336_));
  NAND3_X1   g16144(.A1(new_n16334_), .A2(new_n16336_), .A3(new_n10953_), .ZN(new_n16337_));
  NAND2_X1   g16145(.A1(new_n16337_), .A2(new_n16227_), .ZN(new_n16338_));
  NAND2_X1   g16146(.A1(new_n16334_), .A2(new_n16336_), .ZN(new_n16339_));
  AOI21_X1   g16147(.A1(new_n16339_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n16340_));
  AOI21_X1   g16148(.A1(new_n16340_), .A2(new_n16338_), .B(new_n16329_), .ZN(new_n16341_));
  AOI21_X1   g16149(.A1(new_n16338_), .A2(new_n16319_), .B(new_n10478_), .ZN(new_n16342_));
  OAI21_X1   g16150(.A1(new_n16341_), .A2(new_n16342_), .B(\asqrt[20] ), .ZN(new_n16343_));
  AOI21_X1   g16151(.A1(new_n16325_), .A2(new_n16343_), .B(new_n9590_), .ZN(new_n16344_));
  NOR2_X1    g16152(.A1(new_n16328_), .A2(new_n16344_), .ZN(new_n16345_));
  AOI21_X1   g16153(.A1(new_n16345_), .A2(new_n9177_), .B(new_n16216_), .ZN(new_n16346_));
  OAI21_X1   g16154(.A1(new_n16328_), .A2(new_n16344_), .B(\asqrt[22] ), .ZN(new_n16347_));
  NAND2_X1   g16155(.A1(new_n16347_), .A2(new_n8742_), .ZN(new_n16348_));
  OAI21_X1   g16156(.A1(new_n16346_), .A2(new_n16348_), .B(new_n16212_), .ZN(new_n16349_));
  INV_X1     g16157(.I(new_n16347_), .ZN(new_n16350_));
  OAI21_X1   g16158(.A1(new_n16346_), .A2(new_n16350_), .B(\asqrt[23] ), .ZN(new_n16351_));
  NAND3_X1   g16159(.A1(new_n16349_), .A2(new_n16351_), .A3(new_n8349_), .ZN(new_n16352_));
  NAND2_X1   g16160(.A1(new_n16352_), .A2(new_n16210_), .ZN(new_n16353_));
  NAND2_X1   g16161(.A1(new_n16349_), .A2(new_n16351_), .ZN(new_n16354_));
  AOI21_X1   g16162(.A1(new_n16354_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n16355_));
  AOI21_X1   g16163(.A1(new_n16355_), .A2(new_n16353_), .B(new_n16207_), .ZN(new_n16356_));
  INV_X1     g16164(.I(new_n16212_), .ZN(new_n16357_));
  INV_X1     g16165(.I(new_n16222_), .ZN(new_n16358_));
  NOR2_X1    g16166(.A1(new_n16341_), .A2(new_n16342_), .ZN(new_n16359_));
  AOI21_X1   g16167(.A1(new_n16359_), .A2(new_n10045_), .B(new_n16358_), .ZN(new_n16360_));
  NAND2_X1   g16168(.A1(new_n16343_), .A2(new_n9590_), .ZN(new_n16361_));
  OAI21_X1   g16169(.A1(new_n16360_), .A2(new_n16361_), .B(new_n16218_), .ZN(new_n16362_));
  INV_X1     g16170(.I(new_n16343_), .ZN(new_n16363_));
  OAI21_X1   g16171(.A1(new_n16360_), .A2(new_n16363_), .B(\asqrt[21] ), .ZN(new_n16364_));
  NAND3_X1   g16172(.A1(new_n16362_), .A2(new_n16364_), .A3(new_n9177_), .ZN(new_n16365_));
  NAND2_X1   g16173(.A1(new_n16365_), .A2(new_n16215_), .ZN(new_n16366_));
  NAND2_X1   g16174(.A1(new_n16362_), .A2(new_n16364_), .ZN(new_n16367_));
  AOI21_X1   g16175(.A1(new_n16367_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n16368_));
  AOI21_X1   g16176(.A1(new_n16368_), .A2(new_n16366_), .B(new_n16357_), .ZN(new_n16369_));
  AOI21_X1   g16177(.A1(new_n16366_), .A2(new_n16347_), .B(new_n8742_), .ZN(new_n16370_));
  OAI21_X1   g16178(.A1(new_n16369_), .A2(new_n16370_), .B(\asqrt[24] ), .ZN(new_n16371_));
  AOI21_X1   g16179(.A1(new_n16353_), .A2(new_n16371_), .B(new_n7934_), .ZN(new_n16372_));
  NOR2_X1    g16180(.A1(new_n16356_), .A2(new_n16372_), .ZN(new_n16373_));
  AOI21_X1   g16181(.A1(new_n16373_), .A2(new_n7561_), .B(new_n16204_), .ZN(new_n16374_));
  OAI21_X1   g16182(.A1(new_n16356_), .A2(new_n16372_), .B(\asqrt[26] ), .ZN(new_n16375_));
  NAND2_X1   g16183(.A1(new_n16375_), .A2(new_n7166_), .ZN(new_n16376_));
  OAI21_X1   g16184(.A1(new_n16374_), .A2(new_n16376_), .B(new_n16200_), .ZN(new_n16377_));
  INV_X1     g16185(.I(new_n16375_), .ZN(new_n16378_));
  OAI21_X1   g16186(.A1(new_n16374_), .A2(new_n16378_), .B(\asqrt[27] ), .ZN(new_n16379_));
  NAND3_X1   g16187(.A1(new_n16377_), .A2(new_n16379_), .A3(new_n6813_), .ZN(new_n16380_));
  NAND2_X1   g16188(.A1(new_n16380_), .A2(new_n16198_), .ZN(new_n16381_));
  NAND2_X1   g16189(.A1(new_n16377_), .A2(new_n16379_), .ZN(new_n16382_));
  AOI21_X1   g16190(.A1(new_n16382_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n16383_));
  AOI21_X1   g16191(.A1(new_n16383_), .A2(new_n16381_), .B(new_n16195_), .ZN(new_n16384_));
  INV_X1     g16192(.I(new_n16200_), .ZN(new_n16385_));
  INV_X1     g16193(.I(new_n16210_), .ZN(new_n16386_));
  NOR2_X1    g16194(.A1(new_n16369_), .A2(new_n16370_), .ZN(new_n16387_));
  AOI21_X1   g16195(.A1(new_n16387_), .A2(new_n8349_), .B(new_n16386_), .ZN(new_n16388_));
  NAND2_X1   g16196(.A1(new_n16371_), .A2(new_n7934_), .ZN(new_n16389_));
  OAI21_X1   g16197(.A1(new_n16388_), .A2(new_n16389_), .B(new_n16206_), .ZN(new_n16390_));
  INV_X1     g16198(.I(new_n16371_), .ZN(new_n16391_));
  OAI21_X1   g16199(.A1(new_n16388_), .A2(new_n16391_), .B(\asqrt[25] ), .ZN(new_n16392_));
  NAND3_X1   g16200(.A1(new_n16390_), .A2(new_n16392_), .A3(new_n7561_), .ZN(new_n16393_));
  NAND2_X1   g16201(.A1(new_n16393_), .A2(new_n16203_), .ZN(new_n16394_));
  NAND2_X1   g16202(.A1(new_n16390_), .A2(new_n16392_), .ZN(new_n16395_));
  AOI21_X1   g16203(.A1(new_n16395_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n16396_));
  AOI21_X1   g16204(.A1(new_n16396_), .A2(new_n16394_), .B(new_n16385_), .ZN(new_n16397_));
  AOI21_X1   g16205(.A1(new_n16394_), .A2(new_n16375_), .B(new_n7166_), .ZN(new_n16398_));
  OAI21_X1   g16206(.A1(new_n16397_), .A2(new_n16398_), .B(\asqrt[28] ), .ZN(new_n16399_));
  AOI21_X1   g16207(.A1(new_n16381_), .A2(new_n16399_), .B(new_n6454_), .ZN(new_n16400_));
  NOR2_X1    g16208(.A1(new_n16384_), .A2(new_n16400_), .ZN(new_n16401_));
  AOI21_X1   g16209(.A1(new_n16401_), .A2(new_n6106_), .B(new_n16192_), .ZN(new_n16402_));
  OAI21_X1   g16210(.A1(new_n16384_), .A2(new_n16400_), .B(\asqrt[30] ), .ZN(new_n16403_));
  NAND2_X1   g16211(.A1(new_n16403_), .A2(new_n5750_), .ZN(new_n16404_));
  OAI21_X1   g16212(.A1(new_n16402_), .A2(new_n16404_), .B(new_n16188_), .ZN(new_n16405_));
  INV_X1     g16213(.I(new_n16403_), .ZN(new_n16406_));
  OAI21_X1   g16214(.A1(new_n16402_), .A2(new_n16406_), .B(\asqrt[31] ), .ZN(new_n16407_));
  NAND3_X1   g16215(.A1(new_n16405_), .A2(new_n16407_), .A3(new_n5435_), .ZN(new_n16408_));
  NAND2_X1   g16216(.A1(new_n16408_), .A2(new_n16186_), .ZN(new_n16409_));
  NAND2_X1   g16217(.A1(new_n16405_), .A2(new_n16407_), .ZN(new_n16410_));
  AOI21_X1   g16218(.A1(new_n16410_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n16411_));
  AOI21_X1   g16219(.A1(new_n16411_), .A2(new_n16409_), .B(new_n16183_), .ZN(new_n16412_));
  INV_X1     g16220(.I(new_n16188_), .ZN(new_n16413_));
  INV_X1     g16221(.I(new_n16198_), .ZN(new_n16414_));
  NOR2_X1    g16222(.A1(new_n16397_), .A2(new_n16398_), .ZN(new_n16415_));
  AOI21_X1   g16223(.A1(new_n16415_), .A2(new_n6813_), .B(new_n16414_), .ZN(new_n16416_));
  NAND2_X1   g16224(.A1(new_n16399_), .A2(new_n6454_), .ZN(new_n16417_));
  OAI21_X1   g16225(.A1(new_n16416_), .A2(new_n16417_), .B(new_n16194_), .ZN(new_n16418_));
  INV_X1     g16226(.I(new_n16399_), .ZN(new_n16419_));
  OAI21_X1   g16227(.A1(new_n16416_), .A2(new_n16419_), .B(\asqrt[29] ), .ZN(new_n16420_));
  NAND3_X1   g16228(.A1(new_n16418_), .A2(new_n16420_), .A3(new_n6106_), .ZN(new_n16421_));
  NAND2_X1   g16229(.A1(new_n16421_), .A2(new_n16191_), .ZN(new_n16422_));
  NAND2_X1   g16230(.A1(new_n16418_), .A2(new_n16420_), .ZN(new_n16423_));
  AOI21_X1   g16231(.A1(new_n16423_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n16424_));
  AOI21_X1   g16232(.A1(new_n16424_), .A2(new_n16422_), .B(new_n16413_), .ZN(new_n16425_));
  AOI21_X1   g16233(.A1(new_n16422_), .A2(new_n16403_), .B(new_n5750_), .ZN(new_n16426_));
  OAI21_X1   g16234(.A1(new_n16425_), .A2(new_n16426_), .B(\asqrt[32] ), .ZN(new_n16427_));
  AOI21_X1   g16235(.A1(new_n16409_), .A2(new_n16427_), .B(new_n5110_), .ZN(new_n16428_));
  NOR2_X1    g16236(.A1(new_n16412_), .A2(new_n16428_), .ZN(new_n16429_));
  AOI21_X1   g16237(.A1(new_n16429_), .A2(new_n4810_), .B(new_n16180_), .ZN(new_n16430_));
  OAI21_X1   g16238(.A1(new_n16412_), .A2(new_n16428_), .B(\asqrt[34] ), .ZN(new_n16431_));
  NAND2_X1   g16239(.A1(new_n16431_), .A2(new_n4510_), .ZN(new_n16432_));
  OAI21_X1   g16240(.A1(new_n16430_), .A2(new_n16432_), .B(new_n16176_), .ZN(new_n16433_));
  INV_X1     g16241(.I(new_n16431_), .ZN(new_n16434_));
  OAI21_X1   g16242(.A1(new_n16430_), .A2(new_n16434_), .B(\asqrt[35] ), .ZN(new_n16435_));
  NAND3_X1   g16243(.A1(new_n16433_), .A2(new_n16435_), .A3(new_n4224_), .ZN(new_n16436_));
  NAND2_X1   g16244(.A1(new_n16436_), .A2(new_n16174_), .ZN(new_n16437_));
  NAND2_X1   g16245(.A1(new_n16433_), .A2(new_n16435_), .ZN(new_n16438_));
  AOI21_X1   g16246(.A1(new_n16438_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n16439_));
  AOI21_X1   g16247(.A1(new_n16439_), .A2(new_n16437_), .B(new_n16171_), .ZN(new_n16440_));
  INV_X1     g16248(.I(new_n16176_), .ZN(new_n16441_));
  INV_X1     g16249(.I(new_n16186_), .ZN(new_n16442_));
  NOR2_X1    g16250(.A1(new_n16425_), .A2(new_n16426_), .ZN(new_n16443_));
  AOI21_X1   g16251(.A1(new_n16443_), .A2(new_n5435_), .B(new_n16442_), .ZN(new_n16444_));
  NAND2_X1   g16252(.A1(new_n16427_), .A2(new_n5110_), .ZN(new_n16445_));
  OAI21_X1   g16253(.A1(new_n16444_), .A2(new_n16445_), .B(new_n16182_), .ZN(new_n16446_));
  INV_X1     g16254(.I(new_n16427_), .ZN(new_n16447_));
  OAI21_X1   g16255(.A1(new_n16444_), .A2(new_n16447_), .B(\asqrt[33] ), .ZN(new_n16448_));
  NAND3_X1   g16256(.A1(new_n16446_), .A2(new_n16448_), .A3(new_n4810_), .ZN(new_n16449_));
  NAND2_X1   g16257(.A1(new_n16449_), .A2(new_n16179_), .ZN(new_n16450_));
  NAND2_X1   g16258(.A1(new_n16446_), .A2(new_n16448_), .ZN(new_n16451_));
  AOI21_X1   g16259(.A1(new_n16451_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n16452_));
  AOI21_X1   g16260(.A1(new_n16452_), .A2(new_n16450_), .B(new_n16441_), .ZN(new_n16453_));
  AOI21_X1   g16261(.A1(new_n16450_), .A2(new_n16431_), .B(new_n4510_), .ZN(new_n16454_));
  OAI21_X1   g16262(.A1(new_n16453_), .A2(new_n16454_), .B(\asqrt[36] ), .ZN(new_n16455_));
  AOI21_X1   g16263(.A1(new_n16437_), .A2(new_n16455_), .B(new_n3928_), .ZN(new_n16456_));
  NOR2_X1    g16264(.A1(new_n16440_), .A2(new_n16456_), .ZN(new_n16457_));
  AOI21_X1   g16265(.A1(new_n16457_), .A2(new_n3675_), .B(new_n16168_), .ZN(new_n16458_));
  OAI21_X1   g16266(.A1(new_n16440_), .A2(new_n16456_), .B(\asqrt[38] ), .ZN(new_n16459_));
  NAND2_X1   g16267(.A1(new_n16459_), .A2(new_n3400_), .ZN(new_n16460_));
  OAI21_X1   g16268(.A1(new_n16458_), .A2(new_n16460_), .B(new_n16164_), .ZN(new_n16461_));
  INV_X1     g16269(.I(new_n16459_), .ZN(new_n16462_));
  OAI21_X1   g16270(.A1(new_n16458_), .A2(new_n16462_), .B(\asqrt[39] ), .ZN(new_n16463_));
  NAND3_X1   g16271(.A1(new_n16461_), .A2(new_n16463_), .A3(new_n3167_), .ZN(new_n16464_));
  NAND2_X1   g16272(.A1(new_n16464_), .A2(new_n16162_), .ZN(new_n16465_));
  NAND2_X1   g16273(.A1(new_n16461_), .A2(new_n16463_), .ZN(new_n16466_));
  AOI21_X1   g16274(.A1(new_n16466_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n16467_));
  AOI21_X1   g16275(.A1(new_n16467_), .A2(new_n16465_), .B(new_n16159_), .ZN(new_n16468_));
  INV_X1     g16276(.I(new_n16164_), .ZN(new_n16469_));
  INV_X1     g16277(.I(new_n16174_), .ZN(new_n16470_));
  NOR2_X1    g16278(.A1(new_n16453_), .A2(new_n16454_), .ZN(new_n16471_));
  AOI21_X1   g16279(.A1(new_n16471_), .A2(new_n4224_), .B(new_n16470_), .ZN(new_n16472_));
  NAND2_X1   g16280(.A1(new_n16455_), .A2(new_n3928_), .ZN(new_n16473_));
  OAI21_X1   g16281(.A1(new_n16472_), .A2(new_n16473_), .B(new_n16170_), .ZN(new_n16474_));
  INV_X1     g16282(.I(new_n16455_), .ZN(new_n16475_));
  OAI21_X1   g16283(.A1(new_n16472_), .A2(new_n16475_), .B(\asqrt[37] ), .ZN(new_n16476_));
  NAND3_X1   g16284(.A1(new_n16474_), .A2(new_n16476_), .A3(new_n3675_), .ZN(new_n16477_));
  NAND2_X1   g16285(.A1(new_n16477_), .A2(new_n16167_), .ZN(new_n16478_));
  NAND2_X1   g16286(.A1(new_n16474_), .A2(new_n16476_), .ZN(new_n16479_));
  AOI21_X1   g16287(.A1(new_n16479_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n16480_));
  AOI21_X1   g16288(.A1(new_n16480_), .A2(new_n16478_), .B(new_n16469_), .ZN(new_n16481_));
  AOI21_X1   g16289(.A1(new_n16478_), .A2(new_n16459_), .B(new_n3400_), .ZN(new_n16482_));
  OAI21_X1   g16290(.A1(new_n16481_), .A2(new_n16482_), .B(\asqrt[40] ), .ZN(new_n16483_));
  AOI21_X1   g16291(.A1(new_n16465_), .A2(new_n16483_), .B(new_n2912_), .ZN(new_n16484_));
  NOR2_X1    g16292(.A1(new_n16468_), .A2(new_n16484_), .ZN(new_n16485_));
  AOI21_X1   g16293(.A1(new_n16485_), .A2(new_n2699_), .B(new_n16156_), .ZN(new_n16486_));
  OAI21_X1   g16294(.A1(new_n16468_), .A2(new_n16484_), .B(\asqrt[42] ), .ZN(new_n16487_));
  NAND2_X1   g16295(.A1(new_n16487_), .A2(new_n2464_), .ZN(new_n16488_));
  OAI21_X1   g16296(.A1(new_n16486_), .A2(new_n16488_), .B(new_n16152_), .ZN(new_n16489_));
  INV_X1     g16297(.I(new_n16487_), .ZN(new_n16490_));
  OAI21_X1   g16298(.A1(new_n16486_), .A2(new_n16490_), .B(\asqrt[43] ), .ZN(new_n16491_));
  NAND3_X1   g16299(.A1(new_n16489_), .A2(new_n16491_), .A3(new_n2271_), .ZN(new_n16492_));
  NAND2_X1   g16300(.A1(new_n16492_), .A2(new_n16150_), .ZN(new_n16493_));
  NAND2_X1   g16301(.A1(new_n16489_), .A2(new_n16491_), .ZN(new_n16494_));
  AOI21_X1   g16302(.A1(new_n16494_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n16495_));
  AOI21_X1   g16303(.A1(new_n16495_), .A2(new_n16493_), .B(new_n16147_), .ZN(new_n16496_));
  INV_X1     g16304(.I(new_n16152_), .ZN(new_n16497_));
  INV_X1     g16305(.I(new_n16162_), .ZN(new_n16498_));
  NOR2_X1    g16306(.A1(new_n16481_), .A2(new_n16482_), .ZN(new_n16499_));
  AOI21_X1   g16307(.A1(new_n16499_), .A2(new_n3167_), .B(new_n16498_), .ZN(new_n16500_));
  NAND2_X1   g16308(.A1(new_n16483_), .A2(new_n2912_), .ZN(new_n16501_));
  OAI21_X1   g16309(.A1(new_n16500_), .A2(new_n16501_), .B(new_n16158_), .ZN(new_n16502_));
  INV_X1     g16310(.I(new_n16483_), .ZN(new_n16503_));
  OAI21_X1   g16311(.A1(new_n16500_), .A2(new_n16503_), .B(\asqrt[41] ), .ZN(new_n16504_));
  NAND3_X1   g16312(.A1(new_n16502_), .A2(new_n16504_), .A3(new_n2699_), .ZN(new_n16505_));
  NAND2_X1   g16313(.A1(new_n16505_), .A2(new_n16155_), .ZN(new_n16506_));
  NAND2_X1   g16314(.A1(new_n16502_), .A2(new_n16504_), .ZN(new_n16507_));
  AOI21_X1   g16315(.A1(new_n16507_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n16508_));
  AOI21_X1   g16316(.A1(new_n16508_), .A2(new_n16506_), .B(new_n16497_), .ZN(new_n16509_));
  AOI21_X1   g16317(.A1(new_n16506_), .A2(new_n16487_), .B(new_n2464_), .ZN(new_n16510_));
  OAI21_X1   g16318(.A1(new_n16509_), .A2(new_n16510_), .B(\asqrt[44] ), .ZN(new_n16511_));
  AOI21_X1   g16319(.A1(new_n16493_), .A2(new_n16511_), .B(new_n2072_), .ZN(new_n16512_));
  NOR2_X1    g16320(.A1(new_n16496_), .A2(new_n16512_), .ZN(new_n16513_));
  AOI21_X1   g16321(.A1(new_n16513_), .A2(new_n1884_), .B(new_n16144_), .ZN(new_n16514_));
  OAI21_X1   g16322(.A1(new_n16496_), .A2(new_n16512_), .B(\asqrt[46] ), .ZN(new_n16515_));
  NAND2_X1   g16323(.A1(new_n16515_), .A2(new_n1688_), .ZN(new_n16516_));
  OAI21_X1   g16324(.A1(new_n16514_), .A2(new_n16516_), .B(new_n16140_), .ZN(new_n16517_));
  INV_X1     g16325(.I(new_n16515_), .ZN(new_n16518_));
  OAI21_X1   g16326(.A1(new_n16514_), .A2(new_n16518_), .B(\asqrt[47] ), .ZN(new_n16519_));
  NAND3_X1   g16327(.A1(new_n16517_), .A2(new_n16519_), .A3(new_n1533_), .ZN(new_n16520_));
  NAND2_X1   g16328(.A1(new_n16520_), .A2(new_n16138_), .ZN(new_n16521_));
  NAND2_X1   g16329(.A1(new_n16517_), .A2(new_n16519_), .ZN(new_n16522_));
  AOI21_X1   g16330(.A1(new_n16522_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n16523_));
  AOI21_X1   g16331(.A1(new_n16523_), .A2(new_n16521_), .B(new_n16135_), .ZN(new_n16524_));
  INV_X1     g16332(.I(new_n16140_), .ZN(new_n16525_));
  INV_X1     g16333(.I(new_n16150_), .ZN(new_n16526_));
  NOR2_X1    g16334(.A1(new_n16509_), .A2(new_n16510_), .ZN(new_n16527_));
  AOI21_X1   g16335(.A1(new_n16527_), .A2(new_n2271_), .B(new_n16526_), .ZN(new_n16528_));
  NAND2_X1   g16336(.A1(new_n16511_), .A2(new_n2072_), .ZN(new_n16529_));
  OAI21_X1   g16337(.A1(new_n16528_), .A2(new_n16529_), .B(new_n16146_), .ZN(new_n16530_));
  INV_X1     g16338(.I(new_n16511_), .ZN(new_n16531_));
  OAI21_X1   g16339(.A1(new_n16528_), .A2(new_n16531_), .B(\asqrt[45] ), .ZN(new_n16532_));
  NAND3_X1   g16340(.A1(new_n16530_), .A2(new_n16532_), .A3(new_n1884_), .ZN(new_n16533_));
  NAND2_X1   g16341(.A1(new_n16533_), .A2(new_n16143_), .ZN(new_n16534_));
  NAND2_X1   g16342(.A1(new_n16530_), .A2(new_n16532_), .ZN(new_n16535_));
  AOI21_X1   g16343(.A1(new_n16535_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n16536_));
  AOI21_X1   g16344(.A1(new_n16536_), .A2(new_n16534_), .B(new_n16525_), .ZN(new_n16537_));
  AOI21_X1   g16345(.A1(new_n16534_), .A2(new_n16515_), .B(new_n1688_), .ZN(new_n16538_));
  OAI21_X1   g16346(.A1(new_n16537_), .A2(new_n16538_), .B(\asqrt[48] ), .ZN(new_n16539_));
  AOI21_X1   g16347(.A1(new_n16521_), .A2(new_n16539_), .B(new_n1368_), .ZN(new_n16540_));
  NOR2_X1    g16348(.A1(new_n16524_), .A2(new_n16540_), .ZN(new_n16541_));
  AOI21_X1   g16349(.A1(new_n16541_), .A2(new_n1228_), .B(new_n16132_), .ZN(new_n16542_));
  OAI21_X1   g16350(.A1(new_n16524_), .A2(new_n16540_), .B(\asqrt[50] ), .ZN(new_n16543_));
  NAND2_X1   g16351(.A1(new_n16543_), .A2(new_n1088_), .ZN(new_n16544_));
  OAI21_X1   g16352(.A1(new_n16542_), .A2(new_n16544_), .B(new_n16128_), .ZN(new_n16545_));
  INV_X1     g16353(.I(new_n16543_), .ZN(new_n16546_));
  OAI21_X1   g16354(.A1(new_n16542_), .A2(new_n16546_), .B(\asqrt[51] ), .ZN(new_n16547_));
  NAND3_X1   g16355(.A1(new_n16545_), .A2(new_n16547_), .A3(new_n962_), .ZN(new_n16548_));
  NAND2_X1   g16356(.A1(new_n16548_), .A2(new_n16126_), .ZN(new_n16549_));
  NAND2_X1   g16357(.A1(new_n16545_), .A2(new_n16547_), .ZN(new_n16550_));
  AOI21_X1   g16358(.A1(new_n16550_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n16551_));
  AOI21_X1   g16359(.A1(new_n16551_), .A2(new_n16549_), .B(new_n16123_), .ZN(new_n16552_));
  INV_X1     g16360(.I(new_n16128_), .ZN(new_n16553_));
  INV_X1     g16361(.I(new_n16138_), .ZN(new_n16554_));
  NOR2_X1    g16362(.A1(new_n16537_), .A2(new_n16538_), .ZN(new_n16555_));
  AOI21_X1   g16363(.A1(new_n16555_), .A2(new_n1533_), .B(new_n16554_), .ZN(new_n16556_));
  NAND2_X1   g16364(.A1(new_n16539_), .A2(new_n1368_), .ZN(new_n16557_));
  OAI21_X1   g16365(.A1(new_n16556_), .A2(new_n16557_), .B(new_n16134_), .ZN(new_n16558_));
  INV_X1     g16366(.I(new_n16539_), .ZN(new_n16559_));
  OAI21_X1   g16367(.A1(new_n16556_), .A2(new_n16559_), .B(\asqrt[49] ), .ZN(new_n16560_));
  NAND3_X1   g16368(.A1(new_n16558_), .A2(new_n16560_), .A3(new_n1228_), .ZN(new_n16561_));
  NAND2_X1   g16369(.A1(new_n16561_), .A2(new_n16131_), .ZN(new_n16562_));
  NAND2_X1   g16370(.A1(new_n16558_), .A2(new_n16560_), .ZN(new_n16563_));
  AOI21_X1   g16371(.A1(new_n16563_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n16564_));
  AOI21_X1   g16372(.A1(new_n16564_), .A2(new_n16562_), .B(new_n16553_), .ZN(new_n16565_));
  AOI21_X1   g16373(.A1(new_n16562_), .A2(new_n16543_), .B(new_n1088_), .ZN(new_n16566_));
  OAI21_X1   g16374(.A1(new_n16565_), .A2(new_n16566_), .B(\asqrt[52] ), .ZN(new_n16567_));
  AOI21_X1   g16375(.A1(new_n16549_), .A2(new_n16567_), .B(new_n842_), .ZN(new_n16568_));
  NOR2_X1    g16376(.A1(new_n16552_), .A2(new_n16568_), .ZN(new_n16569_));
  AOI21_X1   g16377(.A1(new_n16569_), .A2(new_n720_), .B(new_n16120_), .ZN(new_n16570_));
  OAI21_X1   g16378(.A1(new_n16552_), .A2(new_n16568_), .B(\asqrt[54] ), .ZN(new_n16571_));
  NAND2_X1   g16379(.A1(new_n16571_), .A2(new_n630_), .ZN(new_n16572_));
  OAI21_X1   g16380(.A1(new_n16570_), .A2(new_n16572_), .B(new_n16116_), .ZN(new_n16573_));
  INV_X1     g16381(.I(new_n16571_), .ZN(new_n16574_));
  OAI21_X1   g16382(.A1(new_n16570_), .A2(new_n16574_), .B(\asqrt[55] ), .ZN(new_n16575_));
  NAND3_X1   g16383(.A1(new_n16573_), .A2(new_n16575_), .A3(new_n545_), .ZN(new_n16576_));
  NAND2_X1   g16384(.A1(new_n16576_), .A2(new_n16114_), .ZN(new_n16577_));
  NAND2_X1   g16385(.A1(new_n16573_), .A2(new_n16575_), .ZN(new_n16578_));
  AOI21_X1   g16386(.A1(new_n16578_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n16579_));
  AOI21_X1   g16387(.A1(new_n16579_), .A2(new_n16577_), .B(new_n16111_), .ZN(new_n16580_));
  INV_X1     g16388(.I(new_n16116_), .ZN(new_n16581_));
  INV_X1     g16389(.I(new_n16126_), .ZN(new_n16582_));
  NOR2_X1    g16390(.A1(new_n16565_), .A2(new_n16566_), .ZN(new_n16583_));
  AOI21_X1   g16391(.A1(new_n16583_), .A2(new_n962_), .B(new_n16582_), .ZN(new_n16584_));
  NAND2_X1   g16392(.A1(new_n16567_), .A2(new_n842_), .ZN(new_n16585_));
  OAI21_X1   g16393(.A1(new_n16584_), .A2(new_n16585_), .B(new_n16122_), .ZN(new_n16586_));
  INV_X1     g16394(.I(new_n16567_), .ZN(new_n16587_));
  OAI21_X1   g16395(.A1(new_n16584_), .A2(new_n16587_), .B(\asqrt[53] ), .ZN(new_n16588_));
  NAND3_X1   g16396(.A1(new_n16586_), .A2(new_n16588_), .A3(new_n720_), .ZN(new_n16589_));
  NAND2_X1   g16397(.A1(new_n16589_), .A2(new_n16119_), .ZN(new_n16590_));
  NAND2_X1   g16398(.A1(new_n16586_), .A2(new_n16588_), .ZN(new_n16591_));
  AOI21_X1   g16399(.A1(new_n16591_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n16592_));
  AOI21_X1   g16400(.A1(new_n16592_), .A2(new_n16590_), .B(new_n16581_), .ZN(new_n16593_));
  AOI21_X1   g16401(.A1(new_n16590_), .A2(new_n16571_), .B(new_n630_), .ZN(new_n16594_));
  OAI21_X1   g16402(.A1(new_n16593_), .A2(new_n16594_), .B(\asqrt[56] ), .ZN(new_n16595_));
  AOI21_X1   g16403(.A1(new_n16577_), .A2(new_n16595_), .B(new_n450_), .ZN(new_n16596_));
  NOR2_X1    g16404(.A1(new_n16580_), .A2(new_n16596_), .ZN(new_n16597_));
  AOI21_X1   g16405(.A1(new_n16597_), .A2(new_n403_), .B(new_n16110_), .ZN(new_n16598_));
  OAI21_X1   g16406(.A1(new_n16580_), .A2(new_n16596_), .B(\asqrt[58] ), .ZN(new_n16599_));
  NAND2_X1   g16407(.A1(new_n16599_), .A2(new_n339_), .ZN(new_n16600_));
  OAI21_X1   g16408(.A1(new_n16598_), .A2(new_n16600_), .B(new_n16106_), .ZN(new_n16601_));
  INV_X1     g16409(.I(new_n16599_), .ZN(new_n16602_));
  OAI21_X1   g16410(.A1(new_n16598_), .A2(new_n16602_), .B(\asqrt[59] ), .ZN(new_n16603_));
  NAND3_X1   g16411(.A1(new_n16601_), .A2(new_n16603_), .A3(new_n288_), .ZN(new_n16604_));
  NAND2_X1   g16412(.A1(new_n16604_), .A2(new_n16104_), .ZN(new_n16605_));
  INV_X1     g16413(.I(new_n16106_), .ZN(new_n16606_));
  INV_X1     g16414(.I(new_n16114_), .ZN(new_n16607_));
  NOR2_X1    g16415(.A1(new_n16593_), .A2(new_n16594_), .ZN(new_n16608_));
  AOI21_X1   g16416(.A1(new_n16608_), .A2(new_n545_), .B(new_n16607_), .ZN(new_n16609_));
  NAND2_X1   g16417(.A1(new_n16595_), .A2(new_n450_), .ZN(new_n16610_));
  OAI21_X1   g16418(.A1(new_n16609_), .A2(new_n16610_), .B(new_n16076_), .ZN(new_n16611_));
  INV_X1     g16419(.I(new_n16595_), .ZN(new_n16612_));
  OAI21_X1   g16420(.A1(new_n16609_), .A2(new_n16612_), .B(\asqrt[57] ), .ZN(new_n16613_));
  NAND3_X1   g16421(.A1(new_n16611_), .A2(new_n16613_), .A3(new_n403_), .ZN(new_n16614_));
  NAND2_X1   g16422(.A1(new_n16614_), .A2(new_n16109_), .ZN(new_n16615_));
  NAND2_X1   g16423(.A1(new_n16611_), .A2(new_n16613_), .ZN(new_n16616_));
  AOI21_X1   g16424(.A1(new_n16616_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n16617_));
  AOI21_X1   g16425(.A1(new_n16617_), .A2(new_n16615_), .B(new_n16606_), .ZN(new_n16618_));
  AOI21_X1   g16426(.A1(new_n16615_), .A2(new_n16599_), .B(new_n339_), .ZN(new_n16619_));
  OAI21_X1   g16427(.A1(new_n16618_), .A2(new_n16619_), .B(\asqrt[60] ), .ZN(new_n16620_));
  AOI21_X1   g16428(.A1(new_n16605_), .A2(new_n16620_), .B(new_n242_), .ZN(new_n16621_));
  NAND3_X1   g16429(.A1(\asqrt[8] ), .A2(new_n16037_), .A3(new_n16052_), .ZN(new_n16622_));
  XOR2_X1    g16430(.A1(new_n16622_), .A2(new_n16077_), .Z(new_n16623_));
  INV_X1     g16431(.I(new_n16623_), .ZN(new_n16624_));
  NAND2_X1   g16432(.A1(new_n16601_), .A2(new_n16603_), .ZN(new_n16625_));
  AOI21_X1   g16433(.A1(new_n16625_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n16626_));
  AOI21_X1   g16434(.A1(new_n16626_), .A2(new_n16605_), .B(new_n16624_), .ZN(new_n16627_));
  OAI21_X1   g16435(.A1(new_n16627_), .A2(new_n16621_), .B(\asqrt[62] ), .ZN(new_n16628_));
  AOI21_X1   g16436(.A1(new_n16038_), .A2(new_n16058_), .B(new_n16053_), .ZN(new_n16629_));
  NAND2_X1   g16437(.A1(\asqrt[8] ), .A2(new_n16629_), .ZN(new_n16630_));
  XOR2_X1    g16438(.A1(new_n16630_), .A2(new_n16056_), .Z(new_n16631_));
  INV_X1     g16439(.I(new_n16104_), .ZN(new_n16632_));
  NOR2_X1    g16440(.A1(new_n16618_), .A2(new_n16619_), .ZN(new_n16633_));
  AOI21_X1   g16441(.A1(new_n16633_), .A2(new_n288_), .B(new_n16632_), .ZN(new_n16634_));
  INV_X1     g16442(.I(new_n16620_), .ZN(new_n16635_));
  OAI21_X1   g16443(.A1(new_n16634_), .A2(new_n16635_), .B(\asqrt[61] ), .ZN(new_n16636_));
  NAND2_X1   g16444(.A1(new_n16620_), .A2(new_n242_), .ZN(new_n16637_));
  OAI21_X1   g16445(.A1(new_n16634_), .A2(new_n16637_), .B(new_n16623_), .ZN(new_n16638_));
  NAND3_X1   g16446(.A1(new_n16638_), .A2(new_n16636_), .A3(new_n234_), .ZN(new_n16639_));
  NAND2_X1   g16447(.A1(new_n16639_), .A2(new_n16631_), .ZN(new_n16640_));
  AOI21_X1   g16448(.A1(new_n16640_), .A2(new_n16628_), .B(new_n16101_), .ZN(new_n16641_));
  AOI21_X1   g16449(.A1(new_n16641_), .A2(new_n16099_), .B(\asqrt[63] ), .ZN(new_n16642_));
  INV_X1     g16450(.I(new_n16628_), .ZN(new_n16643_));
  NOR2_X1    g16451(.A1(new_n16627_), .A2(new_n16621_), .ZN(new_n16644_));
  INV_X1     g16452(.I(new_n16631_), .ZN(new_n16645_));
  AOI21_X1   g16453(.A1(new_n16644_), .A2(new_n234_), .B(new_n16645_), .ZN(new_n16646_));
  NOR3_X1    g16454(.A1(new_n16646_), .A2(new_n16643_), .A3(new_n16099_), .ZN(new_n16647_));
  NOR2_X1    g16455(.A1(\asqrt[8] ), .A2(new_n16088_), .ZN(new_n16648_));
  NOR4_X1    g16456(.A1(new_n16642_), .A2(new_n16096_), .A3(new_n16647_), .A4(new_n16648_), .ZN(new_n16649_));
  OAI21_X1   g16457(.A1(new_n16609_), .A2(new_n16610_), .B(new_n16613_), .ZN(new_n16650_));
  NOR2_X1    g16458(.A1(new_n16649_), .A2(new_n16650_), .ZN(new_n16651_));
  XOR2_X1    g16459(.A1(new_n16651_), .A2(new_n16076_), .Z(new_n16652_));
  INV_X1     g16460(.I(new_n16652_), .ZN(new_n16653_));
  INV_X1     g16461(.I(new_n16096_), .ZN(new_n16654_));
  OAI21_X1   g16462(.A1(new_n16646_), .A2(new_n16643_), .B(new_n16100_), .ZN(new_n16655_));
  OAI21_X1   g16463(.A1(new_n16655_), .A2(new_n16098_), .B(new_n193_), .ZN(new_n16656_));
  INV_X1     g16464(.I(new_n16647_), .ZN(new_n16657_));
  INV_X1     g16465(.I(new_n16648_), .ZN(new_n16658_));
  NAND4_X1   g16466(.A1(new_n16656_), .A2(new_n16654_), .A3(new_n16657_), .A4(new_n16658_), .ZN(\asqrt[7] ));
  NAND3_X1   g16467(.A1(\asqrt[7] ), .A2(new_n16576_), .A3(new_n16595_), .ZN(new_n16660_));
  XOR2_X1    g16468(.A1(new_n16660_), .A2(new_n16607_), .Z(new_n16661_));
  OAI21_X1   g16469(.A1(new_n16570_), .A2(new_n16572_), .B(new_n16575_), .ZN(new_n16662_));
  NOR2_X1    g16470(.A1(new_n16649_), .A2(new_n16662_), .ZN(new_n16663_));
  XOR2_X1    g16471(.A1(new_n16663_), .A2(new_n16116_), .Z(new_n16664_));
  INV_X1     g16472(.I(new_n16664_), .ZN(new_n16665_));
  NAND3_X1   g16473(.A1(\asqrt[7] ), .A2(new_n16589_), .A3(new_n16571_), .ZN(new_n16666_));
  XOR2_X1    g16474(.A1(new_n16666_), .A2(new_n16120_), .Z(new_n16667_));
  INV_X1     g16475(.I(new_n16667_), .ZN(new_n16668_));
  OAI21_X1   g16476(.A1(new_n16584_), .A2(new_n16585_), .B(new_n16588_), .ZN(new_n16669_));
  NOR2_X1    g16477(.A1(new_n16649_), .A2(new_n16669_), .ZN(new_n16670_));
  XOR2_X1    g16478(.A1(new_n16670_), .A2(new_n16122_), .Z(new_n16671_));
  NAND3_X1   g16479(.A1(\asqrt[7] ), .A2(new_n16548_), .A3(new_n16567_), .ZN(new_n16672_));
  XOR2_X1    g16480(.A1(new_n16672_), .A2(new_n16582_), .Z(new_n16673_));
  OAI21_X1   g16481(.A1(new_n16542_), .A2(new_n16544_), .B(new_n16547_), .ZN(new_n16674_));
  NOR2_X1    g16482(.A1(new_n16649_), .A2(new_n16674_), .ZN(new_n16675_));
  XOR2_X1    g16483(.A1(new_n16675_), .A2(new_n16128_), .Z(new_n16676_));
  INV_X1     g16484(.I(new_n16676_), .ZN(new_n16677_));
  NAND3_X1   g16485(.A1(\asqrt[7] ), .A2(new_n16561_), .A3(new_n16543_), .ZN(new_n16678_));
  XOR2_X1    g16486(.A1(new_n16678_), .A2(new_n16132_), .Z(new_n16679_));
  INV_X1     g16487(.I(new_n16679_), .ZN(new_n16680_));
  OAI21_X1   g16488(.A1(new_n16556_), .A2(new_n16557_), .B(new_n16560_), .ZN(new_n16681_));
  NOR2_X1    g16489(.A1(new_n16649_), .A2(new_n16681_), .ZN(new_n16682_));
  XOR2_X1    g16490(.A1(new_n16682_), .A2(new_n16134_), .Z(new_n16683_));
  NAND3_X1   g16491(.A1(\asqrt[7] ), .A2(new_n16520_), .A3(new_n16539_), .ZN(new_n16684_));
  XOR2_X1    g16492(.A1(new_n16684_), .A2(new_n16554_), .Z(new_n16685_));
  OAI21_X1   g16493(.A1(new_n16514_), .A2(new_n16516_), .B(new_n16519_), .ZN(new_n16686_));
  NOR2_X1    g16494(.A1(new_n16649_), .A2(new_n16686_), .ZN(new_n16687_));
  XOR2_X1    g16495(.A1(new_n16687_), .A2(new_n16140_), .Z(new_n16688_));
  INV_X1     g16496(.I(new_n16688_), .ZN(new_n16689_));
  NAND3_X1   g16497(.A1(\asqrt[7] ), .A2(new_n16533_), .A3(new_n16515_), .ZN(new_n16690_));
  XOR2_X1    g16498(.A1(new_n16690_), .A2(new_n16144_), .Z(new_n16691_));
  INV_X1     g16499(.I(new_n16691_), .ZN(new_n16692_));
  OAI21_X1   g16500(.A1(new_n16528_), .A2(new_n16529_), .B(new_n16532_), .ZN(new_n16693_));
  NOR2_X1    g16501(.A1(new_n16649_), .A2(new_n16693_), .ZN(new_n16694_));
  XOR2_X1    g16502(.A1(new_n16694_), .A2(new_n16146_), .Z(new_n16695_));
  NAND3_X1   g16503(.A1(\asqrt[7] ), .A2(new_n16492_), .A3(new_n16511_), .ZN(new_n16696_));
  XOR2_X1    g16504(.A1(new_n16696_), .A2(new_n16526_), .Z(new_n16697_));
  OAI21_X1   g16505(.A1(new_n16486_), .A2(new_n16488_), .B(new_n16491_), .ZN(new_n16698_));
  NOR2_X1    g16506(.A1(new_n16649_), .A2(new_n16698_), .ZN(new_n16699_));
  XOR2_X1    g16507(.A1(new_n16699_), .A2(new_n16152_), .Z(new_n16700_));
  INV_X1     g16508(.I(new_n16700_), .ZN(new_n16701_));
  NAND3_X1   g16509(.A1(\asqrt[7] ), .A2(new_n16505_), .A3(new_n16487_), .ZN(new_n16702_));
  XOR2_X1    g16510(.A1(new_n16702_), .A2(new_n16156_), .Z(new_n16703_));
  INV_X1     g16511(.I(new_n16703_), .ZN(new_n16704_));
  OAI21_X1   g16512(.A1(new_n16500_), .A2(new_n16501_), .B(new_n16504_), .ZN(new_n16705_));
  NOR2_X1    g16513(.A1(new_n16649_), .A2(new_n16705_), .ZN(new_n16706_));
  XOR2_X1    g16514(.A1(new_n16706_), .A2(new_n16158_), .Z(new_n16707_));
  NAND3_X1   g16515(.A1(\asqrt[7] ), .A2(new_n16464_), .A3(new_n16483_), .ZN(new_n16708_));
  XOR2_X1    g16516(.A1(new_n16708_), .A2(new_n16498_), .Z(new_n16709_));
  OAI21_X1   g16517(.A1(new_n16458_), .A2(new_n16460_), .B(new_n16463_), .ZN(new_n16710_));
  NOR2_X1    g16518(.A1(new_n16649_), .A2(new_n16710_), .ZN(new_n16711_));
  XOR2_X1    g16519(.A1(new_n16711_), .A2(new_n16164_), .Z(new_n16712_));
  INV_X1     g16520(.I(new_n16712_), .ZN(new_n16713_));
  NAND3_X1   g16521(.A1(\asqrt[7] ), .A2(new_n16477_), .A3(new_n16459_), .ZN(new_n16714_));
  XOR2_X1    g16522(.A1(new_n16714_), .A2(new_n16168_), .Z(new_n16715_));
  INV_X1     g16523(.I(new_n16715_), .ZN(new_n16716_));
  OAI21_X1   g16524(.A1(new_n16472_), .A2(new_n16473_), .B(new_n16476_), .ZN(new_n16717_));
  NOR2_X1    g16525(.A1(new_n16649_), .A2(new_n16717_), .ZN(new_n16718_));
  XOR2_X1    g16526(.A1(new_n16718_), .A2(new_n16170_), .Z(new_n16719_));
  NAND3_X1   g16527(.A1(\asqrt[7] ), .A2(new_n16436_), .A3(new_n16455_), .ZN(new_n16720_));
  XOR2_X1    g16528(.A1(new_n16720_), .A2(new_n16470_), .Z(new_n16721_));
  OAI21_X1   g16529(.A1(new_n16430_), .A2(new_n16432_), .B(new_n16435_), .ZN(new_n16722_));
  NOR2_X1    g16530(.A1(new_n16649_), .A2(new_n16722_), .ZN(new_n16723_));
  XOR2_X1    g16531(.A1(new_n16723_), .A2(new_n16176_), .Z(new_n16724_));
  INV_X1     g16532(.I(new_n16724_), .ZN(new_n16725_));
  NAND3_X1   g16533(.A1(\asqrt[7] ), .A2(new_n16449_), .A3(new_n16431_), .ZN(new_n16726_));
  XOR2_X1    g16534(.A1(new_n16726_), .A2(new_n16180_), .Z(new_n16727_));
  INV_X1     g16535(.I(new_n16727_), .ZN(new_n16728_));
  OAI21_X1   g16536(.A1(new_n16444_), .A2(new_n16445_), .B(new_n16448_), .ZN(new_n16729_));
  NOR2_X1    g16537(.A1(new_n16649_), .A2(new_n16729_), .ZN(new_n16730_));
  XOR2_X1    g16538(.A1(new_n16730_), .A2(new_n16182_), .Z(new_n16731_));
  NAND3_X1   g16539(.A1(\asqrt[7] ), .A2(new_n16408_), .A3(new_n16427_), .ZN(new_n16732_));
  XOR2_X1    g16540(.A1(new_n16732_), .A2(new_n16442_), .Z(new_n16733_));
  OAI21_X1   g16541(.A1(new_n16402_), .A2(new_n16404_), .B(new_n16407_), .ZN(new_n16734_));
  NOR2_X1    g16542(.A1(new_n16649_), .A2(new_n16734_), .ZN(new_n16735_));
  XOR2_X1    g16543(.A1(new_n16735_), .A2(new_n16188_), .Z(new_n16736_));
  INV_X1     g16544(.I(new_n16736_), .ZN(new_n16737_));
  NAND3_X1   g16545(.A1(\asqrt[7] ), .A2(new_n16421_), .A3(new_n16403_), .ZN(new_n16738_));
  XOR2_X1    g16546(.A1(new_n16738_), .A2(new_n16192_), .Z(new_n16739_));
  INV_X1     g16547(.I(new_n16739_), .ZN(new_n16740_));
  OAI21_X1   g16548(.A1(new_n16416_), .A2(new_n16417_), .B(new_n16420_), .ZN(new_n16741_));
  NOR2_X1    g16549(.A1(new_n16649_), .A2(new_n16741_), .ZN(new_n16742_));
  XOR2_X1    g16550(.A1(new_n16742_), .A2(new_n16194_), .Z(new_n16743_));
  NAND3_X1   g16551(.A1(\asqrt[7] ), .A2(new_n16380_), .A3(new_n16399_), .ZN(new_n16744_));
  XOR2_X1    g16552(.A1(new_n16744_), .A2(new_n16414_), .Z(new_n16745_));
  OAI21_X1   g16553(.A1(new_n16374_), .A2(new_n16376_), .B(new_n16379_), .ZN(new_n16746_));
  NOR2_X1    g16554(.A1(new_n16649_), .A2(new_n16746_), .ZN(new_n16747_));
  XOR2_X1    g16555(.A1(new_n16747_), .A2(new_n16200_), .Z(new_n16748_));
  INV_X1     g16556(.I(new_n16748_), .ZN(new_n16749_));
  NAND3_X1   g16557(.A1(\asqrt[7] ), .A2(new_n16393_), .A3(new_n16375_), .ZN(new_n16750_));
  XOR2_X1    g16558(.A1(new_n16750_), .A2(new_n16204_), .Z(new_n16751_));
  INV_X1     g16559(.I(new_n16751_), .ZN(new_n16752_));
  OAI21_X1   g16560(.A1(new_n16388_), .A2(new_n16389_), .B(new_n16392_), .ZN(new_n16753_));
  NOR2_X1    g16561(.A1(new_n16649_), .A2(new_n16753_), .ZN(new_n16754_));
  XOR2_X1    g16562(.A1(new_n16754_), .A2(new_n16206_), .Z(new_n16755_));
  NAND3_X1   g16563(.A1(\asqrt[7] ), .A2(new_n16352_), .A3(new_n16371_), .ZN(new_n16756_));
  XOR2_X1    g16564(.A1(new_n16756_), .A2(new_n16386_), .Z(new_n16757_));
  OAI21_X1   g16565(.A1(new_n16346_), .A2(new_n16348_), .B(new_n16351_), .ZN(new_n16758_));
  NOR2_X1    g16566(.A1(new_n16649_), .A2(new_n16758_), .ZN(new_n16759_));
  XOR2_X1    g16567(.A1(new_n16759_), .A2(new_n16212_), .Z(new_n16760_));
  INV_X1     g16568(.I(new_n16760_), .ZN(new_n16761_));
  NAND3_X1   g16569(.A1(\asqrt[7] ), .A2(new_n16365_), .A3(new_n16347_), .ZN(new_n16762_));
  XOR2_X1    g16570(.A1(new_n16762_), .A2(new_n16216_), .Z(new_n16763_));
  INV_X1     g16571(.I(new_n16763_), .ZN(new_n16764_));
  OAI21_X1   g16572(.A1(new_n16360_), .A2(new_n16361_), .B(new_n16364_), .ZN(new_n16765_));
  NOR2_X1    g16573(.A1(new_n16649_), .A2(new_n16765_), .ZN(new_n16766_));
  XOR2_X1    g16574(.A1(new_n16766_), .A2(new_n16218_), .Z(new_n16767_));
  NAND3_X1   g16575(.A1(\asqrt[7] ), .A2(new_n16324_), .A3(new_n16343_), .ZN(new_n16768_));
  XOR2_X1    g16576(.A1(new_n16768_), .A2(new_n16358_), .Z(new_n16769_));
  OAI21_X1   g16577(.A1(new_n16318_), .A2(new_n16320_), .B(new_n16323_), .ZN(new_n16770_));
  NOR2_X1    g16578(.A1(new_n16649_), .A2(new_n16770_), .ZN(new_n16771_));
  XOR2_X1    g16579(.A1(new_n16771_), .A2(new_n16224_), .Z(new_n16772_));
  INV_X1     g16580(.I(new_n16772_), .ZN(new_n16773_));
  NAND3_X1   g16581(.A1(\asqrt[7] ), .A2(new_n16337_), .A3(new_n16319_), .ZN(new_n16774_));
  XOR2_X1    g16582(.A1(new_n16774_), .A2(new_n16228_), .Z(new_n16775_));
  INV_X1     g16583(.I(new_n16775_), .ZN(new_n16776_));
  AOI21_X1   g16584(.A1(new_n16284_), .A2(new_n16286_), .B(new_n16316_), .ZN(new_n16777_));
  NAND2_X1   g16585(.A1(\asqrt[7] ), .A2(new_n16777_), .ZN(new_n16778_));
  XOR2_X1    g16586(.A1(new_n16778_), .A2(new_n16231_), .Z(new_n16779_));
  NAND3_X1   g16587(.A1(\asqrt[7] ), .A2(new_n16283_), .A3(new_n16315_), .ZN(new_n16780_));
  XOR2_X1    g16588(.A1(new_n16780_), .A2(new_n16330_), .Z(new_n16781_));
  OAI21_X1   g16589(.A1(new_n16277_), .A2(new_n16279_), .B(new_n16282_), .ZN(new_n16782_));
  NOR2_X1    g16590(.A1(new_n16649_), .A2(new_n16782_), .ZN(new_n16783_));
  XOR2_X1    g16591(.A1(new_n16783_), .A2(new_n16236_), .Z(new_n16784_));
  INV_X1     g16592(.I(new_n16784_), .ZN(new_n16785_));
  NAND3_X1   g16593(.A1(\asqrt[7] ), .A2(new_n16309_), .A3(new_n16278_), .ZN(new_n16786_));
  XOR2_X1    g16594(.A1(new_n16786_), .A2(new_n16240_), .Z(new_n16787_));
  INV_X1     g16595(.I(new_n16787_), .ZN(new_n16788_));
  AOI21_X1   g16596(.A1(new_n16271_), .A2(new_n16272_), .B(new_n16275_), .ZN(new_n16789_));
  NAND2_X1   g16597(.A1(\asqrt[7] ), .A2(new_n16789_), .ZN(new_n16790_));
  XOR2_X1    g16598(.A1(new_n16790_), .A2(new_n16243_), .Z(new_n16791_));
  NOR2_X1    g16599(.A1(new_n16270_), .A2(\asqrt[12] ), .ZN(new_n16792_));
  NOR3_X1    g16600(.A1(new_n16649_), .A2(new_n16792_), .A3(new_n16307_), .ZN(new_n16793_));
  XOR2_X1    g16601(.A1(new_n16793_), .A2(new_n16246_), .Z(new_n16794_));
  NAND3_X1   g16602(.A1(\asqrt[7] ), .A2(new_n16301_), .A3(new_n16269_), .ZN(new_n16795_));
  XOR2_X1    g16603(.A1(new_n16795_), .A2(new_n16268_), .Z(new_n16796_));
  INV_X1     g16604(.I(new_n16796_), .ZN(new_n16797_));
  NAND2_X1   g16605(.A1(new_n16262_), .A2(new_n14985_), .ZN(new_n16798_));
  NAND3_X1   g16606(.A1(\asqrt[7] ), .A2(new_n16798_), .A3(new_n16300_), .ZN(new_n16799_));
  XOR2_X1    g16607(.A1(new_n16799_), .A2(new_n16253_), .Z(new_n16800_));
  INV_X1     g16608(.I(new_n16800_), .ZN(new_n16801_));
  NAND3_X1   g16609(.A1(\asqrt[7] ), .A2(new_n16254_), .A3(new_n16255_), .ZN(new_n16802_));
  NAND4_X1   g16610(.A1(new_n16656_), .A2(\asqrt[8] ), .A3(new_n16657_), .A4(new_n16654_), .ZN(new_n16803_));
  AOI21_X1   g16611(.A1(new_n16802_), .A2(new_n16803_), .B(\a[16] ), .ZN(new_n16804_));
  NOR3_X1    g16612(.A1(new_n16649_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n16805_));
  INV_X1     g16613(.I(new_n16803_), .ZN(new_n16806_));
  NOR3_X1    g16614(.A1(new_n16805_), .A2(new_n15671_), .A3(new_n16806_), .ZN(new_n16807_));
  NOR2_X1    g16615(.A1(new_n16807_), .A2(new_n16804_), .ZN(new_n16808_));
  INV_X1     g16616(.I(\a[12] ), .ZN(new_n16809_));
  INV_X1     g16617(.I(\a[13] ), .ZN(new_n16810_));
  NAND3_X1   g16618(.A1(new_n16809_), .A2(new_n16810_), .A3(new_n16254_), .ZN(new_n16811_));
  OAI21_X1   g16619(.A1(new_n16649_), .A2(new_n16254_), .B(new_n16811_), .ZN(new_n16812_));
  NAND2_X1   g16620(.A1(new_n16812_), .A2(\asqrt[8] ), .ZN(new_n16813_));
  OAI21_X1   g16621(.A1(new_n16649_), .A2(\a[14] ), .B(\a[15] ), .ZN(new_n16814_));
  NAND2_X1   g16622(.A1(new_n16814_), .A2(new_n16802_), .ZN(new_n16815_));
  NOR2_X1    g16623(.A1(new_n16812_), .A2(\asqrt[8] ), .ZN(new_n16816_));
  OAI21_X1   g16624(.A1(new_n16815_), .A2(new_n16816_), .B(new_n16813_), .ZN(new_n16817_));
  OAI21_X1   g16625(.A1(new_n16817_), .A2(\asqrt[9] ), .B(new_n16808_), .ZN(new_n16818_));
  NAND2_X1   g16626(.A1(new_n16817_), .A2(\asqrt[9] ), .ZN(new_n16819_));
  NAND3_X1   g16627(.A1(new_n16818_), .A2(new_n14985_), .A3(new_n16819_), .ZN(new_n16820_));
  NAND3_X1   g16628(.A1(\asqrt[7] ), .A2(new_n16294_), .A3(new_n16261_), .ZN(new_n16821_));
  XOR2_X1    g16629(.A1(new_n16821_), .A2(new_n16296_), .Z(new_n16822_));
  NAND2_X1   g16630(.A1(new_n16820_), .A2(new_n16822_), .ZN(new_n16823_));
  NAND2_X1   g16631(.A1(new_n16818_), .A2(new_n16819_), .ZN(new_n16824_));
  AOI21_X1   g16632(.A1(new_n16824_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n16825_));
  AOI21_X1   g16633(.A1(new_n16825_), .A2(new_n16823_), .B(new_n16801_), .ZN(new_n16826_));
  OAI21_X1   g16634(.A1(new_n16805_), .A2(new_n16806_), .B(new_n15671_), .ZN(new_n16827_));
  NAND3_X1   g16635(.A1(new_n16802_), .A2(\a[16] ), .A3(new_n16803_), .ZN(new_n16828_));
  NAND2_X1   g16636(.A1(new_n16827_), .A2(new_n16828_), .ZN(new_n16829_));
  NAND2_X1   g16637(.A1(\asqrt[7] ), .A2(\a[14] ), .ZN(new_n16830_));
  AOI21_X1   g16638(.A1(new_n16830_), .A2(new_n16811_), .B(new_n16093_), .ZN(new_n16831_));
  AOI21_X1   g16639(.A1(\asqrt[7] ), .A2(new_n16254_), .B(new_n16255_), .ZN(new_n16832_));
  NOR2_X1    g16640(.A1(new_n16805_), .A2(new_n16832_), .ZN(new_n16833_));
  NAND3_X1   g16641(.A1(new_n16830_), .A2(new_n16093_), .A3(new_n16811_), .ZN(new_n16834_));
  AOI21_X1   g16642(.A1(new_n16833_), .A2(new_n16834_), .B(new_n16831_), .ZN(new_n16835_));
  AOI21_X1   g16643(.A1(new_n16835_), .A2(new_n15518_), .B(new_n16829_), .ZN(new_n16836_));
  NOR2_X1    g16644(.A1(new_n16835_), .A2(new_n15518_), .ZN(new_n16837_));
  OAI21_X1   g16645(.A1(new_n16836_), .A2(new_n16837_), .B(\asqrt[10] ), .ZN(new_n16838_));
  AOI21_X1   g16646(.A1(new_n16823_), .A2(new_n16838_), .B(new_n14430_), .ZN(new_n16839_));
  NOR2_X1    g16647(.A1(new_n16826_), .A2(new_n16839_), .ZN(new_n16840_));
  AOI21_X1   g16648(.A1(new_n16840_), .A2(new_n13917_), .B(new_n16797_), .ZN(new_n16841_));
  OAI21_X1   g16649(.A1(new_n16826_), .A2(new_n16839_), .B(\asqrt[12] ), .ZN(new_n16842_));
  NAND2_X1   g16650(.A1(new_n16842_), .A2(new_n13382_), .ZN(new_n16843_));
  OAI21_X1   g16651(.A1(new_n16841_), .A2(new_n16843_), .B(new_n16794_), .ZN(new_n16844_));
  INV_X1     g16652(.I(new_n16842_), .ZN(new_n16845_));
  OAI21_X1   g16653(.A1(new_n16841_), .A2(new_n16845_), .B(\asqrt[13] ), .ZN(new_n16846_));
  NAND3_X1   g16654(.A1(new_n16844_), .A2(new_n16846_), .A3(new_n12889_), .ZN(new_n16847_));
  NAND2_X1   g16655(.A1(new_n16847_), .A2(new_n16791_), .ZN(new_n16848_));
  NAND2_X1   g16656(.A1(new_n16844_), .A2(new_n16846_), .ZN(new_n16849_));
  AOI21_X1   g16657(.A1(new_n16849_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n16850_));
  AOI21_X1   g16658(.A1(new_n16850_), .A2(new_n16848_), .B(new_n16788_), .ZN(new_n16851_));
  INV_X1     g16659(.I(new_n16794_), .ZN(new_n16852_));
  NOR2_X1    g16660(.A1(new_n16836_), .A2(new_n16837_), .ZN(new_n16853_));
  INV_X1     g16661(.I(new_n16822_), .ZN(new_n16854_));
  AOI21_X1   g16662(.A1(new_n16853_), .A2(new_n14985_), .B(new_n16854_), .ZN(new_n16855_));
  NAND2_X1   g16663(.A1(new_n16838_), .A2(new_n14430_), .ZN(new_n16856_));
  OAI21_X1   g16664(.A1(new_n16855_), .A2(new_n16856_), .B(new_n16800_), .ZN(new_n16857_));
  INV_X1     g16665(.I(new_n16838_), .ZN(new_n16858_));
  OAI21_X1   g16666(.A1(new_n16855_), .A2(new_n16858_), .B(\asqrt[11] ), .ZN(new_n16859_));
  NAND3_X1   g16667(.A1(new_n16857_), .A2(new_n16859_), .A3(new_n13917_), .ZN(new_n16860_));
  NAND2_X1   g16668(.A1(new_n16860_), .A2(new_n16796_), .ZN(new_n16861_));
  NAND2_X1   g16669(.A1(new_n16857_), .A2(new_n16859_), .ZN(new_n16862_));
  AOI21_X1   g16670(.A1(new_n16862_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n16863_));
  AOI21_X1   g16671(.A1(new_n16863_), .A2(new_n16861_), .B(new_n16852_), .ZN(new_n16864_));
  AOI21_X1   g16672(.A1(new_n16861_), .A2(new_n16842_), .B(new_n13382_), .ZN(new_n16865_));
  OAI21_X1   g16673(.A1(new_n16864_), .A2(new_n16865_), .B(\asqrt[14] ), .ZN(new_n16866_));
  AOI21_X1   g16674(.A1(new_n16848_), .A2(new_n16866_), .B(new_n12374_), .ZN(new_n16867_));
  NOR2_X1    g16675(.A1(new_n16851_), .A2(new_n16867_), .ZN(new_n16868_));
  AOI21_X1   g16676(.A1(new_n16868_), .A2(new_n11901_), .B(new_n16785_), .ZN(new_n16869_));
  OAI21_X1   g16677(.A1(new_n16851_), .A2(new_n16867_), .B(\asqrt[16] ), .ZN(new_n16870_));
  NAND2_X1   g16678(.A1(new_n16870_), .A2(new_n11406_), .ZN(new_n16871_));
  OAI21_X1   g16679(.A1(new_n16869_), .A2(new_n16871_), .B(new_n16781_), .ZN(new_n16872_));
  INV_X1     g16680(.I(new_n16870_), .ZN(new_n16873_));
  OAI21_X1   g16681(.A1(new_n16869_), .A2(new_n16873_), .B(\asqrt[17] ), .ZN(new_n16874_));
  NAND3_X1   g16682(.A1(new_n16872_), .A2(new_n16874_), .A3(new_n10953_), .ZN(new_n16875_));
  NAND2_X1   g16683(.A1(new_n16875_), .A2(new_n16779_), .ZN(new_n16876_));
  NAND2_X1   g16684(.A1(new_n16872_), .A2(new_n16874_), .ZN(new_n16877_));
  AOI21_X1   g16685(.A1(new_n16877_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n16878_));
  AOI21_X1   g16686(.A1(new_n16878_), .A2(new_n16876_), .B(new_n16776_), .ZN(new_n16879_));
  INV_X1     g16687(.I(new_n16781_), .ZN(new_n16880_));
  INV_X1     g16688(.I(new_n16791_), .ZN(new_n16881_));
  NOR2_X1    g16689(.A1(new_n16864_), .A2(new_n16865_), .ZN(new_n16882_));
  AOI21_X1   g16690(.A1(new_n16882_), .A2(new_n12889_), .B(new_n16881_), .ZN(new_n16883_));
  NAND2_X1   g16691(.A1(new_n16866_), .A2(new_n12374_), .ZN(new_n16884_));
  OAI21_X1   g16692(.A1(new_n16883_), .A2(new_n16884_), .B(new_n16787_), .ZN(new_n16885_));
  INV_X1     g16693(.I(new_n16866_), .ZN(new_n16886_));
  OAI21_X1   g16694(.A1(new_n16883_), .A2(new_n16886_), .B(\asqrt[15] ), .ZN(new_n16887_));
  NAND3_X1   g16695(.A1(new_n16885_), .A2(new_n16887_), .A3(new_n11901_), .ZN(new_n16888_));
  NAND2_X1   g16696(.A1(new_n16888_), .A2(new_n16784_), .ZN(new_n16889_));
  NAND2_X1   g16697(.A1(new_n16885_), .A2(new_n16887_), .ZN(new_n16890_));
  AOI21_X1   g16698(.A1(new_n16890_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n16891_));
  AOI21_X1   g16699(.A1(new_n16891_), .A2(new_n16889_), .B(new_n16880_), .ZN(new_n16892_));
  AOI21_X1   g16700(.A1(new_n16889_), .A2(new_n16870_), .B(new_n11406_), .ZN(new_n16893_));
  OAI21_X1   g16701(.A1(new_n16892_), .A2(new_n16893_), .B(\asqrt[18] ), .ZN(new_n16894_));
  AOI21_X1   g16702(.A1(new_n16876_), .A2(new_n16894_), .B(new_n10478_), .ZN(new_n16895_));
  NOR2_X1    g16703(.A1(new_n16879_), .A2(new_n16895_), .ZN(new_n16896_));
  AOI21_X1   g16704(.A1(new_n16896_), .A2(new_n10045_), .B(new_n16773_), .ZN(new_n16897_));
  OAI21_X1   g16705(.A1(new_n16879_), .A2(new_n16895_), .B(\asqrt[20] ), .ZN(new_n16898_));
  NAND2_X1   g16706(.A1(new_n16898_), .A2(new_n9590_), .ZN(new_n16899_));
  OAI21_X1   g16707(.A1(new_n16897_), .A2(new_n16899_), .B(new_n16769_), .ZN(new_n16900_));
  INV_X1     g16708(.I(new_n16898_), .ZN(new_n16901_));
  OAI21_X1   g16709(.A1(new_n16897_), .A2(new_n16901_), .B(\asqrt[21] ), .ZN(new_n16902_));
  NAND3_X1   g16710(.A1(new_n16900_), .A2(new_n16902_), .A3(new_n9177_), .ZN(new_n16903_));
  NAND2_X1   g16711(.A1(new_n16903_), .A2(new_n16767_), .ZN(new_n16904_));
  NAND2_X1   g16712(.A1(new_n16900_), .A2(new_n16902_), .ZN(new_n16905_));
  AOI21_X1   g16713(.A1(new_n16905_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n16906_));
  AOI21_X1   g16714(.A1(new_n16906_), .A2(new_n16904_), .B(new_n16764_), .ZN(new_n16907_));
  INV_X1     g16715(.I(new_n16769_), .ZN(new_n16908_));
  INV_X1     g16716(.I(new_n16779_), .ZN(new_n16909_));
  NOR2_X1    g16717(.A1(new_n16892_), .A2(new_n16893_), .ZN(new_n16910_));
  AOI21_X1   g16718(.A1(new_n16910_), .A2(new_n10953_), .B(new_n16909_), .ZN(new_n16911_));
  NAND2_X1   g16719(.A1(new_n16894_), .A2(new_n10478_), .ZN(new_n16912_));
  OAI21_X1   g16720(.A1(new_n16911_), .A2(new_n16912_), .B(new_n16775_), .ZN(new_n16913_));
  INV_X1     g16721(.I(new_n16894_), .ZN(new_n16914_));
  OAI21_X1   g16722(.A1(new_n16911_), .A2(new_n16914_), .B(\asqrt[19] ), .ZN(new_n16915_));
  NAND3_X1   g16723(.A1(new_n16913_), .A2(new_n16915_), .A3(new_n10045_), .ZN(new_n16916_));
  NAND2_X1   g16724(.A1(new_n16916_), .A2(new_n16772_), .ZN(new_n16917_));
  NAND2_X1   g16725(.A1(new_n16913_), .A2(new_n16915_), .ZN(new_n16918_));
  AOI21_X1   g16726(.A1(new_n16918_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n16919_));
  AOI21_X1   g16727(.A1(new_n16919_), .A2(new_n16917_), .B(new_n16908_), .ZN(new_n16920_));
  AOI21_X1   g16728(.A1(new_n16917_), .A2(new_n16898_), .B(new_n9590_), .ZN(new_n16921_));
  OAI21_X1   g16729(.A1(new_n16920_), .A2(new_n16921_), .B(\asqrt[22] ), .ZN(new_n16922_));
  AOI21_X1   g16730(.A1(new_n16904_), .A2(new_n16922_), .B(new_n8742_), .ZN(new_n16923_));
  NOR2_X1    g16731(.A1(new_n16907_), .A2(new_n16923_), .ZN(new_n16924_));
  AOI21_X1   g16732(.A1(new_n16924_), .A2(new_n8349_), .B(new_n16761_), .ZN(new_n16925_));
  OAI21_X1   g16733(.A1(new_n16907_), .A2(new_n16923_), .B(\asqrt[24] ), .ZN(new_n16926_));
  NAND2_X1   g16734(.A1(new_n16926_), .A2(new_n7934_), .ZN(new_n16927_));
  OAI21_X1   g16735(.A1(new_n16925_), .A2(new_n16927_), .B(new_n16757_), .ZN(new_n16928_));
  INV_X1     g16736(.I(new_n16926_), .ZN(new_n16929_));
  OAI21_X1   g16737(.A1(new_n16925_), .A2(new_n16929_), .B(\asqrt[25] ), .ZN(new_n16930_));
  NAND3_X1   g16738(.A1(new_n16928_), .A2(new_n16930_), .A3(new_n7561_), .ZN(new_n16931_));
  NAND2_X1   g16739(.A1(new_n16931_), .A2(new_n16755_), .ZN(new_n16932_));
  NAND2_X1   g16740(.A1(new_n16928_), .A2(new_n16930_), .ZN(new_n16933_));
  AOI21_X1   g16741(.A1(new_n16933_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n16934_));
  AOI21_X1   g16742(.A1(new_n16934_), .A2(new_n16932_), .B(new_n16752_), .ZN(new_n16935_));
  INV_X1     g16743(.I(new_n16757_), .ZN(new_n16936_));
  INV_X1     g16744(.I(new_n16767_), .ZN(new_n16937_));
  NOR2_X1    g16745(.A1(new_n16920_), .A2(new_n16921_), .ZN(new_n16938_));
  AOI21_X1   g16746(.A1(new_n16938_), .A2(new_n9177_), .B(new_n16937_), .ZN(new_n16939_));
  NAND2_X1   g16747(.A1(new_n16922_), .A2(new_n8742_), .ZN(new_n16940_));
  OAI21_X1   g16748(.A1(new_n16939_), .A2(new_n16940_), .B(new_n16763_), .ZN(new_n16941_));
  INV_X1     g16749(.I(new_n16922_), .ZN(new_n16942_));
  OAI21_X1   g16750(.A1(new_n16939_), .A2(new_n16942_), .B(\asqrt[23] ), .ZN(new_n16943_));
  NAND3_X1   g16751(.A1(new_n16941_), .A2(new_n16943_), .A3(new_n8349_), .ZN(new_n16944_));
  NAND2_X1   g16752(.A1(new_n16944_), .A2(new_n16760_), .ZN(new_n16945_));
  NAND2_X1   g16753(.A1(new_n16941_), .A2(new_n16943_), .ZN(new_n16946_));
  AOI21_X1   g16754(.A1(new_n16946_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n16947_));
  AOI21_X1   g16755(.A1(new_n16947_), .A2(new_n16945_), .B(new_n16936_), .ZN(new_n16948_));
  AOI21_X1   g16756(.A1(new_n16945_), .A2(new_n16926_), .B(new_n7934_), .ZN(new_n16949_));
  OAI21_X1   g16757(.A1(new_n16948_), .A2(new_n16949_), .B(\asqrt[26] ), .ZN(new_n16950_));
  AOI21_X1   g16758(.A1(new_n16932_), .A2(new_n16950_), .B(new_n7166_), .ZN(new_n16951_));
  NOR2_X1    g16759(.A1(new_n16935_), .A2(new_n16951_), .ZN(new_n16952_));
  AOI21_X1   g16760(.A1(new_n16952_), .A2(new_n6813_), .B(new_n16749_), .ZN(new_n16953_));
  OAI21_X1   g16761(.A1(new_n16935_), .A2(new_n16951_), .B(\asqrt[28] ), .ZN(new_n16954_));
  NAND2_X1   g16762(.A1(new_n16954_), .A2(new_n6454_), .ZN(new_n16955_));
  OAI21_X1   g16763(.A1(new_n16953_), .A2(new_n16955_), .B(new_n16745_), .ZN(new_n16956_));
  INV_X1     g16764(.I(new_n16954_), .ZN(new_n16957_));
  OAI21_X1   g16765(.A1(new_n16953_), .A2(new_n16957_), .B(\asqrt[29] ), .ZN(new_n16958_));
  NAND3_X1   g16766(.A1(new_n16956_), .A2(new_n16958_), .A3(new_n6106_), .ZN(new_n16959_));
  NAND2_X1   g16767(.A1(new_n16959_), .A2(new_n16743_), .ZN(new_n16960_));
  NAND2_X1   g16768(.A1(new_n16956_), .A2(new_n16958_), .ZN(new_n16961_));
  AOI21_X1   g16769(.A1(new_n16961_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n16962_));
  AOI21_X1   g16770(.A1(new_n16962_), .A2(new_n16960_), .B(new_n16740_), .ZN(new_n16963_));
  INV_X1     g16771(.I(new_n16745_), .ZN(new_n16964_));
  INV_X1     g16772(.I(new_n16755_), .ZN(new_n16965_));
  NOR2_X1    g16773(.A1(new_n16948_), .A2(new_n16949_), .ZN(new_n16966_));
  AOI21_X1   g16774(.A1(new_n16966_), .A2(new_n7561_), .B(new_n16965_), .ZN(new_n16967_));
  NAND2_X1   g16775(.A1(new_n16950_), .A2(new_n7166_), .ZN(new_n16968_));
  OAI21_X1   g16776(.A1(new_n16967_), .A2(new_n16968_), .B(new_n16751_), .ZN(new_n16969_));
  INV_X1     g16777(.I(new_n16950_), .ZN(new_n16970_));
  OAI21_X1   g16778(.A1(new_n16967_), .A2(new_n16970_), .B(\asqrt[27] ), .ZN(new_n16971_));
  NAND3_X1   g16779(.A1(new_n16969_), .A2(new_n16971_), .A3(new_n6813_), .ZN(new_n16972_));
  NAND2_X1   g16780(.A1(new_n16972_), .A2(new_n16748_), .ZN(new_n16973_));
  NAND2_X1   g16781(.A1(new_n16969_), .A2(new_n16971_), .ZN(new_n16974_));
  AOI21_X1   g16782(.A1(new_n16974_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n16975_));
  AOI21_X1   g16783(.A1(new_n16975_), .A2(new_n16973_), .B(new_n16964_), .ZN(new_n16976_));
  AOI21_X1   g16784(.A1(new_n16973_), .A2(new_n16954_), .B(new_n6454_), .ZN(new_n16977_));
  OAI21_X1   g16785(.A1(new_n16976_), .A2(new_n16977_), .B(\asqrt[30] ), .ZN(new_n16978_));
  AOI21_X1   g16786(.A1(new_n16960_), .A2(new_n16978_), .B(new_n5750_), .ZN(new_n16979_));
  NOR2_X1    g16787(.A1(new_n16963_), .A2(new_n16979_), .ZN(new_n16980_));
  AOI21_X1   g16788(.A1(new_n16980_), .A2(new_n5435_), .B(new_n16737_), .ZN(new_n16981_));
  OAI21_X1   g16789(.A1(new_n16963_), .A2(new_n16979_), .B(\asqrt[32] ), .ZN(new_n16982_));
  NAND2_X1   g16790(.A1(new_n16982_), .A2(new_n5110_), .ZN(new_n16983_));
  OAI21_X1   g16791(.A1(new_n16981_), .A2(new_n16983_), .B(new_n16733_), .ZN(new_n16984_));
  INV_X1     g16792(.I(new_n16982_), .ZN(new_n16985_));
  OAI21_X1   g16793(.A1(new_n16981_), .A2(new_n16985_), .B(\asqrt[33] ), .ZN(new_n16986_));
  NAND3_X1   g16794(.A1(new_n16984_), .A2(new_n16986_), .A3(new_n4810_), .ZN(new_n16987_));
  NAND2_X1   g16795(.A1(new_n16987_), .A2(new_n16731_), .ZN(new_n16988_));
  NAND2_X1   g16796(.A1(new_n16984_), .A2(new_n16986_), .ZN(new_n16989_));
  AOI21_X1   g16797(.A1(new_n16989_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n16990_));
  AOI21_X1   g16798(.A1(new_n16990_), .A2(new_n16988_), .B(new_n16728_), .ZN(new_n16991_));
  INV_X1     g16799(.I(new_n16733_), .ZN(new_n16992_));
  INV_X1     g16800(.I(new_n16743_), .ZN(new_n16993_));
  NOR2_X1    g16801(.A1(new_n16976_), .A2(new_n16977_), .ZN(new_n16994_));
  AOI21_X1   g16802(.A1(new_n16994_), .A2(new_n6106_), .B(new_n16993_), .ZN(new_n16995_));
  NAND2_X1   g16803(.A1(new_n16978_), .A2(new_n5750_), .ZN(new_n16996_));
  OAI21_X1   g16804(.A1(new_n16995_), .A2(new_n16996_), .B(new_n16739_), .ZN(new_n16997_));
  INV_X1     g16805(.I(new_n16978_), .ZN(new_n16998_));
  OAI21_X1   g16806(.A1(new_n16995_), .A2(new_n16998_), .B(\asqrt[31] ), .ZN(new_n16999_));
  NAND3_X1   g16807(.A1(new_n16997_), .A2(new_n16999_), .A3(new_n5435_), .ZN(new_n17000_));
  NAND2_X1   g16808(.A1(new_n17000_), .A2(new_n16736_), .ZN(new_n17001_));
  NAND2_X1   g16809(.A1(new_n16997_), .A2(new_n16999_), .ZN(new_n17002_));
  AOI21_X1   g16810(.A1(new_n17002_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n17003_));
  AOI21_X1   g16811(.A1(new_n17003_), .A2(new_n17001_), .B(new_n16992_), .ZN(new_n17004_));
  AOI21_X1   g16812(.A1(new_n17001_), .A2(new_n16982_), .B(new_n5110_), .ZN(new_n17005_));
  OAI21_X1   g16813(.A1(new_n17004_), .A2(new_n17005_), .B(\asqrt[34] ), .ZN(new_n17006_));
  AOI21_X1   g16814(.A1(new_n16988_), .A2(new_n17006_), .B(new_n4510_), .ZN(new_n17007_));
  NOR2_X1    g16815(.A1(new_n16991_), .A2(new_n17007_), .ZN(new_n17008_));
  AOI21_X1   g16816(.A1(new_n17008_), .A2(new_n4224_), .B(new_n16725_), .ZN(new_n17009_));
  OAI21_X1   g16817(.A1(new_n16991_), .A2(new_n17007_), .B(\asqrt[36] ), .ZN(new_n17010_));
  NAND2_X1   g16818(.A1(new_n17010_), .A2(new_n3928_), .ZN(new_n17011_));
  OAI21_X1   g16819(.A1(new_n17009_), .A2(new_n17011_), .B(new_n16721_), .ZN(new_n17012_));
  INV_X1     g16820(.I(new_n17010_), .ZN(new_n17013_));
  OAI21_X1   g16821(.A1(new_n17009_), .A2(new_n17013_), .B(\asqrt[37] ), .ZN(new_n17014_));
  NAND3_X1   g16822(.A1(new_n17012_), .A2(new_n17014_), .A3(new_n3675_), .ZN(new_n17015_));
  NAND2_X1   g16823(.A1(new_n17015_), .A2(new_n16719_), .ZN(new_n17016_));
  NAND2_X1   g16824(.A1(new_n17012_), .A2(new_n17014_), .ZN(new_n17017_));
  AOI21_X1   g16825(.A1(new_n17017_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n17018_));
  AOI21_X1   g16826(.A1(new_n17018_), .A2(new_n17016_), .B(new_n16716_), .ZN(new_n17019_));
  INV_X1     g16827(.I(new_n16721_), .ZN(new_n17020_));
  INV_X1     g16828(.I(new_n16731_), .ZN(new_n17021_));
  NOR2_X1    g16829(.A1(new_n17004_), .A2(new_n17005_), .ZN(new_n17022_));
  AOI21_X1   g16830(.A1(new_n17022_), .A2(new_n4810_), .B(new_n17021_), .ZN(new_n17023_));
  NAND2_X1   g16831(.A1(new_n17006_), .A2(new_n4510_), .ZN(new_n17024_));
  OAI21_X1   g16832(.A1(new_n17023_), .A2(new_n17024_), .B(new_n16727_), .ZN(new_n17025_));
  INV_X1     g16833(.I(new_n17006_), .ZN(new_n17026_));
  OAI21_X1   g16834(.A1(new_n17023_), .A2(new_n17026_), .B(\asqrt[35] ), .ZN(new_n17027_));
  NAND3_X1   g16835(.A1(new_n17025_), .A2(new_n17027_), .A3(new_n4224_), .ZN(new_n17028_));
  NAND2_X1   g16836(.A1(new_n17028_), .A2(new_n16724_), .ZN(new_n17029_));
  NAND2_X1   g16837(.A1(new_n17025_), .A2(new_n17027_), .ZN(new_n17030_));
  AOI21_X1   g16838(.A1(new_n17030_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n17031_));
  AOI21_X1   g16839(.A1(new_n17031_), .A2(new_n17029_), .B(new_n17020_), .ZN(new_n17032_));
  AOI21_X1   g16840(.A1(new_n17029_), .A2(new_n17010_), .B(new_n3928_), .ZN(new_n17033_));
  OAI21_X1   g16841(.A1(new_n17032_), .A2(new_n17033_), .B(\asqrt[38] ), .ZN(new_n17034_));
  AOI21_X1   g16842(.A1(new_n17016_), .A2(new_n17034_), .B(new_n3400_), .ZN(new_n17035_));
  NOR2_X1    g16843(.A1(new_n17019_), .A2(new_n17035_), .ZN(new_n17036_));
  AOI21_X1   g16844(.A1(new_n17036_), .A2(new_n3167_), .B(new_n16713_), .ZN(new_n17037_));
  OAI21_X1   g16845(.A1(new_n17019_), .A2(new_n17035_), .B(\asqrt[40] ), .ZN(new_n17038_));
  NAND2_X1   g16846(.A1(new_n17038_), .A2(new_n2912_), .ZN(new_n17039_));
  OAI21_X1   g16847(.A1(new_n17037_), .A2(new_n17039_), .B(new_n16709_), .ZN(new_n17040_));
  INV_X1     g16848(.I(new_n17038_), .ZN(new_n17041_));
  OAI21_X1   g16849(.A1(new_n17037_), .A2(new_n17041_), .B(\asqrt[41] ), .ZN(new_n17042_));
  NAND3_X1   g16850(.A1(new_n17040_), .A2(new_n17042_), .A3(new_n2699_), .ZN(new_n17043_));
  NAND2_X1   g16851(.A1(new_n17043_), .A2(new_n16707_), .ZN(new_n17044_));
  NAND2_X1   g16852(.A1(new_n17040_), .A2(new_n17042_), .ZN(new_n17045_));
  AOI21_X1   g16853(.A1(new_n17045_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n17046_));
  AOI21_X1   g16854(.A1(new_n17046_), .A2(new_n17044_), .B(new_n16704_), .ZN(new_n17047_));
  INV_X1     g16855(.I(new_n16709_), .ZN(new_n17048_));
  INV_X1     g16856(.I(new_n16719_), .ZN(new_n17049_));
  NOR2_X1    g16857(.A1(new_n17032_), .A2(new_n17033_), .ZN(new_n17050_));
  AOI21_X1   g16858(.A1(new_n17050_), .A2(new_n3675_), .B(new_n17049_), .ZN(new_n17051_));
  NAND2_X1   g16859(.A1(new_n17034_), .A2(new_n3400_), .ZN(new_n17052_));
  OAI21_X1   g16860(.A1(new_n17051_), .A2(new_n17052_), .B(new_n16715_), .ZN(new_n17053_));
  INV_X1     g16861(.I(new_n17034_), .ZN(new_n17054_));
  OAI21_X1   g16862(.A1(new_n17051_), .A2(new_n17054_), .B(\asqrt[39] ), .ZN(new_n17055_));
  NAND3_X1   g16863(.A1(new_n17053_), .A2(new_n17055_), .A3(new_n3167_), .ZN(new_n17056_));
  NAND2_X1   g16864(.A1(new_n17056_), .A2(new_n16712_), .ZN(new_n17057_));
  NAND2_X1   g16865(.A1(new_n17053_), .A2(new_n17055_), .ZN(new_n17058_));
  AOI21_X1   g16866(.A1(new_n17058_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n17059_));
  AOI21_X1   g16867(.A1(new_n17059_), .A2(new_n17057_), .B(new_n17048_), .ZN(new_n17060_));
  AOI21_X1   g16868(.A1(new_n17057_), .A2(new_n17038_), .B(new_n2912_), .ZN(new_n17061_));
  OAI21_X1   g16869(.A1(new_n17060_), .A2(new_n17061_), .B(\asqrt[42] ), .ZN(new_n17062_));
  AOI21_X1   g16870(.A1(new_n17044_), .A2(new_n17062_), .B(new_n2464_), .ZN(new_n17063_));
  NOR2_X1    g16871(.A1(new_n17047_), .A2(new_n17063_), .ZN(new_n17064_));
  AOI21_X1   g16872(.A1(new_n17064_), .A2(new_n2271_), .B(new_n16701_), .ZN(new_n17065_));
  OAI21_X1   g16873(.A1(new_n17047_), .A2(new_n17063_), .B(\asqrt[44] ), .ZN(new_n17066_));
  NAND2_X1   g16874(.A1(new_n17066_), .A2(new_n2072_), .ZN(new_n17067_));
  OAI21_X1   g16875(.A1(new_n17065_), .A2(new_n17067_), .B(new_n16697_), .ZN(new_n17068_));
  INV_X1     g16876(.I(new_n17066_), .ZN(new_n17069_));
  OAI21_X1   g16877(.A1(new_n17065_), .A2(new_n17069_), .B(\asqrt[45] ), .ZN(new_n17070_));
  NAND3_X1   g16878(.A1(new_n17068_), .A2(new_n17070_), .A3(new_n1884_), .ZN(new_n17071_));
  NAND2_X1   g16879(.A1(new_n17071_), .A2(new_n16695_), .ZN(new_n17072_));
  NAND2_X1   g16880(.A1(new_n17068_), .A2(new_n17070_), .ZN(new_n17073_));
  AOI21_X1   g16881(.A1(new_n17073_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n17074_));
  AOI21_X1   g16882(.A1(new_n17074_), .A2(new_n17072_), .B(new_n16692_), .ZN(new_n17075_));
  INV_X1     g16883(.I(new_n16697_), .ZN(new_n17076_));
  INV_X1     g16884(.I(new_n16707_), .ZN(new_n17077_));
  NOR2_X1    g16885(.A1(new_n17060_), .A2(new_n17061_), .ZN(new_n17078_));
  AOI21_X1   g16886(.A1(new_n17078_), .A2(new_n2699_), .B(new_n17077_), .ZN(new_n17079_));
  NAND2_X1   g16887(.A1(new_n17062_), .A2(new_n2464_), .ZN(new_n17080_));
  OAI21_X1   g16888(.A1(new_n17079_), .A2(new_n17080_), .B(new_n16703_), .ZN(new_n17081_));
  INV_X1     g16889(.I(new_n17062_), .ZN(new_n17082_));
  OAI21_X1   g16890(.A1(new_n17079_), .A2(new_n17082_), .B(\asqrt[43] ), .ZN(new_n17083_));
  NAND3_X1   g16891(.A1(new_n17081_), .A2(new_n17083_), .A3(new_n2271_), .ZN(new_n17084_));
  NAND2_X1   g16892(.A1(new_n17084_), .A2(new_n16700_), .ZN(new_n17085_));
  NAND2_X1   g16893(.A1(new_n17081_), .A2(new_n17083_), .ZN(new_n17086_));
  AOI21_X1   g16894(.A1(new_n17086_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n17087_));
  AOI21_X1   g16895(.A1(new_n17087_), .A2(new_n17085_), .B(new_n17076_), .ZN(new_n17088_));
  AOI21_X1   g16896(.A1(new_n17085_), .A2(new_n17066_), .B(new_n2072_), .ZN(new_n17089_));
  OAI21_X1   g16897(.A1(new_n17088_), .A2(new_n17089_), .B(\asqrt[46] ), .ZN(new_n17090_));
  AOI21_X1   g16898(.A1(new_n17072_), .A2(new_n17090_), .B(new_n1688_), .ZN(new_n17091_));
  NOR2_X1    g16899(.A1(new_n17075_), .A2(new_n17091_), .ZN(new_n17092_));
  AOI21_X1   g16900(.A1(new_n17092_), .A2(new_n1533_), .B(new_n16689_), .ZN(new_n17093_));
  OAI21_X1   g16901(.A1(new_n17075_), .A2(new_n17091_), .B(\asqrt[48] ), .ZN(new_n17094_));
  NAND2_X1   g16902(.A1(new_n17094_), .A2(new_n1368_), .ZN(new_n17095_));
  OAI21_X1   g16903(.A1(new_n17093_), .A2(new_n17095_), .B(new_n16685_), .ZN(new_n17096_));
  INV_X1     g16904(.I(new_n17094_), .ZN(new_n17097_));
  OAI21_X1   g16905(.A1(new_n17093_), .A2(new_n17097_), .B(\asqrt[49] ), .ZN(new_n17098_));
  NAND3_X1   g16906(.A1(new_n17096_), .A2(new_n17098_), .A3(new_n1228_), .ZN(new_n17099_));
  NAND2_X1   g16907(.A1(new_n17099_), .A2(new_n16683_), .ZN(new_n17100_));
  NAND2_X1   g16908(.A1(new_n17096_), .A2(new_n17098_), .ZN(new_n17101_));
  AOI21_X1   g16909(.A1(new_n17101_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n17102_));
  AOI21_X1   g16910(.A1(new_n17102_), .A2(new_n17100_), .B(new_n16680_), .ZN(new_n17103_));
  INV_X1     g16911(.I(new_n16685_), .ZN(new_n17104_));
  INV_X1     g16912(.I(new_n16695_), .ZN(new_n17105_));
  NOR2_X1    g16913(.A1(new_n17088_), .A2(new_n17089_), .ZN(new_n17106_));
  AOI21_X1   g16914(.A1(new_n17106_), .A2(new_n1884_), .B(new_n17105_), .ZN(new_n17107_));
  NAND2_X1   g16915(.A1(new_n17090_), .A2(new_n1688_), .ZN(new_n17108_));
  OAI21_X1   g16916(.A1(new_n17107_), .A2(new_n17108_), .B(new_n16691_), .ZN(new_n17109_));
  INV_X1     g16917(.I(new_n17090_), .ZN(new_n17110_));
  OAI21_X1   g16918(.A1(new_n17107_), .A2(new_n17110_), .B(\asqrt[47] ), .ZN(new_n17111_));
  NAND3_X1   g16919(.A1(new_n17109_), .A2(new_n17111_), .A3(new_n1533_), .ZN(new_n17112_));
  NAND2_X1   g16920(.A1(new_n17112_), .A2(new_n16688_), .ZN(new_n17113_));
  NAND2_X1   g16921(.A1(new_n17109_), .A2(new_n17111_), .ZN(new_n17114_));
  AOI21_X1   g16922(.A1(new_n17114_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n17115_));
  AOI21_X1   g16923(.A1(new_n17115_), .A2(new_n17113_), .B(new_n17104_), .ZN(new_n17116_));
  AOI21_X1   g16924(.A1(new_n17113_), .A2(new_n17094_), .B(new_n1368_), .ZN(new_n17117_));
  OAI21_X1   g16925(.A1(new_n17116_), .A2(new_n17117_), .B(\asqrt[50] ), .ZN(new_n17118_));
  AOI21_X1   g16926(.A1(new_n17100_), .A2(new_n17118_), .B(new_n1088_), .ZN(new_n17119_));
  NOR2_X1    g16927(.A1(new_n17103_), .A2(new_n17119_), .ZN(new_n17120_));
  AOI21_X1   g16928(.A1(new_n17120_), .A2(new_n962_), .B(new_n16677_), .ZN(new_n17121_));
  OAI21_X1   g16929(.A1(new_n17103_), .A2(new_n17119_), .B(\asqrt[52] ), .ZN(new_n17122_));
  NAND2_X1   g16930(.A1(new_n17122_), .A2(new_n842_), .ZN(new_n17123_));
  OAI21_X1   g16931(.A1(new_n17121_), .A2(new_n17123_), .B(new_n16673_), .ZN(new_n17124_));
  INV_X1     g16932(.I(new_n17122_), .ZN(new_n17125_));
  OAI21_X1   g16933(.A1(new_n17121_), .A2(new_n17125_), .B(\asqrt[53] ), .ZN(new_n17126_));
  NAND3_X1   g16934(.A1(new_n17124_), .A2(new_n17126_), .A3(new_n720_), .ZN(new_n17127_));
  NAND2_X1   g16935(.A1(new_n17127_), .A2(new_n16671_), .ZN(new_n17128_));
  NAND2_X1   g16936(.A1(new_n17124_), .A2(new_n17126_), .ZN(new_n17129_));
  AOI21_X1   g16937(.A1(new_n17129_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n17130_));
  AOI21_X1   g16938(.A1(new_n17130_), .A2(new_n17128_), .B(new_n16668_), .ZN(new_n17131_));
  INV_X1     g16939(.I(new_n16673_), .ZN(new_n17132_));
  INV_X1     g16940(.I(new_n16683_), .ZN(new_n17133_));
  NOR2_X1    g16941(.A1(new_n17116_), .A2(new_n17117_), .ZN(new_n17134_));
  AOI21_X1   g16942(.A1(new_n17134_), .A2(new_n1228_), .B(new_n17133_), .ZN(new_n17135_));
  NAND2_X1   g16943(.A1(new_n17118_), .A2(new_n1088_), .ZN(new_n17136_));
  OAI21_X1   g16944(.A1(new_n17135_), .A2(new_n17136_), .B(new_n16679_), .ZN(new_n17137_));
  INV_X1     g16945(.I(new_n17118_), .ZN(new_n17138_));
  OAI21_X1   g16946(.A1(new_n17135_), .A2(new_n17138_), .B(\asqrt[51] ), .ZN(new_n17139_));
  NAND3_X1   g16947(.A1(new_n17137_), .A2(new_n17139_), .A3(new_n962_), .ZN(new_n17140_));
  NAND2_X1   g16948(.A1(new_n17140_), .A2(new_n16676_), .ZN(new_n17141_));
  NAND2_X1   g16949(.A1(new_n17137_), .A2(new_n17139_), .ZN(new_n17142_));
  AOI21_X1   g16950(.A1(new_n17142_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n17143_));
  AOI21_X1   g16951(.A1(new_n17143_), .A2(new_n17141_), .B(new_n17132_), .ZN(new_n17144_));
  AOI21_X1   g16952(.A1(new_n17141_), .A2(new_n17122_), .B(new_n842_), .ZN(new_n17145_));
  OAI21_X1   g16953(.A1(new_n17144_), .A2(new_n17145_), .B(\asqrt[54] ), .ZN(new_n17146_));
  AOI21_X1   g16954(.A1(new_n17128_), .A2(new_n17146_), .B(new_n630_), .ZN(new_n17147_));
  NOR2_X1    g16955(.A1(new_n17131_), .A2(new_n17147_), .ZN(new_n17148_));
  AOI21_X1   g16956(.A1(new_n17148_), .A2(new_n545_), .B(new_n16665_), .ZN(new_n17149_));
  OAI21_X1   g16957(.A1(new_n17131_), .A2(new_n17147_), .B(\asqrt[56] ), .ZN(new_n17150_));
  NAND2_X1   g16958(.A1(new_n17150_), .A2(new_n450_), .ZN(new_n17151_));
  OAI21_X1   g16959(.A1(new_n17149_), .A2(new_n17151_), .B(new_n16661_), .ZN(new_n17152_));
  INV_X1     g16960(.I(new_n17150_), .ZN(new_n17153_));
  OAI21_X1   g16961(.A1(new_n17149_), .A2(new_n17153_), .B(\asqrt[57] ), .ZN(new_n17154_));
  NAND3_X1   g16962(.A1(new_n17152_), .A2(new_n17154_), .A3(new_n403_), .ZN(new_n17155_));
  INV_X1     g16963(.I(new_n16661_), .ZN(new_n17156_));
  INV_X1     g16964(.I(new_n16671_), .ZN(new_n17157_));
  NOR2_X1    g16965(.A1(new_n17144_), .A2(new_n17145_), .ZN(new_n17158_));
  AOI21_X1   g16966(.A1(new_n17158_), .A2(new_n720_), .B(new_n17157_), .ZN(new_n17159_));
  NAND2_X1   g16967(.A1(new_n17146_), .A2(new_n630_), .ZN(new_n17160_));
  OAI21_X1   g16968(.A1(new_n17159_), .A2(new_n17160_), .B(new_n16667_), .ZN(new_n17161_));
  INV_X1     g16969(.I(new_n17146_), .ZN(new_n17162_));
  OAI21_X1   g16970(.A1(new_n17159_), .A2(new_n17162_), .B(\asqrt[55] ), .ZN(new_n17163_));
  NAND3_X1   g16971(.A1(new_n17161_), .A2(new_n17163_), .A3(new_n545_), .ZN(new_n17164_));
  NAND2_X1   g16972(.A1(new_n17164_), .A2(new_n16664_), .ZN(new_n17165_));
  NAND2_X1   g16973(.A1(new_n17161_), .A2(new_n17163_), .ZN(new_n17166_));
  AOI21_X1   g16974(.A1(new_n17166_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n17167_));
  AOI21_X1   g16975(.A1(new_n17167_), .A2(new_n17165_), .B(new_n17156_), .ZN(new_n17168_));
  AOI21_X1   g16976(.A1(new_n17165_), .A2(new_n17150_), .B(new_n450_), .ZN(new_n17169_));
  OAI21_X1   g16977(.A1(new_n17168_), .A2(new_n17169_), .B(\asqrt[58] ), .ZN(new_n17170_));
  NOR2_X1    g16978(.A1(new_n16646_), .A2(new_n16643_), .ZN(new_n17171_));
  INV_X1     g16979(.I(new_n17171_), .ZN(new_n17172_));
  NAND2_X1   g16980(.A1(new_n17172_), .A2(new_n16098_), .ZN(new_n17173_));
  NOR2_X1    g16981(.A1(new_n16649_), .A2(new_n16098_), .ZN(new_n17174_));
  NAND2_X1   g16982(.A1(new_n17174_), .A2(new_n17171_), .ZN(new_n17175_));
  AOI21_X1   g16983(.A1(new_n17175_), .A2(new_n17173_), .B(new_n193_), .ZN(new_n17176_));
  INV_X1     g16984(.I(new_n17176_), .ZN(new_n17177_));
  NAND3_X1   g16985(.A1(\asqrt[7] ), .A2(new_n16628_), .A3(new_n16639_), .ZN(new_n17178_));
  XOR2_X1    g16986(.A1(new_n17178_), .A2(new_n16645_), .Z(new_n17179_));
  INV_X1     g16987(.I(new_n17179_), .ZN(new_n17180_));
  NAND2_X1   g16988(.A1(new_n17174_), .A2(new_n17172_), .ZN(new_n17181_));
  NAND2_X1   g16989(.A1(new_n17181_), .A2(new_n16657_), .ZN(new_n17182_));
  INV_X1     g16990(.I(new_n17182_), .ZN(new_n17183_));
  OAI21_X1   g16991(.A1(new_n16598_), .A2(new_n16600_), .B(new_n16603_), .ZN(new_n17184_));
  NOR2_X1    g16992(.A1(new_n16649_), .A2(new_n17184_), .ZN(new_n17185_));
  XOR2_X1    g16993(.A1(new_n17185_), .A2(new_n16106_), .Z(new_n17186_));
  NAND3_X1   g16994(.A1(\asqrt[7] ), .A2(new_n16614_), .A3(new_n16599_), .ZN(new_n17187_));
  XOR2_X1    g16995(.A1(new_n17187_), .A2(new_n16110_), .Z(new_n17188_));
  NOR2_X1    g16996(.A1(new_n17168_), .A2(new_n17169_), .ZN(new_n17189_));
  AOI21_X1   g16997(.A1(new_n17189_), .A2(new_n403_), .B(new_n16653_), .ZN(new_n17190_));
  NAND2_X1   g16998(.A1(new_n17170_), .A2(new_n339_), .ZN(new_n17191_));
  OAI21_X1   g16999(.A1(new_n17190_), .A2(new_n17191_), .B(new_n17188_), .ZN(new_n17192_));
  INV_X1     g17000(.I(new_n17170_), .ZN(new_n17193_));
  OAI21_X1   g17001(.A1(new_n17190_), .A2(new_n17193_), .B(\asqrt[59] ), .ZN(new_n17194_));
  NAND3_X1   g17002(.A1(new_n17192_), .A2(new_n17194_), .A3(new_n288_), .ZN(new_n17195_));
  NAND2_X1   g17003(.A1(new_n17195_), .A2(new_n17186_), .ZN(new_n17196_));
  INV_X1     g17004(.I(new_n17188_), .ZN(new_n17197_));
  NAND2_X1   g17005(.A1(new_n17155_), .A2(new_n16652_), .ZN(new_n17198_));
  NAND2_X1   g17006(.A1(new_n17152_), .A2(new_n17154_), .ZN(new_n17199_));
  AOI21_X1   g17007(.A1(new_n17199_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n17200_));
  AOI21_X1   g17008(.A1(new_n17200_), .A2(new_n17198_), .B(new_n17197_), .ZN(new_n17201_));
  AOI21_X1   g17009(.A1(new_n17198_), .A2(new_n17170_), .B(new_n339_), .ZN(new_n17202_));
  OAI21_X1   g17010(.A1(new_n17201_), .A2(new_n17202_), .B(\asqrt[60] ), .ZN(new_n17203_));
  AOI21_X1   g17011(.A1(new_n17196_), .A2(new_n17203_), .B(new_n242_), .ZN(new_n17204_));
  NAND3_X1   g17012(.A1(\asqrt[7] ), .A2(new_n16604_), .A3(new_n16620_), .ZN(new_n17205_));
  XOR2_X1    g17013(.A1(new_n17205_), .A2(new_n16632_), .Z(new_n17206_));
  INV_X1     g17014(.I(new_n17206_), .ZN(new_n17207_));
  NAND2_X1   g17015(.A1(new_n17192_), .A2(new_n17194_), .ZN(new_n17208_));
  AOI21_X1   g17016(.A1(new_n17208_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n17209_));
  AOI21_X1   g17017(.A1(new_n17209_), .A2(new_n17196_), .B(new_n17207_), .ZN(new_n17210_));
  OAI21_X1   g17018(.A1(new_n17210_), .A2(new_n17204_), .B(\asqrt[62] ), .ZN(new_n17211_));
  INV_X1     g17019(.I(new_n17211_), .ZN(new_n17212_));
  NOR2_X1    g17020(.A1(new_n17210_), .A2(new_n17204_), .ZN(new_n17213_));
  AOI21_X1   g17021(.A1(new_n16605_), .A2(new_n16626_), .B(new_n16621_), .ZN(new_n17214_));
  NAND2_X1   g17022(.A1(\asqrt[7] ), .A2(new_n17214_), .ZN(new_n17215_));
  XOR2_X1    g17023(.A1(new_n17215_), .A2(new_n16624_), .Z(new_n17216_));
  INV_X1     g17024(.I(new_n17216_), .ZN(new_n17217_));
  AOI21_X1   g17025(.A1(new_n17213_), .A2(new_n234_), .B(new_n17217_), .ZN(new_n17218_));
  OAI21_X1   g17026(.A1(new_n17218_), .A2(new_n17212_), .B(new_n17183_), .ZN(new_n17219_));
  OAI21_X1   g17027(.A1(new_n17219_), .A2(new_n17180_), .B(new_n193_), .ZN(new_n17220_));
  NOR3_X1    g17028(.A1(new_n17218_), .A2(new_n17212_), .A3(new_n17179_), .ZN(new_n17221_));
  INV_X1     g17029(.I(new_n17221_), .ZN(new_n17222_));
  NOR2_X1    g17030(.A1(\asqrt[7] ), .A2(new_n16099_), .ZN(new_n17223_));
  INV_X1     g17031(.I(new_n17223_), .ZN(new_n17224_));
  NAND4_X1   g17032(.A1(new_n17220_), .A2(new_n17177_), .A3(new_n17222_), .A4(new_n17224_), .ZN(\asqrt[6] ));
  NAND3_X1   g17033(.A1(\asqrt[6] ), .A2(new_n17155_), .A3(new_n17170_), .ZN(new_n17226_));
  XOR2_X1    g17034(.A1(new_n17226_), .A2(new_n16653_), .Z(new_n17227_));
  NOR2_X1    g17035(.A1(new_n17218_), .A2(new_n17212_), .ZN(new_n17228_));
  INV_X1     g17036(.I(new_n17228_), .ZN(new_n17229_));
  NAND2_X1   g17037(.A1(new_n17229_), .A2(new_n17180_), .ZN(new_n17230_));
  INV_X1     g17038(.I(new_n17186_), .ZN(new_n17231_));
  NOR2_X1    g17039(.A1(new_n17201_), .A2(new_n17202_), .ZN(new_n17232_));
  AOI21_X1   g17040(.A1(new_n17232_), .A2(new_n288_), .B(new_n17231_), .ZN(new_n17233_));
  INV_X1     g17041(.I(new_n17203_), .ZN(new_n17234_));
  OAI21_X1   g17042(.A1(new_n17233_), .A2(new_n17234_), .B(\asqrt[61] ), .ZN(new_n17235_));
  NAND2_X1   g17043(.A1(new_n17203_), .A2(new_n242_), .ZN(new_n17236_));
  OAI21_X1   g17044(.A1(new_n17233_), .A2(new_n17236_), .B(new_n17206_), .ZN(new_n17237_));
  NAND3_X1   g17045(.A1(new_n17237_), .A2(new_n17235_), .A3(new_n234_), .ZN(new_n17238_));
  NAND2_X1   g17046(.A1(new_n17238_), .A2(new_n17216_), .ZN(new_n17239_));
  AOI21_X1   g17047(.A1(new_n17239_), .A2(new_n17211_), .B(new_n17182_), .ZN(new_n17240_));
  AOI21_X1   g17048(.A1(new_n17240_), .A2(new_n17179_), .B(\asqrt[63] ), .ZN(new_n17241_));
  NOR4_X1    g17049(.A1(new_n17241_), .A2(new_n17176_), .A3(new_n17221_), .A4(new_n17223_), .ZN(new_n17242_));
  NOR2_X1    g17050(.A1(new_n17242_), .A2(new_n17180_), .ZN(new_n17243_));
  NAND2_X1   g17051(.A1(new_n17243_), .A2(new_n17228_), .ZN(new_n17244_));
  AOI21_X1   g17052(.A1(new_n17244_), .A2(new_n17230_), .B(new_n193_), .ZN(new_n17245_));
  NAND3_X1   g17053(.A1(\asqrt[6] ), .A2(new_n17211_), .A3(new_n17238_), .ZN(new_n17246_));
  XOR2_X1    g17054(.A1(new_n17246_), .A2(new_n17217_), .Z(new_n17247_));
  NAND2_X1   g17055(.A1(new_n17243_), .A2(new_n17229_), .ZN(new_n17248_));
  NAND2_X1   g17056(.A1(new_n17248_), .A2(new_n17222_), .ZN(new_n17249_));
  OAI21_X1   g17057(.A1(new_n17190_), .A2(new_n17191_), .B(new_n17194_), .ZN(new_n17250_));
  NOR2_X1    g17058(.A1(new_n17242_), .A2(new_n17250_), .ZN(new_n17251_));
  XOR2_X1    g17059(.A1(new_n17251_), .A2(new_n17188_), .Z(new_n17252_));
  OAI21_X1   g17060(.A1(new_n17149_), .A2(new_n17151_), .B(new_n17154_), .ZN(new_n17253_));
  NOR2_X1    g17061(.A1(new_n17242_), .A2(new_n17253_), .ZN(new_n17254_));
  XOR2_X1    g17062(.A1(new_n17254_), .A2(new_n16661_), .Z(new_n17255_));
  INV_X1     g17063(.I(new_n17255_), .ZN(new_n17256_));
  NAND3_X1   g17064(.A1(\asqrt[6] ), .A2(new_n17164_), .A3(new_n17150_), .ZN(new_n17257_));
  XOR2_X1    g17065(.A1(new_n17257_), .A2(new_n16665_), .Z(new_n17258_));
  INV_X1     g17066(.I(new_n17258_), .ZN(new_n17259_));
  OAI21_X1   g17067(.A1(new_n17159_), .A2(new_n17160_), .B(new_n17163_), .ZN(new_n17260_));
  NOR2_X1    g17068(.A1(new_n17242_), .A2(new_n17260_), .ZN(new_n17261_));
  XOR2_X1    g17069(.A1(new_n17261_), .A2(new_n16667_), .Z(new_n17262_));
  NAND3_X1   g17070(.A1(\asqrt[6] ), .A2(new_n17127_), .A3(new_n17146_), .ZN(new_n17263_));
  XOR2_X1    g17071(.A1(new_n17263_), .A2(new_n17157_), .Z(new_n17264_));
  OAI21_X1   g17072(.A1(new_n17121_), .A2(new_n17123_), .B(new_n17126_), .ZN(new_n17265_));
  NOR2_X1    g17073(.A1(new_n17242_), .A2(new_n17265_), .ZN(new_n17266_));
  XOR2_X1    g17074(.A1(new_n17266_), .A2(new_n16673_), .Z(new_n17267_));
  INV_X1     g17075(.I(new_n17267_), .ZN(new_n17268_));
  NAND3_X1   g17076(.A1(\asqrt[6] ), .A2(new_n17140_), .A3(new_n17122_), .ZN(new_n17269_));
  XOR2_X1    g17077(.A1(new_n17269_), .A2(new_n16677_), .Z(new_n17270_));
  INV_X1     g17078(.I(new_n17270_), .ZN(new_n17271_));
  OAI21_X1   g17079(.A1(new_n17135_), .A2(new_n17136_), .B(new_n17139_), .ZN(new_n17272_));
  NOR2_X1    g17080(.A1(new_n17242_), .A2(new_n17272_), .ZN(new_n17273_));
  XOR2_X1    g17081(.A1(new_n17273_), .A2(new_n16679_), .Z(new_n17274_));
  NAND3_X1   g17082(.A1(\asqrt[6] ), .A2(new_n17099_), .A3(new_n17118_), .ZN(new_n17275_));
  XOR2_X1    g17083(.A1(new_n17275_), .A2(new_n17133_), .Z(new_n17276_));
  OAI21_X1   g17084(.A1(new_n17093_), .A2(new_n17095_), .B(new_n17098_), .ZN(new_n17277_));
  NOR2_X1    g17085(.A1(new_n17242_), .A2(new_n17277_), .ZN(new_n17278_));
  XOR2_X1    g17086(.A1(new_n17278_), .A2(new_n16685_), .Z(new_n17279_));
  INV_X1     g17087(.I(new_n17279_), .ZN(new_n17280_));
  NAND3_X1   g17088(.A1(\asqrt[6] ), .A2(new_n17112_), .A3(new_n17094_), .ZN(new_n17281_));
  XOR2_X1    g17089(.A1(new_n17281_), .A2(new_n16689_), .Z(new_n17282_));
  INV_X1     g17090(.I(new_n17282_), .ZN(new_n17283_));
  OAI21_X1   g17091(.A1(new_n17107_), .A2(new_n17108_), .B(new_n17111_), .ZN(new_n17284_));
  NOR2_X1    g17092(.A1(new_n17242_), .A2(new_n17284_), .ZN(new_n17285_));
  XOR2_X1    g17093(.A1(new_n17285_), .A2(new_n16691_), .Z(new_n17286_));
  NAND3_X1   g17094(.A1(\asqrt[6] ), .A2(new_n17071_), .A3(new_n17090_), .ZN(new_n17287_));
  XOR2_X1    g17095(.A1(new_n17287_), .A2(new_n17105_), .Z(new_n17288_));
  OAI21_X1   g17096(.A1(new_n17065_), .A2(new_n17067_), .B(new_n17070_), .ZN(new_n17289_));
  NOR2_X1    g17097(.A1(new_n17242_), .A2(new_n17289_), .ZN(new_n17290_));
  XOR2_X1    g17098(.A1(new_n17290_), .A2(new_n16697_), .Z(new_n17291_));
  INV_X1     g17099(.I(new_n17291_), .ZN(new_n17292_));
  NAND3_X1   g17100(.A1(\asqrt[6] ), .A2(new_n17084_), .A3(new_n17066_), .ZN(new_n17293_));
  XOR2_X1    g17101(.A1(new_n17293_), .A2(new_n16701_), .Z(new_n17294_));
  INV_X1     g17102(.I(new_n17294_), .ZN(new_n17295_));
  OAI21_X1   g17103(.A1(new_n17079_), .A2(new_n17080_), .B(new_n17083_), .ZN(new_n17296_));
  NOR2_X1    g17104(.A1(new_n17242_), .A2(new_n17296_), .ZN(new_n17297_));
  XOR2_X1    g17105(.A1(new_n17297_), .A2(new_n16703_), .Z(new_n17298_));
  NAND3_X1   g17106(.A1(\asqrt[6] ), .A2(new_n17043_), .A3(new_n17062_), .ZN(new_n17299_));
  XOR2_X1    g17107(.A1(new_n17299_), .A2(new_n17077_), .Z(new_n17300_));
  OAI21_X1   g17108(.A1(new_n17037_), .A2(new_n17039_), .B(new_n17042_), .ZN(new_n17301_));
  NOR2_X1    g17109(.A1(new_n17242_), .A2(new_n17301_), .ZN(new_n17302_));
  XOR2_X1    g17110(.A1(new_n17302_), .A2(new_n16709_), .Z(new_n17303_));
  INV_X1     g17111(.I(new_n17303_), .ZN(new_n17304_));
  NAND3_X1   g17112(.A1(\asqrt[6] ), .A2(new_n17056_), .A3(new_n17038_), .ZN(new_n17305_));
  XOR2_X1    g17113(.A1(new_n17305_), .A2(new_n16713_), .Z(new_n17306_));
  INV_X1     g17114(.I(new_n17306_), .ZN(new_n17307_));
  OAI21_X1   g17115(.A1(new_n17051_), .A2(new_n17052_), .B(new_n17055_), .ZN(new_n17308_));
  NOR2_X1    g17116(.A1(new_n17242_), .A2(new_n17308_), .ZN(new_n17309_));
  XOR2_X1    g17117(.A1(new_n17309_), .A2(new_n16715_), .Z(new_n17310_));
  NAND3_X1   g17118(.A1(\asqrt[6] ), .A2(new_n17015_), .A3(new_n17034_), .ZN(new_n17311_));
  XOR2_X1    g17119(.A1(new_n17311_), .A2(new_n17049_), .Z(new_n17312_));
  OAI21_X1   g17120(.A1(new_n17009_), .A2(new_n17011_), .B(new_n17014_), .ZN(new_n17313_));
  NOR2_X1    g17121(.A1(new_n17242_), .A2(new_n17313_), .ZN(new_n17314_));
  XOR2_X1    g17122(.A1(new_n17314_), .A2(new_n16721_), .Z(new_n17315_));
  INV_X1     g17123(.I(new_n17315_), .ZN(new_n17316_));
  NAND3_X1   g17124(.A1(\asqrt[6] ), .A2(new_n17028_), .A3(new_n17010_), .ZN(new_n17317_));
  XOR2_X1    g17125(.A1(new_n17317_), .A2(new_n16725_), .Z(new_n17318_));
  INV_X1     g17126(.I(new_n17318_), .ZN(new_n17319_));
  OAI21_X1   g17127(.A1(new_n17023_), .A2(new_n17024_), .B(new_n17027_), .ZN(new_n17320_));
  NOR2_X1    g17128(.A1(new_n17242_), .A2(new_n17320_), .ZN(new_n17321_));
  XOR2_X1    g17129(.A1(new_n17321_), .A2(new_n16727_), .Z(new_n17322_));
  NAND3_X1   g17130(.A1(\asqrt[6] ), .A2(new_n16987_), .A3(new_n17006_), .ZN(new_n17323_));
  XOR2_X1    g17131(.A1(new_n17323_), .A2(new_n17021_), .Z(new_n17324_));
  OAI21_X1   g17132(.A1(new_n16981_), .A2(new_n16983_), .B(new_n16986_), .ZN(new_n17325_));
  NOR2_X1    g17133(.A1(new_n17242_), .A2(new_n17325_), .ZN(new_n17326_));
  XOR2_X1    g17134(.A1(new_n17326_), .A2(new_n16733_), .Z(new_n17327_));
  INV_X1     g17135(.I(new_n17327_), .ZN(new_n17328_));
  NAND3_X1   g17136(.A1(\asqrt[6] ), .A2(new_n17000_), .A3(new_n16982_), .ZN(new_n17329_));
  XOR2_X1    g17137(.A1(new_n17329_), .A2(new_n16737_), .Z(new_n17330_));
  INV_X1     g17138(.I(new_n17330_), .ZN(new_n17331_));
  OAI21_X1   g17139(.A1(new_n16995_), .A2(new_n16996_), .B(new_n16999_), .ZN(new_n17332_));
  NOR2_X1    g17140(.A1(new_n17242_), .A2(new_n17332_), .ZN(new_n17333_));
  XOR2_X1    g17141(.A1(new_n17333_), .A2(new_n16739_), .Z(new_n17334_));
  NAND3_X1   g17142(.A1(\asqrt[6] ), .A2(new_n16959_), .A3(new_n16978_), .ZN(new_n17335_));
  XOR2_X1    g17143(.A1(new_n17335_), .A2(new_n16993_), .Z(new_n17336_));
  OAI21_X1   g17144(.A1(new_n16953_), .A2(new_n16955_), .B(new_n16958_), .ZN(new_n17337_));
  NOR2_X1    g17145(.A1(new_n17242_), .A2(new_n17337_), .ZN(new_n17338_));
  XOR2_X1    g17146(.A1(new_n17338_), .A2(new_n16745_), .Z(new_n17339_));
  INV_X1     g17147(.I(new_n17339_), .ZN(new_n17340_));
  NAND3_X1   g17148(.A1(\asqrt[6] ), .A2(new_n16972_), .A3(new_n16954_), .ZN(new_n17341_));
  XOR2_X1    g17149(.A1(new_n17341_), .A2(new_n16749_), .Z(new_n17342_));
  INV_X1     g17150(.I(new_n17342_), .ZN(new_n17343_));
  OAI21_X1   g17151(.A1(new_n16967_), .A2(new_n16968_), .B(new_n16971_), .ZN(new_n17344_));
  NOR2_X1    g17152(.A1(new_n17242_), .A2(new_n17344_), .ZN(new_n17345_));
  XOR2_X1    g17153(.A1(new_n17345_), .A2(new_n16751_), .Z(new_n17346_));
  NAND3_X1   g17154(.A1(\asqrt[6] ), .A2(new_n16931_), .A3(new_n16950_), .ZN(new_n17347_));
  XOR2_X1    g17155(.A1(new_n17347_), .A2(new_n16965_), .Z(new_n17348_));
  OAI21_X1   g17156(.A1(new_n16925_), .A2(new_n16927_), .B(new_n16930_), .ZN(new_n17349_));
  NOR2_X1    g17157(.A1(new_n17242_), .A2(new_n17349_), .ZN(new_n17350_));
  XOR2_X1    g17158(.A1(new_n17350_), .A2(new_n16757_), .Z(new_n17351_));
  INV_X1     g17159(.I(new_n17351_), .ZN(new_n17352_));
  NAND3_X1   g17160(.A1(\asqrt[6] ), .A2(new_n16944_), .A3(new_n16926_), .ZN(new_n17353_));
  XOR2_X1    g17161(.A1(new_n17353_), .A2(new_n16761_), .Z(new_n17354_));
  INV_X1     g17162(.I(new_n17354_), .ZN(new_n17355_));
  OAI21_X1   g17163(.A1(new_n16939_), .A2(new_n16940_), .B(new_n16943_), .ZN(new_n17356_));
  NOR2_X1    g17164(.A1(new_n17242_), .A2(new_n17356_), .ZN(new_n17357_));
  XOR2_X1    g17165(.A1(new_n17357_), .A2(new_n16763_), .Z(new_n17358_));
  NAND3_X1   g17166(.A1(\asqrt[6] ), .A2(new_n16903_), .A3(new_n16922_), .ZN(new_n17359_));
  XOR2_X1    g17167(.A1(new_n17359_), .A2(new_n16937_), .Z(new_n17360_));
  OAI21_X1   g17168(.A1(new_n16897_), .A2(new_n16899_), .B(new_n16902_), .ZN(new_n17361_));
  NOR2_X1    g17169(.A1(new_n17242_), .A2(new_n17361_), .ZN(new_n17362_));
  XOR2_X1    g17170(.A1(new_n17362_), .A2(new_n16769_), .Z(new_n17363_));
  INV_X1     g17171(.I(new_n17363_), .ZN(new_n17364_));
  NAND3_X1   g17172(.A1(\asqrt[6] ), .A2(new_n16916_), .A3(new_n16898_), .ZN(new_n17365_));
  XOR2_X1    g17173(.A1(new_n17365_), .A2(new_n16773_), .Z(new_n17366_));
  INV_X1     g17174(.I(new_n17366_), .ZN(new_n17367_));
  OAI21_X1   g17175(.A1(new_n16911_), .A2(new_n16912_), .B(new_n16915_), .ZN(new_n17368_));
  NOR2_X1    g17176(.A1(new_n17242_), .A2(new_n17368_), .ZN(new_n17369_));
  XOR2_X1    g17177(.A1(new_n17369_), .A2(new_n16775_), .Z(new_n17370_));
  NAND3_X1   g17178(.A1(\asqrt[6] ), .A2(new_n16875_), .A3(new_n16894_), .ZN(new_n17371_));
  XOR2_X1    g17179(.A1(new_n17371_), .A2(new_n16909_), .Z(new_n17372_));
  OAI21_X1   g17180(.A1(new_n16869_), .A2(new_n16871_), .B(new_n16874_), .ZN(new_n17373_));
  NOR2_X1    g17181(.A1(new_n17242_), .A2(new_n17373_), .ZN(new_n17374_));
  XOR2_X1    g17182(.A1(new_n17374_), .A2(new_n16781_), .Z(new_n17375_));
  INV_X1     g17183(.I(new_n17375_), .ZN(new_n17376_));
  NAND3_X1   g17184(.A1(\asqrt[6] ), .A2(new_n16888_), .A3(new_n16870_), .ZN(new_n17377_));
  XOR2_X1    g17185(.A1(new_n17377_), .A2(new_n16785_), .Z(new_n17378_));
  INV_X1     g17186(.I(new_n17378_), .ZN(new_n17379_));
  OAI21_X1   g17187(.A1(new_n16883_), .A2(new_n16884_), .B(new_n16887_), .ZN(new_n17380_));
  NOR2_X1    g17188(.A1(new_n17242_), .A2(new_n17380_), .ZN(new_n17381_));
  XOR2_X1    g17189(.A1(new_n17381_), .A2(new_n16787_), .Z(new_n17382_));
  NAND3_X1   g17190(.A1(\asqrt[6] ), .A2(new_n16847_), .A3(new_n16866_), .ZN(new_n17383_));
  XOR2_X1    g17191(.A1(new_n17383_), .A2(new_n16881_), .Z(new_n17384_));
  AOI21_X1   g17192(.A1(new_n16861_), .A2(new_n16863_), .B(new_n16865_), .ZN(new_n17385_));
  NAND2_X1   g17193(.A1(\asqrt[6] ), .A2(new_n17385_), .ZN(new_n17386_));
  XOR2_X1    g17194(.A1(new_n17386_), .A2(new_n16852_), .Z(new_n17387_));
  INV_X1     g17195(.I(new_n17387_), .ZN(new_n17388_));
  NAND3_X1   g17196(.A1(\asqrt[6] ), .A2(new_n16860_), .A3(new_n16842_), .ZN(new_n17389_));
  XOR2_X1    g17197(.A1(new_n17389_), .A2(new_n16797_), .Z(new_n17390_));
  INV_X1     g17198(.I(new_n17390_), .ZN(new_n17391_));
  OAI21_X1   g17199(.A1(new_n16855_), .A2(new_n16856_), .B(new_n16859_), .ZN(new_n17392_));
  NOR2_X1    g17200(.A1(new_n17242_), .A2(new_n17392_), .ZN(new_n17393_));
  XOR2_X1    g17201(.A1(new_n17393_), .A2(new_n16800_), .Z(new_n17394_));
  NAND3_X1   g17202(.A1(\asqrt[6] ), .A2(new_n16820_), .A3(new_n16838_), .ZN(new_n17395_));
  XOR2_X1    g17203(.A1(new_n17395_), .A2(new_n16854_), .Z(new_n17396_));
  NAND2_X1   g17204(.A1(new_n16835_), .A2(new_n15518_), .ZN(new_n17397_));
  NAND3_X1   g17205(.A1(\asqrt[6] ), .A2(new_n17397_), .A3(new_n16819_), .ZN(new_n17398_));
  XOR2_X1    g17206(.A1(new_n17398_), .A2(new_n16829_), .Z(new_n17399_));
  INV_X1     g17207(.I(new_n17399_), .ZN(new_n17400_));
  NAND3_X1   g17208(.A1(\asqrt[6] ), .A2(new_n16809_), .A3(new_n16810_), .ZN(new_n17401_));
  NOR4_X1    g17209(.A1(new_n17241_), .A2(new_n16649_), .A3(new_n17176_), .A4(new_n17221_), .ZN(new_n17402_));
  INV_X1     g17210(.I(new_n17402_), .ZN(new_n17403_));
  AOI21_X1   g17211(.A1(new_n17401_), .A2(new_n17403_), .B(\a[14] ), .ZN(new_n17404_));
  NOR3_X1    g17212(.A1(new_n17242_), .A2(\a[12] ), .A3(\a[13] ), .ZN(new_n17405_));
  NOR3_X1    g17213(.A1(new_n17405_), .A2(new_n16254_), .A3(new_n17402_), .ZN(new_n17406_));
  NOR2_X1    g17214(.A1(new_n17406_), .A2(new_n17404_), .ZN(new_n17407_));
  INV_X1     g17215(.I(\a[10] ), .ZN(new_n17408_));
  INV_X1     g17216(.I(\a[11] ), .ZN(new_n17409_));
  NAND3_X1   g17217(.A1(new_n17408_), .A2(new_n17409_), .A3(new_n16809_), .ZN(new_n17410_));
  OAI21_X1   g17218(.A1(new_n17242_), .A2(new_n16809_), .B(new_n17410_), .ZN(new_n17411_));
  NAND2_X1   g17219(.A1(new_n17411_), .A2(\asqrt[7] ), .ZN(new_n17412_));
  OAI21_X1   g17220(.A1(new_n17242_), .A2(\a[12] ), .B(\a[13] ), .ZN(new_n17413_));
  NAND2_X1   g17221(.A1(new_n17413_), .A2(new_n17401_), .ZN(new_n17414_));
  NOR2_X1    g17222(.A1(new_n17411_), .A2(\asqrt[7] ), .ZN(new_n17415_));
  OAI21_X1   g17223(.A1(new_n17414_), .A2(new_n17415_), .B(new_n17412_), .ZN(new_n17416_));
  OAI21_X1   g17224(.A1(new_n17416_), .A2(\asqrt[8] ), .B(new_n17407_), .ZN(new_n17417_));
  NAND2_X1   g17225(.A1(new_n17416_), .A2(\asqrt[8] ), .ZN(new_n17418_));
  NAND3_X1   g17226(.A1(new_n17417_), .A2(new_n15518_), .A3(new_n17418_), .ZN(new_n17419_));
  NAND3_X1   g17227(.A1(\asqrt[6] ), .A2(new_n16813_), .A3(new_n16834_), .ZN(new_n17420_));
  XOR2_X1    g17228(.A1(new_n17420_), .A2(new_n16815_), .Z(new_n17421_));
  AOI21_X1   g17229(.A1(new_n17417_), .A2(new_n17418_), .B(new_n15518_), .ZN(new_n17422_));
  AOI21_X1   g17230(.A1(new_n17419_), .A2(new_n17421_), .B(new_n17422_), .ZN(new_n17423_));
  AOI21_X1   g17231(.A1(new_n17423_), .A2(new_n14985_), .B(new_n17400_), .ZN(new_n17424_));
  OAI21_X1   g17232(.A1(new_n17423_), .A2(new_n14985_), .B(new_n14430_), .ZN(new_n17425_));
  OAI21_X1   g17233(.A1(new_n17424_), .A2(new_n17425_), .B(new_n17396_), .ZN(new_n17426_));
  NOR2_X1    g17234(.A1(new_n17423_), .A2(new_n14985_), .ZN(new_n17427_));
  OAI21_X1   g17235(.A1(new_n17424_), .A2(new_n17427_), .B(\asqrt[11] ), .ZN(new_n17428_));
  NAND3_X1   g17236(.A1(new_n17426_), .A2(new_n17428_), .A3(new_n13917_), .ZN(new_n17429_));
  NAND2_X1   g17237(.A1(new_n17429_), .A2(new_n17394_), .ZN(new_n17430_));
  NAND2_X1   g17238(.A1(new_n17426_), .A2(new_n17428_), .ZN(new_n17431_));
  AOI21_X1   g17239(.A1(new_n17431_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n17432_));
  AOI21_X1   g17240(.A1(new_n17432_), .A2(new_n17430_), .B(new_n17391_), .ZN(new_n17433_));
  INV_X1     g17241(.I(new_n17396_), .ZN(new_n17434_));
  OAI21_X1   g17242(.A1(new_n17405_), .A2(new_n17402_), .B(new_n16254_), .ZN(new_n17435_));
  NAND3_X1   g17243(.A1(new_n17401_), .A2(\a[14] ), .A3(new_n17403_), .ZN(new_n17436_));
  NAND2_X1   g17244(.A1(new_n17435_), .A2(new_n17436_), .ZN(new_n17437_));
  NAND2_X1   g17245(.A1(\asqrt[6] ), .A2(\a[12] ), .ZN(new_n17438_));
  AOI21_X1   g17246(.A1(new_n17438_), .A2(new_n17410_), .B(new_n16649_), .ZN(new_n17439_));
  AOI21_X1   g17247(.A1(\asqrt[6] ), .A2(new_n16809_), .B(new_n16810_), .ZN(new_n17440_));
  NOR2_X1    g17248(.A1(new_n17405_), .A2(new_n17440_), .ZN(new_n17441_));
  NAND3_X1   g17249(.A1(new_n17438_), .A2(new_n16649_), .A3(new_n17410_), .ZN(new_n17442_));
  AOI21_X1   g17250(.A1(new_n17441_), .A2(new_n17442_), .B(new_n17439_), .ZN(new_n17443_));
  AOI21_X1   g17251(.A1(new_n17443_), .A2(new_n16093_), .B(new_n17437_), .ZN(new_n17444_));
  NOR2_X1    g17252(.A1(new_n17443_), .A2(new_n16093_), .ZN(new_n17445_));
  NOR3_X1    g17253(.A1(new_n17444_), .A2(\asqrt[9] ), .A3(new_n17445_), .ZN(new_n17446_));
  INV_X1     g17254(.I(new_n17421_), .ZN(new_n17447_));
  OAI21_X1   g17255(.A1(new_n17444_), .A2(new_n17445_), .B(\asqrt[9] ), .ZN(new_n17448_));
  OAI21_X1   g17256(.A1(new_n17446_), .A2(new_n17447_), .B(new_n17448_), .ZN(new_n17449_));
  OAI21_X1   g17257(.A1(new_n17449_), .A2(\asqrt[10] ), .B(new_n17399_), .ZN(new_n17450_));
  AOI21_X1   g17258(.A1(new_n17449_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n17451_));
  AOI21_X1   g17259(.A1(new_n17451_), .A2(new_n17450_), .B(new_n17434_), .ZN(new_n17452_));
  NAND2_X1   g17260(.A1(new_n17449_), .A2(\asqrt[10] ), .ZN(new_n17453_));
  AOI21_X1   g17261(.A1(new_n17450_), .A2(new_n17453_), .B(new_n14430_), .ZN(new_n17454_));
  OAI21_X1   g17262(.A1(new_n17452_), .A2(new_n17454_), .B(\asqrt[12] ), .ZN(new_n17455_));
  AOI21_X1   g17263(.A1(new_n17430_), .A2(new_n17455_), .B(new_n13382_), .ZN(new_n17456_));
  NOR2_X1    g17264(.A1(new_n17433_), .A2(new_n17456_), .ZN(new_n17457_));
  AOI21_X1   g17265(.A1(new_n17457_), .A2(new_n12889_), .B(new_n17388_), .ZN(new_n17458_));
  OAI21_X1   g17266(.A1(new_n17433_), .A2(new_n17456_), .B(\asqrt[14] ), .ZN(new_n17459_));
  NAND2_X1   g17267(.A1(new_n17459_), .A2(new_n12374_), .ZN(new_n17460_));
  OAI21_X1   g17268(.A1(new_n17458_), .A2(new_n17460_), .B(new_n17384_), .ZN(new_n17461_));
  INV_X1     g17269(.I(new_n17459_), .ZN(new_n17462_));
  OAI21_X1   g17270(.A1(new_n17458_), .A2(new_n17462_), .B(\asqrt[15] ), .ZN(new_n17463_));
  NAND3_X1   g17271(.A1(new_n17461_), .A2(new_n17463_), .A3(new_n11901_), .ZN(new_n17464_));
  NAND2_X1   g17272(.A1(new_n17464_), .A2(new_n17382_), .ZN(new_n17465_));
  NAND2_X1   g17273(.A1(new_n17461_), .A2(new_n17463_), .ZN(new_n17466_));
  AOI21_X1   g17274(.A1(new_n17466_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n17467_));
  AOI21_X1   g17275(.A1(new_n17467_), .A2(new_n17465_), .B(new_n17379_), .ZN(new_n17468_));
  INV_X1     g17276(.I(new_n17384_), .ZN(new_n17469_));
  INV_X1     g17277(.I(new_n17394_), .ZN(new_n17470_));
  NOR2_X1    g17278(.A1(new_n17452_), .A2(new_n17454_), .ZN(new_n17471_));
  AOI21_X1   g17279(.A1(new_n17471_), .A2(new_n13917_), .B(new_n17470_), .ZN(new_n17472_));
  NAND2_X1   g17280(.A1(new_n17455_), .A2(new_n13382_), .ZN(new_n17473_));
  OAI21_X1   g17281(.A1(new_n17472_), .A2(new_n17473_), .B(new_n17390_), .ZN(new_n17474_));
  INV_X1     g17282(.I(new_n17455_), .ZN(new_n17475_));
  OAI21_X1   g17283(.A1(new_n17472_), .A2(new_n17475_), .B(\asqrt[13] ), .ZN(new_n17476_));
  NAND3_X1   g17284(.A1(new_n17474_), .A2(new_n17476_), .A3(new_n12889_), .ZN(new_n17477_));
  NAND2_X1   g17285(.A1(new_n17477_), .A2(new_n17387_), .ZN(new_n17478_));
  NAND2_X1   g17286(.A1(new_n17474_), .A2(new_n17476_), .ZN(new_n17479_));
  AOI21_X1   g17287(.A1(new_n17479_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n17480_));
  AOI21_X1   g17288(.A1(new_n17480_), .A2(new_n17478_), .B(new_n17469_), .ZN(new_n17481_));
  AOI21_X1   g17289(.A1(new_n17478_), .A2(new_n17459_), .B(new_n12374_), .ZN(new_n17482_));
  OAI21_X1   g17290(.A1(new_n17481_), .A2(new_n17482_), .B(\asqrt[16] ), .ZN(new_n17483_));
  AOI21_X1   g17291(.A1(new_n17465_), .A2(new_n17483_), .B(new_n11406_), .ZN(new_n17484_));
  NOR2_X1    g17292(.A1(new_n17468_), .A2(new_n17484_), .ZN(new_n17485_));
  AOI21_X1   g17293(.A1(new_n17485_), .A2(new_n10953_), .B(new_n17376_), .ZN(new_n17486_));
  OAI21_X1   g17294(.A1(new_n17468_), .A2(new_n17484_), .B(\asqrt[18] ), .ZN(new_n17487_));
  NAND2_X1   g17295(.A1(new_n17487_), .A2(new_n10478_), .ZN(new_n17488_));
  OAI21_X1   g17296(.A1(new_n17486_), .A2(new_n17488_), .B(new_n17372_), .ZN(new_n17489_));
  INV_X1     g17297(.I(new_n17487_), .ZN(new_n17490_));
  OAI21_X1   g17298(.A1(new_n17486_), .A2(new_n17490_), .B(\asqrt[19] ), .ZN(new_n17491_));
  NAND3_X1   g17299(.A1(new_n17489_), .A2(new_n17491_), .A3(new_n10045_), .ZN(new_n17492_));
  NAND2_X1   g17300(.A1(new_n17492_), .A2(new_n17370_), .ZN(new_n17493_));
  NAND2_X1   g17301(.A1(new_n17489_), .A2(new_n17491_), .ZN(new_n17494_));
  AOI21_X1   g17302(.A1(new_n17494_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n17495_));
  AOI21_X1   g17303(.A1(new_n17495_), .A2(new_n17493_), .B(new_n17367_), .ZN(new_n17496_));
  INV_X1     g17304(.I(new_n17372_), .ZN(new_n17497_));
  INV_X1     g17305(.I(new_n17382_), .ZN(new_n17498_));
  NOR2_X1    g17306(.A1(new_n17481_), .A2(new_n17482_), .ZN(new_n17499_));
  AOI21_X1   g17307(.A1(new_n17499_), .A2(new_n11901_), .B(new_n17498_), .ZN(new_n17500_));
  NAND2_X1   g17308(.A1(new_n17483_), .A2(new_n11406_), .ZN(new_n17501_));
  OAI21_X1   g17309(.A1(new_n17500_), .A2(new_n17501_), .B(new_n17378_), .ZN(new_n17502_));
  INV_X1     g17310(.I(new_n17483_), .ZN(new_n17503_));
  OAI21_X1   g17311(.A1(new_n17500_), .A2(new_n17503_), .B(\asqrt[17] ), .ZN(new_n17504_));
  NAND3_X1   g17312(.A1(new_n17502_), .A2(new_n17504_), .A3(new_n10953_), .ZN(new_n17505_));
  NAND2_X1   g17313(.A1(new_n17505_), .A2(new_n17375_), .ZN(new_n17506_));
  NAND2_X1   g17314(.A1(new_n17502_), .A2(new_n17504_), .ZN(new_n17507_));
  AOI21_X1   g17315(.A1(new_n17507_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n17508_));
  AOI21_X1   g17316(.A1(new_n17508_), .A2(new_n17506_), .B(new_n17497_), .ZN(new_n17509_));
  AOI21_X1   g17317(.A1(new_n17506_), .A2(new_n17487_), .B(new_n10478_), .ZN(new_n17510_));
  OAI21_X1   g17318(.A1(new_n17509_), .A2(new_n17510_), .B(\asqrt[20] ), .ZN(new_n17511_));
  AOI21_X1   g17319(.A1(new_n17493_), .A2(new_n17511_), .B(new_n9590_), .ZN(new_n17512_));
  NOR2_X1    g17320(.A1(new_n17496_), .A2(new_n17512_), .ZN(new_n17513_));
  AOI21_X1   g17321(.A1(new_n17513_), .A2(new_n9177_), .B(new_n17364_), .ZN(new_n17514_));
  OAI21_X1   g17322(.A1(new_n17496_), .A2(new_n17512_), .B(\asqrt[22] ), .ZN(new_n17515_));
  NAND2_X1   g17323(.A1(new_n17515_), .A2(new_n8742_), .ZN(new_n17516_));
  OAI21_X1   g17324(.A1(new_n17514_), .A2(new_n17516_), .B(new_n17360_), .ZN(new_n17517_));
  INV_X1     g17325(.I(new_n17515_), .ZN(new_n17518_));
  OAI21_X1   g17326(.A1(new_n17514_), .A2(new_n17518_), .B(\asqrt[23] ), .ZN(new_n17519_));
  NAND3_X1   g17327(.A1(new_n17517_), .A2(new_n17519_), .A3(new_n8349_), .ZN(new_n17520_));
  NAND2_X1   g17328(.A1(new_n17520_), .A2(new_n17358_), .ZN(new_n17521_));
  NAND2_X1   g17329(.A1(new_n17517_), .A2(new_n17519_), .ZN(new_n17522_));
  AOI21_X1   g17330(.A1(new_n17522_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n17523_));
  AOI21_X1   g17331(.A1(new_n17523_), .A2(new_n17521_), .B(new_n17355_), .ZN(new_n17524_));
  INV_X1     g17332(.I(new_n17360_), .ZN(new_n17525_));
  INV_X1     g17333(.I(new_n17370_), .ZN(new_n17526_));
  NOR2_X1    g17334(.A1(new_n17509_), .A2(new_n17510_), .ZN(new_n17527_));
  AOI21_X1   g17335(.A1(new_n17527_), .A2(new_n10045_), .B(new_n17526_), .ZN(new_n17528_));
  NAND2_X1   g17336(.A1(new_n17511_), .A2(new_n9590_), .ZN(new_n17529_));
  OAI21_X1   g17337(.A1(new_n17528_), .A2(new_n17529_), .B(new_n17366_), .ZN(new_n17530_));
  INV_X1     g17338(.I(new_n17511_), .ZN(new_n17531_));
  OAI21_X1   g17339(.A1(new_n17528_), .A2(new_n17531_), .B(\asqrt[21] ), .ZN(new_n17532_));
  NAND3_X1   g17340(.A1(new_n17530_), .A2(new_n17532_), .A3(new_n9177_), .ZN(new_n17533_));
  NAND2_X1   g17341(.A1(new_n17533_), .A2(new_n17363_), .ZN(new_n17534_));
  NAND2_X1   g17342(.A1(new_n17530_), .A2(new_n17532_), .ZN(new_n17535_));
  AOI21_X1   g17343(.A1(new_n17535_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n17536_));
  AOI21_X1   g17344(.A1(new_n17536_), .A2(new_n17534_), .B(new_n17525_), .ZN(new_n17537_));
  AOI21_X1   g17345(.A1(new_n17534_), .A2(new_n17515_), .B(new_n8742_), .ZN(new_n17538_));
  OAI21_X1   g17346(.A1(new_n17537_), .A2(new_n17538_), .B(\asqrt[24] ), .ZN(new_n17539_));
  AOI21_X1   g17347(.A1(new_n17521_), .A2(new_n17539_), .B(new_n7934_), .ZN(new_n17540_));
  NOR2_X1    g17348(.A1(new_n17524_), .A2(new_n17540_), .ZN(new_n17541_));
  AOI21_X1   g17349(.A1(new_n17541_), .A2(new_n7561_), .B(new_n17352_), .ZN(new_n17542_));
  OAI21_X1   g17350(.A1(new_n17524_), .A2(new_n17540_), .B(\asqrt[26] ), .ZN(new_n17543_));
  NAND2_X1   g17351(.A1(new_n17543_), .A2(new_n7166_), .ZN(new_n17544_));
  OAI21_X1   g17352(.A1(new_n17542_), .A2(new_n17544_), .B(new_n17348_), .ZN(new_n17545_));
  INV_X1     g17353(.I(new_n17543_), .ZN(new_n17546_));
  OAI21_X1   g17354(.A1(new_n17542_), .A2(new_n17546_), .B(\asqrt[27] ), .ZN(new_n17547_));
  NAND3_X1   g17355(.A1(new_n17545_), .A2(new_n17547_), .A3(new_n6813_), .ZN(new_n17548_));
  NAND2_X1   g17356(.A1(new_n17548_), .A2(new_n17346_), .ZN(new_n17549_));
  NAND2_X1   g17357(.A1(new_n17545_), .A2(new_n17547_), .ZN(new_n17550_));
  AOI21_X1   g17358(.A1(new_n17550_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n17551_));
  AOI21_X1   g17359(.A1(new_n17551_), .A2(new_n17549_), .B(new_n17343_), .ZN(new_n17552_));
  INV_X1     g17360(.I(new_n17348_), .ZN(new_n17553_));
  INV_X1     g17361(.I(new_n17358_), .ZN(new_n17554_));
  NOR2_X1    g17362(.A1(new_n17537_), .A2(new_n17538_), .ZN(new_n17555_));
  AOI21_X1   g17363(.A1(new_n17555_), .A2(new_n8349_), .B(new_n17554_), .ZN(new_n17556_));
  NAND2_X1   g17364(.A1(new_n17539_), .A2(new_n7934_), .ZN(new_n17557_));
  OAI21_X1   g17365(.A1(new_n17556_), .A2(new_n17557_), .B(new_n17354_), .ZN(new_n17558_));
  INV_X1     g17366(.I(new_n17539_), .ZN(new_n17559_));
  OAI21_X1   g17367(.A1(new_n17556_), .A2(new_n17559_), .B(\asqrt[25] ), .ZN(new_n17560_));
  NAND3_X1   g17368(.A1(new_n17558_), .A2(new_n17560_), .A3(new_n7561_), .ZN(new_n17561_));
  NAND2_X1   g17369(.A1(new_n17561_), .A2(new_n17351_), .ZN(new_n17562_));
  NAND2_X1   g17370(.A1(new_n17558_), .A2(new_n17560_), .ZN(new_n17563_));
  AOI21_X1   g17371(.A1(new_n17563_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n17564_));
  AOI21_X1   g17372(.A1(new_n17564_), .A2(new_n17562_), .B(new_n17553_), .ZN(new_n17565_));
  AOI21_X1   g17373(.A1(new_n17562_), .A2(new_n17543_), .B(new_n7166_), .ZN(new_n17566_));
  OAI21_X1   g17374(.A1(new_n17565_), .A2(new_n17566_), .B(\asqrt[28] ), .ZN(new_n17567_));
  AOI21_X1   g17375(.A1(new_n17549_), .A2(new_n17567_), .B(new_n6454_), .ZN(new_n17568_));
  NOR2_X1    g17376(.A1(new_n17552_), .A2(new_n17568_), .ZN(new_n17569_));
  AOI21_X1   g17377(.A1(new_n17569_), .A2(new_n6106_), .B(new_n17340_), .ZN(new_n17570_));
  OAI21_X1   g17378(.A1(new_n17552_), .A2(new_n17568_), .B(\asqrt[30] ), .ZN(new_n17571_));
  NAND2_X1   g17379(.A1(new_n17571_), .A2(new_n5750_), .ZN(new_n17572_));
  OAI21_X1   g17380(.A1(new_n17570_), .A2(new_n17572_), .B(new_n17336_), .ZN(new_n17573_));
  INV_X1     g17381(.I(new_n17571_), .ZN(new_n17574_));
  OAI21_X1   g17382(.A1(new_n17570_), .A2(new_n17574_), .B(\asqrt[31] ), .ZN(new_n17575_));
  NAND3_X1   g17383(.A1(new_n17573_), .A2(new_n17575_), .A3(new_n5435_), .ZN(new_n17576_));
  NAND2_X1   g17384(.A1(new_n17576_), .A2(new_n17334_), .ZN(new_n17577_));
  NAND2_X1   g17385(.A1(new_n17573_), .A2(new_n17575_), .ZN(new_n17578_));
  AOI21_X1   g17386(.A1(new_n17578_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n17579_));
  AOI21_X1   g17387(.A1(new_n17579_), .A2(new_n17577_), .B(new_n17331_), .ZN(new_n17580_));
  INV_X1     g17388(.I(new_n17336_), .ZN(new_n17581_));
  INV_X1     g17389(.I(new_n17346_), .ZN(new_n17582_));
  NOR2_X1    g17390(.A1(new_n17565_), .A2(new_n17566_), .ZN(new_n17583_));
  AOI21_X1   g17391(.A1(new_n17583_), .A2(new_n6813_), .B(new_n17582_), .ZN(new_n17584_));
  NAND2_X1   g17392(.A1(new_n17567_), .A2(new_n6454_), .ZN(new_n17585_));
  OAI21_X1   g17393(.A1(new_n17584_), .A2(new_n17585_), .B(new_n17342_), .ZN(new_n17586_));
  INV_X1     g17394(.I(new_n17567_), .ZN(new_n17587_));
  OAI21_X1   g17395(.A1(new_n17584_), .A2(new_n17587_), .B(\asqrt[29] ), .ZN(new_n17588_));
  NAND3_X1   g17396(.A1(new_n17586_), .A2(new_n17588_), .A3(new_n6106_), .ZN(new_n17589_));
  NAND2_X1   g17397(.A1(new_n17589_), .A2(new_n17339_), .ZN(new_n17590_));
  NAND2_X1   g17398(.A1(new_n17586_), .A2(new_n17588_), .ZN(new_n17591_));
  AOI21_X1   g17399(.A1(new_n17591_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n17592_));
  AOI21_X1   g17400(.A1(new_n17592_), .A2(new_n17590_), .B(new_n17581_), .ZN(new_n17593_));
  AOI21_X1   g17401(.A1(new_n17590_), .A2(new_n17571_), .B(new_n5750_), .ZN(new_n17594_));
  OAI21_X1   g17402(.A1(new_n17593_), .A2(new_n17594_), .B(\asqrt[32] ), .ZN(new_n17595_));
  AOI21_X1   g17403(.A1(new_n17577_), .A2(new_n17595_), .B(new_n5110_), .ZN(new_n17596_));
  NOR2_X1    g17404(.A1(new_n17580_), .A2(new_n17596_), .ZN(new_n17597_));
  AOI21_X1   g17405(.A1(new_n17597_), .A2(new_n4810_), .B(new_n17328_), .ZN(new_n17598_));
  OAI21_X1   g17406(.A1(new_n17580_), .A2(new_n17596_), .B(\asqrt[34] ), .ZN(new_n17599_));
  NAND2_X1   g17407(.A1(new_n17599_), .A2(new_n4510_), .ZN(new_n17600_));
  OAI21_X1   g17408(.A1(new_n17598_), .A2(new_n17600_), .B(new_n17324_), .ZN(new_n17601_));
  INV_X1     g17409(.I(new_n17599_), .ZN(new_n17602_));
  OAI21_X1   g17410(.A1(new_n17598_), .A2(new_n17602_), .B(\asqrt[35] ), .ZN(new_n17603_));
  NAND3_X1   g17411(.A1(new_n17601_), .A2(new_n17603_), .A3(new_n4224_), .ZN(new_n17604_));
  NAND2_X1   g17412(.A1(new_n17604_), .A2(new_n17322_), .ZN(new_n17605_));
  NAND2_X1   g17413(.A1(new_n17601_), .A2(new_n17603_), .ZN(new_n17606_));
  AOI21_X1   g17414(.A1(new_n17606_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n17607_));
  AOI21_X1   g17415(.A1(new_n17607_), .A2(new_n17605_), .B(new_n17319_), .ZN(new_n17608_));
  INV_X1     g17416(.I(new_n17324_), .ZN(new_n17609_));
  INV_X1     g17417(.I(new_n17334_), .ZN(new_n17610_));
  NOR2_X1    g17418(.A1(new_n17593_), .A2(new_n17594_), .ZN(new_n17611_));
  AOI21_X1   g17419(.A1(new_n17611_), .A2(new_n5435_), .B(new_n17610_), .ZN(new_n17612_));
  NAND2_X1   g17420(.A1(new_n17595_), .A2(new_n5110_), .ZN(new_n17613_));
  OAI21_X1   g17421(.A1(new_n17612_), .A2(new_n17613_), .B(new_n17330_), .ZN(new_n17614_));
  INV_X1     g17422(.I(new_n17595_), .ZN(new_n17615_));
  OAI21_X1   g17423(.A1(new_n17612_), .A2(new_n17615_), .B(\asqrt[33] ), .ZN(new_n17616_));
  NAND3_X1   g17424(.A1(new_n17614_), .A2(new_n17616_), .A3(new_n4810_), .ZN(new_n17617_));
  NAND2_X1   g17425(.A1(new_n17617_), .A2(new_n17327_), .ZN(new_n17618_));
  NAND2_X1   g17426(.A1(new_n17614_), .A2(new_n17616_), .ZN(new_n17619_));
  AOI21_X1   g17427(.A1(new_n17619_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n17620_));
  AOI21_X1   g17428(.A1(new_n17620_), .A2(new_n17618_), .B(new_n17609_), .ZN(new_n17621_));
  AOI21_X1   g17429(.A1(new_n17618_), .A2(new_n17599_), .B(new_n4510_), .ZN(new_n17622_));
  OAI21_X1   g17430(.A1(new_n17621_), .A2(new_n17622_), .B(\asqrt[36] ), .ZN(new_n17623_));
  AOI21_X1   g17431(.A1(new_n17605_), .A2(new_n17623_), .B(new_n3928_), .ZN(new_n17624_));
  NOR2_X1    g17432(.A1(new_n17608_), .A2(new_n17624_), .ZN(new_n17625_));
  AOI21_X1   g17433(.A1(new_n17625_), .A2(new_n3675_), .B(new_n17316_), .ZN(new_n17626_));
  OAI21_X1   g17434(.A1(new_n17608_), .A2(new_n17624_), .B(\asqrt[38] ), .ZN(new_n17627_));
  NAND2_X1   g17435(.A1(new_n17627_), .A2(new_n3400_), .ZN(new_n17628_));
  OAI21_X1   g17436(.A1(new_n17626_), .A2(new_n17628_), .B(new_n17312_), .ZN(new_n17629_));
  INV_X1     g17437(.I(new_n17627_), .ZN(new_n17630_));
  OAI21_X1   g17438(.A1(new_n17626_), .A2(new_n17630_), .B(\asqrt[39] ), .ZN(new_n17631_));
  NAND3_X1   g17439(.A1(new_n17629_), .A2(new_n17631_), .A3(new_n3167_), .ZN(new_n17632_));
  NAND2_X1   g17440(.A1(new_n17632_), .A2(new_n17310_), .ZN(new_n17633_));
  NAND2_X1   g17441(.A1(new_n17629_), .A2(new_n17631_), .ZN(new_n17634_));
  AOI21_X1   g17442(.A1(new_n17634_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n17635_));
  AOI21_X1   g17443(.A1(new_n17635_), .A2(new_n17633_), .B(new_n17307_), .ZN(new_n17636_));
  INV_X1     g17444(.I(new_n17312_), .ZN(new_n17637_));
  INV_X1     g17445(.I(new_n17322_), .ZN(new_n17638_));
  NOR2_X1    g17446(.A1(new_n17621_), .A2(new_n17622_), .ZN(new_n17639_));
  AOI21_X1   g17447(.A1(new_n17639_), .A2(new_n4224_), .B(new_n17638_), .ZN(new_n17640_));
  NAND2_X1   g17448(.A1(new_n17623_), .A2(new_n3928_), .ZN(new_n17641_));
  OAI21_X1   g17449(.A1(new_n17640_), .A2(new_n17641_), .B(new_n17318_), .ZN(new_n17642_));
  INV_X1     g17450(.I(new_n17623_), .ZN(new_n17643_));
  OAI21_X1   g17451(.A1(new_n17640_), .A2(new_n17643_), .B(\asqrt[37] ), .ZN(new_n17644_));
  NAND3_X1   g17452(.A1(new_n17642_), .A2(new_n17644_), .A3(new_n3675_), .ZN(new_n17645_));
  NAND2_X1   g17453(.A1(new_n17645_), .A2(new_n17315_), .ZN(new_n17646_));
  NAND2_X1   g17454(.A1(new_n17642_), .A2(new_n17644_), .ZN(new_n17647_));
  AOI21_X1   g17455(.A1(new_n17647_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n17648_));
  AOI21_X1   g17456(.A1(new_n17648_), .A2(new_n17646_), .B(new_n17637_), .ZN(new_n17649_));
  AOI21_X1   g17457(.A1(new_n17646_), .A2(new_n17627_), .B(new_n3400_), .ZN(new_n17650_));
  OAI21_X1   g17458(.A1(new_n17649_), .A2(new_n17650_), .B(\asqrt[40] ), .ZN(new_n17651_));
  AOI21_X1   g17459(.A1(new_n17633_), .A2(new_n17651_), .B(new_n2912_), .ZN(new_n17652_));
  NOR2_X1    g17460(.A1(new_n17636_), .A2(new_n17652_), .ZN(new_n17653_));
  AOI21_X1   g17461(.A1(new_n17653_), .A2(new_n2699_), .B(new_n17304_), .ZN(new_n17654_));
  OAI21_X1   g17462(.A1(new_n17636_), .A2(new_n17652_), .B(\asqrt[42] ), .ZN(new_n17655_));
  NAND2_X1   g17463(.A1(new_n17655_), .A2(new_n2464_), .ZN(new_n17656_));
  OAI21_X1   g17464(.A1(new_n17654_), .A2(new_n17656_), .B(new_n17300_), .ZN(new_n17657_));
  INV_X1     g17465(.I(new_n17655_), .ZN(new_n17658_));
  OAI21_X1   g17466(.A1(new_n17654_), .A2(new_n17658_), .B(\asqrt[43] ), .ZN(new_n17659_));
  NAND3_X1   g17467(.A1(new_n17657_), .A2(new_n17659_), .A3(new_n2271_), .ZN(new_n17660_));
  NAND2_X1   g17468(.A1(new_n17660_), .A2(new_n17298_), .ZN(new_n17661_));
  NAND2_X1   g17469(.A1(new_n17657_), .A2(new_n17659_), .ZN(new_n17662_));
  AOI21_X1   g17470(.A1(new_n17662_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n17663_));
  AOI21_X1   g17471(.A1(new_n17663_), .A2(new_n17661_), .B(new_n17295_), .ZN(new_n17664_));
  INV_X1     g17472(.I(new_n17300_), .ZN(new_n17665_));
  INV_X1     g17473(.I(new_n17310_), .ZN(new_n17666_));
  NOR2_X1    g17474(.A1(new_n17649_), .A2(new_n17650_), .ZN(new_n17667_));
  AOI21_X1   g17475(.A1(new_n17667_), .A2(new_n3167_), .B(new_n17666_), .ZN(new_n17668_));
  NAND2_X1   g17476(.A1(new_n17651_), .A2(new_n2912_), .ZN(new_n17669_));
  OAI21_X1   g17477(.A1(new_n17668_), .A2(new_n17669_), .B(new_n17306_), .ZN(new_n17670_));
  INV_X1     g17478(.I(new_n17651_), .ZN(new_n17671_));
  OAI21_X1   g17479(.A1(new_n17668_), .A2(new_n17671_), .B(\asqrt[41] ), .ZN(new_n17672_));
  NAND3_X1   g17480(.A1(new_n17670_), .A2(new_n17672_), .A3(new_n2699_), .ZN(new_n17673_));
  NAND2_X1   g17481(.A1(new_n17673_), .A2(new_n17303_), .ZN(new_n17674_));
  NAND2_X1   g17482(.A1(new_n17670_), .A2(new_n17672_), .ZN(new_n17675_));
  AOI21_X1   g17483(.A1(new_n17675_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n17676_));
  AOI21_X1   g17484(.A1(new_n17676_), .A2(new_n17674_), .B(new_n17665_), .ZN(new_n17677_));
  AOI21_X1   g17485(.A1(new_n17674_), .A2(new_n17655_), .B(new_n2464_), .ZN(new_n17678_));
  OAI21_X1   g17486(.A1(new_n17677_), .A2(new_n17678_), .B(\asqrt[44] ), .ZN(new_n17679_));
  AOI21_X1   g17487(.A1(new_n17661_), .A2(new_n17679_), .B(new_n2072_), .ZN(new_n17680_));
  NOR2_X1    g17488(.A1(new_n17664_), .A2(new_n17680_), .ZN(new_n17681_));
  AOI21_X1   g17489(.A1(new_n17681_), .A2(new_n1884_), .B(new_n17292_), .ZN(new_n17682_));
  OAI21_X1   g17490(.A1(new_n17664_), .A2(new_n17680_), .B(\asqrt[46] ), .ZN(new_n17683_));
  NAND2_X1   g17491(.A1(new_n17683_), .A2(new_n1688_), .ZN(new_n17684_));
  OAI21_X1   g17492(.A1(new_n17682_), .A2(new_n17684_), .B(new_n17288_), .ZN(new_n17685_));
  INV_X1     g17493(.I(new_n17683_), .ZN(new_n17686_));
  OAI21_X1   g17494(.A1(new_n17682_), .A2(new_n17686_), .B(\asqrt[47] ), .ZN(new_n17687_));
  NAND3_X1   g17495(.A1(new_n17685_), .A2(new_n17687_), .A3(new_n1533_), .ZN(new_n17688_));
  NAND2_X1   g17496(.A1(new_n17688_), .A2(new_n17286_), .ZN(new_n17689_));
  NAND2_X1   g17497(.A1(new_n17685_), .A2(new_n17687_), .ZN(new_n17690_));
  AOI21_X1   g17498(.A1(new_n17690_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n17691_));
  AOI21_X1   g17499(.A1(new_n17691_), .A2(new_n17689_), .B(new_n17283_), .ZN(new_n17692_));
  INV_X1     g17500(.I(new_n17288_), .ZN(new_n17693_));
  INV_X1     g17501(.I(new_n17298_), .ZN(new_n17694_));
  NOR2_X1    g17502(.A1(new_n17677_), .A2(new_n17678_), .ZN(new_n17695_));
  AOI21_X1   g17503(.A1(new_n17695_), .A2(new_n2271_), .B(new_n17694_), .ZN(new_n17696_));
  NAND2_X1   g17504(.A1(new_n17679_), .A2(new_n2072_), .ZN(new_n17697_));
  OAI21_X1   g17505(.A1(new_n17696_), .A2(new_n17697_), .B(new_n17294_), .ZN(new_n17698_));
  INV_X1     g17506(.I(new_n17679_), .ZN(new_n17699_));
  OAI21_X1   g17507(.A1(new_n17696_), .A2(new_n17699_), .B(\asqrt[45] ), .ZN(new_n17700_));
  NAND3_X1   g17508(.A1(new_n17698_), .A2(new_n17700_), .A3(new_n1884_), .ZN(new_n17701_));
  NAND2_X1   g17509(.A1(new_n17701_), .A2(new_n17291_), .ZN(new_n17702_));
  NAND2_X1   g17510(.A1(new_n17698_), .A2(new_n17700_), .ZN(new_n17703_));
  AOI21_X1   g17511(.A1(new_n17703_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n17704_));
  AOI21_X1   g17512(.A1(new_n17704_), .A2(new_n17702_), .B(new_n17693_), .ZN(new_n17705_));
  AOI21_X1   g17513(.A1(new_n17702_), .A2(new_n17683_), .B(new_n1688_), .ZN(new_n17706_));
  OAI21_X1   g17514(.A1(new_n17705_), .A2(new_n17706_), .B(\asqrt[48] ), .ZN(new_n17707_));
  AOI21_X1   g17515(.A1(new_n17689_), .A2(new_n17707_), .B(new_n1368_), .ZN(new_n17708_));
  NOR2_X1    g17516(.A1(new_n17692_), .A2(new_n17708_), .ZN(new_n17709_));
  AOI21_X1   g17517(.A1(new_n17709_), .A2(new_n1228_), .B(new_n17280_), .ZN(new_n17710_));
  OAI21_X1   g17518(.A1(new_n17692_), .A2(new_n17708_), .B(\asqrt[50] ), .ZN(new_n17711_));
  NAND2_X1   g17519(.A1(new_n17711_), .A2(new_n1088_), .ZN(new_n17712_));
  OAI21_X1   g17520(.A1(new_n17710_), .A2(new_n17712_), .B(new_n17276_), .ZN(new_n17713_));
  INV_X1     g17521(.I(new_n17711_), .ZN(new_n17714_));
  OAI21_X1   g17522(.A1(new_n17710_), .A2(new_n17714_), .B(\asqrt[51] ), .ZN(new_n17715_));
  NAND3_X1   g17523(.A1(new_n17713_), .A2(new_n17715_), .A3(new_n962_), .ZN(new_n17716_));
  NAND2_X1   g17524(.A1(new_n17716_), .A2(new_n17274_), .ZN(new_n17717_));
  NAND2_X1   g17525(.A1(new_n17713_), .A2(new_n17715_), .ZN(new_n17718_));
  AOI21_X1   g17526(.A1(new_n17718_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n17719_));
  AOI21_X1   g17527(.A1(new_n17719_), .A2(new_n17717_), .B(new_n17271_), .ZN(new_n17720_));
  INV_X1     g17528(.I(new_n17276_), .ZN(new_n17721_));
  INV_X1     g17529(.I(new_n17286_), .ZN(new_n17722_));
  NOR2_X1    g17530(.A1(new_n17705_), .A2(new_n17706_), .ZN(new_n17723_));
  AOI21_X1   g17531(.A1(new_n17723_), .A2(new_n1533_), .B(new_n17722_), .ZN(new_n17724_));
  NAND2_X1   g17532(.A1(new_n17707_), .A2(new_n1368_), .ZN(new_n17725_));
  OAI21_X1   g17533(.A1(new_n17724_), .A2(new_n17725_), .B(new_n17282_), .ZN(new_n17726_));
  INV_X1     g17534(.I(new_n17707_), .ZN(new_n17727_));
  OAI21_X1   g17535(.A1(new_n17724_), .A2(new_n17727_), .B(\asqrt[49] ), .ZN(new_n17728_));
  NAND3_X1   g17536(.A1(new_n17726_), .A2(new_n17728_), .A3(new_n1228_), .ZN(new_n17729_));
  NAND2_X1   g17537(.A1(new_n17729_), .A2(new_n17279_), .ZN(new_n17730_));
  NAND2_X1   g17538(.A1(new_n17726_), .A2(new_n17728_), .ZN(new_n17731_));
  AOI21_X1   g17539(.A1(new_n17731_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n17732_));
  AOI21_X1   g17540(.A1(new_n17732_), .A2(new_n17730_), .B(new_n17721_), .ZN(new_n17733_));
  AOI21_X1   g17541(.A1(new_n17730_), .A2(new_n17711_), .B(new_n1088_), .ZN(new_n17734_));
  OAI21_X1   g17542(.A1(new_n17733_), .A2(new_n17734_), .B(\asqrt[52] ), .ZN(new_n17735_));
  AOI21_X1   g17543(.A1(new_n17717_), .A2(new_n17735_), .B(new_n842_), .ZN(new_n17736_));
  NOR2_X1    g17544(.A1(new_n17720_), .A2(new_n17736_), .ZN(new_n17737_));
  AOI21_X1   g17545(.A1(new_n17737_), .A2(new_n720_), .B(new_n17268_), .ZN(new_n17738_));
  OAI21_X1   g17546(.A1(new_n17720_), .A2(new_n17736_), .B(\asqrt[54] ), .ZN(new_n17739_));
  NAND2_X1   g17547(.A1(new_n17739_), .A2(new_n630_), .ZN(new_n17740_));
  OAI21_X1   g17548(.A1(new_n17738_), .A2(new_n17740_), .B(new_n17264_), .ZN(new_n17741_));
  INV_X1     g17549(.I(new_n17739_), .ZN(new_n17742_));
  OAI21_X1   g17550(.A1(new_n17738_), .A2(new_n17742_), .B(\asqrt[55] ), .ZN(new_n17743_));
  NAND3_X1   g17551(.A1(new_n17741_), .A2(new_n17743_), .A3(new_n545_), .ZN(new_n17744_));
  NAND2_X1   g17552(.A1(new_n17744_), .A2(new_n17262_), .ZN(new_n17745_));
  NAND2_X1   g17553(.A1(new_n17741_), .A2(new_n17743_), .ZN(new_n17746_));
  AOI21_X1   g17554(.A1(new_n17746_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n17747_));
  AOI21_X1   g17555(.A1(new_n17747_), .A2(new_n17745_), .B(new_n17259_), .ZN(new_n17748_));
  INV_X1     g17556(.I(new_n17264_), .ZN(new_n17749_));
  INV_X1     g17557(.I(new_n17274_), .ZN(new_n17750_));
  NOR2_X1    g17558(.A1(new_n17733_), .A2(new_n17734_), .ZN(new_n17751_));
  AOI21_X1   g17559(.A1(new_n17751_), .A2(new_n962_), .B(new_n17750_), .ZN(new_n17752_));
  NAND2_X1   g17560(.A1(new_n17735_), .A2(new_n842_), .ZN(new_n17753_));
  OAI21_X1   g17561(.A1(new_n17752_), .A2(new_n17753_), .B(new_n17270_), .ZN(new_n17754_));
  INV_X1     g17562(.I(new_n17735_), .ZN(new_n17755_));
  OAI21_X1   g17563(.A1(new_n17752_), .A2(new_n17755_), .B(\asqrt[53] ), .ZN(new_n17756_));
  NAND3_X1   g17564(.A1(new_n17754_), .A2(new_n17756_), .A3(new_n720_), .ZN(new_n17757_));
  NAND2_X1   g17565(.A1(new_n17757_), .A2(new_n17267_), .ZN(new_n17758_));
  NAND2_X1   g17566(.A1(new_n17754_), .A2(new_n17756_), .ZN(new_n17759_));
  AOI21_X1   g17567(.A1(new_n17759_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n17760_));
  AOI21_X1   g17568(.A1(new_n17760_), .A2(new_n17758_), .B(new_n17749_), .ZN(new_n17761_));
  AOI21_X1   g17569(.A1(new_n17758_), .A2(new_n17739_), .B(new_n630_), .ZN(new_n17762_));
  OAI21_X1   g17570(.A1(new_n17761_), .A2(new_n17762_), .B(\asqrt[56] ), .ZN(new_n17763_));
  AOI21_X1   g17571(.A1(new_n17745_), .A2(new_n17763_), .B(new_n450_), .ZN(new_n17764_));
  NOR2_X1    g17572(.A1(new_n17748_), .A2(new_n17764_), .ZN(new_n17765_));
  AOI21_X1   g17573(.A1(new_n17765_), .A2(new_n403_), .B(new_n17256_), .ZN(new_n17766_));
  OAI21_X1   g17574(.A1(new_n17748_), .A2(new_n17764_), .B(\asqrt[58] ), .ZN(new_n17767_));
  NAND2_X1   g17575(.A1(new_n17767_), .A2(new_n339_), .ZN(new_n17768_));
  OAI21_X1   g17576(.A1(new_n17766_), .A2(new_n17768_), .B(new_n17227_), .ZN(new_n17769_));
  INV_X1     g17577(.I(new_n17767_), .ZN(new_n17770_));
  OAI21_X1   g17578(.A1(new_n17766_), .A2(new_n17770_), .B(\asqrt[59] ), .ZN(new_n17771_));
  NAND3_X1   g17579(.A1(new_n17769_), .A2(new_n17771_), .A3(new_n288_), .ZN(new_n17772_));
  NAND2_X1   g17580(.A1(new_n17772_), .A2(new_n17252_), .ZN(new_n17773_));
  INV_X1     g17581(.I(new_n17227_), .ZN(new_n17774_));
  INV_X1     g17582(.I(new_n17262_), .ZN(new_n17775_));
  NOR2_X1    g17583(.A1(new_n17761_), .A2(new_n17762_), .ZN(new_n17776_));
  AOI21_X1   g17584(.A1(new_n17776_), .A2(new_n545_), .B(new_n17775_), .ZN(new_n17777_));
  NAND2_X1   g17585(.A1(new_n17763_), .A2(new_n450_), .ZN(new_n17778_));
  OAI21_X1   g17586(.A1(new_n17777_), .A2(new_n17778_), .B(new_n17258_), .ZN(new_n17779_));
  INV_X1     g17587(.I(new_n17763_), .ZN(new_n17780_));
  OAI21_X1   g17588(.A1(new_n17777_), .A2(new_n17780_), .B(\asqrt[57] ), .ZN(new_n17781_));
  NAND3_X1   g17589(.A1(new_n17779_), .A2(new_n17781_), .A3(new_n403_), .ZN(new_n17782_));
  NAND2_X1   g17590(.A1(new_n17782_), .A2(new_n17255_), .ZN(new_n17783_));
  NAND2_X1   g17591(.A1(new_n17779_), .A2(new_n17781_), .ZN(new_n17784_));
  AOI21_X1   g17592(.A1(new_n17784_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n17785_));
  AOI21_X1   g17593(.A1(new_n17785_), .A2(new_n17783_), .B(new_n17774_), .ZN(new_n17786_));
  AOI21_X1   g17594(.A1(new_n17783_), .A2(new_n17767_), .B(new_n339_), .ZN(new_n17787_));
  OAI21_X1   g17595(.A1(new_n17786_), .A2(new_n17787_), .B(\asqrt[60] ), .ZN(new_n17788_));
  AOI21_X1   g17596(.A1(new_n17773_), .A2(new_n17788_), .B(new_n242_), .ZN(new_n17789_));
  NAND3_X1   g17597(.A1(\asqrt[6] ), .A2(new_n17195_), .A3(new_n17203_), .ZN(new_n17790_));
  XOR2_X1    g17598(.A1(new_n17790_), .A2(new_n17231_), .Z(new_n17791_));
  INV_X1     g17599(.I(new_n17791_), .ZN(new_n17792_));
  NAND2_X1   g17600(.A1(new_n17769_), .A2(new_n17771_), .ZN(new_n17793_));
  AOI21_X1   g17601(.A1(new_n17793_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n17794_));
  AOI21_X1   g17602(.A1(new_n17794_), .A2(new_n17773_), .B(new_n17792_), .ZN(new_n17795_));
  OAI21_X1   g17603(.A1(new_n17795_), .A2(new_n17789_), .B(\asqrt[62] ), .ZN(new_n17796_));
  AOI21_X1   g17604(.A1(new_n17196_), .A2(new_n17209_), .B(new_n17204_), .ZN(new_n17797_));
  NAND2_X1   g17605(.A1(\asqrt[6] ), .A2(new_n17797_), .ZN(new_n17798_));
  XOR2_X1    g17606(.A1(new_n17798_), .A2(new_n17207_), .Z(new_n17799_));
  INV_X1     g17607(.I(new_n17252_), .ZN(new_n17800_));
  NOR2_X1    g17608(.A1(new_n17786_), .A2(new_n17787_), .ZN(new_n17801_));
  AOI21_X1   g17609(.A1(new_n17801_), .A2(new_n288_), .B(new_n17800_), .ZN(new_n17802_));
  INV_X1     g17610(.I(new_n17788_), .ZN(new_n17803_));
  OAI21_X1   g17611(.A1(new_n17802_), .A2(new_n17803_), .B(\asqrt[61] ), .ZN(new_n17804_));
  NAND2_X1   g17612(.A1(new_n17788_), .A2(new_n242_), .ZN(new_n17805_));
  OAI21_X1   g17613(.A1(new_n17802_), .A2(new_n17805_), .B(new_n17791_), .ZN(new_n17806_));
  NAND3_X1   g17614(.A1(new_n17806_), .A2(new_n17804_), .A3(new_n234_), .ZN(new_n17807_));
  NAND2_X1   g17615(.A1(new_n17807_), .A2(new_n17799_), .ZN(new_n17808_));
  AOI21_X1   g17616(.A1(new_n17808_), .A2(new_n17796_), .B(new_n17249_), .ZN(new_n17809_));
  AOI21_X1   g17617(.A1(new_n17809_), .A2(new_n17247_), .B(\asqrt[63] ), .ZN(new_n17810_));
  AOI21_X1   g17618(.A1(new_n17806_), .A2(new_n17804_), .B(new_n234_), .ZN(new_n17811_));
  INV_X1     g17619(.I(new_n17799_), .ZN(new_n17812_));
  NOR3_X1    g17620(.A1(new_n17795_), .A2(new_n17789_), .A3(\asqrt[62] ), .ZN(new_n17813_));
  NOR2_X1    g17621(.A1(new_n17813_), .A2(new_n17812_), .ZN(new_n17814_));
  NOR3_X1    g17622(.A1(new_n17814_), .A2(new_n17247_), .A3(new_n17811_), .ZN(new_n17815_));
  NOR3_X1    g17623(.A1(new_n17810_), .A2(new_n17245_), .A3(new_n17815_), .ZN(new_n17816_));
  OAI21_X1   g17624(.A1(new_n17766_), .A2(new_n17768_), .B(new_n17771_), .ZN(new_n17817_));
  NOR2_X1    g17625(.A1(new_n17816_), .A2(new_n17817_), .ZN(new_n17818_));
  XOR2_X1    g17626(.A1(new_n17818_), .A2(new_n17227_), .Z(new_n17819_));
  INV_X1     g17627(.I(new_n17819_), .ZN(new_n17820_));
  INV_X1     g17628(.I(new_n17245_), .ZN(new_n17821_));
  INV_X1     g17629(.I(new_n17247_), .ZN(new_n17822_));
  INV_X1     g17630(.I(new_n17249_), .ZN(new_n17823_));
  OAI21_X1   g17631(.A1(new_n17814_), .A2(new_n17811_), .B(new_n17823_), .ZN(new_n17824_));
  OAI21_X1   g17632(.A1(new_n17824_), .A2(new_n17822_), .B(new_n193_), .ZN(new_n17825_));
  AOI21_X1   g17633(.A1(new_n17799_), .A2(new_n17807_), .B(new_n17811_), .ZN(new_n17826_));
  NAND2_X1   g17634(.A1(new_n17826_), .A2(new_n17822_), .ZN(new_n17827_));
  NAND3_X1   g17635(.A1(new_n17825_), .A2(new_n17821_), .A3(new_n17827_), .ZN(\asqrt[5] ));
  NAND3_X1   g17636(.A1(\asqrt[5] ), .A2(new_n17782_), .A3(new_n17767_), .ZN(new_n17829_));
  XOR2_X1    g17637(.A1(new_n17829_), .A2(new_n17256_), .Z(new_n17830_));
  OAI21_X1   g17638(.A1(new_n17777_), .A2(new_n17778_), .B(new_n17781_), .ZN(new_n17831_));
  NOR2_X1    g17639(.A1(new_n17816_), .A2(new_n17831_), .ZN(new_n17832_));
  XOR2_X1    g17640(.A1(new_n17832_), .A2(new_n17258_), .Z(new_n17833_));
  INV_X1     g17641(.I(new_n17833_), .ZN(new_n17834_));
  NAND3_X1   g17642(.A1(\asqrt[5] ), .A2(new_n17744_), .A3(new_n17763_), .ZN(new_n17835_));
  XOR2_X1    g17643(.A1(new_n17835_), .A2(new_n17775_), .Z(new_n17836_));
  INV_X1     g17644(.I(new_n17836_), .ZN(new_n17837_));
  OAI21_X1   g17645(.A1(new_n17738_), .A2(new_n17740_), .B(new_n17743_), .ZN(new_n17838_));
  NOR2_X1    g17646(.A1(new_n17816_), .A2(new_n17838_), .ZN(new_n17839_));
  XOR2_X1    g17647(.A1(new_n17839_), .A2(new_n17264_), .Z(new_n17840_));
  NAND3_X1   g17648(.A1(\asqrt[5] ), .A2(new_n17757_), .A3(new_n17739_), .ZN(new_n17841_));
  XOR2_X1    g17649(.A1(new_n17841_), .A2(new_n17268_), .Z(new_n17842_));
  OAI21_X1   g17650(.A1(new_n17752_), .A2(new_n17753_), .B(new_n17756_), .ZN(new_n17843_));
  NOR2_X1    g17651(.A1(new_n17816_), .A2(new_n17843_), .ZN(new_n17844_));
  XOR2_X1    g17652(.A1(new_n17844_), .A2(new_n17270_), .Z(new_n17845_));
  INV_X1     g17653(.I(new_n17845_), .ZN(new_n17846_));
  NAND3_X1   g17654(.A1(\asqrt[5] ), .A2(new_n17716_), .A3(new_n17735_), .ZN(new_n17847_));
  XOR2_X1    g17655(.A1(new_n17847_), .A2(new_n17750_), .Z(new_n17848_));
  INV_X1     g17656(.I(new_n17848_), .ZN(new_n17849_));
  OAI21_X1   g17657(.A1(new_n17710_), .A2(new_n17712_), .B(new_n17715_), .ZN(new_n17850_));
  NOR2_X1    g17658(.A1(new_n17816_), .A2(new_n17850_), .ZN(new_n17851_));
  XOR2_X1    g17659(.A1(new_n17851_), .A2(new_n17276_), .Z(new_n17852_));
  NAND3_X1   g17660(.A1(\asqrt[5] ), .A2(new_n17729_), .A3(new_n17711_), .ZN(new_n17853_));
  XOR2_X1    g17661(.A1(new_n17853_), .A2(new_n17280_), .Z(new_n17854_));
  OAI21_X1   g17662(.A1(new_n17724_), .A2(new_n17725_), .B(new_n17728_), .ZN(new_n17855_));
  NOR2_X1    g17663(.A1(new_n17816_), .A2(new_n17855_), .ZN(new_n17856_));
  XOR2_X1    g17664(.A1(new_n17856_), .A2(new_n17282_), .Z(new_n17857_));
  INV_X1     g17665(.I(new_n17857_), .ZN(new_n17858_));
  NAND3_X1   g17666(.A1(\asqrt[5] ), .A2(new_n17688_), .A3(new_n17707_), .ZN(new_n17859_));
  XOR2_X1    g17667(.A1(new_n17859_), .A2(new_n17722_), .Z(new_n17860_));
  INV_X1     g17668(.I(new_n17860_), .ZN(new_n17861_));
  OAI21_X1   g17669(.A1(new_n17682_), .A2(new_n17684_), .B(new_n17687_), .ZN(new_n17862_));
  NOR2_X1    g17670(.A1(new_n17816_), .A2(new_n17862_), .ZN(new_n17863_));
  XOR2_X1    g17671(.A1(new_n17863_), .A2(new_n17288_), .Z(new_n17864_));
  NAND3_X1   g17672(.A1(\asqrt[5] ), .A2(new_n17701_), .A3(new_n17683_), .ZN(new_n17865_));
  XOR2_X1    g17673(.A1(new_n17865_), .A2(new_n17292_), .Z(new_n17866_));
  OAI21_X1   g17674(.A1(new_n17696_), .A2(new_n17697_), .B(new_n17700_), .ZN(new_n17867_));
  NOR2_X1    g17675(.A1(new_n17816_), .A2(new_n17867_), .ZN(new_n17868_));
  XOR2_X1    g17676(.A1(new_n17868_), .A2(new_n17294_), .Z(new_n17869_));
  INV_X1     g17677(.I(new_n17869_), .ZN(new_n17870_));
  NAND3_X1   g17678(.A1(\asqrt[5] ), .A2(new_n17660_), .A3(new_n17679_), .ZN(new_n17871_));
  XOR2_X1    g17679(.A1(new_n17871_), .A2(new_n17694_), .Z(new_n17872_));
  INV_X1     g17680(.I(new_n17872_), .ZN(new_n17873_));
  OAI21_X1   g17681(.A1(new_n17654_), .A2(new_n17656_), .B(new_n17659_), .ZN(new_n17874_));
  NOR2_X1    g17682(.A1(new_n17816_), .A2(new_n17874_), .ZN(new_n17875_));
  XOR2_X1    g17683(.A1(new_n17875_), .A2(new_n17300_), .Z(new_n17876_));
  NAND3_X1   g17684(.A1(\asqrt[5] ), .A2(new_n17673_), .A3(new_n17655_), .ZN(new_n17877_));
  XOR2_X1    g17685(.A1(new_n17877_), .A2(new_n17304_), .Z(new_n17878_));
  OAI21_X1   g17686(.A1(new_n17668_), .A2(new_n17669_), .B(new_n17672_), .ZN(new_n17879_));
  NOR2_X1    g17687(.A1(new_n17816_), .A2(new_n17879_), .ZN(new_n17880_));
  XOR2_X1    g17688(.A1(new_n17880_), .A2(new_n17306_), .Z(new_n17881_));
  INV_X1     g17689(.I(new_n17881_), .ZN(new_n17882_));
  NAND3_X1   g17690(.A1(\asqrt[5] ), .A2(new_n17632_), .A3(new_n17651_), .ZN(new_n17883_));
  XOR2_X1    g17691(.A1(new_n17883_), .A2(new_n17666_), .Z(new_n17884_));
  INV_X1     g17692(.I(new_n17884_), .ZN(new_n17885_));
  OAI21_X1   g17693(.A1(new_n17626_), .A2(new_n17628_), .B(new_n17631_), .ZN(new_n17886_));
  NOR2_X1    g17694(.A1(new_n17816_), .A2(new_n17886_), .ZN(new_n17887_));
  XOR2_X1    g17695(.A1(new_n17887_), .A2(new_n17312_), .Z(new_n17888_));
  NAND3_X1   g17696(.A1(\asqrt[5] ), .A2(new_n17645_), .A3(new_n17627_), .ZN(new_n17889_));
  XOR2_X1    g17697(.A1(new_n17889_), .A2(new_n17316_), .Z(new_n17890_));
  OAI21_X1   g17698(.A1(new_n17640_), .A2(new_n17641_), .B(new_n17644_), .ZN(new_n17891_));
  NOR2_X1    g17699(.A1(new_n17816_), .A2(new_n17891_), .ZN(new_n17892_));
  XOR2_X1    g17700(.A1(new_n17892_), .A2(new_n17318_), .Z(new_n17893_));
  INV_X1     g17701(.I(new_n17893_), .ZN(new_n17894_));
  NAND3_X1   g17702(.A1(\asqrt[5] ), .A2(new_n17604_), .A3(new_n17623_), .ZN(new_n17895_));
  XOR2_X1    g17703(.A1(new_n17895_), .A2(new_n17638_), .Z(new_n17896_));
  INV_X1     g17704(.I(new_n17896_), .ZN(new_n17897_));
  OAI21_X1   g17705(.A1(new_n17598_), .A2(new_n17600_), .B(new_n17603_), .ZN(new_n17898_));
  NOR2_X1    g17706(.A1(new_n17816_), .A2(new_n17898_), .ZN(new_n17899_));
  XOR2_X1    g17707(.A1(new_n17899_), .A2(new_n17324_), .Z(new_n17900_));
  NAND3_X1   g17708(.A1(\asqrt[5] ), .A2(new_n17617_), .A3(new_n17599_), .ZN(new_n17901_));
  XOR2_X1    g17709(.A1(new_n17901_), .A2(new_n17328_), .Z(new_n17902_));
  OAI21_X1   g17710(.A1(new_n17612_), .A2(new_n17613_), .B(new_n17616_), .ZN(new_n17903_));
  NOR2_X1    g17711(.A1(new_n17816_), .A2(new_n17903_), .ZN(new_n17904_));
  XOR2_X1    g17712(.A1(new_n17904_), .A2(new_n17330_), .Z(new_n17905_));
  INV_X1     g17713(.I(new_n17905_), .ZN(new_n17906_));
  NAND3_X1   g17714(.A1(\asqrt[5] ), .A2(new_n17576_), .A3(new_n17595_), .ZN(new_n17907_));
  XOR2_X1    g17715(.A1(new_n17907_), .A2(new_n17610_), .Z(new_n17908_));
  INV_X1     g17716(.I(new_n17908_), .ZN(new_n17909_));
  OAI21_X1   g17717(.A1(new_n17570_), .A2(new_n17572_), .B(new_n17575_), .ZN(new_n17910_));
  NOR2_X1    g17718(.A1(new_n17816_), .A2(new_n17910_), .ZN(new_n17911_));
  XOR2_X1    g17719(.A1(new_n17911_), .A2(new_n17336_), .Z(new_n17912_));
  NAND3_X1   g17720(.A1(\asqrt[5] ), .A2(new_n17589_), .A3(new_n17571_), .ZN(new_n17913_));
  XOR2_X1    g17721(.A1(new_n17913_), .A2(new_n17340_), .Z(new_n17914_));
  OAI21_X1   g17722(.A1(new_n17584_), .A2(new_n17585_), .B(new_n17588_), .ZN(new_n17915_));
  NOR2_X1    g17723(.A1(new_n17816_), .A2(new_n17915_), .ZN(new_n17916_));
  XOR2_X1    g17724(.A1(new_n17916_), .A2(new_n17342_), .Z(new_n17917_));
  INV_X1     g17725(.I(new_n17917_), .ZN(new_n17918_));
  NAND3_X1   g17726(.A1(\asqrt[5] ), .A2(new_n17548_), .A3(new_n17567_), .ZN(new_n17919_));
  XOR2_X1    g17727(.A1(new_n17919_), .A2(new_n17582_), .Z(new_n17920_));
  INV_X1     g17728(.I(new_n17920_), .ZN(new_n17921_));
  OAI21_X1   g17729(.A1(new_n17542_), .A2(new_n17544_), .B(new_n17547_), .ZN(new_n17922_));
  NOR2_X1    g17730(.A1(new_n17816_), .A2(new_n17922_), .ZN(new_n17923_));
  XOR2_X1    g17731(.A1(new_n17923_), .A2(new_n17348_), .Z(new_n17924_));
  NAND3_X1   g17732(.A1(\asqrt[5] ), .A2(new_n17561_), .A3(new_n17543_), .ZN(new_n17925_));
  XOR2_X1    g17733(.A1(new_n17925_), .A2(new_n17352_), .Z(new_n17926_));
  OAI21_X1   g17734(.A1(new_n17556_), .A2(new_n17557_), .B(new_n17560_), .ZN(new_n17927_));
  NOR2_X1    g17735(.A1(new_n17816_), .A2(new_n17927_), .ZN(new_n17928_));
  XOR2_X1    g17736(.A1(new_n17928_), .A2(new_n17354_), .Z(new_n17929_));
  INV_X1     g17737(.I(new_n17929_), .ZN(new_n17930_));
  NAND3_X1   g17738(.A1(\asqrt[5] ), .A2(new_n17520_), .A3(new_n17539_), .ZN(new_n17931_));
  XOR2_X1    g17739(.A1(new_n17931_), .A2(new_n17554_), .Z(new_n17932_));
  INV_X1     g17740(.I(new_n17932_), .ZN(new_n17933_));
  AOI21_X1   g17741(.A1(new_n17534_), .A2(new_n17536_), .B(new_n17538_), .ZN(new_n17934_));
  NAND2_X1   g17742(.A1(\asqrt[5] ), .A2(new_n17934_), .ZN(new_n17935_));
  XOR2_X1    g17743(.A1(new_n17935_), .A2(new_n17525_), .Z(new_n17936_));
  NAND3_X1   g17744(.A1(\asqrt[5] ), .A2(new_n17533_), .A3(new_n17515_), .ZN(new_n17937_));
  XOR2_X1    g17745(.A1(new_n17937_), .A2(new_n17364_), .Z(new_n17938_));
  OAI21_X1   g17746(.A1(new_n17528_), .A2(new_n17529_), .B(new_n17532_), .ZN(new_n17939_));
  NOR2_X1    g17747(.A1(new_n17816_), .A2(new_n17939_), .ZN(new_n17940_));
  XOR2_X1    g17748(.A1(new_n17940_), .A2(new_n17366_), .Z(new_n17941_));
  INV_X1     g17749(.I(new_n17941_), .ZN(new_n17942_));
  NAND3_X1   g17750(.A1(\asqrt[5] ), .A2(new_n17492_), .A3(new_n17511_), .ZN(new_n17943_));
  XOR2_X1    g17751(.A1(new_n17943_), .A2(new_n17526_), .Z(new_n17944_));
  INV_X1     g17752(.I(new_n17944_), .ZN(new_n17945_));
  AOI21_X1   g17753(.A1(new_n17506_), .A2(new_n17508_), .B(new_n17510_), .ZN(new_n17946_));
  NAND2_X1   g17754(.A1(\asqrt[5] ), .A2(new_n17946_), .ZN(new_n17947_));
  XOR2_X1    g17755(.A1(new_n17947_), .A2(new_n17497_), .Z(new_n17948_));
  NAND3_X1   g17756(.A1(\asqrt[5] ), .A2(new_n17505_), .A3(new_n17487_), .ZN(new_n17949_));
  XOR2_X1    g17757(.A1(new_n17949_), .A2(new_n17376_), .Z(new_n17950_));
  OAI21_X1   g17758(.A1(new_n17500_), .A2(new_n17501_), .B(new_n17504_), .ZN(new_n17951_));
  NOR2_X1    g17759(.A1(new_n17816_), .A2(new_n17951_), .ZN(new_n17952_));
  XOR2_X1    g17760(.A1(new_n17952_), .A2(new_n17378_), .Z(new_n17953_));
  INV_X1     g17761(.I(new_n17953_), .ZN(new_n17954_));
  NAND3_X1   g17762(.A1(\asqrt[5] ), .A2(new_n17464_), .A3(new_n17483_), .ZN(new_n17955_));
  XOR2_X1    g17763(.A1(new_n17955_), .A2(new_n17498_), .Z(new_n17956_));
  INV_X1     g17764(.I(new_n17956_), .ZN(new_n17957_));
  AOI21_X1   g17765(.A1(new_n17478_), .A2(new_n17480_), .B(new_n17482_), .ZN(new_n17958_));
  NAND2_X1   g17766(.A1(\asqrt[5] ), .A2(new_n17958_), .ZN(new_n17959_));
  XOR2_X1    g17767(.A1(new_n17959_), .A2(new_n17469_), .Z(new_n17960_));
  NAND3_X1   g17768(.A1(\asqrt[5] ), .A2(new_n17477_), .A3(new_n17459_), .ZN(new_n17961_));
  XOR2_X1    g17769(.A1(new_n17961_), .A2(new_n17388_), .Z(new_n17962_));
  OAI21_X1   g17770(.A1(new_n17472_), .A2(new_n17473_), .B(new_n17476_), .ZN(new_n17963_));
  NOR2_X1    g17771(.A1(new_n17816_), .A2(new_n17963_), .ZN(new_n17964_));
  XOR2_X1    g17772(.A1(new_n17964_), .A2(new_n17390_), .Z(new_n17965_));
  INV_X1     g17773(.I(new_n17965_), .ZN(new_n17966_));
  NAND3_X1   g17774(.A1(\asqrt[5] ), .A2(new_n17429_), .A3(new_n17455_), .ZN(new_n17967_));
  XOR2_X1    g17775(.A1(new_n17967_), .A2(new_n17470_), .Z(new_n17968_));
  INV_X1     g17776(.I(new_n17968_), .ZN(new_n17969_));
  AOI21_X1   g17777(.A1(new_n17450_), .A2(new_n17451_), .B(new_n17454_), .ZN(new_n17970_));
  NAND2_X1   g17778(.A1(\asqrt[5] ), .A2(new_n17970_), .ZN(new_n17971_));
  XOR2_X1    g17779(.A1(new_n17971_), .A2(new_n17434_), .Z(new_n17972_));
  NOR2_X1    g17780(.A1(new_n17449_), .A2(\asqrt[10] ), .ZN(new_n17973_));
  NOR3_X1    g17781(.A1(new_n17816_), .A2(new_n17973_), .A3(new_n17427_), .ZN(new_n17974_));
  XOR2_X1    g17782(.A1(new_n17974_), .A2(new_n17399_), .Z(new_n17975_));
  NAND3_X1   g17783(.A1(\asqrt[5] ), .A2(new_n17419_), .A3(new_n17448_), .ZN(new_n17976_));
  XOR2_X1    g17784(.A1(new_n17976_), .A2(new_n17447_), .Z(new_n17977_));
  INV_X1     g17785(.I(new_n17977_), .ZN(new_n17978_));
  NAND2_X1   g17786(.A1(new_n17443_), .A2(new_n16093_), .ZN(new_n17979_));
  NAND3_X1   g17787(.A1(\asqrt[5] ), .A2(new_n17979_), .A3(new_n17418_), .ZN(new_n17980_));
  XOR2_X1    g17788(.A1(new_n17980_), .A2(new_n17437_), .Z(new_n17981_));
  INV_X1     g17789(.I(new_n17981_), .ZN(new_n17982_));
  NAND2_X1   g17790(.A1(new_n17816_), .A2(\asqrt[6] ), .ZN(new_n17983_));
  NAND3_X1   g17791(.A1(\asqrt[5] ), .A2(new_n17408_), .A3(new_n17409_), .ZN(new_n17984_));
  AOI21_X1   g17792(.A1(new_n17984_), .A2(new_n17983_), .B(\a[12] ), .ZN(new_n17985_));
  NOR2_X1    g17793(.A1(\asqrt[5] ), .A2(new_n17242_), .ZN(new_n17986_));
  NOR3_X1    g17794(.A1(new_n17816_), .A2(\a[10] ), .A3(\a[11] ), .ZN(new_n17987_));
  NOR3_X1    g17795(.A1(new_n17987_), .A2(new_n17986_), .A3(new_n16809_), .ZN(new_n17988_));
  OR2_X2     g17796(.A1(new_n17988_), .A2(new_n17985_), .Z(new_n17989_));
  NOR3_X1    g17797(.A1(\a[8] ), .A2(\a[9] ), .A3(\a[10] ), .ZN(new_n17990_));
  INV_X1     g17798(.I(new_n17990_), .ZN(new_n17991_));
  NOR3_X1    g17799(.A1(new_n17826_), .A2(new_n17822_), .A3(new_n17249_), .ZN(new_n17992_));
  OAI21_X1   g17800(.A1(new_n17992_), .A2(\asqrt[63] ), .B(new_n17827_), .ZN(new_n17993_));
  OAI21_X1   g17801(.A1(new_n17993_), .A2(new_n17245_), .B(\a[10] ), .ZN(new_n17994_));
  AOI21_X1   g17802(.A1(new_n17994_), .A2(new_n17991_), .B(new_n17242_), .ZN(new_n17995_));
  AOI21_X1   g17803(.A1(\asqrt[5] ), .A2(new_n17408_), .B(new_n17409_), .ZN(new_n17996_));
  OAI21_X1   g17804(.A1(new_n17812_), .A2(new_n17813_), .B(new_n17796_), .ZN(new_n17997_));
  NAND3_X1   g17805(.A1(new_n17997_), .A2(new_n17247_), .A3(new_n17823_), .ZN(new_n17998_));
  AOI21_X1   g17806(.A1(new_n17998_), .A2(new_n193_), .B(new_n17815_), .ZN(new_n17999_));
  AOI21_X1   g17807(.A1(new_n17999_), .A2(new_n17821_), .B(new_n17408_), .ZN(new_n18000_));
  NOR3_X1    g17808(.A1(new_n18000_), .A2(\asqrt[6] ), .A3(new_n17990_), .ZN(new_n18001_));
  NOR3_X1    g17809(.A1(new_n18001_), .A2(new_n17987_), .A3(new_n17996_), .ZN(new_n18002_));
  NOR3_X1    g17810(.A1(new_n18002_), .A2(\asqrt[7] ), .A3(new_n17995_), .ZN(new_n18003_));
  OAI21_X1   g17811(.A1(new_n18002_), .A2(new_n17995_), .B(\asqrt[7] ), .ZN(new_n18004_));
  OAI21_X1   g17812(.A1(new_n17989_), .A2(new_n18003_), .B(new_n18004_), .ZN(new_n18005_));
  NAND3_X1   g17813(.A1(\asqrt[5] ), .A2(new_n17412_), .A3(new_n17442_), .ZN(new_n18006_));
  XOR2_X1    g17814(.A1(new_n18006_), .A2(new_n17414_), .Z(new_n18007_));
  OAI21_X1   g17815(.A1(new_n18005_), .A2(\asqrt[8] ), .B(new_n18007_), .ZN(new_n18008_));
  AOI21_X1   g17816(.A1(new_n18005_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n18009_));
  AOI21_X1   g17817(.A1(new_n18009_), .A2(new_n18008_), .B(new_n17982_), .ZN(new_n18010_));
  NAND2_X1   g17818(.A1(new_n18005_), .A2(\asqrt[8] ), .ZN(new_n18011_));
  AOI21_X1   g17819(.A1(new_n18008_), .A2(new_n18011_), .B(new_n15518_), .ZN(new_n18012_));
  NOR2_X1    g17820(.A1(new_n18010_), .A2(new_n18012_), .ZN(new_n18013_));
  AOI21_X1   g17821(.A1(new_n18013_), .A2(new_n14985_), .B(new_n17978_), .ZN(new_n18014_));
  OAI21_X1   g17822(.A1(new_n18010_), .A2(new_n18012_), .B(\asqrt[10] ), .ZN(new_n18015_));
  NAND2_X1   g17823(.A1(new_n18015_), .A2(new_n14430_), .ZN(new_n18016_));
  OAI21_X1   g17824(.A1(new_n18014_), .A2(new_n18016_), .B(new_n17975_), .ZN(new_n18017_));
  INV_X1     g17825(.I(new_n18015_), .ZN(new_n18018_));
  OAI21_X1   g17826(.A1(new_n18014_), .A2(new_n18018_), .B(\asqrt[11] ), .ZN(new_n18019_));
  NAND3_X1   g17827(.A1(new_n18017_), .A2(new_n18019_), .A3(new_n13917_), .ZN(new_n18020_));
  NAND2_X1   g17828(.A1(new_n18020_), .A2(new_n17972_), .ZN(new_n18021_));
  NAND2_X1   g17829(.A1(new_n18017_), .A2(new_n18019_), .ZN(new_n18022_));
  AOI21_X1   g17830(.A1(new_n18022_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n18023_));
  AOI21_X1   g17831(.A1(new_n18023_), .A2(new_n18021_), .B(new_n17969_), .ZN(new_n18024_));
  INV_X1     g17832(.I(new_n17975_), .ZN(new_n18025_));
  NOR2_X1    g17833(.A1(new_n17988_), .A2(new_n17985_), .ZN(new_n18026_));
  INV_X1     g17834(.I(new_n17995_), .ZN(new_n18027_));
  OAI21_X1   g17835(.A1(new_n17816_), .A2(\a[10] ), .B(\a[11] ), .ZN(new_n18028_));
  NAND3_X1   g17836(.A1(new_n17994_), .A2(new_n17242_), .A3(new_n17991_), .ZN(new_n18029_));
  NAND3_X1   g17837(.A1(new_n18029_), .A2(new_n17984_), .A3(new_n18028_), .ZN(new_n18030_));
  NAND3_X1   g17838(.A1(new_n18030_), .A2(new_n16649_), .A3(new_n18027_), .ZN(new_n18031_));
  AOI21_X1   g17839(.A1(new_n18030_), .A2(new_n18027_), .B(new_n16649_), .ZN(new_n18032_));
  AOI21_X1   g17840(.A1(new_n18026_), .A2(new_n18031_), .B(new_n18032_), .ZN(new_n18033_));
  INV_X1     g17841(.I(new_n18007_), .ZN(new_n18034_));
  AOI21_X1   g17842(.A1(new_n18033_), .A2(new_n16093_), .B(new_n18034_), .ZN(new_n18035_));
  OAI21_X1   g17843(.A1(new_n18033_), .A2(new_n16093_), .B(new_n15518_), .ZN(new_n18036_));
  OAI21_X1   g17844(.A1(new_n18035_), .A2(new_n18036_), .B(new_n17981_), .ZN(new_n18037_));
  NOR2_X1    g17845(.A1(new_n18033_), .A2(new_n16093_), .ZN(new_n18038_));
  OAI21_X1   g17846(.A1(new_n18035_), .A2(new_n18038_), .B(\asqrt[9] ), .ZN(new_n18039_));
  NAND3_X1   g17847(.A1(new_n18037_), .A2(new_n18039_), .A3(new_n14985_), .ZN(new_n18040_));
  NAND2_X1   g17848(.A1(new_n18040_), .A2(new_n17977_), .ZN(new_n18041_));
  NAND2_X1   g17849(.A1(new_n18037_), .A2(new_n18039_), .ZN(new_n18042_));
  AOI21_X1   g17850(.A1(new_n18042_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n18043_));
  AOI21_X1   g17851(.A1(new_n18043_), .A2(new_n18041_), .B(new_n18025_), .ZN(new_n18044_));
  AOI21_X1   g17852(.A1(new_n18041_), .A2(new_n18015_), .B(new_n14430_), .ZN(new_n18045_));
  OAI21_X1   g17853(.A1(new_n18044_), .A2(new_n18045_), .B(\asqrt[12] ), .ZN(new_n18046_));
  AOI21_X1   g17854(.A1(new_n18021_), .A2(new_n18046_), .B(new_n13382_), .ZN(new_n18047_));
  NOR2_X1    g17855(.A1(new_n18024_), .A2(new_n18047_), .ZN(new_n18048_));
  AOI21_X1   g17856(.A1(new_n18048_), .A2(new_n12889_), .B(new_n17966_), .ZN(new_n18049_));
  OAI21_X1   g17857(.A1(new_n18024_), .A2(new_n18047_), .B(\asqrt[14] ), .ZN(new_n18050_));
  NAND2_X1   g17858(.A1(new_n18050_), .A2(new_n12374_), .ZN(new_n18051_));
  OAI21_X1   g17859(.A1(new_n18049_), .A2(new_n18051_), .B(new_n17962_), .ZN(new_n18052_));
  INV_X1     g17860(.I(new_n18050_), .ZN(new_n18053_));
  OAI21_X1   g17861(.A1(new_n18049_), .A2(new_n18053_), .B(\asqrt[15] ), .ZN(new_n18054_));
  NAND3_X1   g17862(.A1(new_n18052_), .A2(new_n18054_), .A3(new_n11901_), .ZN(new_n18055_));
  NAND2_X1   g17863(.A1(new_n18055_), .A2(new_n17960_), .ZN(new_n18056_));
  NAND2_X1   g17864(.A1(new_n18052_), .A2(new_n18054_), .ZN(new_n18057_));
  AOI21_X1   g17865(.A1(new_n18057_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n18058_));
  AOI21_X1   g17866(.A1(new_n18058_), .A2(new_n18056_), .B(new_n17957_), .ZN(new_n18059_));
  INV_X1     g17867(.I(new_n17962_), .ZN(new_n18060_));
  INV_X1     g17868(.I(new_n17972_), .ZN(new_n18061_));
  NOR2_X1    g17869(.A1(new_n18044_), .A2(new_n18045_), .ZN(new_n18062_));
  AOI21_X1   g17870(.A1(new_n18062_), .A2(new_n13917_), .B(new_n18061_), .ZN(new_n18063_));
  NAND2_X1   g17871(.A1(new_n18046_), .A2(new_n13382_), .ZN(new_n18064_));
  OAI21_X1   g17872(.A1(new_n18063_), .A2(new_n18064_), .B(new_n17968_), .ZN(new_n18065_));
  INV_X1     g17873(.I(new_n18046_), .ZN(new_n18066_));
  OAI21_X1   g17874(.A1(new_n18063_), .A2(new_n18066_), .B(\asqrt[13] ), .ZN(new_n18067_));
  NAND3_X1   g17875(.A1(new_n18065_), .A2(new_n18067_), .A3(new_n12889_), .ZN(new_n18068_));
  NAND2_X1   g17876(.A1(new_n18068_), .A2(new_n17965_), .ZN(new_n18069_));
  NAND2_X1   g17877(.A1(new_n18065_), .A2(new_n18067_), .ZN(new_n18070_));
  AOI21_X1   g17878(.A1(new_n18070_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n18071_));
  AOI21_X1   g17879(.A1(new_n18071_), .A2(new_n18069_), .B(new_n18060_), .ZN(new_n18072_));
  AOI21_X1   g17880(.A1(new_n18069_), .A2(new_n18050_), .B(new_n12374_), .ZN(new_n18073_));
  OAI21_X1   g17881(.A1(new_n18072_), .A2(new_n18073_), .B(\asqrt[16] ), .ZN(new_n18074_));
  AOI21_X1   g17882(.A1(new_n18056_), .A2(new_n18074_), .B(new_n11406_), .ZN(new_n18075_));
  NOR2_X1    g17883(.A1(new_n18059_), .A2(new_n18075_), .ZN(new_n18076_));
  AOI21_X1   g17884(.A1(new_n18076_), .A2(new_n10953_), .B(new_n17954_), .ZN(new_n18077_));
  OAI21_X1   g17885(.A1(new_n18059_), .A2(new_n18075_), .B(\asqrt[18] ), .ZN(new_n18078_));
  NAND2_X1   g17886(.A1(new_n18078_), .A2(new_n10478_), .ZN(new_n18079_));
  OAI21_X1   g17887(.A1(new_n18077_), .A2(new_n18079_), .B(new_n17950_), .ZN(new_n18080_));
  INV_X1     g17888(.I(new_n18078_), .ZN(new_n18081_));
  OAI21_X1   g17889(.A1(new_n18077_), .A2(new_n18081_), .B(\asqrt[19] ), .ZN(new_n18082_));
  NAND3_X1   g17890(.A1(new_n18080_), .A2(new_n18082_), .A3(new_n10045_), .ZN(new_n18083_));
  NAND2_X1   g17891(.A1(new_n18083_), .A2(new_n17948_), .ZN(new_n18084_));
  NAND2_X1   g17892(.A1(new_n18080_), .A2(new_n18082_), .ZN(new_n18085_));
  AOI21_X1   g17893(.A1(new_n18085_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n18086_));
  AOI21_X1   g17894(.A1(new_n18086_), .A2(new_n18084_), .B(new_n17945_), .ZN(new_n18087_));
  INV_X1     g17895(.I(new_n17950_), .ZN(new_n18088_));
  INV_X1     g17896(.I(new_n17960_), .ZN(new_n18089_));
  NOR2_X1    g17897(.A1(new_n18072_), .A2(new_n18073_), .ZN(new_n18090_));
  AOI21_X1   g17898(.A1(new_n18090_), .A2(new_n11901_), .B(new_n18089_), .ZN(new_n18091_));
  NAND2_X1   g17899(.A1(new_n18074_), .A2(new_n11406_), .ZN(new_n18092_));
  OAI21_X1   g17900(.A1(new_n18091_), .A2(new_n18092_), .B(new_n17956_), .ZN(new_n18093_));
  INV_X1     g17901(.I(new_n18074_), .ZN(new_n18094_));
  OAI21_X1   g17902(.A1(new_n18091_), .A2(new_n18094_), .B(\asqrt[17] ), .ZN(new_n18095_));
  NAND3_X1   g17903(.A1(new_n18093_), .A2(new_n18095_), .A3(new_n10953_), .ZN(new_n18096_));
  NAND2_X1   g17904(.A1(new_n18096_), .A2(new_n17953_), .ZN(new_n18097_));
  NAND2_X1   g17905(.A1(new_n18093_), .A2(new_n18095_), .ZN(new_n18098_));
  AOI21_X1   g17906(.A1(new_n18098_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n18099_));
  AOI21_X1   g17907(.A1(new_n18099_), .A2(new_n18097_), .B(new_n18088_), .ZN(new_n18100_));
  AOI21_X1   g17908(.A1(new_n18097_), .A2(new_n18078_), .B(new_n10478_), .ZN(new_n18101_));
  OAI21_X1   g17909(.A1(new_n18100_), .A2(new_n18101_), .B(\asqrt[20] ), .ZN(new_n18102_));
  AOI21_X1   g17910(.A1(new_n18084_), .A2(new_n18102_), .B(new_n9590_), .ZN(new_n18103_));
  NOR2_X1    g17911(.A1(new_n18087_), .A2(new_n18103_), .ZN(new_n18104_));
  AOI21_X1   g17912(.A1(new_n18104_), .A2(new_n9177_), .B(new_n17942_), .ZN(new_n18105_));
  OAI21_X1   g17913(.A1(new_n18087_), .A2(new_n18103_), .B(\asqrt[22] ), .ZN(new_n18106_));
  NAND2_X1   g17914(.A1(new_n18106_), .A2(new_n8742_), .ZN(new_n18107_));
  OAI21_X1   g17915(.A1(new_n18105_), .A2(new_n18107_), .B(new_n17938_), .ZN(new_n18108_));
  INV_X1     g17916(.I(new_n18106_), .ZN(new_n18109_));
  OAI21_X1   g17917(.A1(new_n18105_), .A2(new_n18109_), .B(\asqrt[23] ), .ZN(new_n18110_));
  NAND3_X1   g17918(.A1(new_n18108_), .A2(new_n18110_), .A3(new_n8349_), .ZN(new_n18111_));
  NAND2_X1   g17919(.A1(new_n18111_), .A2(new_n17936_), .ZN(new_n18112_));
  NAND2_X1   g17920(.A1(new_n18108_), .A2(new_n18110_), .ZN(new_n18113_));
  AOI21_X1   g17921(.A1(new_n18113_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n18114_));
  AOI21_X1   g17922(.A1(new_n18114_), .A2(new_n18112_), .B(new_n17933_), .ZN(new_n18115_));
  INV_X1     g17923(.I(new_n17938_), .ZN(new_n18116_));
  INV_X1     g17924(.I(new_n17948_), .ZN(new_n18117_));
  NOR2_X1    g17925(.A1(new_n18100_), .A2(new_n18101_), .ZN(new_n18118_));
  AOI21_X1   g17926(.A1(new_n18118_), .A2(new_n10045_), .B(new_n18117_), .ZN(new_n18119_));
  NAND2_X1   g17927(.A1(new_n18102_), .A2(new_n9590_), .ZN(new_n18120_));
  OAI21_X1   g17928(.A1(new_n18119_), .A2(new_n18120_), .B(new_n17944_), .ZN(new_n18121_));
  INV_X1     g17929(.I(new_n18102_), .ZN(new_n18122_));
  OAI21_X1   g17930(.A1(new_n18119_), .A2(new_n18122_), .B(\asqrt[21] ), .ZN(new_n18123_));
  NAND3_X1   g17931(.A1(new_n18121_), .A2(new_n18123_), .A3(new_n9177_), .ZN(new_n18124_));
  NAND2_X1   g17932(.A1(new_n18124_), .A2(new_n17941_), .ZN(new_n18125_));
  NAND2_X1   g17933(.A1(new_n18121_), .A2(new_n18123_), .ZN(new_n18126_));
  AOI21_X1   g17934(.A1(new_n18126_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n18127_));
  AOI21_X1   g17935(.A1(new_n18127_), .A2(new_n18125_), .B(new_n18116_), .ZN(new_n18128_));
  AOI21_X1   g17936(.A1(new_n18125_), .A2(new_n18106_), .B(new_n8742_), .ZN(new_n18129_));
  OAI21_X1   g17937(.A1(new_n18128_), .A2(new_n18129_), .B(\asqrt[24] ), .ZN(new_n18130_));
  AOI21_X1   g17938(.A1(new_n18112_), .A2(new_n18130_), .B(new_n7934_), .ZN(new_n18131_));
  NOR2_X1    g17939(.A1(new_n18115_), .A2(new_n18131_), .ZN(new_n18132_));
  AOI21_X1   g17940(.A1(new_n18132_), .A2(new_n7561_), .B(new_n17930_), .ZN(new_n18133_));
  OAI21_X1   g17941(.A1(new_n18115_), .A2(new_n18131_), .B(\asqrt[26] ), .ZN(new_n18134_));
  NAND2_X1   g17942(.A1(new_n18134_), .A2(new_n7166_), .ZN(new_n18135_));
  OAI21_X1   g17943(.A1(new_n18133_), .A2(new_n18135_), .B(new_n17926_), .ZN(new_n18136_));
  INV_X1     g17944(.I(new_n18134_), .ZN(new_n18137_));
  OAI21_X1   g17945(.A1(new_n18133_), .A2(new_n18137_), .B(\asqrt[27] ), .ZN(new_n18138_));
  NAND3_X1   g17946(.A1(new_n18136_), .A2(new_n18138_), .A3(new_n6813_), .ZN(new_n18139_));
  NAND2_X1   g17947(.A1(new_n18139_), .A2(new_n17924_), .ZN(new_n18140_));
  NAND2_X1   g17948(.A1(new_n18136_), .A2(new_n18138_), .ZN(new_n18141_));
  AOI21_X1   g17949(.A1(new_n18141_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n18142_));
  AOI21_X1   g17950(.A1(new_n18142_), .A2(new_n18140_), .B(new_n17921_), .ZN(new_n18143_));
  INV_X1     g17951(.I(new_n17926_), .ZN(new_n18144_));
  INV_X1     g17952(.I(new_n17936_), .ZN(new_n18145_));
  NOR2_X1    g17953(.A1(new_n18128_), .A2(new_n18129_), .ZN(new_n18146_));
  AOI21_X1   g17954(.A1(new_n18146_), .A2(new_n8349_), .B(new_n18145_), .ZN(new_n18147_));
  NAND2_X1   g17955(.A1(new_n18130_), .A2(new_n7934_), .ZN(new_n18148_));
  OAI21_X1   g17956(.A1(new_n18147_), .A2(new_n18148_), .B(new_n17932_), .ZN(new_n18149_));
  INV_X1     g17957(.I(new_n18130_), .ZN(new_n18150_));
  OAI21_X1   g17958(.A1(new_n18147_), .A2(new_n18150_), .B(\asqrt[25] ), .ZN(new_n18151_));
  NAND3_X1   g17959(.A1(new_n18149_), .A2(new_n18151_), .A3(new_n7561_), .ZN(new_n18152_));
  NAND2_X1   g17960(.A1(new_n18152_), .A2(new_n17929_), .ZN(new_n18153_));
  NAND2_X1   g17961(.A1(new_n18149_), .A2(new_n18151_), .ZN(new_n18154_));
  AOI21_X1   g17962(.A1(new_n18154_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n18155_));
  AOI21_X1   g17963(.A1(new_n18155_), .A2(new_n18153_), .B(new_n18144_), .ZN(new_n18156_));
  AOI21_X1   g17964(.A1(new_n18153_), .A2(new_n18134_), .B(new_n7166_), .ZN(new_n18157_));
  OAI21_X1   g17965(.A1(new_n18156_), .A2(new_n18157_), .B(\asqrt[28] ), .ZN(new_n18158_));
  AOI21_X1   g17966(.A1(new_n18140_), .A2(new_n18158_), .B(new_n6454_), .ZN(new_n18159_));
  NOR2_X1    g17967(.A1(new_n18143_), .A2(new_n18159_), .ZN(new_n18160_));
  AOI21_X1   g17968(.A1(new_n18160_), .A2(new_n6106_), .B(new_n17918_), .ZN(new_n18161_));
  OAI21_X1   g17969(.A1(new_n18143_), .A2(new_n18159_), .B(\asqrt[30] ), .ZN(new_n18162_));
  NAND2_X1   g17970(.A1(new_n18162_), .A2(new_n5750_), .ZN(new_n18163_));
  OAI21_X1   g17971(.A1(new_n18161_), .A2(new_n18163_), .B(new_n17914_), .ZN(new_n18164_));
  INV_X1     g17972(.I(new_n18162_), .ZN(new_n18165_));
  OAI21_X1   g17973(.A1(new_n18161_), .A2(new_n18165_), .B(\asqrt[31] ), .ZN(new_n18166_));
  NAND3_X1   g17974(.A1(new_n18164_), .A2(new_n18166_), .A3(new_n5435_), .ZN(new_n18167_));
  NAND2_X1   g17975(.A1(new_n18167_), .A2(new_n17912_), .ZN(new_n18168_));
  NAND2_X1   g17976(.A1(new_n18164_), .A2(new_n18166_), .ZN(new_n18169_));
  AOI21_X1   g17977(.A1(new_n18169_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n18170_));
  AOI21_X1   g17978(.A1(new_n18170_), .A2(new_n18168_), .B(new_n17909_), .ZN(new_n18171_));
  INV_X1     g17979(.I(new_n17914_), .ZN(new_n18172_));
  INV_X1     g17980(.I(new_n17924_), .ZN(new_n18173_));
  NOR2_X1    g17981(.A1(new_n18156_), .A2(new_n18157_), .ZN(new_n18174_));
  AOI21_X1   g17982(.A1(new_n18174_), .A2(new_n6813_), .B(new_n18173_), .ZN(new_n18175_));
  NAND2_X1   g17983(.A1(new_n18158_), .A2(new_n6454_), .ZN(new_n18176_));
  OAI21_X1   g17984(.A1(new_n18175_), .A2(new_n18176_), .B(new_n17920_), .ZN(new_n18177_));
  INV_X1     g17985(.I(new_n18158_), .ZN(new_n18178_));
  OAI21_X1   g17986(.A1(new_n18175_), .A2(new_n18178_), .B(\asqrt[29] ), .ZN(new_n18179_));
  NAND3_X1   g17987(.A1(new_n18177_), .A2(new_n18179_), .A3(new_n6106_), .ZN(new_n18180_));
  NAND2_X1   g17988(.A1(new_n18180_), .A2(new_n17917_), .ZN(new_n18181_));
  NAND2_X1   g17989(.A1(new_n18177_), .A2(new_n18179_), .ZN(new_n18182_));
  AOI21_X1   g17990(.A1(new_n18182_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n18183_));
  AOI21_X1   g17991(.A1(new_n18183_), .A2(new_n18181_), .B(new_n18172_), .ZN(new_n18184_));
  AOI21_X1   g17992(.A1(new_n18181_), .A2(new_n18162_), .B(new_n5750_), .ZN(new_n18185_));
  OAI21_X1   g17993(.A1(new_n18184_), .A2(new_n18185_), .B(\asqrt[32] ), .ZN(new_n18186_));
  AOI21_X1   g17994(.A1(new_n18168_), .A2(new_n18186_), .B(new_n5110_), .ZN(new_n18187_));
  NOR2_X1    g17995(.A1(new_n18171_), .A2(new_n18187_), .ZN(new_n18188_));
  AOI21_X1   g17996(.A1(new_n18188_), .A2(new_n4810_), .B(new_n17906_), .ZN(new_n18189_));
  OAI21_X1   g17997(.A1(new_n18171_), .A2(new_n18187_), .B(\asqrt[34] ), .ZN(new_n18190_));
  NAND2_X1   g17998(.A1(new_n18190_), .A2(new_n4510_), .ZN(new_n18191_));
  OAI21_X1   g17999(.A1(new_n18189_), .A2(new_n18191_), .B(new_n17902_), .ZN(new_n18192_));
  INV_X1     g18000(.I(new_n18190_), .ZN(new_n18193_));
  OAI21_X1   g18001(.A1(new_n18189_), .A2(new_n18193_), .B(\asqrt[35] ), .ZN(new_n18194_));
  NAND3_X1   g18002(.A1(new_n18192_), .A2(new_n18194_), .A3(new_n4224_), .ZN(new_n18195_));
  NAND2_X1   g18003(.A1(new_n18195_), .A2(new_n17900_), .ZN(new_n18196_));
  NAND2_X1   g18004(.A1(new_n18192_), .A2(new_n18194_), .ZN(new_n18197_));
  AOI21_X1   g18005(.A1(new_n18197_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n18198_));
  AOI21_X1   g18006(.A1(new_n18198_), .A2(new_n18196_), .B(new_n17897_), .ZN(new_n18199_));
  INV_X1     g18007(.I(new_n17902_), .ZN(new_n18200_));
  INV_X1     g18008(.I(new_n17912_), .ZN(new_n18201_));
  NOR2_X1    g18009(.A1(new_n18184_), .A2(new_n18185_), .ZN(new_n18202_));
  AOI21_X1   g18010(.A1(new_n18202_), .A2(new_n5435_), .B(new_n18201_), .ZN(new_n18203_));
  NAND2_X1   g18011(.A1(new_n18186_), .A2(new_n5110_), .ZN(new_n18204_));
  OAI21_X1   g18012(.A1(new_n18203_), .A2(new_n18204_), .B(new_n17908_), .ZN(new_n18205_));
  INV_X1     g18013(.I(new_n18186_), .ZN(new_n18206_));
  OAI21_X1   g18014(.A1(new_n18203_), .A2(new_n18206_), .B(\asqrt[33] ), .ZN(new_n18207_));
  NAND3_X1   g18015(.A1(new_n18205_), .A2(new_n18207_), .A3(new_n4810_), .ZN(new_n18208_));
  NAND2_X1   g18016(.A1(new_n18208_), .A2(new_n17905_), .ZN(new_n18209_));
  NAND2_X1   g18017(.A1(new_n18205_), .A2(new_n18207_), .ZN(new_n18210_));
  AOI21_X1   g18018(.A1(new_n18210_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n18211_));
  AOI21_X1   g18019(.A1(new_n18211_), .A2(new_n18209_), .B(new_n18200_), .ZN(new_n18212_));
  AOI21_X1   g18020(.A1(new_n18209_), .A2(new_n18190_), .B(new_n4510_), .ZN(new_n18213_));
  OAI21_X1   g18021(.A1(new_n18212_), .A2(new_n18213_), .B(\asqrt[36] ), .ZN(new_n18214_));
  AOI21_X1   g18022(.A1(new_n18196_), .A2(new_n18214_), .B(new_n3928_), .ZN(new_n18215_));
  NOR2_X1    g18023(.A1(new_n18199_), .A2(new_n18215_), .ZN(new_n18216_));
  AOI21_X1   g18024(.A1(new_n18216_), .A2(new_n3675_), .B(new_n17894_), .ZN(new_n18217_));
  OAI21_X1   g18025(.A1(new_n18199_), .A2(new_n18215_), .B(\asqrt[38] ), .ZN(new_n18218_));
  NAND2_X1   g18026(.A1(new_n18218_), .A2(new_n3400_), .ZN(new_n18219_));
  OAI21_X1   g18027(.A1(new_n18217_), .A2(new_n18219_), .B(new_n17890_), .ZN(new_n18220_));
  INV_X1     g18028(.I(new_n18218_), .ZN(new_n18221_));
  OAI21_X1   g18029(.A1(new_n18217_), .A2(new_n18221_), .B(\asqrt[39] ), .ZN(new_n18222_));
  NAND3_X1   g18030(.A1(new_n18220_), .A2(new_n18222_), .A3(new_n3167_), .ZN(new_n18223_));
  NAND2_X1   g18031(.A1(new_n18223_), .A2(new_n17888_), .ZN(new_n18224_));
  NAND2_X1   g18032(.A1(new_n18220_), .A2(new_n18222_), .ZN(new_n18225_));
  AOI21_X1   g18033(.A1(new_n18225_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n18226_));
  AOI21_X1   g18034(.A1(new_n18226_), .A2(new_n18224_), .B(new_n17885_), .ZN(new_n18227_));
  INV_X1     g18035(.I(new_n17890_), .ZN(new_n18228_));
  INV_X1     g18036(.I(new_n17900_), .ZN(new_n18229_));
  NOR2_X1    g18037(.A1(new_n18212_), .A2(new_n18213_), .ZN(new_n18230_));
  AOI21_X1   g18038(.A1(new_n18230_), .A2(new_n4224_), .B(new_n18229_), .ZN(new_n18231_));
  NAND2_X1   g18039(.A1(new_n18214_), .A2(new_n3928_), .ZN(new_n18232_));
  OAI21_X1   g18040(.A1(new_n18231_), .A2(new_n18232_), .B(new_n17896_), .ZN(new_n18233_));
  INV_X1     g18041(.I(new_n18214_), .ZN(new_n18234_));
  OAI21_X1   g18042(.A1(new_n18231_), .A2(new_n18234_), .B(\asqrt[37] ), .ZN(new_n18235_));
  NAND3_X1   g18043(.A1(new_n18233_), .A2(new_n18235_), .A3(new_n3675_), .ZN(new_n18236_));
  NAND2_X1   g18044(.A1(new_n18236_), .A2(new_n17893_), .ZN(new_n18237_));
  NAND2_X1   g18045(.A1(new_n18233_), .A2(new_n18235_), .ZN(new_n18238_));
  AOI21_X1   g18046(.A1(new_n18238_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n18239_));
  AOI21_X1   g18047(.A1(new_n18239_), .A2(new_n18237_), .B(new_n18228_), .ZN(new_n18240_));
  AOI21_X1   g18048(.A1(new_n18237_), .A2(new_n18218_), .B(new_n3400_), .ZN(new_n18241_));
  OAI21_X1   g18049(.A1(new_n18240_), .A2(new_n18241_), .B(\asqrt[40] ), .ZN(new_n18242_));
  AOI21_X1   g18050(.A1(new_n18224_), .A2(new_n18242_), .B(new_n2912_), .ZN(new_n18243_));
  NOR2_X1    g18051(.A1(new_n18227_), .A2(new_n18243_), .ZN(new_n18244_));
  AOI21_X1   g18052(.A1(new_n18244_), .A2(new_n2699_), .B(new_n17882_), .ZN(new_n18245_));
  OAI21_X1   g18053(.A1(new_n18227_), .A2(new_n18243_), .B(\asqrt[42] ), .ZN(new_n18246_));
  NAND2_X1   g18054(.A1(new_n18246_), .A2(new_n2464_), .ZN(new_n18247_));
  OAI21_X1   g18055(.A1(new_n18245_), .A2(new_n18247_), .B(new_n17878_), .ZN(new_n18248_));
  INV_X1     g18056(.I(new_n18246_), .ZN(new_n18249_));
  OAI21_X1   g18057(.A1(new_n18245_), .A2(new_n18249_), .B(\asqrt[43] ), .ZN(new_n18250_));
  NAND3_X1   g18058(.A1(new_n18248_), .A2(new_n18250_), .A3(new_n2271_), .ZN(new_n18251_));
  NAND2_X1   g18059(.A1(new_n18251_), .A2(new_n17876_), .ZN(new_n18252_));
  NAND2_X1   g18060(.A1(new_n18248_), .A2(new_n18250_), .ZN(new_n18253_));
  AOI21_X1   g18061(.A1(new_n18253_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n18254_));
  AOI21_X1   g18062(.A1(new_n18254_), .A2(new_n18252_), .B(new_n17873_), .ZN(new_n18255_));
  INV_X1     g18063(.I(new_n17878_), .ZN(new_n18256_));
  INV_X1     g18064(.I(new_n17888_), .ZN(new_n18257_));
  NOR2_X1    g18065(.A1(new_n18240_), .A2(new_n18241_), .ZN(new_n18258_));
  AOI21_X1   g18066(.A1(new_n18258_), .A2(new_n3167_), .B(new_n18257_), .ZN(new_n18259_));
  NAND2_X1   g18067(.A1(new_n18242_), .A2(new_n2912_), .ZN(new_n18260_));
  OAI21_X1   g18068(.A1(new_n18259_), .A2(new_n18260_), .B(new_n17884_), .ZN(new_n18261_));
  INV_X1     g18069(.I(new_n18242_), .ZN(new_n18262_));
  OAI21_X1   g18070(.A1(new_n18259_), .A2(new_n18262_), .B(\asqrt[41] ), .ZN(new_n18263_));
  NAND3_X1   g18071(.A1(new_n18261_), .A2(new_n18263_), .A3(new_n2699_), .ZN(new_n18264_));
  NAND2_X1   g18072(.A1(new_n18264_), .A2(new_n17881_), .ZN(new_n18265_));
  NAND2_X1   g18073(.A1(new_n18261_), .A2(new_n18263_), .ZN(new_n18266_));
  AOI21_X1   g18074(.A1(new_n18266_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n18267_));
  AOI21_X1   g18075(.A1(new_n18267_), .A2(new_n18265_), .B(new_n18256_), .ZN(new_n18268_));
  AOI21_X1   g18076(.A1(new_n18265_), .A2(new_n18246_), .B(new_n2464_), .ZN(new_n18269_));
  OAI21_X1   g18077(.A1(new_n18268_), .A2(new_n18269_), .B(\asqrt[44] ), .ZN(new_n18270_));
  AOI21_X1   g18078(.A1(new_n18252_), .A2(new_n18270_), .B(new_n2072_), .ZN(new_n18271_));
  NOR2_X1    g18079(.A1(new_n18255_), .A2(new_n18271_), .ZN(new_n18272_));
  AOI21_X1   g18080(.A1(new_n18272_), .A2(new_n1884_), .B(new_n17870_), .ZN(new_n18273_));
  OAI21_X1   g18081(.A1(new_n18255_), .A2(new_n18271_), .B(\asqrt[46] ), .ZN(new_n18274_));
  NAND2_X1   g18082(.A1(new_n18274_), .A2(new_n1688_), .ZN(new_n18275_));
  OAI21_X1   g18083(.A1(new_n18273_), .A2(new_n18275_), .B(new_n17866_), .ZN(new_n18276_));
  INV_X1     g18084(.I(new_n18274_), .ZN(new_n18277_));
  OAI21_X1   g18085(.A1(new_n18273_), .A2(new_n18277_), .B(\asqrt[47] ), .ZN(new_n18278_));
  NAND3_X1   g18086(.A1(new_n18276_), .A2(new_n18278_), .A3(new_n1533_), .ZN(new_n18279_));
  NAND2_X1   g18087(.A1(new_n18279_), .A2(new_n17864_), .ZN(new_n18280_));
  NAND2_X1   g18088(.A1(new_n18276_), .A2(new_n18278_), .ZN(new_n18281_));
  AOI21_X1   g18089(.A1(new_n18281_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n18282_));
  AOI21_X1   g18090(.A1(new_n18282_), .A2(new_n18280_), .B(new_n17861_), .ZN(new_n18283_));
  INV_X1     g18091(.I(new_n17866_), .ZN(new_n18284_));
  INV_X1     g18092(.I(new_n17876_), .ZN(new_n18285_));
  NOR2_X1    g18093(.A1(new_n18268_), .A2(new_n18269_), .ZN(new_n18286_));
  AOI21_X1   g18094(.A1(new_n18286_), .A2(new_n2271_), .B(new_n18285_), .ZN(new_n18287_));
  NAND2_X1   g18095(.A1(new_n18270_), .A2(new_n2072_), .ZN(new_n18288_));
  OAI21_X1   g18096(.A1(new_n18287_), .A2(new_n18288_), .B(new_n17872_), .ZN(new_n18289_));
  INV_X1     g18097(.I(new_n18270_), .ZN(new_n18290_));
  OAI21_X1   g18098(.A1(new_n18287_), .A2(new_n18290_), .B(\asqrt[45] ), .ZN(new_n18291_));
  NAND3_X1   g18099(.A1(new_n18289_), .A2(new_n18291_), .A3(new_n1884_), .ZN(new_n18292_));
  NAND2_X1   g18100(.A1(new_n18292_), .A2(new_n17869_), .ZN(new_n18293_));
  NAND2_X1   g18101(.A1(new_n18289_), .A2(new_n18291_), .ZN(new_n18294_));
  AOI21_X1   g18102(.A1(new_n18294_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n18295_));
  AOI21_X1   g18103(.A1(new_n18295_), .A2(new_n18293_), .B(new_n18284_), .ZN(new_n18296_));
  AOI21_X1   g18104(.A1(new_n18293_), .A2(new_n18274_), .B(new_n1688_), .ZN(new_n18297_));
  OAI21_X1   g18105(.A1(new_n18296_), .A2(new_n18297_), .B(\asqrt[48] ), .ZN(new_n18298_));
  AOI21_X1   g18106(.A1(new_n18280_), .A2(new_n18298_), .B(new_n1368_), .ZN(new_n18299_));
  NOR2_X1    g18107(.A1(new_n18283_), .A2(new_n18299_), .ZN(new_n18300_));
  AOI21_X1   g18108(.A1(new_n18300_), .A2(new_n1228_), .B(new_n17858_), .ZN(new_n18301_));
  OAI21_X1   g18109(.A1(new_n18283_), .A2(new_n18299_), .B(\asqrt[50] ), .ZN(new_n18302_));
  NAND2_X1   g18110(.A1(new_n18302_), .A2(new_n1088_), .ZN(new_n18303_));
  OAI21_X1   g18111(.A1(new_n18301_), .A2(new_n18303_), .B(new_n17854_), .ZN(new_n18304_));
  INV_X1     g18112(.I(new_n18302_), .ZN(new_n18305_));
  OAI21_X1   g18113(.A1(new_n18301_), .A2(new_n18305_), .B(\asqrt[51] ), .ZN(new_n18306_));
  NAND3_X1   g18114(.A1(new_n18304_), .A2(new_n18306_), .A3(new_n962_), .ZN(new_n18307_));
  NAND2_X1   g18115(.A1(new_n18307_), .A2(new_n17852_), .ZN(new_n18308_));
  NAND2_X1   g18116(.A1(new_n18304_), .A2(new_n18306_), .ZN(new_n18309_));
  AOI21_X1   g18117(.A1(new_n18309_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n18310_));
  AOI21_X1   g18118(.A1(new_n18310_), .A2(new_n18308_), .B(new_n17849_), .ZN(new_n18311_));
  INV_X1     g18119(.I(new_n17854_), .ZN(new_n18312_));
  INV_X1     g18120(.I(new_n17864_), .ZN(new_n18313_));
  NOR2_X1    g18121(.A1(new_n18296_), .A2(new_n18297_), .ZN(new_n18314_));
  AOI21_X1   g18122(.A1(new_n18314_), .A2(new_n1533_), .B(new_n18313_), .ZN(new_n18315_));
  NAND2_X1   g18123(.A1(new_n18298_), .A2(new_n1368_), .ZN(new_n18316_));
  OAI21_X1   g18124(.A1(new_n18315_), .A2(new_n18316_), .B(new_n17860_), .ZN(new_n18317_));
  INV_X1     g18125(.I(new_n18298_), .ZN(new_n18318_));
  OAI21_X1   g18126(.A1(new_n18315_), .A2(new_n18318_), .B(\asqrt[49] ), .ZN(new_n18319_));
  NAND3_X1   g18127(.A1(new_n18317_), .A2(new_n18319_), .A3(new_n1228_), .ZN(new_n18320_));
  NAND2_X1   g18128(.A1(new_n18320_), .A2(new_n17857_), .ZN(new_n18321_));
  NAND2_X1   g18129(.A1(new_n18317_), .A2(new_n18319_), .ZN(new_n18322_));
  AOI21_X1   g18130(.A1(new_n18322_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n18323_));
  AOI21_X1   g18131(.A1(new_n18323_), .A2(new_n18321_), .B(new_n18312_), .ZN(new_n18324_));
  AOI21_X1   g18132(.A1(new_n18321_), .A2(new_n18302_), .B(new_n1088_), .ZN(new_n18325_));
  OAI21_X1   g18133(.A1(new_n18324_), .A2(new_n18325_), .B(\asqrt[52] ), .ZN(new_n18326_));
  AOI21_X1   g18134(.A1(new_n18308_), .A2(new_n18326_), .B(new_n842_), .ZN(new_n18327_));
  NOR2_X1    g18135(.A1(new_n18311_), .A2(new_n18327_), .ZN(new_n18328_));
  AOI21_X1   g18136(.A1(new_n18328_), .A2(new_n720_), .B(new_n17846_), .ZN(new_n18329_));
  OAI21_X1   g18137(.A1(new_n18311_), .A2(new_n18327_), .B(\asqrt[54] ), .ZN(new_n18330_));
  NAND2_X1   g18138(.A1(new_n18330_), .A2(new_n630_), .ZN(new_n18331_));
  OAI21_X1   g18139(.A1(new_n18329_), .A2(new_n18331_), .B(new_n17842_), .ZN(new_n18332_));
  INV_X1     g18140(.I(new_n18330_), .ZN(new_n18333_));
  OAI21_X1   g18141(.A1(new_n18329_), .A2(new_n18333_), .B(\asqrt[55] ), .ZN(new_n18334_));
  NAND3_X1   g18142(.A1(new_n18332_), .A2(new_n18334_), .A3(new_n545_), .ZN(new_n18335_));
  NAND2_X1   g18143(.A1(new_n18335_), .A2(new_n17840_), .ZN(new_n18336_));
  NAND2_X1   g18144(.A1(new_n18332_), .A2(new_n18334_), .ZN(new_n18337_));
  AOI21_X1   g18145(.A1(new_n18337_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n18338_));
  AOI21_X1   g18146(.A1(new_n18338_), .A2(new_n18336_), .B(new_n17837_), .ZN(new_n18339_));
  INV_X1     g18147(.I(new_n17842_), .ZN(new_n18340_));
  INV_X1     g18148(.I(new_n17852_), .ZN(new_n18341_));
  NOR2_X1    g18149(.A1(new_n18324_), .A2(new_n18325_), .ZN(new_n18342_));
  AOI21_X1   g18150(.A1(new_n18342_), .A2(new_n962_), .B(new_n18341_), .ZN(new_n18343_));
  NAND2_X1   g18151(.A1(new_n18326_), .A2(new_n842_), .ZN(new_n18344_));
  OAI21_X1   g18152(.A1(new_n18343_), .A2(new_n18344_), .B(new_n17848_), .ZN(new_n18345_));
  INV_X1     g18153(.I(new_n18326_), .ZN(new_n18346_));
  OAI21_X1   g18154(.A1(new_n18343_), .A2(new_n18346_), .B(\asqrt[53] ), .ZN(new_n18347_));
  NAND3_X1   g18155(.A1(new_n18345_), .A2(new_n18347_), .A3(new_n720_), .ZN(new_n18348_));
  NAND2_X1   g18156(.A1(new_n18348_), .A2(new_n17845_), .ZN(new_n18349_));
  NAND2_X1   g18157(.A1(new_n18345_), .A2(new_n18347_), .ZN(new_n18350_));
  AOI21_X1   g18158(.A1(new_n18350_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n18351_));
  AOI21_X1   g18159(.A1(new_n18351_), .A2(new_n18349_), .B(new_n18340_), .ZN(new_n18352_));
  AOI21_X1   g18160(.A1(new_n18349_), .A2(new_n18330_), .B(new_n630_), .ZN(new_n18353_));
  OAI21_X1   g18161(.A1(new_n18352_), .A2(new_n18353_), .B(\asqrt[56] ), .ZN(new_n18354_));
  AOI21_X1   g18162(.A1(new_n18336_), .A2(new_n18354_), .B(new_n450_), .ZN(new_n18355_));
  NOR2_X1    g18163(.A1(new_n18339_), .A2(new_n18355_), .ZN(new_n18356_));
  AOI21_X1   g18164(.A1(new_n18356_), .A2(new_n403_), .B(new_n17834_), .ZN(new_n18357_));
  OAI21_X1   g18165(.A1(new_n18339_), .A2(new_n18355_), .B(\asqrt[58] ), .ZN(new_n18358_));
  NAND2_X1   g18166(.A1(new_n18358_), .A2(new_n339_), .ZN(new_n18359_));
  OAI21_X1   g18167(.A1(new_n18357_), .A2(new_n18359_), .B(new_n17830_), .ZN(new_n18360_));
  INV_X1     g18168(.I(new_n18358_), .ZN(new_n18361_));
  OAI21_X1   g18169(.A1(new_n18357_), .A2(new_n18361_), .B(\asqrt[59] ), .ZN(new_n18362_));
  NAND3_X1   g18170(.A1(new_n18360_), .A2(new_n18362_), .A3(new_n288_), .ZN(new_n18363_));
  INV_X1     g18171(.I(new_n17830_), .ZN(new_n18364_));
  INV_X1     g18172(.I(new_n17840_), .ZN(new_n18365_));
  NOR2_X1    g18173(.A1(new_n18352_), .A2(new_n18353_), .ZN(new_n18366_));
  AOI21_X1   g18174(.A1(new_n18366_), .A2(new_n545_), .B(new_n18365_), .ZN(new_n18367_));
  NAND2_X1   g18175(.A1(new_n18354_), .A2(new_n450_), .ZN(new_n18368_));
  OAI21_X1   g18176(.A1(new_n18367_), .A2(new_n18368_), .B(new_n17836_), .ZN(new_n18369_));
  INV_X1     g18177(.I(new_n18354_), .ZN(new_n18370_));
  OAI21_X1   g18178(.A1(new_n18367_), .A2(new_n18370_), .B(\asqrt[57] ), .ZN(new_n18371_));
  NAND3_X1   g18179(.A1(new_n18369_), .A2(new_n18371_), .A3(new_n403_), .ZN(new_n18372_));
  NAND2_X1   g18180(.A1(new_n18372_), .A2(new_n17833_), .ZN(new_n18373_));
  NAND2_X1   g18181(.A1(new_n18369_), .A2(new_n18371_), .ZN(new_n18374_));
  AOI21_X1   g18182(.A1(new_n18374_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n18375_));
  AOI21_X1   g18183(.A1(new_n18375_), .A2(new_n18373_), .B(new_n18364_), .ZN(new_n18376_));
  AOI21_X1   g18184(.A1(new_n18373_), .A2(new_n18358_), .B(new_n339_), .ZN(new_n18377_));
  OAI21_X1   g18185(.A1(new_n18376_), .A2(new_n18377_), .B(\asqrt[60] ), .ZN(new_n18378_));
  NOR2_X1    g18186(.A1(new_n17826_), .A2(new_n17247_), .ZN(new_n18379_));
  NOR2_X1    g18187(.A1(new_n17816_), .A2(new_n17822_), .ZN(new_n18380_));
  AOI21_X1   g18188(.A1(new_n18380_), .A2(new_n17826_), .B(new_n18379_), .ZN(new_n18381_));
  NOR2_X1    g18189(.A1(new_n18381_), .A2(new_n193_), .ZN(new_n18382_));
  INV_X1     g18190(.I(new_n18382_), .ZN(new_n18383_));
  NAND3_X1   g18191(.A1(\asqrt[5] ), .A2(new_n17796_), .A3(new_n17807_), .ZN(new_n18384_));
  XOR2_X1    g18192(.A1(new_n18384_), .A2(new_n17812_), .Z(new_n18385_));
  INV_X1     g18193(.I(new_n18385_), .ZN(new_n18386_));
  AOI21_X1   g18194(.A1(new_n18380_), .A2(new_n17997_), .B(new_n17815_), .ZN(new_n18387_));
  NAND2_X1   g18195(.A1(new_n18363_), .A2(new_n17819_), .ZN(new_n18388_));
  AOI21_X1   g18196(.A1(new_n18388_), .A2(new_n18378_), .B(new_n242_), .ZN(new_n18389_));
  NAND3_X1   g18197(.A1(\asqrt[5] ), .A2(new_n17772_), .A3(new_n17788_), .ZN(new_n18390_));
  XOR2_X1    g18198(.A1(new_n18390_), .A2(new_n17800_), .Z(new_n18391_));
  INV_X1     g18199(.I(new_n18391_), .ZN(new_n18392_));
  NAND2_X1   g18200(.A1(new_n18360_), .A2(new_n18362_), .ZN(new_n18393_));
  AOI21_X1   g18201(.A1(new_n18393_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n18394_));
  AOI21_X1   g18202(.A1(new_n18394_), .A2(new_n18388_), .B(new_n18392_), .ZN(new_n18395_));
  OAI21_X1   g18203(.A1(new_n18395_), .A2(new_n18389_), .B(\asqrt[62] ), .ZN(new_n18396_));
  INV_X1     g18204(.I(new_n18396_), .ZN(new_n18397_));
  NOR2_X1    g18205(.A1(new_n18395_), .A2(new_n18389_), .ZN(new_n18398_));
  AOI21_X1   g18206(.A1(new_n17773_), .A2(new_n17794_), .B(new_n17789_), .ZN(new_n18399_));
  NAND2_X1   g18207(.A1(\asqrt[5] ), .A2(new_n18399_), .ZN(new_n18400_));
  XOR2_X1    g18208(.A1(new_n18400_), .A2(new_n17792_), .Z(new_n18401_));
  INV_X1     g18209(.I(new_n18401_), .ZN(new_n18402_));
  AOI21_X1   g18210(.A1(new_n18398_), .A2(new_n234_), .B(new_n18402_), .ZN(new_n18403_));
  OAI21_X1   g18211(.A1(new_n18403_), .A2(new_n18397_), .B(new_n18387_), .ZN(new_n18404_));
  OAI21_X1   g18212(.A1(new_n18404_), .A2(new_n18386_), .B(new_n193_), .ZN(new_n18405_));
  NOR3_X1    g18213(.A1(new_n18403_), .A2(new_n18397_), .A3(new_n18385_), .ZN(new_n18406_));
  INV_X1     g18214(.I(new_n18406_), .ZN(new_n18407_));
  NAND3_X1   g18215(.A1(new_n18405_), .A2(new_n18383_), .A3(new_n18407_), .ZN(\asqrt[4] ));
  NAND3_X1   g18216(.A1(\asqrt[4] ), .A2(new_n18363_), .A3(new_n18378_), .ZN(new_n18409_));
  XOR2_X1    g18217(.A1(new_n18409_), .A2(new_n17820_), .Z(new_n18410_));
  INV_X1     g18218(.I(new_n18410_), .ZN(new_n18411_));
  NOR2_X1    g18219(.A1(new_n18376_), .A2(new_n18377_), .ZN(new_n18412_));
  AOI21_X1   g18220(.A1(new_n18412_), .A2(new_n288_), .B(new_n17820_), .ZN(new_n18413_));
  INV_X1     g18221(.I(new_n18378_), .ZN(new_n18414_));
  OAI21_X1   g18222(.A1(new_n18413_), .A2(new_n18414_), .B(\asqrt[61] ), .ZN(new_n18415_));
  NAND2_X1   g18223(.A1(new_n18378_), .A2(new_n242_), .ZN(new_n18416_));
  OAI21_X1   g18224(.A1(new_n18413_), .A2(new_n18416_), .B(new_n18391_), .ZN(new_n18417_));
  NAND3_X1   g18225(.A1(new_n18417_), .A2(new_n18415_), .A3(new_n234_), .ZN(new_n18418_));
  NAND2_X1   g18226(.A1(new_n18418_), .A2(new_n18401_), .ZN(new_n18419_));
  NAND2_X1   g18227(.A1(new_n18419_), .A2(new_n18396_), .ZN(new_n18420_));
  INV_X1     g18228(.I(new_n18387_), .ZN(new_n18421_));
  AOI21_X1   g18229(.A1(new_n18419_), .A2(new_n18396_), .B(new_n18421_), .ZN(new_n18422_));
  AOI21_X1   g18230(.A1(new_n18422_), .A2(new_n18385_), .B(\asqrt[63] ), .ZN(new_n18423_));
  NOR3_X1    g18231(.A1(new_n18423_), .A2(new_n18382_), .A3(new_n18406_), .ZN(new_n18424_));
  NOR3_X1    g18232(.A1(new_n18424_), .A2(new_n18386_), .A3(new_n18420_), .ZN(new_n18425_));
  AOI21_X1   g18233(.A1(new_n18386_), .A2(new_n18420_), .B(new_n18425_), .ZN(new_n18426_));
  NOR2_X1    g18234(.A1(new_n18426_), .A2(new_n193_), .ZN(new_n18427_));
  INV_X1     g18235(.I(new_n18427_), .ZN(new_n18428_));
  NAND3_X1   g18236(.A1(\asqrt[4] ), .A2(new_n18396_), .A3(new_n18418_), .ZN(new_n18429_));
  XOR2_X1    g18237(.A1(new_n18429_), .A2(new_n18402_), .Z(new_n18430_));
  NOR2_X1    g18238(.A1(new_n18424_), .A2(new_n18386_), .ZN(new_n18431_));
  AOI21_X1   g18239(.A1(new_n18431_), .A2(new_n18420_), .B(new_n18406_), .ZN(new_n18432_));
  OAI21_X1   g18240(.A1(new_n18357_), .A2(new_n18359_), .B(new_n18362_), .ZN(new_n18433_));
  NOR2_X1    g18241(.A1(new_n18424_), .A2(new_n18433_), .ZN(new_n18434_));
  XOR2_X1    g18242(.A1(new_n18434_), .A2(new_n17830_), .Z(new_n18435_));
  NAND3_X1   g18243(.A1(\asqrt[4] ), .A2(new_n18372_), .A3(new_n18358_), .ZN(new_n18436_));
  XOR2_X1    g18244(.A1(new_n18436_), .A2(new_n17834_), .Z(new_n18437_));
  OAI21_X1   g18245(.A1(new_n18367_), .A2(new_n18368_), .B(new_n18371_), .ZN(new_n18438_));
  NOR2_X1    g18246(.A1(new_n18424_), .A2(new_n18438_), .ZN(new_n18439_));
  XOR2_X1    g18247(.A1(new_n18439_), .A2(new_n17836_), .Z(new_n18440_));
  INV_X1     g18248(.I(new_n18440_), .ZN(new_n18441_));
  NAND3_X1   g18249(.A1(\asqrt[4] ), .A2(new_n18335_), .A3(new_n18354_), .ZN(new_n18442_));
  XOR2_X1    g18250(.A1(new_n18442_), .A2(new_n18365_), .Z(new_n18443_));
  INV_X1     g18251(.I(new_n18443_), .ZN(new_n18444_));
  OAI21_X1   g18252(.A1(new_n18329_), .A2(new_n18331_), .B(new_n18334_), .ZN(new_n18445_));
  NOR2_X1    g18253(.A1(new_n18424_), .A2(new_n18445_), .ZN(new_n18446_));
  XOR2_X1    g18254(.A1(new_n18446_), .A2(new_n17842_), .Z(new_n18447_));
  NAND3_X1   g18255(.A1(\asqrt[4] ), .A2(new_n18348_), .A3(new_n18330_), .ZN(new_n18448_));
  XOR2_X1    g18256(.A1(new_n18448_), .A2(new_n17846_), .Z(new_n18449_));
  OAI21_X1   g18257(.A1(new_n18343_), .A2(new_n18344_), .B(new_n18347_), .ZN(new_n18450_));
  NOR2_X1    g18258(.A1(new_n18424_), .A2(new_n18450_), .ZN(new_n18451_));
  XOR2_X1    g18259(.A1(new_n18451_), .A2(new_n17848_), .Z(new_n18452_));
  INV_X1     g18260(.I(new_n18452_), .ZN(new_n18453_));
  NAND3_X1   g18261(.A1(\asqrt[4] ), .A2(new_n18307_), .A3(new_n18326_), .ZN(new_n18454_));
  XOR2_X1    g18262(.A1(new_n18454_), .A2(new_n18341_), .Z(new_n18455_));
  INV_X1     g18263(.I(new_n18455_), .ZN(new_n18456_));
  OAI21_X1   g18264(.A1(new_n18301_), .A2(new_n18303_), .B(new_n18306_), .ZN(new_n18457_));
  NOR2_X1    g18265(.A1(new_n18424_), .A2(new_n18457_), .ZN(new_n18458_));
  XOR2_X1    g18266(.A1(new_n18458_), .A2(new_n17854_), .Z(new_n18459_));
  NAND3_X1   g18267(.A1(\asqrt[4] ), .A2(new_n18320_), .A3(new_n18302_), .ZN(new_n18460_));
  XOR2_X1    g18268(.A1(new_n18460_), .A2(new_n17858_), .Z(new_n18461_));
  OAI21_X1   g18269(.A1(new_n18315_), .A2(new_n18316_), .B(new_n18319_), .ZN(new_n18462_));
  NOR2_X1    g18270(.A1(new_n18424_), .A2(new_n18462_), .ZN(new_n18463_));
  XOR2_X1    g18271(.A1(new_n18463_), .A2(new_n17860_), .Z(new_n18464_));
  INV_X1     g18272(.I(new_n18464_), .ZN(new_n18465_));
  NAND3_X1   g18273(.A1(\asqrt[4] ), .A2(new_n18279_), .A3(new_n18298_), .ZN(new_n18466_));
  XOR2_X1    g18274(.A1(new_n18466_), .A2(new_n18313_), .Z(new_n18467_));
  INV_X1     g18275(.I(new_n18467_), .ZN(new_n18468_));
  OAI21_X1   g18276(.A1(new_n18273_), .A2(new_n18275_), .B(new_n18278_), .ZN(new_n18469_));
  NOR2_X1    g18277(.A1(new_n18424_), .A2(new_n18469_), .ZN(new_n18470_));
  XOR2_X1    g18278(.A1(new_n18470_), .A2(new_n17866_), .Z(new_n18471_));
  NAND3_X1   g18279(.A1(\asqrt[4] ), .A2(new_n18292_), .A3(new_n18274_), .ZN(new_n18472_));
  XOR2_X1    g18280(.A1(new_n18472_), .A2(new_n17870_), .Z(new_n18473_));
  OAI21_X1   g18281(.A1(new_n18287_), .A2(new_n18288_), .B(new_n18291_), .ZN(new_n18474_));
  NOR2_X1    g18282(.A1(new_n18424_), .A2(new_n18474_), .ZN(new_n18475_));
  XOR2_X1    g18283(.A1(new_n18475_), .A2(new_n17872_), .Z(new_n18476_));
  INV_X1     g18284(.I(new_n18476_), .ZN(new_n18477_));
  NAND3_X1   g18285(.A1(\asqrt[4] ), .A2(new_n18251_), .A3(new_n18270_), .ZN(new_n18478_));
  XOR2_X1    g18286(.A1(new_n18478_), .A2(new_n18285_), .Z(new_n18479_));
  INV_X1     g18287(.I(new_n18479_), .ZN(new_n18480_));
  OAI21_X1   g18288(.A1(new_n18245_), .A2(new_n18247_), .B(new_n18250_), .ZN(new_n18481_));
  NOR2_X1    g18289(.A1(new_n18424_), .A2(new_n18481_), .ZN(new_n18482_));
  XOR2_X1    g18290(.A1(new_n18482_), .A2(new_n17878_), .Z(new_n18483_));
  NAND3_X1   g18291(.A1(\asqrt[4] ), .A2(new_n18264_), .A3(new_n18246_), .ZN(new_n18484_));
  XOR2_X1    g18292(.A1(new_n18484_), .A2(new_n17882_), .Z(new_n18485_));
  OAI21_X1   g18293(.A1(new_n18259_), .A2(new_n18260_), .B(new_n18263_), .ZN(new_n18486_));
  NOR2_X1    g18294(.A1(new_n18424_), .A2(new_n18486_), .ZN(new_n18487_));
  XOR2_X1    g18295(.A1(new_n18487_), .A2(new_n17884_), .Z(new_n18488_));
  INV_X1     g18296(.I(new_n18488_), .ZN(new_n18489_));
  NAND3_X1   g18297(.A1(\asqrt[4] ), .A2(new_n18223_), .A3(new_n18242_), .ZN(new_n18490_));
  XOR2_X1    g18298(.A1(new_n18490_), .A2(new_n18257_), .Z(new_n18491_));
  INV_X1     g18299(.I(new_n18491_), .ZN(new_n18492_));
  OAI21_X1   g18300(.A1(new_n18217_), .A2(new_n18219_), .B(new_n18222_), .ZN(new_n18493_));
  NOR2_X1    g18301(.A1(new_n18424_), .A2(new_n18493_), .ZN(new_n18494_));
  XOR2_X1    g18302(.A1(new_n18494_), .A2(new_n17890_), .Z(new_n18495_));
  NAND3_X1   g18303(.A1(\asqrt[4] ), .A2(new_n18236_), .A3(new_n18218_), .ZN(new_n18496_));
  XOR2_X1    g18304(.A1(new_n18496_), .A2(new_n17894_), .Z(new_n18497_));
  OAI21_X1   g18305(.A1(new_n18231_), .A2(new_n18232_), .B(new_n18235_), .ZN(new_n18498_));
  NOR2_X1    g18306(.A1(new_n18424_), .A2(new_n18498_), .ZN(new_n18499_));
  XOR2_X1    g18307(.A1(new_n18499_), .A2(new_n17896_), .Z(new_n18500_));
  INV_X1     g18308(.I(new_n18500_), .ZN(new_n18501_));
  NAND3_X1   g18309(.A1(\asqrt[4] ), .A2(new_n18195_), .A3(new_n18214_), .ZN(new_n18502_));
  XOR2_X1    g18310(.A1(new_n18502_), .A2(new_n18229_), .Z(new_n18503_));
  INV_X1     g18311(.I(new_n18503_), .ZN(new_n18504_));
  OAI21_X1   g18312(.A1(new_n18189_), .A2(new_n18191_), .B(new_n18194_), .ZN(new_n18505_));
  NOR2_X1    g18313(.A1(new_n18424_), .A2(new_n18505_), .ZN(new_n18506_));
  XOR2_X1    g18314(.A1(new_n18506_), .A2(new_n17902_), .Z(new_n18507_));
  NAND3_X1   g18315(.A1(\asqrt[4] ), .A2(new_n18208_), .A3(new_n18190_), .ZN(new_n18508_));
  XOR2_X1    g18316(.A1(new_n18508_), .A2(new_n17906_), .Z(new_n18509_));
  OAI21_X1   g18317(.A1(new_n18203_), .A2(new_n18204_), .B(new_n18207_), .ZN(new_n18510_));
  NOR2_X1    g18318(.A1(new_n18424_), .A2(new_n18510_), .ZN(new_n18511_));
  XOR2_X1    g18319(.A1(new_n18511_), .A2(new_n17908_), .Z(new_n18512_));
  INV_X1     g18320(.I(new_n18512_), .ZN(new_n18513_));
  NAND3_X1   g18321(.A1(\asqrt[4] ), .A2(new_n18167_), .A3(new_n18186_), .ZN(new_n18514_));
  XOR2_X1    g18322(.A1(new_n18514_), .A2(new_n18201_), .Z(new_n18515_));
  INV_X1     g18323(.I(new_n18515_), .ZN(new_n18516_));
  OAI21_X1   g18324(.A1(new_n18161_), .A2(new_n18163_), .B(new_n18166_), .ZN(new_n18517_));
  NOR2_X1    g18325(.A1(new_n18424_), .A2(new_n18517_), .ZN(new_n18518_));
  XOR2_X1    g18326(.A1(new_n18518_), .A2(new_n17914_), .Z(new_n18519_));
  NAND3_X1   g18327(.A1(\asqrt[4] ), .A2(new_n18180_), .A3(new_n18162_), .ZN(new_n18520_));
  XOR2_X1    g18328(.A1(new_n18520_), .A2(new_n17918_), .Z(new_n18521_));
  OAI21_X1   g18329(.A1(new_n18175_), .A2(new_n18176_), .B(new_n18179_), .ZN(new_n18522_));
  NOR2_X1    g18330(.A1(new_n18424_), .A2(new_n18522_), .ZN(new_n18523_));
  XOR2_X1    g18331(.A1(new_n18523_), .A2(new_n17920_), .Z(new_n18524_));
  INV_X1     g18332(.I(new_n18524_), .ZN(new_n18525_));
  NAND3_X1   g18333(.A1(\asqrt[4] ), .A2(new_n18139_), .A3(new_n18158_), .ZN(new_n18526_));
  XOR2_X1    g18334(.A1(new_n18526_), .A2(new_n18173_), .Z(new_n18527_));
  INV_X1     g18335(.I(new_n18527_), .ZN(new_n18528_));
  OAI21_X1   g18336(.A1(new_n18133_), .A2(new_n18135_), .B(new_n18138_), .ZN(new_n18529_));
  NOR2_X1    g18337(.A1(new_n18424_), .A2(new_n18529_), .ZN(new_n18530_));
  XOR2_X1    g18338(.A1(new_n18530_), .A2(new_n17926_), .Z(new_n18531_));
  NAND3_X1   g18339(.A1(\asqrt[4] ), .A2(new_n18152_), .A3(new_n18134_), .ZN(new_n18532_));
  XOR2_X1    g18340(.A1(new_n18532_), .A2(new_n17930_), .Z(new_n18533_));
  OAI21_X1   g18341(.A1(new_n18147_), .A2(new_n18148_), .B(new_n18151_), .ZN(new_n18534_));
  NOR2_X1    g18342(.A1(new_n18424_), .A2(new_n18534_), .ZN(new_n18535_));
  XOR2_X1    g18343(.A1(new_n18535_), .A2(new_n17932_), .Z(new_n18536_));
  INV_X1     g18344(.I(new_n18536_), .ZN(new_n18537_));
  NAND3_X1   g18345(.A1(\asqrt[4] ), .A2(new_n18111_), .A3(new_n18130_), .ZN(new_n18538_));
  XOR2_X1    g18346(.A1(new_n18538_), .A2(new_n18145_), .Z(new_n18539_));
  INV_X1     g18347(.I(new_n18539_), .ZN(new_n18540_));
  OAI21_X1   g18348(.A1(new_n18105_), .A2(new_n18107_), .B(new_n18110_), .ZN(new_n18541_));
  NOR2_X1    g18349(.A1(new_n18424_), .A2(new_n18541_), .ZN(new_n18542_));
  XOR2_X1    g18350(.A1(new_n18542_), .A2(new_n17938_), .Z(new_n18543_));
  NAND3_X1   g18351(.A1(\asqrt[4] ), .A2(new_n18124_), .A3(new_n18106_), .ZN(new_n18544_));
  XOR2_X1    g18352(.A1(new_n18544_), .A2(new_n17942_), .Z(new_n18545_));
  OAI21_X1   g18353(.A1(new_n18119_), .A2(new_n18120_), .B(new_n18123_), .ZN(new_n18546_));
  NOR2_X1    g18354(.A1(new_n18424_), .A2(new_n18546_), .ZN(new_n18547_));
  XOR2_X1    g18355(.A1(new_n18547_), .A2(new_n17944_), .Z(new_n18548_));
  INV_X1     g18356(.I(new_n18548_), .ZN(new_n18549_));
  NAND3_X1   g18357(.A1(\asqrt[4] ), .A2(new_n18083_), .A3(new_n18102_), .ZN(new_n18550_));
  XOR2_X1    g18358(.A1(new_n18550_), .A2(new_n18117_), .Z(new_n18551_));
  INV_X1     g18359(.I(new_n18551_), .ZN(new_n18552_));
  OAI21_X1   g18360(.A1(new_n18077_), .A2(new_n18079_), .B(new_n18082_), .ZN(new_n18553_));
  NOR2_X1    g18361(.A1(new_n18424_), .A2(new_n18553_), .ZN(new_n18554_));
  XOR2_X1    g18362(.A1(new_n18554_), .A2(new_n17950_), .Z(new_n18555_));
  NAND3_X1   g18363(.A1(\asqrt[4] ), .A2(new_n18096_), .A3(new_n18078_), .ZN(new_n18556_));
  XOR2_X1    g18364(.A1(new_n18556_), .A2(new_n17954_), .Z(new_n18557_));
  AOI21_X1   g18365(.A1(new_n18056_), .A2(new_n18058_), .B(new_n18075_), .ZN(new_n18558_));
  NAND2_X1   g18366(.A1(\asqrt[4] ), .A2(new_n18558_), .ZN(new_n18559_));
  XOR2_X1    g18367(.A1(new_n18559_), .A2(new_n17957_), .Z(new_n18560_));
  INV_X1     g18368(.I(new_n18560_), .ZN(new_n18561_));
  NAND3_X1   g18369(.A1(\asqrt[4] ), .A2(new_n18055_), .A3(new_n18074_), .ZN(new_n18562_));
  XOR2_X1    g18370(.A1(new_n18562_), .A2(new_n18089_), .Z(new_n18563_));
  INV_X1     g18371(.I(new_n18563_), .ZN(new_n18564_));
  OAI21_X1   g18372(.A1(new_n18049_), .A2(new_n18051_), .B(new_n18054_), .ZN(new_n18565_));
  NOR2_X1    g18373(.A1(new_n18424_), .A2(new_n18565_), .ZN(new_n18566_));
  XOR2_X1    g18374(.A1(new_n18566_), .A2(new_n17962_), .Z(new_n18567_));
  NAND3_X1   g18375(.A1(\asqrt[4] ), .A2(new_n18068_), .A3(new_n18050_), .ZN(new_n18568_));
  XOR2_X1    g18376(.A1(new_n18568_), .A2(new_n17966_), .Z(new_n18569_));
  AOI21_X1   g18377(.A1(new_n18021_), .A2(new_n18023_), .B(new_n18047_), .ZN(new_n18570_));
  NAND2_X1   g18378(.A1(\asqrt[4] ), .A2(new_n18570_), .ZN(new_n18571_));
  XOR2_X1    g18379(.A1(new_n18571_), .A2(new_n17969_), .Z(new_n18572_));
  INV_X1     g18380(.I(new_n18572_), .ZN(new_n18573_));
  NAND3_X1   g18381(.A1(\asqrt[4] ), .A2(new_n18020_), .A3(new_n18046_), .ZN(new_n18574_));
  XOR2_X1    g18382(.A1(new_n18574_), .A2(new_n18061_), .Z(new_n18575_));
  INV_X1     g18383(.I(new_n18575_), .ZN(new_n18576_));
  OAI21_X1   g18384(.A1(new_n18014_), .A2(new_n18016_), .B(new_n18019_), .ZN(new_n18577_));
  NOR2_X1    g18385(.A1(new_n18424_), .A2(new_n18577_), .ZN(new_n18578_));
  XOR2_X1    g18386(.A1(new_n18578_), .A2(new_n17975_), .Z(new_n18579_));
  NAND3_X1   g18387(.A1(\asqrt[4] ), .A2(new_n18040_), .A3(new_n18015_), .ZN(new_n18580_));
  XOR2_X1    g18388(.A1(new_n18580_), .A2(new_n17978_), .Z(new_n18581_));
  OAI21_X1   g18389(.A1(new_n18035_), .A2(new_n18036_), .B(new_n18039_), .ZN(new_n18582_));
  NOR2_X1    g18390(.A1(new_n18424_), .A2(new_n18582_), .ZN(new_n18583_));
  XOR2_X1    g18391(.A1(new_n18583_), .A2(new_n17981_), .Z(new_n18584_));
  INV_X1     g18392(.I(new_n18584_), .ZN(new_n18585_));
  NAND2_X1   g18393(.A1(new_n18033_), .A2(new_n16093_), .ZN(new_n18586_));
  NAND3_X1   g18394(.A1(\asqrt[4] ), .A2(new_n18586_), .A3(new_n18011_), .ZN(new_n18587_));
  XOR2_X1    g18395(.A1(new_n18587_), .A2(new_n18034_), .Z(new_n18588_));
  INV_X1     g18396(.I(new_n18588_), .ZN(new_n18589_));
  NAND3_X1   g18397(.A1(\asqrt[4] ), .A2(new_n18031_), .A3(new_n18004_), .ZN(new_n18590_));
  XOR2_X1    g18398(.A1(new_n18590_), .A2(new_n17989_), .Z(new_n18591_));
  NAND4_X1   g18399(.A1(new_n18405_), .A2(\asqrt[5] ), .A3(new_n18407_), .A4(new_n18383_), .ZN(new_n18592_));
  INV_X1     g18400(.I(new_n18592_), .ZN(new_n18593_));
  NOR3_X1    g18401(.A1(new_n18424_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n18594_));
  OAI21_X1   g18402(.A1(new_n18594_), .A2(new_n18593_), .B(new_n17408_), .ZN(new_n18595_));
  INV_X1     g18403(.I(\a[8] ), .ZN(new_n18596_));
  INV_X1     g18404(.I(\a[9] ), .ZN(new_n18597_));
  NAND3_X1   g18405(.A1(\asqrt[4] ), .A2(new_n18596_), .A3(new_n18597_), .ZN(new_n18598_));
  NAND3_X1   g18406(.A1(new_n18598_), .A2(\a[10] ), .A3(new_n18592_), .ZN(new_n18599_));
  NAND2_X1   g18407(.A1(new_n18595_), .A2(new_n18599_), .ZN(new_n18600_));
  NOR3_X1    g18408(.A1(\a[6] ), .A2(\a[7] ), .A3(\a[8] ), .ZN(new_n18601_));
  AOI21_X1   g18409(.A1(\asqrt[4] ), .A2(\a[8] ), .B(new_n18601_), .ZN(new_n18602_));
  NOR2_X1    g18410(.A1(new_n18602_), .A2(new_n17816_), .ZN(new_n18603_));
  AOI21_X1   g18411(.A1(\asqrt[4] ), .A2(new_n18596_), .B(new_n18597_), .ZN(new_n18604_));
  NOR2_X1    g18412(.A1(new_n18594_), .A2(new_n18604_), .ZN(new_n18605_));
  NAND2_X1   g18413(.A1(new_n18602_), .A2(new_n17816_), .ZN(new_n18606_));
  AOI21_X1   g18414(.A1(new_n18605_), .A2(new_n18606_), .B(new_n18603_), .ZN(new_n18607_));
  AOI21_X1   g18415(.A1(new_n18607_), .A2(new_n17242_), .B(new_n18600_), .ZN(new_n18608_));
  NOR2_X1    g18416(.A1(new_n18607_), .A2(new_n17242_), .ZN(new_n18609_));
  NOR3_X1    g18417(.A1(new_n18608_), .A2(new_n18609_), .A3(\asqrt[7] ), .ZN(new_n18610_));
  NOR2_X1    g18418(.A1(new_n17996_), .A2(new_n17987_), .ZN(new_n18611_));
  NAND3_X1   g18419(.A1(\asqrt[4] ), .A2(new_n18027_), .A3(new_n18029_), .ZN(new_n18612_));
  XNOR2_X1   g18420(.A1(new_n18612_), .A2(new_n18611_), .ZN(new_n18613_));
  INV_X1     g18421(.I(new_n18613_), .ZN(new_n18614_));
  OAI21_X1   g18422(.A1(new_n18608_), .A2(new_n18609_), .B(\asqrt[7] ), .ZN(new_n18615_));
  OAI21_X1   g18423(.A1(new_n18610_), .A2(new_n18614_), .B(new_n18615_), .ZN(new_n18616_));
  OAI21_X1   g18424(.A1(new_n18616_), .A2(\asqrt[8] ), .B(new_n18591_), .ZN(new_n18617_));
  AOI21_X1   g18425(.A1(new_n18616_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n18618_));
  AOI21_X1   g18426(.A1(new_n18618_), .A2(new_n18617_), .B(new_n18589_), .ZN(new_n18619_));
  NAND2_X1   g18427(.A1(new_n18616_), .A2(\asqrt[8] ), .ZN(new_n18620_));
  AOI21_X1   g18428(.A1(new_n18617_), .A2(new_n18620_), .B(new_n15518_), .ZN(new_n18621_));
  NOR2_X1    g18429(.A1(new_n18619_), .A2(new_n18621_), .ZN(new_n18622_));
  AOI21_X1   g18430(.A1(new_n18622_), .A2(new_n14985_), .B(new_n18585_), .ZN(new_n18623_));
  OAI21_X1   g18431(.A1(new_n18619_), .A2(new_n18621_), .B(\asqrt[10] ), .ZN(new_n18624_));
  NAND2_X1   g18432(.A1(new_n18624_), .A2(new_n14430_), .ZN(new_n18625_));
  OAI21_X1   g18433(.A1(new_n18623_), .A2(new_n18625_), .B(new_n18581_), .ZN(new_n18626_));
  INV_X1     g18434(.I(new_n18624_), .ZN(new_n18627_));
  OAI21_X1   g18435(.A1(new_n18623_), .A2(new_n18627_), .B(\asqrt[11] ), .ZN(new_n18628_));
  NAND3_X1   g18436(.A1(new_n18626_), .A2(new_n18628_), .A3(new_n13917_), .ZN(new_n18629_));
  NAND2_X1   g18437(.A1(new_n18629_), .A2(new_n18579_), .ZN(new_n18630_));
  NAND2_X1   g18438(.A1(new_n18626_), .A2(new_n18628_), .ZN(new_n18631_));
  AOI21_X1   g18439(.A1(new_n18631_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n18632_));
  AOI21_X1   g18440(.A1(new_n18632_), .A2(new_n18630_), .B(new_n18576_), .ZN(new_n18633_));
  INV_X1     g18441(.I(new_n18581_), .ZN(new_n18634_));
  INV_X1     g18442(.I(new_n18591_), .ZN(new_n18635_));
  AOI21_X1   g18443(.A1(new_n18598_), .A2(new_n18592_), .B(\a[10] ), .ZN(new_n18636_));
  NOR3_X1    g18444(.A1(new_n18594_), .A2(new_n18593_), .A3(new_n17408_), .ZN(new_n18637_));
  NOR2_X1    g18445(.A1(new_n18637_), .A2(new_n18636_), .ZN(new_n18638_));
  NAND3_X1   g18446(.A1(new_n18420_), .A2(new_n18385_), .A3(new_n18387_), .ZN(new_n18639_));
  AOI21_X1   g18447(.A1(new_n18639_), .A2(new_n193_), .B(new_n18406_), .ZN(new_n18640_));
  AOI21_X1   g18448(.A1(new_n18640_), .A2(new_n18383_), .B(new_n18596_), .ZN(new_n18641_));
  OAI21_X1   g18449(.A1(new_n18641_), .A2(new_n18601_), .B(\asqrt[5] ), .ZN(new_n18642_));
  OAI21_X1   g18450(.A1(new_n18424_), .A2(\a[8] ), .B(\a[9] ), .ZN(new_n18643_));
  NAND2_X1   g18451(.A1(new_n18643_), .A2(new_n18598_), .ZN(new_n18644_));
  NOR3_X1    g18452(.A1(new_n18641_), .A2(\asqrt[5] ), .A3(new_n18601_), .ZN(new_n18645_));
  OAI21_X1   g18453(.A1(new_n18644_), .A2(new_n18645_), .B(new_n18642_), .ZN(new_n18646_));
  OAI21_X1   g18454(.A1(\asqrt[6] ), .A2(new_n18646_), .B(new_n18638_), .ZN(new_n18647_));
  NAND2_X1   g18455(.A1(new_n18646_), .A2(\asqrt[6] ), .ZN(new_n18648_));
  NAND3_X1   g18456(.A1(new_n18647_), .A2(new_n16649_), .A3(new_n18648_), .ZN(new_n18649_));
  AOI21_X1   g18457(.A1(new_n18647_), .A2(new_n18648_), .B(new_n16649_), .ZN(new_n18650_));
  AOI21_X1   g18458(.A1(new_n18649_), .A2(new_n18613_), .B(new_n18650_), .ZN(new_n18651_));
  AOI21_X1   g18459(.A1(new_n18651_), .A2(new_n16093_), .B(new_n18635_), .ZN(new_n18652_));
  OAI21_X1   g18460(.A1(new_n18651_), .A2(new_n16093_), .B(new_n15518_), .ZN(new_n18653_));
  OAI21_X1   g18461(.A1(new_n18652_), .A2(new_n18653_), .B(new_n18588_), .ZN(new_n18654_));
  NOR2_X1    g18462(.A1(new_n18651_), .A2(new_n16093_), .ZN(new_n18655_));
  OAI21_X1   g18463(.A1(new_n18652_), .A2(new_n18655_), .B(\asqrt[9] ), .ZN(new_n18656_));
  NAND3_X1   g18464(.A1(new_n18654_), .A2(new_n18656_), .A3(new_n14985_), .ZN(new_n18657_));
  NAND2_X1   g18465(.A1(new_n18657_), .A2(new_n18584_), .ZN(new_n18658_));
  NAND2_X1   g18466(.A1(new_n18654_), .A2(new_n18656_), .ZN(new_n18659_));
  AOI21_X1   g18467(.A1(new_n18659_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n18660_));
  AOI21_X1   g18468(.A1(new_n18660_), .A2(new_n18658_), .B(new_n18634_), .ZN(new_n18661_));
  AOI21_X1   g18469(.A1(new_n18658_), .A2(new_n18624_), .B(new_n14430_), .ZN(new_n18662_));
  OAI21_X1   g18470(.A1(new_n18661_), .A2(new_n18662_), .B(\asqrt[12] ), .ZN(new_n18663_));
  AOI21_X1   g18471(.A1(new_n18630_), .A2(new_n18663_), .B(new_n13382_), .ZN(new_n18664_));
  NOR2_X1    g18472(.A1(new_n18633_), .A2(new_n18664_), .ZN(new_n18665_));
  AOI21_X1   g18473(.A1(new_n18665_), .A2(new_n12889_), .B(new_n18573_), .ZN(new_n18666_));
  OAI21_X1   g18474(.A1(new_n18633_), .A2(new_n18664_), .B(\asqrt[14] ), .ZN(new_n18667_));
  NAND2_X1   g18475(.A1(new_n18667_), .A2(new_n12374_), .ZN(new_n18668_));
  OAI21_X1   g18476(.A1(new_n18666_), .A2(new_n18668_), .B(new_n18569_), .ZN(new_n18669_));
  INV_X1     g18477(.I(new_n18667_), .ZN(new_n18670_));
  OAI21_X1   g18478(.A1(new_n18666_), .A2(new_n18670_), .B(\asqrt[15] ), .ZN(new_n18671_));
  NAND3_X1   g18479(.A1(new_n18669_), .A2(new_n18671_), .A3(new_n11901_), .ZN(new_n18672_));
  NAND2_X1   g18480(.A1(new_n18672_), .A2(new_n18567_), .ZN(new_n18673_));
  NAND2_X1   g18481(.A1(new_n18669_), .A2(new_n18671_), .ZN(new_n18674_));
  AOI21_X1   g18482(.A1(new_n18674_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n18675_));
  AOI21_X1   g18483(.A1(new_n18675_), .A2(new_n18673_), .B(new_n18564_), .ZN(new_n18676_));
  INV_X1     g18484(.I(new_n18569_), .ZN(new_n18677_));
  INV_X1     g18485(.I(new_n18579_), .ZN(new_n18678_));
  NOR2_X1    g18486(.A1(new_n18661_), .A2(new_n18662_), .ZN(new_n18679_));
  AOI21_X1   g18487(.A1(new_n18679_), .A2(new_n13917_), .B(new_n18678_), .ZN(new_n18680_));
  NAND2_X1   g18488(.A1(new_n18663_), .A2(new_n13382_), .ZN(new_n18681_));
  OAI21_X1   g18489(.A1(new_n18680_), .A2(new_n18681_), .B(new_n18575_), .ZN(new_n18682_));
  INV_X1     g18490(.I(new_n18663_), .ZN(new_n18683_));
  OAI21_X1   g18491(.A1(new_n18680_), .A2(new_n18683_), .B(\asqrt[13] ), .ZN(new_n18684_));
  NAND3_X1   g18492(.A1(new_n18682_), .A2(new_n18684_), .A3(new_n12889_), .ZN(new_n18685_));
  NAND2_X1   g18493(.A1(new_n18685_), .A2(new_n18572_), .ZN(new_n18686_));
  NAND2_X1   g18494(.A1(new_n18682_), .A2(new_n18684_), .ZN(new_n18687_));
  AOI21_X1   g18495(.A1(new_n18687_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n18688_));
  AOI21_X1   g18496(.A1(new_n18688_), .A2(new_n18686_), .B(new_n18677_), .ZN(new_n18689_));
  AOI21_X1   g18497(.A1(new_n18686_), .A2(new_n18667_), .B(new_n12374_), .ZN(new_n18690_));
  OAI21_X1   g18498(.A1(new_n18689_), .A2(new_n18690_), .B(\asqrt[16] ), .ZN(new_n18691_));
  AOI21_X1   g18499(.A1(new_n18673_), .A2(new_n18691_), .B(new_n11406_), .ZN(new_n18692_));
  NOR2_X1    g18500(.A1(new_n18676_), .A2(new_n18692_), .ZN(new_n18693_));
  AOI21_X1   g18501(.A1(new_n18693_), .A2(new_n10953_), .B(new_n18561_), .ZN(new_n18694_));
  OAI21_X1   g18502(.A1(new_n18676_), .A2(new_n18692_), .B(\asqrt[18] ), .ZN(new_n18695_));
  NAND2_X1   g18503(.A1(new_n18695_), .A2(new_n10478_), .ZN(new_n18696_));
  OAI21_X1   g18504(.A1(new_n18694_), .A2(new_n18696_), .B(new_n18557_), .ZN(new_n18697_));
  INV_X1     g18505(.I(new_n18695_), .ZN(new_n18698_));
  OAI21_X1   g18506(.A1(new_n18694_), .A2(new_n18698_), .B(\asqrt[19] ), .ZN(new_n18699_));
  NAND3_X1   g18507(.A1(new_n18697_), .A2(new_n18699_), .A3(new_n10045_), .ZN(new_n18700_));
  NAND2_X1   g18508(.A1(new_n18700_), .A2(new_n18555_), .ZN(new_n18701_));
  NAND2_X1   g18509(.A1(new_n18697_), .A2(new_n18699_), .ZN(new_n18702_));
  AOI21_X1   g18510(.A1(new_n18702_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n18703_));
  AOI21_X1   g18511(.A1(new_n18703_), .A2(new_n18701_), .B(new_n18552_), .ZN(new_n18704_));
  INV_X1     g18512(.I(new_n18557_), .ZN(new_n18705_));
  INV_X1     g18513(.I(new_n18567_), .ZN(new_n18706_));
  NOR2_X1    g18514(.A1(new_n18689_), .A2(new_n18690_), .ZN(new_n18707_));
  AOI21_X1   g18515(.A1(new_n18707_), .A2(new_n11901_), .B(new_n18706_), .ZN(new_n18708_));
  NAND2_X1   g18516(.A1(new_n18691_), .A2(new_n11406_), .ZN(new_n18709_));
  OAI21_X1   g18517(.A1(new_n18708_), .A2(new_n18709_), .B(new_n18563_), .ZN(new_n18710_));
  INV_X1     g18518(.I(new_n18691_), .ZN(new_n18711_));
  OAI21_X1   g18519(.A1(new_n18708_), .A2(new_n18711_), .B(\asqrt[17] ), .ZN(new_n18712_));
  NAND3_X1   g18520(.A1(new_n18710_), .A2(new_n18712_), .A3(new_n10953_), .ZN(new_n18713_));
  NAND2_X1   g18521(.A1(new_n18713_), .A2(new_n18560_), .ZN(new_n18714_));
  NAND2_X1   g18522(.A1(new_n18710_), .A2(new_n18712_), .ZN(new_n18715_));
  AOI21_X1   g18523(.A1(new_n18715_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n18716_));
  AOI21_X1   g18524(.A1(new_n18716_), .A2(new_n18714_), .B(new_n18705_), .ZN(new_n18717_));
  AOI21_X1   g18525(.A1(new_n18714_), .A2(new_n18695_), .B(new_n10478_), .ZN(new_n18718_));
  OAI21_X1   g18526(.A1(new_n18717_), .A2(new_n18718_), .B(\asqrt[20] ), .ZN(new_n18719_));
  AOI21_X1   g18527(.A1(new_n18701_), .A2(new_n18719_), .B(new_n9590_), .ZN(new_n18720_));
  NOR2_X1    g18528(.A1(new_n18704_), .A2(new_n18720_), .ZN(new_n18721_));
  AOI21_X1   g18529(.A1(new_n18721_), .A2(new_n9177_), .B(new_n18549_), .ZN(new_n18722_));
  OAI21_X1   g18530(.A1(new_n18704_), .A2(new_n18720_), .B(\asqrt[22] ), .ZN(new_n18723_));
  NAND2_X1   g18531(.A1(new_n18723_), .A2(new_n8742_), .ZN(new_n18724_));
  OAI21_X1   g18532(.A1(new_n18722_), .A2(new_n18724_), .B(new_n18545_), .ZN(new_n18725_));
  INV_X1     g18533(.I(new_n18723_), .ZN(new_n18726_));
  OAI21_X1   g18534(.A1(new_n18722_), .A2(new_n18726_), .B(\asqrt[23] ), .ZN(new_n18727_));
  NAND3_X1   g18535(.A1(new_n18725_), .A2(new_n18727_), .A3(new_n8349_), .ZN(new_n18728_));
  NAND2_X1   g18536(.A1(new_n18728_), .A2(new_n18543_), .ZN(new_n18729_));
  NAND2_X1   g18537(.A1(new_n18725_), .A2(new_n18727_), .ZN(new_n18730_));
  AOI21_X1   g18538(.A1(new_n18730_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n18731_));
  AOI21_X1   g18539(.A1(new_n18731_), .A2(new_n18729_), .B(new_n18540_), .ZN(new_n18732_));
  INV_X1     g18540(.I(new_n18545_), .ZN(new_n18733_));
  INV_X1     g18541(.I(new_n18555_), .ZN(new_n18734_));
  NOR2_X1    g18542(.A1(new_n18717_), .A2(new_n18718_), .ZN(new_n18735_));
  AOI21_X1   g18543(.A1(new_n18735_), .A2(new_n10045_), .B(new_n18734_), .ZN(new_n18736_));
  NAND2_X1   g18544(.A1(new_n18719_), .A2(new_n9590_), .ZN(new_n18737_));
  OAI21_X1   g18545(.A1(new_n18736_), .A2(new_n18737_), .B(new_n18551_), .ZN(new_n18738_));
  INV_X1     g18546(.I(new_n18719_), .ZN(new_n18739_));
  OAI21_X1   g18547(.A1(new_n18736_), .A2(new_n18739_), .B(\asqrt[21] ), .ZN(new_n18740_));
  NAND3_X1   g18548(.A1(new_n18738_), .A2(new_n18740_), .A3(new_n9177_), .ZN(new_n18741_));
  NAND2_X1   g18549(.A1(new_n18741_), .A2(new_n18548_), .ZN(new_n18742_));
  NAND2_X1   g18550(.A1(new_n18738_), .A2(new_n18740_), .ZN(new_n18743_));
  AOI21_X1   g18551(.A1(new_n18743_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n18744_));
  AOI21_X1   g18552(.A1(new_n18744_), .A2(new_n18742_), .B(new_n18733_), .ZN(new_n18745_));
  AOI21_X1   g18553(.A1(new_n18742_), .A2(new_n18723_), .B(new_n8742_), .ZN(new_n18746_));
  OAI21_X1   g18554(.A1(new_n18745_), .A2(new_n18746_), .B(\asqrt[24] ), .ZN(new_n18747_));
  AOI21_X1   g18555(.A1(new_n18729_), .A2(new_n18747_), .B(new_n7934_), .ZN(new_n18748_));
  NOR2_X1    g18556(.A1(new_n18732_), .A2(new_n18748_), .ZN(new_n18749_));
  AOI21_X1   g18557(.A1(new_n18749_), .A2(new_n7561_), .B(new_n18537_), .ZN(new_n18750_));
  OAI21_X1   g18558(.A1(new_n18732_), .A2(new_n18748_), .B(\asqrt[26] ), .ZN(new_n18751_));
  NAND2_X1   g18559(.A1(new_n18751_), .A2(new_n7166_), .ZN(new_n18752_));
  OAI21_X1   g18560(.A1(new_n18750_), .A2(new_n18752_), .B(new_n18533_), .ZN(new_n18753_));
  INV_X1     g18561(.I(new_n18751_), .ZN(new_n18754_));
  OAI21_X1   g18562(.A1(new_n18750_), .A2(new_n18754_), .B(\asqrt[27] ), .ZN(new_n18755_));
  NAND3_X1   g18563(.A1(new_n18753_), .A2(new_n18755_), .A3(new_n6813_), .ZN(new_n18756_));
  NAND2_X1   g18564(.A1(new_n18756_), .A2(new_n18531_), .ZN(new_n18757_));
  NAND2_X1   g18565(.A1(new_n18753_), .A2(new_n18755_), .ZN(new_n18758_));
  AOI21_X1   g18566(.A1(new_n18758_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n18759_));
  AOI21_X1   g18567(.A1(new_n18759_), .A2(new_n18757_), .B(new_n18528_), .ZN(new_n18760_));
  INV_X1     g18568(.I(new_n18533_), .ZN(new_n18761_));
  INV_X1     g18569(.I(new_n18543_), .ZN(new_n18762_));
  NOR2_X1    g18570(.A1(new_n18745_), .A2(new_n18746_), .ZN(new_n18763_));
  AOI21_X1   g18571(.A1(new_n18763_), .A2(new_n8349_), .B(new_n18762_), .ZN(new_n18764_));
  NAND2_X1   g18572(.A1(new_n18747_), .A2(new_n7934_), .ZN(new_n18765_));
  OAI21_X1   g18573(.A1(new_n18764_), .A2(new_n18765_), .B(new_n18539_), .ZN(new_n18766_));
  INV_X1     g18574(.I(new_n18747_), .ZN(new_n18767_));
  OAI21_X1   g18575(.A1(new_n18764_), .A2(new_n18767_), .B(\asqrt[25] ), .ZN(new_n18768_));
  NAND3_X1   g18576(.A1(new_n18766_), .A2(new_n18768_), .A3(new_n7561_), .ZN(new_n18769_));
  NAND2_X1   g18577(.A1(new_n18769_), .A2(new_n18536_), .ZN(new_n18770_));
  NAND2_X1   g18578(.A1(new_n18766_), .A2(new_n18768_), .ZN(new_n18771_));
  AOI21_X1   g18579(.A1(new_n18771_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n18772_));
  AOI21_X1   g18580(.A1(new_n18772_), .A2(new_n18770_), .B(new_n18761_), .ZN(new_n18773_));
  AOI21_X1   g18581(.A1(new_n18770_), .A2(new_n18751_), .B(new_n7166_), .ZN(new_n18774_));
  OAI21_X1   g18582(.A1(new_n18773_), .A2(new_n18774_), .B(\asqrt[28] ), .ZN(new_n18775_));
  AOI21_X1   g18583(.A1(new_n18757_), .A2(new_n18775_), .B(new_n6454_), .ZN(new_n18776_));
  NOR2_X1    g18584(.A1(new_n18760_), .A2(new_n18776_), .ZN(new_n18777_));
  AOI21_X1   g18585(.A1(new_n18777_), .A2(new_n6106_), .B(new_n18525_), .ZN(new_n18778_));
  OAI21_X1   g18586(.A1(new_n18760_), .A2(new_n18776_), .B(\asqrt[30] ), .ZN(new_n18779_));
  NAND2_X1   g18587(.A1(new_n18779_), .A2(new_n5750_), .ZN(new_n18780_));
  OAI21_X1   g18588(.A1(new_n18778_), .A2(new_n18780_), .B(new_n18521_), .ZN(new_n18781_));
  INV_X1     g18589(.I(new_n18779_), .ZN(new_n18782_));
  OAI21_X1   g18590(.A1(new_n18778_), .A2(new_n18782_), .B(\asqrt[31] ), .ZN(new_n18783_));
  NAND3_X1   g18591(.A1(new_n18781_), .A2(new_n18783_), .A3(new_n5435_), .ZN(new_n18784_));
  NAND2_X1   g18592(.A1(new_n18784_), .A2(new_n18519_), .ZN(new_n18785_));
  NAND2_X1   g18593(.A1(new_n18781_), .A2(new_n18783_), .ZN(new_n18786_));
  AOI21_X1   g18594(.A1(new_n18786_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n18787_));
  AOI21_X1   g18595(.A1(new_n18787_), .A2(new_n18785_), .B(new_n18516_), .ZN(new_n18788_));
  INV_X1     g18596(.I(new_n18521_), .ZN(new_n18789_));
  INV_X1     g18597(.I(new_n18531_), .ZN(new_n18790_));
  NOR2_X1    g18598(.A1(new_n18773_), .A2(new_n18774_), .ZN(new_n18791_));
  AOI21_X1   g18599(.A1(new_n18791_), .A2(new_n6813_), .B(new_n18790_), .ZN(new_n18792_));
  NAND2_X1   g18600(.A1(new_n18775_), .A2(new_n6454_), .ZN(new_n18793_));
  OAI21_X1   g18601(.A1(new_n18792_), .A2(new_n18793_), .B(new_n18527_), .ZN(new_n18794_));
  INV_X1     g18602(.I(new_n18775_), .ZN(new_n18795_));
  OAI21_X1   g18603(.A1(new_n18792_), .A2(new_n18795_), .B(\asqrt[29] ), .ZN(new_n18796_));
  NAND3_X1   g18604(.A1(new_n18794_), .A2(new_n18796_), .A3(new_n6106_), .ZN(new_n18797_));
  NAND2_X1   g18605(.A1(new_n18797_), .A2(new_n18524_), .ZN(new_n18798_));
  NAND2_X1   g18606(.A1(new_n18794_), .A2(new_n18796_), .ZN(new_n18799_));
  AOI21_X1   g18607(.A1(new_n18799_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n18800_));
  AOI21_X1   g18608(.A1(new_n18800_), .A2(new_n18798_), .B(new_n18789_), .ZN(new_n18801_));
  AOI21_X1   g18609(.A1(new_n18798_), .A2(new_n18779_), .B(new_n5750_), .ZN(new_n18802_));
  OAI21_X1   g18610(.A1(new_n18801_), .A2(new_n18802_), .B(\asqrt[32] ), .ZN(new_n18803_));
  AOI21_X1   g18611(.A1(new_n18785_), .A2(new_n18803_), .B(new_n5110_), .ZN(new_n18804_));
  NOR2_X1    g18612(.A1(new_n18788_), .A2(new_n18804_), .ZN(new_n18805_));
  AOI21_X1   g18613(.A1(new_n18805_), .A2(new_n4810_), .B(new_n18513_), .ZN(new_n18806_));
  OAI21_X1   g18614(.A1(new_n18788_), .A2(new_n18804_), .B(\asqrt[34] ), .ZN(new_n18807_));
  NAND2_X1   g18615(.A1(new_n18807_), .A2(new_n4510_), .ZN(new_n18808_));
  OAI21_X1   g18616(.A1(new_n18806_), .A2(new_n18808_), .B(new_n18509_), .ZN(new_n18809_));
  INV_X1     g18617(.I(new_n18807_), .ZN(new_n18810_));
  OAI21_X1   g18618(.A1(new_n18806_), .A2(new_n18810_), .B(\asqrt[35] ), .ZN(new_n18811_));
  NAND3_X1   g18619(.A1(new_n18809_), .A2(new_n18811_), .A3(new_n4224_), .ZN(new_n18812_));
  NAND2_X1   g18620(.A1(new_n18812_), .A2(new_n18507_), .ZN(new_n18813_));
  NAND2_X1   g18621(.A1(new_n18809_), .A2(new_n18811_), .ZN(new_n18814_));
  AOI21_X1   g18622(.A1(new_n18814_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n18815_));
  AOI21_X1   g18623(.A1(new_n18815_), .A2(new_n18813_), .B(new_n18504_), .ZN(new_n18816_));
  INV_X1     g18624(.I(new_n18509_), .ZN(new_n18817_));
  INV_X1     g18625(.I(new_n18519_), .ZN(new_n18818_));
  NOR2_X1    g18626(.A1(new_n18801_), .A2(new_n18802_), .ZN(new_n18819_));
  AOI21_X1   g18627(.A1(new_n18819_), .A2(new_n5435_), .B(new_n18818_), .ZN(new_n18820_));
  NAND2_X1   g18628(.A1(new_n18803_), .A2(new_n5110_), .ZN(new_n18821_));
  OAI21_X1   g18629(.A1(new_n18820_), .A2(new_n18821_), .B(new_n18515_), .ZN(new_n18822_));
  INV_X1     g18630(.I(new_n18803_), .ZN(new_n18823_));
  OAI21_X1   g18631(.A1(new_n18820_), .A2(new_n18823_), .B(\asqrt[33] ), .ZN(new_n18824_));
  NAND3_X1   g18632(.A1(new_n18822_), .A2(new_n18824_), .A3(new_n4810_), .ZN(new_n18825_));
  NAND2_X1   g18633(.A1(new_n18825_), .A2(new_n18512_), .ZN(new_n18826_));
  NAND2_X1   g18634(.A1(new_n18822_), .A2(new_n18824_), .ZN(new_n18827_));
  AOI21_X1   g18635(.A1(new_n18827_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n18828_));
  AOI21_X1   g18636(.A1(new_n18828_), .A2(new_n18826_), .B(new_n18817_), .ZN(new_n18829_));
  AOI21_X1   g18637(.A1(new_n18826_), .A2(new_n18807_), .B(new_n4510_), .ZN(new_n18830_));
  OAI21_X1   g18638(.A1(new_n18829_), .A2(new_n18830_), .B(\asqrt[36] ), .ZN(new_n18831_));
  AOI21_X1   g18639(.A1(new_n18813_), .A2(new_n18831_), .B(new_n3928_), .ZN(new_n18832_));
  NOR2_X1    g18640(.A1(new_n18816_), .A2(new_n18832_), .ZN(new_n18833_));
  AOI21_X1   g18641(.A1(new_n18833_), .A2(new_n3675_), .B(new_n18501_), .ZN(new_n18834_));
  OAI21_X1   g18642(.A1(new_n18816_), .A2(new_n18832_), .B(\asqrt[38] ), .ZN(new_n18835_));
  NAND2_X1   g18643(.A1(new_n18835_), .A2(new_n3400_), .ZN(new_n18836_));
  OAI21_X1   g18644(.A1(new_n18834_), .A2(new_n18836_), .B(new_n18497_), .ZN(new_n18837_));
  INV_X1     g18645(.I(new_n18835_), .ZN(new_n18838_));
  OAI21_X1   g18646(.A1(new_n18834_), .A2(new_n18838_), .B(\asqrt[39] ), .ZN(new_n18839_));
  NAND3_X1   g18647(.A1(new_n18837_), .A2(new_n18839_), .A3(new_n3167_), .ZN(new_n18840_));
  NAND2_X1   g18648(.A1(new_n18840_), .A2(new_n18495_), .ZN(new_n18841_));
  NAND2_X1   g18649(.A1(new_n18837_), .A2(new_n18839_), .ZN(new_n18842_));
  AOI21_X1   g18650(.A1(new_n18842_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n18843_));
  AOI21_X1   g18651(.A1(new_n18843_), .A2(new_n18841_), .B(new_n18492_), .ZN(new_n18844_));
  INV_X1     g18652(.I(new_n18497_), .ZN(new_n18845_));
  INV_X1     g18653(.I(new_n18507_), .ZN(new_n18846_));
  NOR2_X1    g18654(.A1(new_n18829_), .A2(new_n18830_), .ZN(new_n18847_));
  AOI21_X1   g18655(.A1(new_n18847_), .A2(new_n4224_), .B(new_n18846_), .ZN(new_n18848_));
  NAND2_X1   g18656(.A1(new_n18831_), .A2(new_n3928_), .ZN(new_n18849_));
  OAI21_X1   g18657(.A1(new_n18848_), .A2(new_n18849_), .B(new_n18503_), .ZN(new_n18850_));
  INV_X1     g18658(.I(new_n18831_), .ZN(new_n18851_));
  OAI21_X1   g18659(.A1(new_n18848_), .A2(new_n18851_), .B(\asqrt[37] ), .ZN(new_n18852_));
  NAND3_X1   g18660(.A1(new_n18850_), .A2(new_n18852_), .A3(new_n3675_), .ZN(new_n18853_));
  NAND2_X1   g18661(.A1(new_n18853_), .A2(new_n18500_), .ZN(new_n18854_));
  NAND2_X1   g18662(.A1(new_n18850_), .A2(new_n18852_), .ZN(new_n18855_));
  AOI21_X1   g18663(.A1(new_n18855_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n18856_));
  AOI21_X1   g18664(.A1(new_n18856_), .A2(new_n18854_), .B(new_n18845_), .ZN(new_n18857_));
  AOI21_X1   g18665(.A1(new_n18854_), .A2(new_n18835_), .B(new_n3400_), .ZN(new_n18858_));
  OAI21_X1   g18666(.A1(new_n18857_), .A2(new_n18858_), .B(\asqrt[40] ), .ZN(new_n18859_));
  AOI21_X1   g18667(.A1(new_n18841_), .A2(new_n18859_), .B(new_n2912_), .ZN(new_n18860_));
  NOR2_X1    g18668(.A1(new_n18844_), .A2(new_n18860_), .ZN(new_n18861_));
  AOI21_X1   g18669(.A1(new_n18861_), .A2(new_n2699_), .B(new_n18489_), .ZN(new_n18862_));
  OAI21_X1   g18670(.A1(new_n18844_), .A2(new_n18860_), .B(\asqrt[42] ), .ZN(new_n18863_));
  NAND2_X1   g18671(.A1(new_n18863_), .A2(new_n2464_), .ZN(new_n18864_));
  OAI21_X1   g18672(.A1(new_n18862_), .A2(new_n18864_), .B(new_n18485_), .ZN(new_n18865_));
  INV_X1     g18673(.I(new_n18863_), .ZN(new_n18866_));
  OAI21_X1   g18674(.A1(new_n18862_), .A2(new_n18866_), .B(\asqrt[43] ), .ZN(new_n18867_));
  NAND3_X1   g18675(.A1(new_n18865_), .A2(new_n18867_), .A3(new_n2271_), .ZN(new_n18868_));
  NAND2_X1   g18676(.A1(new_n18868_), .A2(new_n18483_), .ZN(new_n18869_));
  NAND2_X1   g18677(.A1(new_n18865_), .A2(new_n18867_), .ZN(new_n18870_));
  AOI21_X1   g18678(.A1(new_n18870_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n18871_));
  AOI21_X1   g18679(.A1(new_n18871_), .A2(new_n18869_), .B(new_n18480_), .ZN(new_n18872_));
  INV_X1     g18680(.I(new_n18485_), .ZN(new_n18873_));
  INV_X1     g18681(.I(new_n18495_), .ZN(new_n18874_));
  NOR2_X1    g18682(.A1(new_n18857_), .A2(new_n18858_), .ZN(new_n18875_));
  AOI21_X1   g18683(.A1(new_n18875_), .A2(new_n3167_), .B(new_n18874_), .ZN(new_n18876_));
  NAND2_X1   g18684(.A1(new_n18859_), .A2(new_n2912_), .ZN(new_n18877_));
  OAI21_X1   g18685(.A1(new_n18876_), .A2(new_n18877_), .B(new_n18491_), .ZN(new_n18878_));
  INV_X1     g18686(.I(new_n18859_), .ZN(new_n18879_));
  OAI21_X1   g18687(.A1(new_n18876_), .A2(new_n18879_), .B(\asqrt[41] ), .ZN(new_n18880_));
  NAND3_X1   g18688(.A1(new_n18878_), .A2(new_n18880_), .A3(new_n2699_), .ZN(new_n18881_));
  NAND2_X1   g18689(.A1(new_n18881_), .A2(new_n18488_), .ZN(new_n18882_));
  NAND2_X1   g18690(.A1(new_n18878_), .A2(new_n18880_), .ZN(new_n18883_));
  AOI21_X1   g18691(.A1(new_n18883_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n18884_));
  AOI21_X1   g18692(.A1(new_n18884_), .A2(new_n18882_), .B(new_n18873_), .ZN(new_n18885_));
  AOI21_X1   g18693(.A1(new_n18882_), .A2(new_n18863_), .B(new_n2464_), .ZN(new_n18886_));
  OAI21_X1   g18694(.A1(new_n18885_), .A2(new_n18886_), .B(\asqrt[44] ), .ZN(new_n18887_));
  AOI21_X1   g18695(.A1(new_n18869_), .A2(new_n18887_), .B(new_n2072_), .ZN(new_n18888_));
  NOR2_X1    g18696(.A1(new_n18872_), .A2(new_n18888_), .ZN(new_n18889_));
  AOI21_X1   g18697(.A1(new_n18889_), .A2(new_n1884_), .B(new_n18477_), .ZN(new_n18890_));
  OAI21_X1   g18698(.A1(new_n18872_), .A2(new_n18888_), .B(\asqrt[46] ), .ZN(new_n18891_));
  NAND2_X1   g18699(.A1(new_n18891_), .A2(new_n1688_), .ZN(new_n18892_));
  OAI21_X1   g18700(.A1(new_n18890_), .A2(new_n18892_), .B(new_n18473_), .ZN(new_n18893_));
  INV_X1     g18701(.I(new_n18891_), .ZN(new_n18894_));
  OAI21_X1   g18702(.A1(new_n18890_), .A2(new_n18894_), .B(\asqrt[47] ), .ZN(new_n18895_));
  NAND3_X1   g18703(.A1(new_n18893_), .A2(new_n18895_), .A3(new_n1533_), .ZN(new_n18896_));
  NAND2_X1   g18704(.A1(new_n18896_), .A2(new_n18471_), .ZN(new_n18897_));
  NAND2_X1   g18705(.A1(new_n18893_), .A2(new_n18895_), .ZN(new_n18898_));
  AOI21_X1   g18706(.A1(new_n18898_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n18899_));
  AOI21_X1   g18707(.A1(new_n18899_), .A2(new_n18897_), .B(new_n18468_), .ZN(new_n18900_));
  INV_X1     g18708(.I(new_n18473_), .ZN(new_n18901_));
  INV_X1     g18709(.I(new_n18483_), .ZN(new_n18902_));
  NOR2_X1    g18710(.A1(new_n18885_), .A2(new_n18886_), .ZN(new_n18903_));
  AOI21_X1   g18711(.A1(new_n18903_), .A2(new_n2271_), .B(new_n18902_), .ZN(new_n18904_));
  NAND2_X1   g18712(.A1(new_n18887_), .A2(new_n2072_), .ZN(new_n18905_));
  OAI21_X1   g18713(.A1(new_n18904_), .A2(new_n18905_), .B(new_n18479_), .ZN(new_n18906_));
  INV_X1     g18714(.I(new_n18887_), .ZN(new_n18907_));
  OAI21_X1   g18715(.A1(new_n18904_), .A2(new_n18907_), .B(\asqrt[45] ), .ZN(new_n18908_));
  NAND3_X1   g18716(.A1(new_n18906_), .A2(new_n18908_), .A3(new_n1884_), .ZN(new_n18909_));
  NAND2_X1   g18717(.A1(new_n18909_), .A2(new_n18476_), .ZN(new_n18910_));
  NAND2_X1   g18718(.A1(new_n18906_), .A2(new_n18908_), .ZN(new_n18911_));
  AOI21_X1   g18719(.A1(new_n18911_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n18912_));
  AOI21_X1   g18720(.A1(new_n18912_), .A2(new_n18910_), .B(new_n18901_), .ZN(new_n18913_));
  AOI21_X1   g18721(.A1(new_n18910_), .A2(new_n18891_), .B(new_n1688_), .ZN(new_n18914_));
  OAI21_X1   g18722(.A1(new_n18913_), .A2(new_n18914_), .B(\asqrt[48] ), .ZN(new_n18915_));
  AOI21_X1   g18723(.A1(new_n18897_), .A2(new_n18915_), .B(new_n1368_), .ZN(new_n18916_));
  NOR2_X1    g18724(.A1(new_n18900_), .A2(new_n18916_), .ZN(new_n18917_));
  AOI21_X1   g18725(.A1(new_n18917_), .A2(new_n1228_), .B(new_n18465_), .ZN(new_n18918_));
  OAI21_X1   g18726(.A1(new_n18900_), .A2(new_n18916_), .B(\asqrt[50] ), .ZN(new_n18919_));
  NAND2_X1   g18727(.A1(new_n18919_), .A2(new_n1088_), .ZN(new_n18920_));
  OAI21_X1   g18728(.A1(new_n18918_), .A2(new_n18920_), .B(new_n18461_), .ZN(new_n18921_));
  INV_X1     g18729(.I(new_n18919_), .ZN(new_n18922_));
  OAI21_X1   g18730(.A1(new_n18918_), .A2(new_n18922_), .B(\asqrt[51] ), .ZN(new_n18923_));
  NAND3_X1   g18731(.A1(new_n18921_), .A2(new_n18923_), .A3(new_n962_), .ZN(new_n18924_));
  NAND2_X1   g18732(.A1(new_n18924_), .A2(new_n18459_), .ZN(new_n18925_));
  NAND2_X1   g18733(.A1(new_n18921_), .A2(new_n18923_), .ZN(new_n18926_));
  AOI21_X1   g18734(.A1(new_n18926_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n18927_));
  AOI21_X1   g18735(.A1(new_n18927_), .A2(new_n18925_), .B(new_n18456_), .ZN(new_n18928_));
  INV_X1     g18736(.I(new_n18461_), .ZN(new_n18929_));
  INV_X1     g18737(.I(new_n18471_), .ZN(new_n18930_));
  NOR2_X1    g18738(.A1(new_n18913_), .A2(new_n18914_), .ZN(new_n18931_));
  AOI21_X1   g18739(.A1(new_n18931_), .A2(new_n1533_), .B(new_n18930_), .ZN(new_n18932_));
  NAND2_X1   g18740(.A1(new_n18915_), .A2(new_n1368_), .ZN(new_n18933_));
  OAI21_X1   g18741(.A1(new_n18932_), .A2(new_n18933_), .B(new_n18467_), .ZN(new_n18934_));
  INV_X1     g18742(.I(new_n18915_), .ZN(new_n18935_));
  OAI21_X1   g18743(.A1(new_n18932_), .A2(new_n18935_), .B(\asqrt[49] ), .ZN(new_n18936_));
  NAND3_X1   g18744(.A1(new_n18934_), .A2(new_n18936_), .A3(new_n1228_), .ZN(new_n18937_));
  NAND2_X1   g18745(.A1(new_n18937_), .A2(new_n18464_), .ZN(new_n18938_));
  NAND2_X1   g18746(.A1(new_n18934_), .A2(new_n18936_), .ZN(new_n18939_));
  AOI21_X1   g18747(.A1(new_n18939_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n18940_));
  AOI21_X1   g18748(.A1(new_n18940_), .A2(new_n18938_), .B(new_n18929_), .ZN(new_n18941_));
  AOI21_X1   g18749(.A1(new_n18938_), .A2(new_n18919_), .B(new_n1088_), .ZN(new_n18942_));
  OAI21_X1   g18750(.A1(new_n18941_), .A2(new_n18942_), .B(\asqrt[52] ), .ZN(new_n18943_));
  AOI21_X1   g18751(.A1(new_n18925_), .A2(new_n18943_), .B(new_n842_), .ZN(new_n18944_));
  NOR2_X1    g18752(.A1(new_n18928_), .A2(new_n18944_), .ZN(new_n18945_));
  AOI21_X1   g18753(.A1(new_n18945_), .A2(new_n720_), .B(new_n18453_), .ZN(new_n18946_));
  OAI21_X1   g18754(.A1(new_n18928_), .A2(new_n18944_), .B(\asqrt[54] ), .ZN(new_n18947_));
  NAND2_X1   g18755(.A1(new_n18947_), .A2(new_n630_), .ZN(new_n18948_));
  OAI21_X1   g18756(.A1(new_n18946_), .A2(new_n18948_), .B(new_n18449_), .ZN(new_n18949_));
  INV_X1     g18757(.I(new_n18947_), .ZN(new_n18950_));
  OAI21_X1   g18758(.A1(new_n18946_), .A2(new_n18950_), .B(\asqrt[55] ), .ZN(new_n18951_));
  NAND3_X1   g18759(.A1(new_n18949_), .A2(new_n18951_), .A3(new_n545_), .ZN(new_n18952_));
  NAND2_X1   g18760(.A1(new_n18952_), .A2(new_n18447_), .ZN(new_n18953_));
  NAND2_X1   g18761(.A1(new_n18949_), .A2(new_n18951_), .ZN(new_n18954_));
  AOI21_X1   g18762(.A1(new_n18954_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n18955_));
  AOI21_X1   g18763(.A1(new_n18955_), .A2(new_n18953_), .B(new_n18444_), .ZN(new_n18956_));
  INV_X1     g18764(.I(new_n18449_), .ZN(new_n18957_));
  INV_X1     g18765(.I(new_n18459_), .ZN(new_n18958_));
  NOR2_X1    g18766(.A1(new_n18941_), .A2(new_n18942_), .ZN(new_n18959_));
  AOI21_X1   g18767(.A1(new_n18959_), .A2(new_n962_), .B(new_n18958_), .ZN(new_n18960_));
  NAND2_X1   g18768(.A1(new_n18943_), .A2(new_n842_), .ZN(new_n18961_));
  OAI21_X1   g18769(.A1(new_n18960_), .A2(new_n18961_), .B(new_n18455_), .ZN(new_n18962_));
  INV_X1     g18770(.I(new_n18943_), .ZN(new_n18963_));
  OAI21_X1   g18771(.A1(new_n18960_), .A2(new_n18963_), .B(\asqrt[53] ), .ZN(new_n18964_));
  NAND3_X1   g18772(.A1(new_n18962_), .A2(new_n18964_), .A3(new_n720_), .ZN(new_n18965_));
  NAND2_X1   g18773(.A1(new_n18965_), .A2(new_n18452_), .ZN(new_n18966_));
  NAND2_X1   g18774(.A1(new_n18962_), .A2(new_n18964_), .ZN(new_n18967_));
  AOI21_X1   g18775(.A1(new_n18967_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n18968_));
  AOI21_X1   g18776(.A1(new_n18968_), .A2(new_n18966_), .B(new_n18957_), .ZN(new_n18969_));
  AOI21_X1   g18777(.A1(new_n18966_), .A2(new_n18947_), .B(new_n630_), .ZN(new_n18970_));
  OAI21_X1   g18778(.A1(new_n18969_), .A2(new_n18970_), .B(\asqrt[56] ), .ZN(new_n18971_));
  AOI21_X1   g18779(.A1(new_n18953_), .A2(new_n18971_), .B(new_n450_), .ZN(new_n18972_));
  NOR2_X1    g18780(.A1(new_n18956_), .A2(new_n18972_), .ZN(new_n18973_));
  AOI21_X1   g18781(.A1(new_n18973_), .A2(new_n403_), .B(new_n18441_), .ZN(new_n18974_));
  OAI21_X1   g18782(.A1(new_n18956_), .A2(new_n18972_), .B(\asqrt[58] ), .ZN(new_n18975_));
  NAND2_X1   g18783(.A1(new_n18975_), .A2(new_n339_), .ZN(new_n18976_));
  OAI21_X1   g18784(.A1(new_n18974_), .A2(new_n18976_), .B(new_n18437_), .ZN(new_n18977_));
  INV_X1     g18785(.I(new_n18975_), .ZN(new_n18978_));
  OAI21_X1   g18786(.A1(new_n18974_), .A2(new_n18978_), .B(\asqrt[59] ), .ZN(new_n18979_));
  NAND3_X1   g18787(.A1(new_n18977_), .A2(new_n18979_), .A3(new_n288_), .ZN(new_n18980_));
  NAND2_X1   g18788(.A1(new_n18980_), .A2(new_n18435_), .ZN(new_n18981_));
  INV_X1     g18789(.I(new_n18437_), .ZN(new_n18982_));
  INV_X1     g18790(.I(new_n18447_), .ZN(new_n18983_));
  NOR2_X1    g18791(.A1(new_n18969_), .A2(new_n18970_), .ZN(new_n18984_));
  AOI21_X1   g18792(.A1(new_n18984_), .A2(new_n545_), .B(new_n18983_), .ZN(new_n18985_));
  NAND2_X1   g18793(.A1(new_n18971_), .A2(new_n450_), .ZN(new_n18986_));
  OAI21_X1   g18794(.A1(new_n18985_), .A2(new_n18986_), .B(new_n18443_), .ZN(new_n18987_));
  INV_X1     g18795(.I(new_n18971_), .ZN(new_n18988_));
  OAI21_X1   g18796(.A1(new_n18985_), .A2(new_n18988_), .B(\asqrt[57] ), .ZN(new_n18989_));
  NAND3_X1   g18797(.A1(new_n18987_), .A2(new_n18989_), .A3(new_n403_), .ZN(new_n18990_));
  NAND2_X1   g18798(.A1(new_n18990_), .A2(new_n18440_), .ZN(new_n18991_));
  NAND2_X1   g18799(.A1(new_n18987_), .A2(new_n18989_), .ZN(new_n18992_));
  AOI21_X1   g18800(.A1(new_n18992_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n18993_));
  AOI21_X1   g18801(.A1(new_n18993_), .A2(new_n18991_), .B(new_n18982_), .ZN(new_n18994_));
  AOI21_X1   g18802(.A1(new_n18991_), .A2(new_n18975_), .B(new_n339_), .ZN(new_n18995_));
  OAI21_X1   g18803(.A1(new_n18994_), .A2(new_n18995_), .B(\asqrt[60] ), .ZN(new_n18996_));
  AOI21_X1   g18804(.A1(new_n18981_), .A2(new_n18996_), .B(new_n242_), .ZN(new_n18997_));
  NAND2_X1   g18805(.A1(new_n18977_), .A2(new_n18979_), .ZN(new_n18998_));
  AOI21_X1   g18806(.A1(new_n18998_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n18999_));
  AOI21_X1   g18807(.A1(new_n18999_), .A2(new_n18981_), .B(new_n18411_), .ZN(new_n19000_));
  OAI21_X1   g18808(.A1(new_n19000_), .A2(new_n18997_), .B(\asqrt[62] ), .ZN(new_n19001_));
  AOI21_X1   g18809(.A1(new_n18388_), .A2(new_n18394_), .B(new_n18389_), .ZN(new_n19002_));
  NAND2_X1   g18810(.A1(\asqrt[4] ), .A2(new_n19002_), .ZN(new_n19003_));
  XOR2_X1    g18811(.A1(new_n19003_), .A2(new_n18392_), .Z(new_n19004_));
  INV_X1     g18812(.I(new_n19004_), .ZN(new_n19005_));
  NOR3_X1    g18813(.A1(new_n19000_), .A2(new_n18997_), .A3(\asqrt[62] ), .ZN(new_n19006_));
  OAI21_X1   g18814(.A1(new_n19005_), .A2(new_n19006_), .B(new_n19001_), .ZN(new_n19007_));
  NAND3_X1   g18815(.A1(new_n19007_), .A2(new_n18430_), .A3(new_n18432_), .ZN(new_n19008_));
  INV_X1     g18816(.I(new_n18435_), .ZN(new_n19009_));
  NOR2_X1    g18817(.A1(new_n18994_), .A2(new_n18995_), .ZN(new_n19010_));
  AOI21_X1   g18818(.A1(new_n19010_), .A2(new_n288_), .B(new_n19009_), .ZN(new_n19011_));
  INV_X1     g18819(.I(new_n18996_), .ZN(new_n19012_));
  OAI21_X1   g18820(.A1(new_n19011_), .A2(new_n19012_), .B(\asqrt[61] ), .ZN(new_n19013_));
  NAND2_X1   g18821(.A1(new_n18996_), .A2(new_n242_), .ZN(new_n19014_));
  OAI21_X1   g18822(.A1(new_n19011_), .A2(new_n19014_), .B(new_n18410_), .ZN(new_n19015_));
  AOI21_X1   g18823(.A1(new_n19015_), .A2(new_n19013_), .B(new_n234_), .ZN(new_n19016_));
  NOR2_X1    g18824(.A1(new_n19006_), .A2(new_n19005_), .ZN(new_n19017_));
  NOR3_X1    g18825(.A1(new_n19017_), .A2(new_n18430_), .A3(new_n19016_), .ZN(new_n19018_));
  AOI21_X1   g18826(.A1(new_n19008_), .A2(new_n193_), .B(new_n19018_), .ZN(new_n19019_));
  NAND2_X1   g18827(.A1(new_n19019_), .A2(new_n18428_), .ZN(\asqrt[3] ));
  AOI21_X1   g18828(.A1(new_n18981_), .A2(new_n18999_), .B(new_n18997_), .ZN(new_n19021_));
  NAND2_X1   g18829(.A1(\asqrt[3] ), .A2(new_n19021_), .ZN(new_n19022_));
  XOR2_X1    g18830(.A1(new_n19022_), .A2(new_n18411_), .Z(new_n19023_));
  AOI21_X1   g18831(.A1(new_n18991_), .A2(new_n18993_), .B(new_n18995_), .ZN(new_n19024_));
  NAND2_X1   g18832(.A1(\asqrt[3] ), .A2(new_n19024_), .ZN(new_n19025_));
  XOR2_X1    g18833(.A1(new_n19025_), .A2(new_n18982_), .Z(new_n19026_));
  NAND3_X1   g18834(.A1(\asqrt[3] ), .A2(new_n18990_), .A3(new_n18975_), .ZN(new_n19027_));
  XOR2_X1    g18835(.A1(new_n19027_), .A2(new_n18441_), .Z(new_n19028_));
  AOI21_X1   g18836(.A1(new_n18953_), .A2(new_n18955_), .B(new_n18972_), .ZN(new_n19029_));
  NAND2_X1   g18837(.A1(\asqrt[3] ), .A2(new_n19029_), .ZN(new_n19030_));
  XOR2_X1    g18838(.A1(new_n19030_), .A2(new_n18444_), .Z(new_n19031_));
  INV_X1     g18839(.I(new_n19031_), .ZN(new_n19032_));
  NAND3_X1   g18840(.A1(\asqrt[3] ), .A2(new_n18952_), .A3(new_n18971_), .ZN(new_n19033_));
  XOR2_X1    g18841(.A1(new_n19033_), .A2(new_n18983_), .Z(new_n19034_));
  INV_X1     g18842(.I(new_n19034_), .ZN(new_n19035_));
  AOI21_X1   g18843(.A1(new_n18966_), .A2(new_n18968_), .B(new_n18970_), .ZN(new_n19036_));
  NAND2_X1   g18844(.A1(\asqrt[3] ), .A2(new_n19036_), .ZN(new_n19037_));
  XOR2_X1    g18845(.A1(new_n19037_), .A2(new_n18957_), .Z(new_n19038_));
  NAND3_X1   g18846(.A1(\asqrt[3] ), .A2(new_n18965_), .A3(new_n18947_), .ZN(new_n19039_));
  XOR2_X1    g18847(.A1(new_n19039_), .A2(new_n18453_), .Z(new_n19040_));
  AOI21_X1   g18848(.A1(new_n18925_), .A2(new_n18927_), .B(new_n18944_), .ZN(new_n19041_));
  NAND2_X1   g18849(.A1(\asqrt[3] ), .A2(new_n19041_), .ZN(new_n19042_));
  XOR2_X1    g18850(.A1(new_n19042_), .A2(new_n18456_), .Z(new_n19043_));
  INV_X1     g18851(.I(new_n19043_), .ZN(new_n19044_));
  NAND3_X1   g18852(.A1(\asqrt[3] ), .A2(new_n18924_), .A3(new_n18943_), .ZN(new_n19045_));
  XOR2_X1    g18853(.A1(new_n19045_), .A2(new_n18958_), .Z(new_n19046_));
  INV_X1     g18854(.I(new_n19046_), .ZN(new_n19047_));
  AOI21_X1   g18855(.A1(new_n18938_), .A2(new_n18940_), .B(new_n18942_), .ZN(new_n19048_));
  NAND2_X1   g18856(.A1(\asqrt[3] ), .A2(new_n19048_), .ZN(new_n19049_));
  XOR2_X1    g18857(.A1(new_n19049_), .A2(new_n18929_), .Z(new_n19050_));
  NAND3_X1   g18858(.A1(\asqrt[3] ), .A2(new_n18937_), .A3(new_n18919_), .ZN(new_n19051_));
  XOR2_X1    g18859(.A1(new_n19051_), .A2(new_n18465_), .Z(new_n19052_));
  AOI21_X1   g18860(.A1(new_n18897_), .A2(new_n18899_), .B(new_n18916_), .ZN(new_n19053_));
  NAND2_X1   g18861(.A1(\asqrt[3] ), .A2(new_n19053_), .ZN(new_n19054_));
  XOR2_X1    g18862(.A1(new_n19054_), .A2(new_n18468_), .Z(new_n19055_));
  INV_X1     g18863(.I(new_n19055_), .ZN(new_n19056_));
  NAND3_X1   g18864(.A1(\asqrt[3] ), .A2(new_n18896_), .A3(new_n18915_), .ZN(new_n19057_));
  XOR2_X1    g18865(.A1(new_n19057_), .A2(new_n18930_), .Z(new_n19058_));
  INV_X1     g18866(.I(new_n19058_), .ZN(new_n19059_));
  AOI21_X1   g18867(.A1(new_n18910_), .A2(new_n18912_), .B(new_n18914_), .ZN(new_n19060_));
  NAND2_X1   g18868(.A1(\asqrt[3] ), .A2(new_n19060_), .ZN(new_n19061_));
  XOR2_X1    g18869(.A1(new_n19061_), .A2(new_n18901_), .Z(new_n19062_));
  NAND3_X1   g18870(.A1(\asqrt[3] ), .A2(new_n18909_), .A3(new_n18891_), .ZN(new_n19063_));
  XOR2_X1    g18871(.A1(new_n19063_), .A2(new_n18477_), .Z(new_n19064_));
  AOI21_X1   g18872(.A1(new_n18869_), .A2(new_n18871_), .B(new_n18888_), .ZN(new_n19065_));
  NAND2_X1   g18873(.A1(\asqrt[3] ), .A2(new_n19065_), .ZN(new_n19066_));
  XOR2_X1    g18874(.A1(new_n19066_), .A2(new_n18480_), .Z(new_n19067_));
  INV_X1     g18875(.I(new_n19067_), .ZN(new_n19068_));
  NAND3_X1   g18876(.A1(\asqrt[3] ), .A2(new_n18868_), .A3(new_n18887_), .ZN(new_n19069_));
  XOR2_X1    g18877(.A1(new_n19069_), .A2(new_n18902_), .Z(new_n19070_));
  INV_X1     g18878(.I(new_n19070_), .ZN(new_n19071_));
  AOI21_X1   g18879(.A1(new_n18882_), .A2(new_n18884_), .B(new_n18886_), .ZN(new_n19072_));
  NAND2_X1   g18880(.A1(\asqrt[3] ), .A2(new_n19072_), .ZN(new_n19073_));
  XOR2_X1    g18881(.A1(new_n19073_), .A2(new_n18873_), .Z(new_n19074_));
  NAND3_X1   g18882(.A1(\asqrt[3] ), .A2(new_n18881_), .A3(new_n18863_), .ZN(new_n19075_));
  XOR2_X1    g18883(.A1(new_n19075_), .A2(new_n18489_), .Z(new_n19076_));
  AOI21_X1   g18884(.A1(new_n18841_), .A2(new_n18843_), .B(new_n18860_), .ZN(new_n19077_));
  NAND2_X1   g18885(.A1(\asqrt[3] ), .A2(new_n19077_), .ZN(new_n19078_));
  XOR2_X1    g18886(.A1(new_n19078_), .A2(new_n18492_), .Z(new_n19079_));
  INV_X1     g18887(.I(new_n19079_), .ZN(new_n19080_));
  NAND3_X1   g18888(.A1(\asqrt[3] ), .A2(new_n18840_), .A3(new_n18859_), .ZN(new_n19081_));
  XOR2_X1    g18889(.A1(new_n19081_), .A2(new_n18874_), .Z(new_n19082_));
  INV_X1     g18890(.I(new_n19082_), .ZN(new_n19083_));
  AOI21_X1   g18891(.A1(new_n18854_), .A2(new_n18856_), .B(new_n18858_), .ZN(new_n19084_));
  NAND2_X1   g18892(.A1(\asqrt[3] ), .A2(new_n19084_), .ZN(new_n19085_));
  XOR2_X1    g18893(.A1(new_n19085_), .A2(new_n18845_), .Z(new_n19086_));
  NAND3_X1   g18894(.A1(\asqrt[3] ), .A2(new_n18853_), .A3(new_n18835_), .ZN(new_n19087_));
  XOR2_X1    g18895(.A1(new_n19087_), .A2(new_n18501_), .Z(new_n19088_));
  AOI21_X1   g18896(.A1(new_n18813_), .A2(new_n18815_), .B(new_n18832_), .ZN(new_n19089_));
  NAND2_X1   g18897(.A1(\asqrt[3] ), .A2(new_n19089_), .ZN(new_n19090_));
  XOR2_X1    g18898(.A1(new_n19090_), .A2(new_n18504_), .Z(new_n19091_));
  INV_X1     g18899(.I(new_n19091_), .ZN(new_n19092_));
  NAND3_X1   g18900(.A1(\asqrt[3] ), .A2(new_n18812_), .A3(new_n18831_), .ZN(new_n19093_));
  XOR2_X1    g18901(.A1(new_n19093_), .A2(new_n18846_), .Z(new_n19094_));
  INV_X1     g18902(.I(new_n19094_), .ZN(new_n19095_));
  AOI21_X1   g18903(.A1(new_n18826_), .A2(new_n18828_), .B(new_n18830_), .ZN(new_n19096_));
  NAND2_X1   g18904(.A1(\asqrt[3] ), .A2(new_n19096_), .ZN(new_n19097_));
  XOR2_X1    g18905(.A1(new_n19097_), .A2(new_n18817_), .Z(new_n19098_));
  NAND3_X1   g18906(.A1(\asqrt[3] ), .A2(new_n18825_), .A3(new_n18807_), .ZN(new_n19099_));
  XOR2_X1    g18907(.A1(new_n19099_), .A2(new_n18513_), .Z(new_n19100_));
  AOI21_X1   g18908(.A1(new_n18785_), .A2(new_n18787_), .B(new_n18804_), .ZN(new_n19101_));
  NAND2_X1   g18909(.A1(\asqrt[3] ), .A2(new_n19101_), .ZN(new_n19102_));
  XOR2_X1    g18910(.A1(new_n19102_), .A2(new_n18516_), .Z(new_n19103_));
  INV_X1     g18911(.I(new_n19103_), .ZN(new_n19104_));
  NAND3_X1   g18912(.A1(\asqrt[3] ), .A2(new_n18784_), .A3(new_n18803_), .ZN(new_n19105_));
  XOR2_X1    g18913(.A1(new_n19105_), .A2(new_n18818_), .Z(new_n19106_));
  INV_X1     g18914(.I(new_n19106_), .ZN(new_n19107_));
  AOI21_X1   g18915(.A1(new_n18798_), .A2(new_n18800_), .B(new_n18802_), .ZN(new_n19108_));
  NAND2_X1   g18916(.A1(\asqrt[3] ), .A2(new_n19108_), .ZN(new_n19109_));
  XOR2_X1    g18917(.A1(new_n19109_), .A2(new_n18789_), .Z(new_n19110_));
  NAND3_X1   g18918(.A1(\asqrt[3] ), .A2(new_n18797_), .A3(new_n18779_), .ZN(new_n19111_));
  XOR2_X1    g18919(.A1(new_n19111_), .A2(new_n18525_), .Z(new_n19112_));
  AOI21_X1   g18920(.A1(new_n18757_), .A2(new_n18759_), .B(new_n18776_), .ZN(new_n19113_));
  NAND2_X1   g18921(.A1(\asqrt[3] ), .A2(new_n19113_), .ZN(new_n19114_));
  XOR2_X1    g18922(.A1(new_n19114_), .A2(new_n18528_), .Z(new_n19115_));
  INV_X1     g18923(.I(new_n19115_), .ZN(new_n19116_));
  NAND3_X1   g18924(.A1(\asqrt[3] ), .A2(new_n18756_), .A3(new_n18775_), .ZN(new_n19117_));
  XOR2_X1    g18925(.A1(new_n19117_), .A2(new_n18790_), .Z(new_n19118_));
  INV_X1     g18926(.I(new_n19118_), .ZN(new_n19119_));
  AOI21_X1   g18927(.A1(new_n18770_), .A2(new_n18772_), .B(new_n18774_), .ZN(new_n19120_));
  NAND2_X1   g18928(.A1(\asqrt[3] ), .A2(new_n19120_), .ZN(new_n19121_));
  XOR2_X1    g18929(.A1(new_n19121_), .A2(new_n18761_), .Z(new_n19122_));
  NAND3_X1   g18930(.A1(\asqrt[3] ), .A2(new_n18769_), .A3(new_n18751_), .ZN(new_n19123_));
  XOR2_X1    g18931(.A1(new_n19123_), .A2(new_n18537_), .Z(new_n19124_));
  AOI21_X1   g18932(.A1(new_n18729_), .A2(new_n18731_), .B(new_n18748_), .ZN(new_n19125_));
  NAND2_X1   g18933(.A1(\asqrt[3] ), .A2(new_n19125_), .ZN(new_n19126_));
  XOR2_X1    g18934(.A1(new_n19126_), .A2(new_n18540_), .Z(new_n19127_));
  INV_X1     g18935(.I(new_n19127_), .ZN(new_n19128_));
  NAND3_X1   g18936(.A1(\asqrt[3] ), .A2(new_n18728_), .A3(new_n18747_), .ZN(new_n19129_));
  XOR2_X1    g18937(.A1(new_n19129_), .A2(new_n18762_), .Z(new_n19130_));
  INV_X1     g18938(.I(new_n19130_), .ZN(new_n19131_));
  AOI21_X1   g18939(.A1(new_n18742_), .A2(new_n18744_), .B(new_n18746_), .ZN(new_n19132_));
  NAND2_X1   g18940(.A1(\asqrt[3] ), .A2(new_n19132_), .ZN(new_n19133_));
  XOR2_X1    g18941(.A1(new_n19133_), .A2(new_n18733_), .Z(new_n19134_));
  NAND3_X1   g18942(.A1(\asqrt[3] ), .A2(new_n18741_), .A3(new_n18723_), .ZN(new_n19135_));
  XOR2_X1    g18943(.A1(new_n19135_), .A2(new_n18549_), .Z(new_n19136_));
  AOI21_X1   g18944(.A1(new_n18701_), .A2(new_n18703_), .B(new_n18720_), .ZN(new_n19137_));
  NAND2_X1   g18945(.A1(\asqrt[3] ), .A2(new_n19137_), .ZN(new_n19138_));
  XOR2_X1    g18946(.A1(new_n19138_), .A2(new_n18552_), .Z(new_n19139_));
  INV_X1     g18947(.I(new_n19139_), .ZN(new_n19140_));
  NAND3_X1   g18948(.A1(\asqrt[3] ), .A2(new_n18700_), .A3(new_n18719_), .ZN(new_n19141_));
  XOR2_X1    g18949(.A1(new_n19141_), .A2(new_n18734_), .Z(new_n19142_));
  INV_X1     g18950(.I(new_n19142_), .ZN(new_n19143_));
  AOI21_X1   g18951(.A1(new_n18714_), .A2(new_n18716_), .B(new_n18718_), .ZN(new_n19144_));
  NAND2_X1   g18952(.A1(\asqrt[3] ), .A2(new_n19144_), .ZN(new_n19145_));
  XOR2_X1    g18953(.A1(new_n19145_), .A2(new_n18705_), .Z(new_n19146_));
  NAND3_X1   g18954(.A1(\asqrt[3] ), .A2(new_n18713_), .A3(new_n18695_), .ZN(new_n19147_));
  XOR2_X1    g18955(.A1(new_n19147_), .A2(new_n18561_), .Z(new_n19148_));
  AOI21_X1   g18956(.A1(new_n18673_), .A2(new_n18675_), .B(new_n18692_), .ZN(new_n19149_));
  NAND2_X1   g18957(.A1(\asqrt[3] ), .A2(new_n19149_), .ZN(new_n19150_));
  XOR2_X1    g18958(.A1(new_n19150_), .A2(new_n18564_), .Z(new_n19151_));
  INV_X1     g18959(.I(new_n19151_), .ZN(new_n19152_));
  NAND3_X1   g18960(.A1(\asqrt[3] ), .A2(new_n18672_), .A3(new_n18691_), .ZN(new_n19153_));
  XOR2_X1    g18961(.A1(new_n19153_), .A2(new_n18706_), .Z(new_n19154_));
  INV_X1     g18962(.I(new_n19154_), .ZN(new_n19155_));
  AOI21_X1   g18963(.A1(new_n18686_), .A2(new_n18688_), .B(new_n18690_), .ZN(new_n19156_));
  NAND2_X1   g18964(.A1(\asqrt[3] ), .A2(new_n19156_), .ZN(new_n19157_));
  XOR2_X1    g18965(.A1(new_n19157_), .A2(new_n18677_), .Z(new_n19158_));
  NAND3_X1   g18966(.A1(\asqrt[3] ), .A2(new_n18685_), .A3(new_n18667_), .ZN(new_n19159_));
  XOR2_X1    g18967(.A1(new_n19159_), .A2(new_n18573_), .Z(new_n19160_));
  AOI21_X1   g18968(.A1(new_n18630_), .A2(new_n18632_), .B(new_n18664_), .ZN(new_n19161_));
  NAND2_X1   g18969(.A1(\asqrt[3] ), .A2(new_n19161_), .ZN(new_n19162_));
  XOR2_X1    g18970(.A1(new_n19162_), .A2(new_n18576_), .Z(new_n19163_));
  INV_X1     g18971(.I(new_n19163_), .ZN(new_n19164_));
  NAND3_X1   g18972(.A1(\asqrt[3] ), .A2(new_n18629_), .A3(new_n18663_), .ZN(new_n19165_));
  XOR2_X1    g18973(.A1(new_n19165_), .A2(new_n18678_), .Z(new_n19166_));
  INV_X1     g18974(.I(new_n19166_), .ZN(new_n19167_));
  INV_X1     g18975(.I(new_n18432_), .ZN(new_n19168_));
  NAND3_X1   g18976(.A1(new_n19015_), .A2(new_n19013_), .A3(new_n234_), .ZN(new_n19169_));
  NAND2_X1   g18977(.A1(new_n19169_), .A2(new_n19004_), .ZN(new_n19170_));
  AOI21_X1   g18978(.A1(new_n19170_), .A2(new_n19001_), .B(new_n19168_), .ZN(new_n19171_));
  AOI21_X1   g18979(.A1(new_n19171_), .A2(new_n18430_), .B(\asqrt[63] ), .ZN(new_n19172_));
  NOR3_X1    g18980(.A1(new_n19172_), .A2(new_n18427_), .A3(new_n19018_), .ZN(new_n19173_));
  OAI21_X1   g18981(.A1(new_n18623_), .A2(new_n18625_), .B(new_n18628_), .ZN(new_n19174_));
  NOR2_X1    g18982(.A1(new_n19173_), .A2(new_n19174_), .ZN(new_n19175_));
  XOR2_X1    g18983(.A1(new_n19175_), .A2(new_n18581_), .Z(new_n19176_));
  NAND3_X1   g18984(.A1(\asqrt[3] ), .A2(new_n18657_), .A3(new_n18624_), .ZN(new_n19177_));
  XOR2_X1    g18985(.A1(new_n19177_), .A2(new_n18585_), .Z(new_n19178_));
  AOI21_X1   g18986(.A1(new_n18617_), .A2(new_n18618_), .B(new_n18621_), .ZN(new_n19179_));
  NAND2_X1   g18987(.A1(\asqrt[3] ), .A2(new_n19179_), .ZN(new_n19180_));
  XOR2_X1    g18988(.A1(new_n19180_), .A2(new_n18589_), .Z(new_n19181_));
  INV_X1     g18989(.I(new_n19181_), .ZN(new_n19182_));
  NAND2_X1   g18990(.A1(new_n18651_), .A2(new_n16093_), .ZN(new_n19183_));
  NAND3_X1   g18991(.A1(\asqrt[3] ), .A2(new_n19183_), .A3(new_n18620_), .ZN(new_n19184_));
  XOR2_X1    g18992(.A1(new_n19184_), .A2(new_n18635_), .Z(new_n19185_));
  INV_X1     g18993(.I(new_n19185_), .ZN(new_n19186_));
  NAND3_X1   g18994(.A1(\asqrt[3] ), .A2(new_n18649_), .A3(new_n18615_), .ZN(new_n19187_));
  XOR2_X1    g18995(.A1(new_n19187_), .A2(new_n18614_), .Z(new_n19188_));
  NOR2_X1    g18996(.A1(new_n18646_), .A2(\asqrt[6] ), .ZN(new_n19189_));
  OR3_X2     g18997(.A1(new_n19173_), .A2(new_n19189_), .A3(new_n18609_), .Z(new_n19190_));
  XOR2_X1    g18998(.A1(new_n19190_), .A2(new_n18600_), .Z(new_n19191_));
  NOR2_X1    g18999(.A1(\asqrt[3] ), .A2(new_n18424_), .ZN(new_n19192_));
  NOR3_X1    g19000(.A1(new_n19173_), .A2(\a[6] ), .A3(\a[7] ), .ZN(new_n19193_));
  OAI21_X1   g19001(.A1(new_n19193_), .A2(new_n19192_), .B(new_n18596_), .ZN(new_n19194_));
  NAND2_X1   g19002(.A1(new_n19173_), .A2(\asqrt[4] ), .ZN(new_n19195_));
  INV_X1     g19003(.I(\a[6] ), .ZN(new_n19196_));
  INV_X1     g19004(.I(\a[7] ), .ZN(new_n19197_));
  NAND3_X1   g19005(.A1(\asqrt[3] ), .A2(new_n19196_), .A3(new_n19197_), .ZN(new_n19198_));
  NAND3_X1   g19006(.A1(new_n19198_), .A2(\a[8] ), .A3(new_n19195_), .ZN(new_n19199_));
  AND2_X2    g19007(.A1(new_n19194_), .A2(new_n19199_), .Z(new_n19200_));
  NOR3_X1    g19008(.A1(\a[4] ), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n19201_));
  INV_X1     g19009(.I(new_n19201_), .ZN(new_n19202_));
  INV_X1     g19010(.I(new_n18430_), .ZN(new_n19203_));
  AOI21_X1   g19011(.A1(new_n19004_), .A2(new_n19169_), .B(new_n19016_), .ZN(new_n19204_));
  NOR3_X1    g19012(.A1(new_n19204_), .A2(new_n19203_), .A3(new_n19168_), .ZN(new_n19205_));
  NAND3_X1   g19013(.A1(new_n19170_), .A2(new_n19203_), .A3(new_n19001_), .ZN(new_n19206_));
  OAI21_X1   g19014(.A1(new_n19205_), .A2(\asqrt[63] ), .B(new_n19206_), .ZN(new_n19207_));
  OAI21_X1   g19015(.A1(new_n19207_), .A2(new_n18427_), .B(\a[6] ), .ZN(new_n19208_));
  AOI21_X1   g19016(.A1(new_n19208_), .A2(new_n19202_), .B(new_n18424_), .ZN(new_n19209_));
  INV_X1     g19017(.I(new_n19209_), .ZN(new_n19210_));
  OAI21_X1   g19018(.A1(new_n19173_), .A2(\a[6] ), .B(\a[7] ), .ZN(new_n19211_));
  NAND3_X1   g19019(.A1(new_n19208_), .A2(new_n18424_), .A3(new_n19202_), .ZN(new_n19212_));
  NAND3_X1   g19020(.A1(new_n19212_), .A2(new_n19198_), .A3(new_n19211_), .ZN(new_n19213_));
  NAND3_X1   g19021(.A1(new_n19213_), .A2(new_n17816_), .A3(new_n19210_), .ZN(new_n19214_));
  AOI21_X1   g19022(.A1(new_n19213_), .A2(new_n19210_), .B(new_n17816_), .ZN(new_n19215_));
  AOI21_X1   g19023(.A1(new_n19200_), .A2(new_n19214_), .B(new_n19215_), .ZN(new_n19216_));
  NAND3_X1   g19024(.A1(\asqrt[3] ), .A2(new_n18642_), .A3(new_n18606_), .ZN(new_n19217_));
  XOR2_X1    g19025(.A1(new_n19217_), .A2(new_n18644_), .Z(new_n19218_));
  INV_X1     g19026(.I(new_n19218_), .ZN(new_n19219_));
  AOI21_X1   g19027(.A1(new_n19216_), .A2(new_n17242_), .B(new_n19219_), .ZN(new_n19220_));
  OAI21_X1   g19028(.A1(new_n19216_), .A2(new_n17242_), .B(new_n16649_), .ZN(new_n19221_));
  OAI21_X1   g19029(.A1(new_n19220_), .A2(new_n19221_), .B(new_n19191_), .ZN(new_n19222_));
  NOR2_X1    g19030(.A1(new_n19216_), .A2(new_n17242_), .ZN(new_n19223_));
  OAI21_X1   g19031(.A1(new_n19220_), .A2(new_n19223_), .B(\asqrt[7] ), .ZN(new_n19224_));
  NAND3_X1   g19032(.A1(new_n19222_), .A2(new_n19224_), .A3(new_n16093_), .ZN(new_n19225_));
  NAND2_X1   g19033(.A1(new_n19225_), .A2(new_n19188_), .ZN(new_n19226_));
  NAND2_X1   g19034(.A1(new_n19222_), .A2(new_n19224_), .ZN(new_n19227_));
  AOI21_X1   g19035(.A1(new_n19227_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n19228_));
  AOI21_X1   g19036(.A1(new_n19228_), .A2(new_n19226_), .B(new_n19186_), .ZN(new_n19229_));
  INV_X1     g19037(.I(new_n19191_), .ZN(new_n19230_));
  NAND2_X1   g19038(.A1(new_n19194_), .A2(new_n19199_), .ZN(new_n19231_));
  AOI21_X1   g19039(.A1(\asqrt[3] ), .A2(new_n19196_), .B(new_n19197_), .ZN(new_n19232_));
  AOI21_X1   g19040(.A1(new_n19019_), .A2(new_n18428_), .B(new_n19196_), .ZN(new_n19233_));
  NOR3_X1    g19041(.A1(new_n19233_), .A2(\asqrt[4] ), .A3(new_n19201_), .ZN(new_n19234_));
  NOR3_X1    g19042(.A1(new_n19234_), .A2(new_n19232_), .A3(new_n19193_), .ZN(new_n19235_));
  NOR3_X1    g19043(.A1(new_n19235_), .A2(\asqrt[5] ), .A3(new_n19209_), .ZN(new_n19236_));
  OAI21_X1   g19044(.A1(new_n19235_), .A2(new_n19209_), .B(\asqrt[5] ), .ZN(new_n19237_));
  OAI21_X1   g19045(.A1(new_n19231_), .A2(new_n19236_), .B(new_n19237_), .ZN(new_n19238_));
  OAI21_X1   g19046(.A1(new_n19238_), .A2(\asqrt[6] ), .B(new_n19218_), .ZN(new_n19239_));
  AOI21_X1   g19047(.A1(new_n19238_), .A2(\asqrt[6] ), .B(\asqrt[7] ), .ZN(new_n19240_));
  AOI21_X1   g19048(.A1(new_n19240_), .A2(new_n19239_), .B(new_n19230_), .ZN(new_n19241_));
  NAND2_X1   g19049(.A1(new_n19238_), .A2(\asqrt[6] ), .ZN(new_n19242_));
  AOI21_X1   g19050(.A1(new_n19239_), .A2(new_n19242_), .B(new_n16649_), .ZN(new_n19243_));
  OAI21_X1   g19051(.A1(new_n19241_), .A2(new_n19243_), .B(\asqrt[8] ), .ZN(new_n19244_));
  AOI21_X1   g19052(.A1(new_n19226_), .A2(new_n19244_), .B(new_n15518_), .ZN(new_n19245_));
  NOR2_X1    g19053(.A1(new_n19229_), .A2(new_n19245_), .ZN(new_n19246_));
  AOI21_X1   g19054(.A1(new_n19246_), .A2(new_n14985_), .B(new_n19182_), .ZN(new_n19247_));
  OAI21_X1   g19055(.A1(new_n19229_), .A2(new_n19245_), .B(\asqrt[10] ), .ZN(new_n19248_));
  NAND2_X1   g19056(.A1(new_n19248_), .A2(new_n14430_), .ZN(new_n19249_));
  OAI21_X1   g19057(.A1(new_n19247_), .A2(new_n19249_), .B(new_n19178_), .ZN(new_n19250_));
  INV_X1     g19058(.I(new_n19248_), .ZN(new_n19251_));
  OAI21_X1   g19059(.A1(new_n19247_), .A2(new_n19251_), .B(\asqrt[11] ), .ZN(new_n19252_));
  NAND3_X1   g19060(.A1(new_n19250_), .A2(new_n19252_), .A3(new_n13917_), .ZN(new_n19253_));
  NAND2_X1   g19061(.A1(new_n19253_), .A2(new_n19176_), .ZN(new_n19254_));
  NAND2_X1   g19062(.A1(new_n19250_), .A2(new_n19252_), .ZN(new_n19255_));
  AOI21_X1   g19063(.A1(new_n19255_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n19256_));
  AOI21_X1   g19064(.A1(new_n19256_), .A2(new_n19254_), .B(new_n19167_), .ZN(new_n19257_));
  INV_X1     g19065(.I(new_n19178_), .ZN(new_n19258_));
  INV_X1     g19066(.I(new_n19188_), .ZN(new_n19259_));
  NOR2_X1    g19067(.A1(new_n19241_), .A2(new_n19243_), .ZN(new_n19260_));
  AOI21_X1   g19068(.A1(new_n19260_), .A2(new_n16093_), .B(new_n19259_), .ZN(new_n19261_));
  NAND2_X1   g19069(.A1(new_n19244_), .A2(new_n15518_), .ZN(new_n19262_));
  OAI21_X1   g19070(.A1(new_n19261_), .A2(new_n19262_), .B(new_n19185_), .ZN(new_n19263_));
  INV_X1     g19071(.I(new_n19244_), .ZN(new_n19264_));
  OAI21_X1   g19072(.A1(new_n19261_), .A2(new_n19264_), .B(\asqrt[9] ), .ZN(new_n19265_));
  NAND3_X1   g19073(.A1(new_n19263_), .A2(new_n19265_), .A3(new_n14985_), .ZN(new_n19266_));
  NAND2_X1   g19074(.A1(new_n19266_), .A2(new_n19181_), .ZN(new_n19267_));
  NAND2_X1   g19075(.A1(new_n19263_), .A2(new_n19265_), .ZN(new_n19268_));
  AOI21_X1   g19076(.A1(new_n19268_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n19269_));
  AOI21_X1   g19077(.A1(new_n19269_), .A2(new_n19267_), .B(new_n19258_), .ZN(new_n19270_));
  AOI21_X1   g19078(.A1(new_n19267_), .A2(new_n19248_), .B(new_n14430_), .ZN(new_n19271_));
  OAI21_X1   g19079(.A1(new_n19270_), .A2(new_n19271_), .B(\asqrt[12] ), .ZN(new_n19272_));
  AOI21_X1   g19080(.A1(new_n19254_), .A2(new_n19272_), .B(new_n13382_), .ZN(new_n19273_));
  NOR2_X1    g19081(.A1(new_n19257_), .A2(new_n19273_), .ZN(new_n19274_));
  AOI21_X1   g19082(.A1(new_n19274_), .A2(new_n12889_), .B(new_n19164_), .ZN(new_n19275_));
  OAI21_X1   g19083(.A1(new_n19257_), .A2(new_n19273_), .B(\asqrt[14] ), .ZN(new_n19276_));
  NAND2_X1   g19084(.A1(new_n19276_), .A2(new_n12374_), .ZN(new_n19277_));
  OAI21_X1   g19085(.A1(new_n19275_), .A2(new_n19277_), .B(new_n19160_), .ZN(new_n19278_));
  INV_X1     g19086(.I(new_n19276_), .ZN(new_n19279_));
  OAI21_X1   g19087(.A1(new_n19275_), .A2(new_n19279_), .B(\asqrt[15] ), .ZN(new_n19280_));
  NAND3_X1   g19088(.A1(new_n19278_), .A2(new_n19280_), .A3(new_n11901_), .ZN(new_n19281_));
  NAND2_X1   g19089(.A1(new_n19281_), .A2(new_n19158_), .ZN(new_n19282_));
  NAND2_X1   g19090(.A1(new_n19278_), .A2(new_n19280_), .ZN(new_n19283_));
  AOI21_X1   g19091(.A1(new_n19283_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n19284_));
  AOI21_X1   g19092(.A1(new_n19284_), .A2(new_n19282_), .B(new_n19155_), .ZN(new_n19285_));
  INV_X1     g19093(.I(new_n19160_), .ZN(new_n19286_));
  INV_X1     g19094(.I(new_n19176_), .ZN(new_n19287_));
  NOR2_X1    g19095(.A1(new_n19270_), .A2(new_n19271_), .ZN(new_n19288_));
  AOI21_X1   g19096(.A1(new_n19288_), .A2(new_n13917_), .B(new_n19287_), .ZN(new_n19289_));
  NAND2_X1   g19097(.A1(new_n19272_), .A2(new_n13382_), .ZN(new_n19290_));
  OAI21_X1   g19098(.A1(new_n19289_), .A2(new_n19290_), .B(new_n19166_), .ZN(new_n19291_));
  INV_X1     g19099(.I(new_n19272_), .ZN(new_n19292_));
  OAI21_X1   g19100(.A1(new_n19289_), .A2(new_n19292_), .B(\asqrt[13] ), .ZN(new_n19293_));
  NAND3_X1   g19101(.A1(new_n19291_), .A2(new_n19293_), .A3(new_n12889_), .ZN(new_n19294_));
  NAND2_X1   g19102(.A1(new_n19294_), .A2(new_n19163_), .ZN(new_n19295_));
  NAND2_X1   g19103(.A1(new_n19291_), .A2(new_n19293_), .ZN(new_n19296_));
  AOI21_X1   g19104(.A1(new_n19296_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n19297_));
  AOI21_X1   g19105(.A1(new_n19297_), .A2(new_n19295_), .B(new_n19286_), .ZN(new_n19298_));
  AOI21_X1   g19106(.A1(new_n19295_), .A2(new_n19276_), .B(new_n12374_), .ZN(new_n19299_));
  OAI21_X1   g19107(.A1(new_n19298_), .A2(new_n19299_), .B(\asqrt[16] ), .ZN(new_n19300_));
  AOI21_X1   g19108(.A1(new_n19282_), .A2(new_n19300_), .B(new_n11406_), .ZN(new_n19301_));
  NOR2_X1    g19109(.A1(new_n19285_), .A2(new_n19301_), .ZN(new_n19302_));
  AOI21_X1   g19110(.A1(new_n19302_), .A2(new_n10953_), .B(new_n19152_), .ZN(new_n19303_));
  OAI21_X1   g19111(.A1(new_n19285_), .A2(new_n19301_), .B(\asqrt[18] ), .ZN(new_n19304_));
  NAND2_X1   g19112(.A1(new_n19304_), .A2(new_n10478_), .ZN(new_n19305_));
  OAI21_X1   g19113(.A1(new_n19303_), .A2(new_n19305_), .B(new_n19148_), .ZN(new_n19306_));
  INV_X1     g19114(.I(new_n19304_), .ZN(new_n19307_));
  OAI21_X1   g19115(.A1(new_n19303_), .A2(new_n19307_), .B(\asqrt[19] ), .ZN(new_n19308_));
  NAND3_X1   g19116(.A1(new_n19306_), .A2(new_n19308_), .A3(new_n10045_), .ZN(new_n19309_));
  NAND2_X1   g19117(.A1(new_n19309_), .A2(new_n19146_), .ZN(new_n19310_));
  NAND2_X1   g19118(.A1(new_n19306_), .A2(new_n19308_), .ZN(new_n19311_));
  AOI21_X1   g19119(.A1(new_n19311_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n19312_));
  AOI21_X1   g19120(.A1(new_n19312_), .A2(new_n19310_), .B(new_n19143_), .ZN(new_n19313_));
  INV_X1     g19121(.I(new_n19148_), .ZN(new_n19314_));
  INV_X1     g19122(.I(new_n19158_), .ZN(new_n19315_));
  NOR2_X1    g19123(.A1(new_n19298_), .A2(new_n19299_), .ZN(new_n19316_));
  AOI21_X1   g19124(.A1(new_n19316_), .A2(new_n11901_), .B(new_n19315_), .ZN(new_n19317_));
  NAND2_X1   g19125(.A1(new_n19300_), .A2(new_n11406_), .ZN(new_n19318_));
  OAI21_X1   g19126(.A1(new_n19317_), .A2(new_n19318_), .B(new_n19154_), .ZN(new_n19319_));
  INV_X1     g19127(.I(new_n19300_), .ZN(new_n19320_));
  OAI21_X1   g19128(.A1(new_n19317_), .A2(new_n19320_), .B(\asqrt[17] ), .ZN(new_n19321_));
  NAND3_X1   g19129(.A1(new_n19319_), .A2(new_n19321_), .A3(new_n10953_), .ZN(new_n19322_));
  NAND2_X1   g19130(.A1(new_n19322_), .A2(new_n19151_), .ZN(new_n19323_));
  NAND2_X1   g19131(.A1(new_n19319_), .A2(new_n19321_), .ZN(new_n19324_));
  AOI21_X1   g19132(.A1(new_n19324_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n19325_));
  AOI21_X1   g19133(.A1(new_n19325_), .A2(new_n19323_), .B(new_n19314_), .ZN(new_n19326_));
  AOI21_X1   g19134(.A1(new_n19323_), .A2(new_n19304_), .B(new_n10478_), .ZN(new_n19327_));
  OAI21_X1   g19135(.A1(new_n19326_), .A2(new_n19327_), .B(\asqrt[20] ), .ZN(new_n19328_));
  AOI21_X1   g19136(.A1(new_n19310_), .A2(new_n19328_), .B(new_n9590_), .ZN(new_n19329_));
  NOR2_X1    g19137(.A1(new_n19313_), .A2(new_n19329_), .ZN(new_n19330_));
  AOI21_X1   g19138(.A1(new_n19330_), .A2(new_n9177_), .B(new_n19140_), .ZN(new_n19331_));
  OAI21_X1   g19139(.A1(new_n19313_), .A2(new_n19329_), .B(\asqrt[22] ), .ZN(new_n19332_));
  NAND2_X1   g19140(.A1(new_n19332_), .A2(new_n8742_), .ZN(new_n19333_));
  OAI21_X1   g19141(.A1(new_n19331_), .A2(new_n19333_), .B(new_n19136_), .ZN(new_n19334_));
  INV_X1     g19142(.I(new_n19332_), .ZN(new_n19335_));
  OAI21_X1   g19143(.A1(new_n19331_), .A2(new_n19335_), .B(\asqrt[23] ), .ZN(new_n19336_));
  NAND3_X1   g19144(.A1(new_n19334_), .A2(new_n19336_), .A3(new_n8349_), .ZN(new_n19337_));
  NAND2_X1   g19145(.A1(new_n19337_), .A2(new_n19134_), .ZN(new_n19338_));
  NAND2_X1   g19146(.A1(new_n19334_), .A2(new_n19336_), .ZN(new_n19339_));
  AOI21_X1   g19147(.A1(new_n19339_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n19340_));
  AOI21_X1   g19148(.A1(new_n19340_), .A2(new_n19338_), .B(new_n19131_), .ZN(new_n19341_));
  INV_X1     g19149(.I(new_n19136_), .ZN(new_n19342_));
  INV_X1     g19150(.I(new_n19146_), .ZN(new_n19343_));
  NOR2_X1    g19151(.A1(new_n19326_), .A2(new_n19327_), .ZN(new_n19344_));
  AOI21_X1   g19152(.A1(new_n19344_), .A2(new_n10045_), .B(new_n19343_), .ZN(new_n19345_));
  NAND2_X1   g19153(.A1(new_n19328_), .A2(new_n9590_), .ZN(new_n19346_));
  OAI21_X1   g19154(.A1(new_n19345_), .A2(new_n19346_), .B(new_n19142_), .ZN(new_n19347_));
  INV_X1     g19155(.I(new_n19328_), .ZN(new_n19348_));
  OAI21_X1   g19156(.A1(new_n19345_), .A2(new_n19348_), .B(\asqrt[21] ), .ZN(new_n19349_));
  NAND3_X1   g19157(.A1(new_n19347_), .A2(new_n19349_), .A3(new_n9177_), .ZN(new_n19350_));
  NAND2_X1   g19158(.A1(new_n19350_), .A2(new_n19139_), .ZN(new_n19351_));
  NAND2_X1   g19159(.A1(new_n19347_), .A2(new_n19349_), .ZN(new_n19352_));
  AOI21_X1   g19160(.A1(new_n19352_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n19353_));
  AOI21_X1   g19161(.A1(new_n19353_), .A2(new_n19351_), .B(new_n19342_), .ZN(new_n19354_));
  AOI21_X1   g19162(.A1(new_n19351_), .A2(new_n19332_), .B(new_n8742_), .ZN(new_n19355_));
  OAI21_X1   g19163(.A1(new_n19354_), .A2(new_n19355_), .B(\asqrt[24] ), .ZN(new_n19356_));
  AOI21_X1   g19164(.A1(new_n19338_), .A2(new_n19356_), .B(new_n7934_), .ZN(new_n19357_));
  NOR2_X1    g19165(.A1(new_n19341_), .A2(new_n19357_), .ZN(new_n19358_));
  AOI21_X1   g19166(.A1(new_n19358_), .A2(new_n7561_), .B(new_n19128_), .ZN(new_n19359_));
  OAI21_X1   g19167(.A1(new_n19341_), .A2(new_n19357_), .B(\asqrt[26] ), .ZN(new_n19360_));
  NAND2_X1   g19168(.A1(new_n19360_), .A2(new_n7166_), .ZN(new_n19361_));
  OAI21_X1   g19169(.A1(new_n19359_), .A2(new_n19361_), .B(new_n19124_), .ZN(new_n19362_));
  INV_X1     g19170(.I(new_n19360_), .ZN(new_n19363_));
  OAI21_X1   g19171(.A1(new_n19359_), .A2(new_n19363_), .B(\asqrt[27] ), .ZN(new_n19364_));
  NAND3_X1   g19172(.A1(new_n19362_), .A2(new_n19364_), .A3(new_n6813_), .ZN(new_n19365_));
  NAND2_X1   g19173(.A1(new_n19365_), .A2(new_n19122_), .ZN(new_n19366_));
  NAND2_X1   g19174(.A1(new_n19362_), .A2(new_n19364_), .ZN(new_n19367_));
  AOI21_X1   g19175(.A1(new_n19367_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n19368_));
  AOI21_X1   g19176(.A1(new_n19368_), .A2(new_n19366_), .B(new_n19119_), .ZN(new_n19369_));
  INV_X1     g19177(.I(new_n19124_), .ZN(new_n19370_));
  INV_X1     g19178(.I(new_n19134_), .ZN(new_n19371_));
  NOR2_X1    g19179(.A1(new_n19354_), .A2(new_n19355_), .ZN(new_n19372_));
  AOI21_X1   g19180(.A1(new_n19372_), .A2(new_n8349_), .B(new_n19371_), .ZN(new_n19373_));
  NAND2_X1   g19181(.A1(new_n19356_), .A2(new_n7934_), .ZN(new_n19374_));
  OAI21_X1   g19182(.A1(new_n19373_), .A2(new_n19374_), .B(new_n19130_), .ZN(new_n19375_));
  INV_X1     g19183(.I(new_n19356_), .ZN(new_n19376_));
  OAI21_X1   g19184(.A1(new_n19373_), .A2(new_n19376_), .B(\asqrt[25] ), .ZN(new_n19377_));
  NAND3_X1   g19185(.A1(new_n19375_), .A2(new_n19377_), .A3(new_n7561_), .ZN(new_n19378_));
  NAND2_X1   g19186(.A1(new_n19378_), .A2(new_n19127_), .ZN(new_n19379_));
  NAND2_X1   g19187(.A1(new_n19375_), .A2(new_n19377_), .ZN(new_n19380_));
  AOI21_X1   g19188(.A1(new_n19380_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n19381_));
  AOI21_X1   g19189(.A1(new_n19381_), .A2(new_n19379_), .B(new_n19370_), .ZN(new_n19382_));
  AOI21_X1   g19190(.A1(new_n19379_), .A2(new_n19360_), .B(new_n7166_), .ZN(new_n19383_));
  OAI21_X1   g19191(.A1(new_n19382_), .A2(new_n19383_), .B(\asqrt[28] ), .ZN(new_n19384_));
  AOI21_X1   g19192(.A1(new_n19366_), .A2(new_n19384_), .B(new_n6454_), .ZN(new_n19385_));
  NOR2_X1    g19193(.A1(new_n19369_), .A2(new_n19385_), .ZN(new_n19386_));
  AOI21_X1   g19194(.A1(new_n19386_), .A2(new_n6106_), .B(new_n19116_), .ZN(new_n19387_));
  OAI21_X1   g19195(.A1(new_n19369_), .A2(new_n19385_), .B(\asqrt[30] ), .ZN(new_n19388_));
  NAND2_X1   g19196(.A1(new_n19388_), .A2(new_n5750_), .ZN(new_n19389_));
  OAI21_X1   g19197(.A1(new_n19387_), .A2(new_n19389_), .B(new_n19112_), .ZN(new_n19390_));
  INV_X1     g19198(.I(new_n19388_), .ZN(new_n19391_));
  OAI21_X1   g19199(.A1(new_n19387_), .A2(new_n19391_), .B(\asqrt[31] ), .ZN(new_n19392_));
  NAND3_X1   g19200(.A1(new_n19390_), .A2(new_n19392_), .A3(new_n5435_), .ZN(new_n19393_));
  NAND2_X1   g19201(.A1(new_n19393_), .A2(new_n19110_), .ZN(new_n19394_));
  NAND2_X1   g19202(.A1(new_n19390_), .A2(new_n19392_), .ZN(new_n19395_));
  AOI21_X1   g19203(.A1(new_n19395_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n19396_));
  AOI21_X1   g19204(.A1(new_n19396_), .A2(new_n19394_), .B(new_n19107_), .ZN(new_n19397_));
  INV_X1     g19205(.I(new_n19112_), .ZN(new_n19398_));
  INV_X1     g19206(.I(new_n19122_), .ZN(new_n19399_));
  NOR2_X1    g19207(.A1(new_n19382_), .A2(new_n19383_), .ZN(new_n19400_));
  AOI21_X1   g19208(.A1(new_n19400_), .A2(new_n6813_), .B(new_n19399_), .ZN(new_n19401_));
  NAND2_X1   g19209(.A1(new_n19384_), .A2(new_n6454_), .ZN(new_n19402_));
  OAI21_X1   g19210(.A1(new_n19401_), .A2(new_n19402_), .B(new_n19118_), .ZN(new_n19403_));
  INV_X1     g19211(.I(new_n19384_), .ZN(new_n19404_));
  OAI21_X1   g19212(.A1(new_n19401_), .A2(new_n19404_), .B(\asqrt[29] ), .ZN(new_n19405_));
  NAND3_X1   g19213(.A1(new_n19403_), .A2(new_n19405_), .A3(new_n6106_), .ZN(new_n19406_));
  NAND2_X1   g19214(.A1(new_n19406_), .A2(new_n19115_), .ZN(new_n19407_));
  NAND2_X1   g19215(.A1(new_n19403_), .A2(new_n19405_), .ZN(new_n19408_));
  AOI21_X1   g19216(.A1(new_n19408_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n19409_));
  AOI21_X1   g19217(.A1(new_n19409_), .A2(new_n19407_), .B(new_n19398_), .ZN(new_n19410_));
  AOI21_X1   g19218(.A1(new_n19407_), .A2(new_n19388_), .B(new_n5750_), .ZN(new_n19411_));
  OAI21_X1   g19219(.A1(new_n19410_), .A2(new_n19411_), .B(\asqrt[32] ), .ZN(new_n19412_));
  AOI21_X1   g19220(.A1(new_n19394_), .A2(new_n19412_), .B(new_n5110_), .ZN(new_n19413_));
  NOR2_X1    g19221(.A1(new_n19397_), .A2(new_n19413_), .ZN(new_n19414_));
  AOI21_X1   g19222(.A1(new_n19414_), .A2(new_n4810_), .B(new_n19104_), .ZN(new_n19415_));
  OAI21_X1   g19223(.A1(new_n19397_), .A2(new_n19413_), .B(\asqrt[34] ), .ZN(new_n19416_));
  NAND2_X1   g19224(.A1(new_n19416_), .A2(new_n4510_), .ZN(new_n19417_));
  OAI21_X1   g19225(.A1(new_n19415_), .A2(new_n19417_), .B(new_n19100_), .ZN(new_n19418_));
  INV_X1     g19226(.I(new_n19416_), .ZN(new_n19419_));
  OAI21_X1   g19227(.A1(new_n19415_), .A2(new_n19419_), .B(\asqrt[35] ), .ZN(new_n19420_));
  NAND3_X1   g19228(.A1(new_n19418_), .A2(new_n19420_), .A3(new_n4224_), .ZN(new_n19421_));
  NAND2_X1   g19229(.A1(new_n19421_), .A2(new_n19098_), .ZN(new_n19422_));
  NAND2_X1   g19230(.A1(new_n19418_), .A2(new_n19420_), .ZN(new_n19423_));
  AOI21_X1   g19231(.A1(new_n19423_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n19424_));
  AOI21_X1   g19232(.A1(new_n19424_), .A2(new_n19422_), .B(new_n19095_), .ZN(new_n19425_));
  INV_X1     g19233(.I(new_n19100_), .ZN(new_n19426_));
  INV_X1     g19234(.I(new_n19110_), .ZN(new_n19427_));
  NOR2_X1    g19235(.A1(new_n19410_), .A2(new_n19411_), .ZN(new_n19428_));
  AOI21_X1   g19236(.A1(new_n19428_), .A2(new_n5435_), .B(new_n19427_), .ZN(new_n19429_));
  NAND2_X1   g19237(.A1(new_n19412_), .A2(new_n5110_), .ZN(new_n19430_));
  OAI21_X1   g19238(.A1(new_n19429_), .A2(new_n19430_), .B(new_n19106_), .ZN(new_n19431_));
  INV_X1     g19239(.I(new_n19412_), .ZN(new_n19432_));
  OAI21_X1   g19240(.A1(new_n19429_), .A2(new_n19432_), .B(\asqrt[33] ), .ZN(new_n19433_));
  NAND3_X1   g19241(.A1(new_n19431_), .A2(new_n19433_), .A3(new_n4810_), .ZN(new_n19434_));
  NAND2_X1   g19242(.A1(new_n19434_), .A2(new_n19103_), .ZN(new_n19435_));
  NAND2_X1   g19243(.A1(new_n19431_), .A2(new_n19433_), .ZN(new_n19436_));
  AOI21_X1   g19244(.A1(new_n19436_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n19437_));
  AOI21_X1   g19245(.A1(new_n19437_), .A2(new_n19435_), .B(new_n19426_), .ZN(new_n19438_));
  AOI21_X1   g19246(.A1(new_n19435_), .A2(new_n19416_), .B(new_n4510_), .ZN(new_n19439_));
  OAI21_X1   g19247(.A1(new_n19438_), .A2(new_n19439_), .B(\asqrt[36] ), .ZN(new_n19440_));
  AOI21_X1   g19248(.A1(new_n19422_), .A2(new_n19440_), .B(new_n3928_), .ZN(new_n19441_));
  NOR2_X1    g19249(.A1(new_n19425_), .A2(new_n19441_), .ZN(new_n19442_));
  AOI21_X1   g19250(.A1(new_n19442_), .A2(new_n3675_), .B(new_n19092_), .ZN(new_n19443_));
  OAI21_X1   g19251(.A1(new_n19425_), .A2(new_n19441_), .B(\asqrt[38] ), .ZN(new_n19444_));
  NAND2_X1   g19252(.A1(new_n19444_), .A2(new_n3400_), .ZN(new_n19445_));
  OAI21_X1   g19253(.A1(new_n19443_), .A2(new_n19445_), .B(new_n19088_), .ZN(new_n19446_));
  INV_X1     g19254(.I(new_n19444_), .ZN(new_n19447_));
  OAI21_X1   g19255(.A1(new_n19443_), .A2(new_n19447_), .B(\asqrt[39] ), .ZN(new_n19448_));
  NAND3_X1   g19256(.A1(new_n19446_), .A2(new_n19448_), .A3(new_n3167_), .ZN(new_n19449_));
  NAND2_X1   g19257(.A1(new_n19449_), .A2(new_n19086_), .ZN(new_n19450_));
  NAND2_X1   g19258(.A1(new_n19446_), .A2(new_n19448_), .ZN(new_n19451_));
  AOI21_X1   g19259(.A1(new_n19451_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n19452_));
  AOI21_X1   g19260(.A1(new_n19452_), .A2(new_n19450_), .B(new_n19083_), .ZN(new_n19453_));
  INV_X1     g19261(.I(new_n19088_), .ZN(new_n19454_));
  INV_X1     g19262(.I(new_n19098_), .ZN(new_n19455_));
  NOR2_X1    g19263(.A1(new_n19438_), .A2(new_n19439_), .ZN(new_n19456_));
  AOI21_X1   g19264(.A1(new_n19456_), .A2(new_n4224_), .B(new_n19455_), .ZN(new_n19457_));
  NAND2_X1   g19265(.A1(new_n19440_), .A2(new_n3928_), .ZN(new_n19458_));
  OAI21_X1   g19266(.A1(new_n19457_), .A2(new_n19458_), .B(new_n19094_), .ZN(new_n19459_));
  INV_X1     g19267(.I(new_n19440_), .ZN(new_n19460_));
  OAI21_X1   g19268(.A1(new_n19457_), .A2(new_n19460_), .B(\asqrt[37] ), .ZN(new_n19461_));
  NAND3_X1   g19269(.A1(new_n19459_), .A2(new_n19461_), .A3(new_n3675_), .ZN(new_n19462_));
  NAND2_X1   g19270(.A1(new_n19462_), .A2(new_n19091_), .ZN(new_n19463_));
  NAND2_X1   g19271(.A1(new_n19459_), .A2(new_n19461_), .ZN(new_n19464_));
  AOI21_X1   g19272(.A1(new_n19464_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n19465_));
  AOI21_X1   g19273(.A1(new_n19465_), .A2(new_n19463_), .B(new_n19454_), .ZN(new_n19466_));
  AOI21_X1   g19274(.A1(new_n19463_), .A2(new_n19444_), .B(new_n3400_), .ZN(new_n19467_));
  OAI21_X1   g19275(.A1(new_n19466_), .A2(new_n19467_), .B(\asqrt[40] ), .ZN(new_n19468_));
  AOI21_X1   g19276(.A1(new_n19450_), .A2(new_n19468_), .B(new_n2912_), .ZN(new_n19469_));
  NOR2_X1    g19277(.A1(new_n19453_), .A2(new_n19469_), .ZN(new_n19470_));
  AOI21_X1   g19278(.A1(new_n19470_), .A2(new_n2699_), .B(new_n19080_), .ZN(new_n19471_));
  OAI21_X1   g19279(.A1(new_n19453_), .A2(new_n19469_), .B(\asqrt[42] ), .ZN(new_n19472_));
  NAND2_X1   g19280(.A1(new_n19472_), .A2(new_n2464_), .ZN(new_n19473_));
  OAI21_X1   g19281(.A1(new_n19471_), .A2(new_n19473_), .B(new_n19076_), .ZN(new_n19474_));
  INV_X1     g19282(.I(new_n19472_), .ZN(new_n19475_));
  OAI21_X1   g19283(.A1(new_n19471_), .A2(new_n19475_), .B(\asqrt[43] ), .ZN(new_n19476_));
  NAND3_X1   g19284(.A1(new_n19474_), .A2(new_n19476_), .A3(new_n2271_), .ZN(new_n19477_));
  NAND2_X1   g19285(.A1(new_n19477_), .A2(new_n19074_), .ZN(new_n19478_));
  NAND2_X1   g19286(.A1(new_n19474_), .A2(new_n19476_), .ZN(new_n19479_));
  AOI21_X1   g19287(.A1(new_n19479_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n19480_));
  AOI21_X1   g19288(.A1(new_n19480_), .A2(new_n19478_), .B(new_n19071_), .ZN(new_n19481_));
  INV_X1     g19289(.I(new_n19076_), .ZN(new_n19482_));
  INV_X1     g19290(.I(new_n19086_), .ZN(new_n19483_));
  NOR2_X1    g19291(.A1(new_n19466_), .A2(new_n19467_), .ZN(new_n19484_));
  AOI21_X1   g19292(.A1(new_n19484_), .A2(new_n3167_), .B(new_n19483_), .ZN(new_n19485_));
  NAND2_X1   g19293(.A1(new_n19468_), .A2(new_n2912_), .ZN(new_n19486_));
  OAI21_X1   g19294(.A1(new_n19485_), .A2(new_n19486_), .B(new_n19082_), .ZN(new_n19487_));
  INV_X1     g19295(.I(new_n19468_), .ZN(new_n19488_));
  OAI21_X1   g19296(.A1(new_n19485_), .A2(new_n19488_), .B(\asqrt[41] ), .ZN(new_n19489_));
  NAND3_X1   g19297(.A1(new_n19487_), .A2(new_n19489_), .A3(new_n2699_), .ZN(new_n19490_));
  NAND2_X1   g19298(.A1(new_n19490_), .A2(new_n19079_), .ZN(new_n19491_));
  NAND2_X1   g19299(.A1(new_n19487_), .A2(new_n19489_), .ZN(new_n19492_));
  AOI21_X1   g19300(.A1(new_n19492_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n19493_));
  AOI21_X1   g19301(.A1(new_n19493_), .A2(new_n19491_), .B(new_n19482_), .ZN(new_n19494_));
  AOI21_X1   g19302(.A1(new_n19491_), .A2(new_n19472_), .B(new_n2464_), .ZN(new_n19495_));
  OAI21_X1   g19303(.A1(new_n19494_), .A2(new_n19495_), .B(\asqrt[44] ), .ZN(new_n19496_));
  AOI21_X1   g19304(.A1(new_n19478_), .A2(new_n19496_), .B(new_n2072_), .ZN(new_n19497_));
  NOR2_X1    g19305(.A1(new_n19481_), .A2(new_n19497_), .ZN(new_n19498_));
  AOI21_X1   g19306(.A1(new_n19498_), .A2(new_n1884_), .B(new_n19068_), .ZN(new_n19499_));
  OAI21_X1   g19307(.A1(new_n19481_), .A2(new_n19497_), .B(\asqrt[46] ), .ZN(new_n19500_));
  NAND2_X1   g19308(.A1(new_n19500_), .A2(new_n1688_), .ZN(new_n19501_));
  OAI21_X1   g19309(.A1(new_n19499_), .A2(new_n19501_), .B(new_n19064_), .ZN(new_n19502_));
  INV_X1     g19310(.I(new_n19500_), .ZN(new_n19503_));
  OAI21_X1   g19311(.A1(new_n19499_), .A2(new_n19503_), .B(\asqrt[47] ), .ZN(new_n19504_));
  NAND3_X1   g19312(.A1(new_n19502_), .A2(new_n19504_), .A3(new_n1533_), .ZN(new_n19505_));
  NAND2_X1   g19313(.A1(new_n19505_), .A2(new_n19062_), .ZN(new_n19506_));
  NAND2_X1   g19314(.A1(new_n19502_), .A2(new_n19504_), .ZN(new_n19507_));
  AOI21_X1   g19315(.A1(new_n19507_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n19508_));
  AOI21_X1   g19316(.A1(new_n19508_), .A2(new_n19506_), .B(new_n19059_), .ZN(new_n19509_));
  INV_X1     g19317(.I(new_n19064_), .ZN(new_n19510_));
  INV_X1     g19318(.I(new_n19074_), .ZN(new_n19511_));
  NOR2_X1    g19319(.A1(new_n19494_), .A2(new_n19495_), .ZN(new_n19512_));
  AOI21_X1   g19320(.A1(new_n19512_), .A2(new_n2271_), .B(new_n19511_), .ZN(new_n19513_));
  NAND2_X1   g19321(.A1(new_n19496_), .A2(new_n2072_), .ZN(new_n19514_));
  OAI21_X1   g19322(.A1(new_n19513_), .A2(new_n19514_), .B(new_n19070_), .ZN(new_n19515_));
  INV_X1     g19323(.I(new_n19496_), .ZN(new_n19516_));
  OAI21_X1   g19324(.A1(new_n19513_), .A2(new_n19516_), .B(\asqrt[45] ), .ZN(new_n19517_));
  NAND3_X1   g19325(.A1(new_n19515_), .A2(new_n19517_), .A3(new_n1884_), .ZN(new_n19518_));
  NAND2_X1   g19326(.A1(new_n19518_), .A2(new_n19067_), .ZN(new_n19519_));
  NAND2_X1   g19327(.A1(new_n19515_), .A2(new_n19517_), .ZN(new_n19520_));
  AOI21_X1   g19328(.A1(new_n19520_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n19521_));
  AOI21_X1   g19329(.A1(new_n19521_), .A2(new_n19519_), .B(new_n19510_), .ZN(new_n19522_));
  AOI21_X1   g19330(.A1(new_n19519_), .A2(new_n19500_), .B(new_n1688_), .ZN(new_n19523_));
  OAI21_X1   g19331(.A1(new_n19522_), .A2(new_n19523_), .B(\asqrt[48] ), .ZN(new_n19524_));
  AOI21_X1   g19332(.A1(new_n19506_), .A2(new_n19524_), .B(new_n1368_), .ZN(new_n19525_));
  NOR2_X1    g19333(.A1(new_n19509_), .A2(new_n19525_), .ZN(new_n19526_));
  AOI21_X1   g19334(.A1(new_n19526_), .A2(new_n1228_), .B(new_n19056_), .ZN(new_n19527_));
  OAI21_X1   g19335(.A1(new_n19509_), .A2(new_n19525_), .B(\asqrt[50] ), .ZN(new_n19528_));
  NAND2_X1   g19336(.A1(new_n19528_), .A2(new_n1088_), .ZN(new_n19529_));
  OAI21_X1   g19337(.A1(new_n19527_), .A2(new_n19529_), .B(new_n19052_), .ZN(new_n19530_));
  INV_X1     g19338(.I(new_n19528_), .ZN(new_n19531_));
  OAI21_X1   g19339(.A1(new_n19527_), .A2(new_n19531_), .B(\asqrt[51] ), .ZN(new_n19532_));
  NAND3_X1   g19340(.A1(new_n19530_), .A2(new_n19532_), .A3(new_n962_), .ZN(new_n19533_));
  NAND2_X1   g19341(.A1(new_n19533_), .A2(new_n19050_), .ZN(new_n19534_));
  NAND2_X1   g19342(.A1(new_n19530_), .A2(new_n19532_), .ZN(new_n19535_));
  AOI21_X1   g19343(.A1(new_n19535_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n19536_));
  AOI21_X1   g19344(.A1(new_n19536_), .A2(new_n19534_), .B(new_n19047_), .ZN(new_n19537_));
  INV_X1     g19345(.I(new_n19052_), .ZN(new_n19538_));
  INV_X1     g19346(.I(new_n19062_), .ZN(new_n19539_));
  NOR2_X1    g19347(.A1(new_n19522_), .A2(new_n19523_), .ZN(new_n19540_));
  AOI21_X1   g19348(.A1(new_n19540_), .A2(new_n1533_), .B(new_n19539_), .ZN(new_n19541_));
  NAND2_X1   g19349(.A1(new_n19524_), .A2(new_n1368_), .ZN(new_n19542_));
  OAI21_X1   g19350(.A1(new_n19541_), .A2(new_n19542_), .B(new_n19058_), .ZN(new_n19543_));
  INV_X1     g19351(.I(new_n19524_), .ZN(new_n19544_));
  OAI21_X1   g19352(.A1(new_n19541_), .A2(new_n19544_), .B(\asqrt[49] ), .ZN(new_n19545_));
  NAND3_X1   g19353(.A1(new_n19543_), .A2(new_n19545_), .A3(new_n1228_), .ZN(new_n19546_));
  NAND2_X1   g19354(.A1(new_n19546_), .A2(new_n19055_), .ZN(new_n19547_));
  NAND2_X1   g19355(.A1(new_n19543_), .A2(new_n19545_), .ZN(new_n19548_));
  AOI21_X1   g19356(.A1(new_n19548_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n19549_));
  AOI21_X1   g19357(.A1(new_n19549_), .A2(new_n19547_), .B(new_n19538_), .ZN(new_n19550_));
  AOI21_X1   g19358(.A1(new_n19547_), .A2(new_n19528_), .B(new_n1088_), .ZN(new_n19551_));
  OAI21_X1   g19359(.A1(new_n19550_), .A2(new_n19551_), .B(\asqrt[52] ), .ZN(new_n19552_));
  AOI21_X1   g19360(.A1(new_n19534_), .A2(new_n19552_), .B(new_n842_), .ZN(new_n19553_));
  NOR2_X1    g19361(.A1(new_n19537_), .A2(new_n19553_), .ZN(new_n19554_));
  AOI21_X1   g19362(.A1(new_n19554_), .A2(new_n720_), .B(new_n19044_), .ZN(new_n19555_));
  OAI21_X1   g19363(.A1(new_n19537_), .A2(new_n19553_), .B(\asqrt[54] ), .ZN(new_n19556_));
  NAND2_X1   g19364(.A1(new_n19556_), .A2(new_n630_), .ZN(new_n19557_));
  OAI21_X1   g19365(.A1(new_n19555_), .A2(new_n19557_), .B(new_n19040_), .ZN(new_n19558_));
  INV_X1     g19366(.I(new_n19556_), .ZN(new_n19559_));
  OAI21_X1   g19367(.A1(new_n19555_), .A2(new_n19559_), .B(\asqrt[55] ), .ZN(new_n19560_));
  NAND3_X1   g19368(.A1(new_n19558_), .A2(new_n19560_), .A3(new_n545_), .ZN(new_n19561_));
  NAND2_X1   g19369(.A1(new_n19561_), .A2(new_n19038_), .ZN(new_n19562_));
  NAND2_X1   g19370(.A1(new_n19558_), .A2(new_n19560_), .ZN(new_n19563_));
  AOI21_X1   g19371(.A1(new_n19563_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n19564_));
  AOI21_X1   g19372(.A1(new_n19564_), .A2(new_n19562_), .B(new_n19035_), .ZN(new_n19565_));
  INV_X1     g19373(.I(new_n19040_), .ZN(new_n19566_));
  INV_X1     g19374(.I(new_n19050_), .ZN(new_n19567_));
  NOR2_X1    g19375(.A1(new_n19550_), .A2(new_n19551_), .ZN(new_n19568_));
  AOI21_X1   g19376(.A1(new_n19568_), .A2(new_n962_), .B(new_n19567_), .ZN(new_n19569_));
  NAND2_X1   g19377(.A1(new_n19552_), .A2(new_n842_), .ZN(new_n19570_));
  OAI21_X1   g19378(.A1(new_n19569_), .A2(new_n19570_), .B(new_n19046_), .ZN(new_n19571_));
  INV_X1     g19379(.I(new_n19552_), .ZN(new_n19572_));
  OAI21_X1   g19380(.A1(new_n19569_), .A2(new_n19572_), .B(\asqrt[53] ), .ZN(new_n19573_));
  NAND3_X1   g19381(.A1(new_n19571_), .A2(new_n19573_), .A3(new_n720_), .ZN(new_n19574_));
  NAND2_X1   g19382(.A1(new_n19574_), .A2(new_n19043_), .ZN(new_n19575_));
  NAND2_X1   g19383(.A1(new_n19571_), .A2(new_n19573_), .ZN(new_n19576_));
  AOI21_X1   g19384(.A1(new_n19576_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n19577_));
  AOI21_X1   g19385(.A1(new_n19577_), .A2(new_n19575_), .B(new_n19566_), .ZN(new_n19578_));
  AOI21_X1   g19386(.A1(new_n19575_), .A2(new_n19556_), .B(new_n630_), .ZN(new_n19579_));
  OAI21_X1   g19387(.A1(new_n19578_), .A2(new_n19579_), .B(\asqrt[56] ), .ZN(new_n19580_));
  AOI21_X1   g19388(.A1(new_n19562_), .A2(new_n19580_), .B(new_n450_), .ZN(new_n19581_));
  NOR2_X1    g19389(.A1(new_n19565_), .A2(new_n19581_), .ZN(new_n19582_));
  AOI21_X1   g19390(.A1(new_n19582_), .A2(new_n403_), .B(new_n19032_), .ZN(new_n19583_));
  OAI21_X1   g19391(.A1(new_n19565_), .A2(new_n19581_), .B(\asqrt[58] ), .ZN(new_n19584_));
  NAND2_X1   g19392(.A1(new_n19584_), .A2(new_n339_), .ZN(new_n19585_));
  OAI21_X1   g19393(.A1(new_n19583_), .A2(new_n19585_), .B(new_n19028_), .ZN(new_n19586_));
  INV_X1     g19394(.I(new_n19584_), .ZN(new_n19587_));
  OAI21_X1   g19395(.A1(new_n19583_), .A2(new_n19587_), .B(\asqrt[59] ), .ZN(new_n19588_));
  NAND3_X1   g19396(.A1(new_n19586_), .A2(new_n19588_), .A3(new_n288_), .ZN(new_n19589_));
  NAND2_X1   g19397(.A1(new_n19589_), .A2(new_n19026_), .ZN(new_n19590_));
  INV_X1     g19398(.I(new_n19028_), .ZN(new_n19591_));
  INV_X1     g19399(.I(new_n19038_), .ZN(new_n19592_));
  NOR2_X1    g19400(.A1(new_n19578_), .A2(new_n19579_), .ZN(new_n19593_));
  AOI21_X1   g19401(.A1(new_n19593_), .A2(new_n545_), .B(new_n19592_), .ZN(new_n19594_));
  NAND2_X1   g19402(.A1(new_n19580_), .A2(new_n450_), .ZN(new_n19595_));
  OAI21_X1   g19403(.A1(new_n19594_), .A2(new_n19595_), .B(new_n19034_), .ZN(new_n19596_));
  INV_X1     g19404(.I(new_n19580_), .ZN(new_n19597_));
  OAI21_X1   g19405(.A1(new_n19594_), .A2(new_n19597_), .B(\asqrt[57] ), .ZN(new_n19598_));
  NAND3_X1   g19406(.A1(new_n19596_), .A2(new_n19598_), .A3(new_n403_), .ZN(new_n19599_));
  NAND2_X1   g19407(.A1(new_n19599_), .A2(new_n19031_), .ZN(new_n19600_));
  NAND2_X1   g19408(.A1(new_n19596_), .A2(new_n19598_), .ZN(new_n19601_));
  AOI21_X1   g19409(.A1(new_n19601_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n19602_));
  AOI21_X1   g19410(.A1(new_n19602_), .A2(new_n19600_), .B(new_n19591_), .ZN(new_n19603_));
  AOI21_X1   g19411(.A1(new_n19600_), .A2(new_n19584_), .B(new_n339_), .ZN(new_n19604_));
  OAI21_X1   g19412(.A1(new_n19603_), .A2(new_n19604_), .B(\asqrt[60] ), .ZN(new_n19605_));
  AOI21_X1   g19413(.A1(new_n19590_), .A2(new_n19605_), .B(new_n242_), .ZN(new_n19606_));
  NAND3_X1   g19414(.A1(\asqrt[3] ), .A2(new_n18980_), .A3(new_n18996_), .ZN(new_n19607_));
  XOR2_X1    g19415(.A1(new_n19607_), .A2(new_n19009_), .Z(new_n19608_));
  INV_X1     g19416(.I(new_n19608_), .ZN(new_n19609_));
  NAND2_X1   g19417(.A1(new_n19586_), .A2(new_n19588_), .ZN(new_n19610_));
  AOI21_X1   g19418(.A1(new_n19610_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n19611_));
  AOI21_X1   g19419(.A1(new_n19611_), .A2(new_n19590_), .B(new_n19609_), .ZN(new_n19612_));
  OAI21_X1   g19420(.A1(new_n19612_), .A2(new_n19606_), .B(\asqrt[62] ), .ZN(new_n19613_));
  INV_X1     g19421(.I(new_n19026_), .ZN(new_n19614_));
  NOR2_X1    g19422(.A1(new_n19603_), .A2(new_n19604_), .ZN(new_n19615_));
  AOI21_X1   g19423(.A1(new_n19615_), .A2(new_n288_), .B(new_n19614_), .ZN(new_n19616_));
  INV_X1     g19424(.I(new_n19605_), .ZN(new_n19617_));
  OAI21_X1   g19425(.A1(new_n19616_), .A2(new_n19617_), .B(\asqrt[61] ), .ZN(new_n19618_));
  NAND2_X1   g19426(.A1(new_n19605_), .A2(new_n242_), .ZN(new_n19619_));
  OAI21_X1   g19427(.A1(new_n19616_), .A2(new_n19619_), .B(new_n19608_), .ZN(new_n19620_));
  NAND3_X1   g19428(.A1(new_n19620_), .A2(new_n19618_), .A3(new_n234_), .ZN(new_n19621_));
  NOR2_X1    g19429(.A1(new_n19204_), .A2(new_n18430_), .ZN(new_n19622_));
  NOR2_X1    g19430(.A1(new_n19173_), .A2(new_n19203_), .ZN(new_n19623_));
  AOI21_X1   g19431(.A1(new_n19623_), .A2(new_n19204_), .B(new_n19622_), .ZN(new_n19624_));
  NOR2_X1    g19432(.A1(new_n19624_), .A2(new_n193_), .ZN(new_n19625_));
  INV_X1     g19433(.I(new_n19625_), .ZN(new_n19626_));
  NAND3_X1   g19434(.A1(\asqrt[3] ), .A2(new_n19001_), .A3(new_n19169_), .ZN(new_n19627_));
  XOR2_X1    g19435(.A1(new_n19627_), .A2(new_n19005_), .Z(new_n19628_));
  INV_X1     g19436(.I(new_n19628_), .ZN(new_n19629_));
  AOI21_X1   g19437(.A1(new_n19623_), .A2(new_n19007_), .B(new_n19018_), .ZN(new_n19630_));
  AOI21_X1   g19438(.A1(new_n19620_), .A2(new_n19618_), .B(new_n234_), .ZN(new_n19631_));
  INV_X1     g19439(.I(new_n19023_), .ZN(new_n19632_));
  NOR2_X1    g19440(.A1(new_n19612_), .A2(new_n19606_), .ZN(new_n19633_));
  AOI21_X1   g19441(.A1(new_n19633_), .A2(new_n234_), .B(new_n19632_), .ZN(new_n19634_));
  OAI21_X1   g19442(.A1(new_n19634_), .A2(new_n19631_), .B(new_n19630_), .ZN(new_n19635_));
  OAI21_X1   g19443(.A1(new_n19635_), .A2(new_n19629_), .B(new_n193_), .ZN(new_n19636_));
  AOI21_X1   g19444(.A1(new_n19023_), .A2(new_n19621_), .B(new_n19631_), .ZN(new_n19637_));
  NAND2_X1   g19445(.A1(new_n19637_), .A2(new_n19629_), .ZN(new_n19638_));
  NAND3_X1   g19446(.A1(new_n19636_), .A2(new_n19626_), .A3(new_n19638_), .ZN(\asqrt[2] ));
  AND3_X2    g19447(.A1(\asqrt[2] ), .A2(new_n19613_), .A3(new_n19621_), .Z(new_n19640_));
  XOR2_X1    g19448(.A1(new_n19640_), .A2(new_n19023_), .Z(new_n19641_));
  AOI21_X1   g19449(.A1(new_n19590_), .A2(new_n19611_), .B(new_n19606_), .ZN(new_n19642_));
  NAND2_X1   g19450(.A1(\asqrt[2] ), .A2(new_n19642_), .ZN(new_n19643_));
  XOR2_X1    g19451(.A1(new_n19643_), .A2(new_n19609_), .Z(new_n19644_));
  NAND3_X1   g19452(.A1(\asqrt[2] ), .A2(new_n19589_), .A3(new_n19605_), .ZN(new_n19645_));
  XOR2_X1    g19453(.A1(new_n19645_), .A2(new_n19614_), .Z(new_n19646_));
  INV_X1     g19454(.I(new_n19630_), .ZN(new_n19647_));
  NAND2_X1   g19455(.A1(new_n19621_), .A2(new_n19023_), .ZN(new_n19648_));
  AOI21_X1   g19456(.A1(new_n19648_), .A2(new_n19613_), .B(new_n19647_), .ZN(new_n19649_));
  AOI21_X1   g19457(.A1(new_n19649_), .A2(new_n19628_), .B(\asqrt[63] ), .ZN(new_n19650_));
  NAND2_X1   g19458(.A1(new_n19648_), .A2(new_n19613_), .ZN(new_n19651_));
  NOR2_X1    g19459(.A1(new_n19651_), .A2(new_n19628_), .ZN(new_n19652_));
  NOR3_X1    g19460(.A1(new_n19650_), .A2(new_n19625_), .A3(new_n19652_), .ZN(new_n19653_));
  OAI21_X1   g19461(.A1(new_n19583_), .A2(new_n19585_), .B(new_n19588_), .ZN(new_n19654_));
  NOR2_X1    g19462(.A1(new_n19653_), .A2(new_n19654_), .ZN(new_n19655_));
  XOR2_X1    g19463(.A1(new_n19655_), .A2(new_n19028_), .Z(new_n19656_));
  INV_X1     g19464(.I(new_n19656_), .ZN(new_n19657_));
  NAND3_X1   g19465(.A1(\asqrt[2] ), .A2(new_n19599_), .A3(new_n19584_), .ZN(new_n19658_));
  XOR2_X1    g19466(.A1(new_n19658_), .A2(new_n19032_), .Z(new_n19659_));
  INV_X1     g19467(.I(new_n19659_), .ZN(new_n19660_));
  OAI21_X1   g19468(.A1(new_n19594_), .A2(new_n19595_), .B(new_n19598_), .ZN(new_n19661_));
  NOR2_X1    g19469(.A1(new_n19653_), .A2(new_n19661_), .ZN(new_n19662_));
  XOR2_X1    g19470(.A1(new_n19662_), .A2(new_n19034_), .Z(new_n19663_));
  NAND3_X1   g19471(.A1(\asqrt[2] ), .A2(new_n19561_), .A3(new_n19580_), .ZN(new_n19664_));
  XOR2_X1    g19472(.A1(new_n19664_), .A2(new_n19592_), .Z(new_n19665_));
  OAI21_X1   g19473(.A1(new_n19555_), .A2(new_n19557_), .B(new_n19560_), .ZN(new_n19666_));
  NOR2_X1    g19474(.A1(new_n19653_), .A2(new_n19666_), .ZN(new_n19667_));
  XOR2_X1    g19475(.A1(new_n19667_), .A2(new_n19040_), .Z(new_n19668_));
  INV_X1     g19476(.I(new_n19668_), .ZN(new_n19669_));
  NAND3_X1   g19477(.A1(\asqrt[2] ), .A2(new_n19574_), .A3(new_n19556_), .ZN(new_n19670_));
  XOR2_X1    g19478(.A1(new_n19670_), .A2(new_n19044_), .Z(new_n19671_));
  INV_X1     g19479(.I(new_n19671_), .ZN(new_n19672_));
  OAI21_X1   g19480(.A1(new_n19569_), .A2(new_n19570_), .B(new_n19573_), .ZN(new_n19673_));
  NOR2_X1    g19481(.A1(new_n19653_), .A2(new_n19673_), .ZN(new_n19674_));
  XOR2_X1    g19482(.A1(new_n19674_), .A2(new_n19046_), .Z(new_n19675_));
  NAND3_X1   g19483(.A1(\asqrt[2] ), .A2(new_n19533_), .A3(new_n19552_), .ZN(new_n19676_));
  XOR2_X1    g19484(.A1(new_n19676_), .A2(new_n19567_), .Z(new_n19677_));
  OAI21_X1   g19485(.A1(new_n19527_), .A2(new_n19529_), .B(new_n19532_), .ZN(new_n19678_));
  NOR2_X1    g19486(.A1(new_n19653_), .A2(new_n19678_), .ZN(new_n19679_));
  XOR2_X1    g19487(.A1(new_n19679_), .A2(new_n19052_), .Z(new_n19680_));
  INV_X1     g19488(.I(new_n19680_), .ZN(new_n19681_));
  NAND3_X1   g19489(.A1(\asqrt[2] ), .A2(new_n19546_), .A3(new_n19528_), .ZN(new_n19682_));
  XOR2_X1    g19490(.A1(new_n19682_), .A2(new_n19056_), .Z(new_n19683_));
  INV_X1     g19491(.I(new_n19683_), .ZN(new_n19684_));
  OAI21_X1   g19492(.A1(new_n19541_), .A2(new_n19542_), .B(new_n19545_), .ZN(new_n19685_));
  NOR2_X1    g19493(.A1(new_n19653_), .A2(new_n19685_), .ZN(new_n19686_));
  XOR2_X1    g19494(.A1(new_n19686_), .A2(new_n19058_), .Z(new_n19687_));
  NAND3_X1   g19495(.A1(\asqrt[2] ), .A2(new_n19505_), .A3(new_n19524_), .ZN(new_n19688_));
  XOR2_X1    g19496(.A1(new_n19688_), .A2(new_n19539_), .Z(new_n19689_));
  OAI21_X1   g19497(.A1(new_n19499_), .A2(new_n19501_), .B(new_n19504_), .ZN(new_n19690_));
  NOR2_X1    g19498(.A1(new_n19653_), .A2(new_n19690_), .ZN(new_n19691_));
  XOR2_X1    g19499(.A1(new_n19691_), .A2(new_n19064_), .Z(new_n19692_));
  INV_X1     g19500(.I(new_n19692_), .ZN(new_n19693_));
  NAND3_X1   g19501(.A1(\asqrt[2] ), .A2(new_n19518_), .A3(new_n19500_), .ZN(new_n19694_));
  XOR2_X1    g19502(.A1(new_n19694_), .A2(new_n19068_), .Z(new_n19695_));
  INV_X1     g19503(.I(new_n19695_), .ZN(new_n19696_));
  OAI21_X1   g19504(.A1(new_n19513_), .A2(new_n19514_), .B(new_n19517_), .ZN(new_n19697_));
  NOR2_X1    g19505(.A1(new_n19653_), .A2(new_n19697_), .ZN(new_n19698_));
  XOR2_X1    g19506(.A1(new_n19698_), .A2(new_n19070_), .Z(new_n19699_));
  NAND3_X1   g19507(.A1(\asqrt[2] ), .A2(new_n19477_), .A3(new_n19496_), .ZN(new_n19700_));
  XOR2_X1    g19508(.A1(new_n19700_), .A2(new_n19511_), .Z(new_n19701_));
  OAI21_X1   g19509(.A1(new_n19471_), .A2(new_n19473_), .B(new_n19476_), .ZN(new_n19702_));
  NOR2_X1    g19510(.A1(new_n19653_), .A2(new_n19702_), .ZN(new_n19703_));
  XOR2_X1    g19511(.A1(new_n19703_), .A2(new_n19076_), .Z(new_n19704_));
  INV_X1     g19512(.I(new_n19704_), .ZN(new_n19705_));
  NAND3_X1   g19513(.A1(\asqrt[2] ), .A2(new_n19490_), .A3(new_n19472_), .ZN(new_n19706_));
  XOR2_X1    g19514(.A1(new_n19706_), .A2(new_n19080_), .Z(new_n19707_));
  INV_X1     g19515(.I(new_n19707_), .ZN(new_n19708_));
  OAI21_X1   g19516(.A1(new_n19485_), .A2(new_n19486_), .B(new_n19489_), .ZN(new_n19709_));
  NOR2_X1    g19517(.A1(new_n19653_), .A2(new_n19709_), .ZN(new_n19710_));
  XOR2_X1    g19518(.A1(new_n19710_), .A2(new_n19082_), .Z(new_n19711_));
  NAND3_X1   g19519(.A1(\asqrt[2] ), .A2(new_n19449_), .A3(new_n19468_), .ZN(new_n19712_));
  XOR2_X1    g19520(.A1(new_n19712_), .A2(new_n19483_), .Z(new_n19713_));
  OAI21_X1   g19521(.A1(new_n19443_), .A2(new_n19445_), .B(new_n19448_), .ZN(new_n19714_));
  NOR2_X1    g19522(.A1(new_n19653_), .A2(new_n19714_), .ZN(new_n19715_));
  XOR2_X1    g19523(.A1(new_n19715_), .A2(new_n19088_), .Z(new_n19716_));
  INV_X1     g19524(.I(new_n19716_), .ZN(new_n19717_));
  NAND3_X1   g19525(.A1(\asqrt[2] ), .A2(new_n19462_), .A3(new_n19444_), .ZN(new_n19718_));
  XOR2_X1    g19526(.A1(new_n19718_), .A2(new_n19092_), .Z(new_n19719_));
  INV_X1     g19527(.I(new_n19719_), .ZN(new_n19720_));
  OAI21_X1   g19528(.A1(new_n19457_), .A2(new_n19458_), .B(new_n19461_), .ZN(new_n19721_));
  NOR2_X1    g19529(.A1(new_n19653_), .A2(new_n19721_), .ZN(new_n19722_));
  XOR2_X1    g19530(.A1(new_n19722_), .A2(new_n19094_), .Z(new_n19723_));
  NAND3_X1   g19531(.A1(\asqrt[2] ), .A2(new_n19421_), .A3(new_n19440_), .ZN(new_n19724_));
  XOR2_X1    g19532(.A1(new_n19724_), .A2(new_n19455_), .Z(new_n19725_));
  OAI21_X1   g19533(.A1(new_n19415_), .A2(new_n19417_), .B(new_n19420_), .ZN(new_n19726_));
  NOR2_X1    g19534(.A1(new_n19653_), .A2(new_n19726_), .ZN(new_n19727_));
  XOR2_X1    g19535(.A1(new_n19727_), .A2(new_n19100_), .Z(new_n19728_));
  INV_X1     g19536(.I(new_n19728_), .ZN(new_n19729_));
  NAND3_X1   g19537(.A1(\asqrt[2] ), .A2(new_n19434_), .A3(new_n19416_), .ZN(new_n19730_));
  XOR2_X1    g19538(.A1(new_n19730_), .A2(new_n19104_), .Z(new_n19731_));
  INV_X1     g19539(.I(new_n19731_), .ZN(new_n19732_));
  OAI21_X1   g19540(.A1(new_n19429_), .A2(new_n19430_), .B(new_n19433_), .ZN(new_n19733_));
  NOR2_X1    g19541(.A1(new_n19653_), .A2(new_n19733_), .ZN(new_n19734_));
  XOR2_X1    g19542(.A1(new_n19734_), .A2(new_n19106_), .Z(new_n19735_));
  NAND3_X1   g19543(.A1(\asqrt[2] ), .A2(new_n19393_), .A3(new_n19412_), .ZN(new_n19736_));
  XOR2_X1    g19544(.A1(new_n19736_), .A2(new_n19427_), .Z(new_n19737_));
  OAI21_X1   g19545(.A1(new_n19387_), .A2(new_n19389_), .B(new_n19392_), .ZN(new_n19738_));
  NOR2_X1    g19546(.A1(new_n19653_), .A2(new_n19738_), .ZN(new_n19739_));
  XOR2_X1    g19547(.A1(new_n19739_), .A2(new_n19112_), .Z(new_n19740_));
  INV_X1     g19548(.I(new_n19740_), .ZN(new_n19741_));
  NAND3_X1   g19549(.A1(\asqrt[2] ), .A2(new_n19406_), .A3(new_n19388_), .ZN(new_n19742_));
  XOR2_X1    g19550(.A1(new_n19742_), .A2(new_n19116_), .Z(new_n19743_));
  INV_X1     g19551(.I(new_n19743_), .ZN(new_n19744_));
  OAI21_X1   g19552(.A1(new_n19401_), .A2(new_n19402_), .B(new_n19405_), .ZN(new_n19745_));
  NOR2_X1    g19553(.A1(new_n19653_), .A2(new_n19745_), .ZN(new_n19746_));
  XOR2_X1    g19554(.A1(new_n19746_), .A2(new_n19118_), .Z(new_n19747_));
  NAND3_X1   g19555(.A1(\asqrt[2] ), .A2(new_n19365_), .A3(new_n19384_), .ZN(new_n19748_));
  XOR2_X1    g19556(.A1(new_n19748_), .A2(new_n19399_), .Z(new_n19749_));
  OAI21_X1   g19557(.A1(new_n19359_), .A2(new_n19361_), .B(new_n19364_), .ZN(new_n19750_));
  NOR2_X1    g19558(.A1(new_n19653_), .A2(new_n19750_), .ZN(new_n19751_));
  XOR2_X1    g19559(.A1(new_n19751_), .A2(new_n19124_), .Z(new_n19752_));
  INV_X1     g19560(.I(new_n19752_), .ZN(new_n19753_));
  NAND3_X1   g19561(.A1(\asqrt[2] ), .A2(new_n19378_), .A3(new_n19360_), .ZN(new_n19754_));
  XOR2_X1    g19562(.A1(new_n19754_), .A2(new_n19128_), .Z(new_n19755_));
  INV_X1     g19563(.I(new_n19755_), .ZN(new_n19756_));
  OAI21_X1   g19564(.A1(new_n19373_), .A2(new_n19374_), .B(new_n19377_), .ZN(new_n19757_));
  NOR2_X1    g19565(.A1(new_n19653_), .A2(new_n19757_), .ZN(new_n19758_));
  XOR2_X1    g19566(.A1(new_n19758_), .A2(new_n19130_), .Z(new_n19759_));
  NAND3_X1   g19567(.A1(\asqrt[2] ), .A2(new_n19337_), .A3(new_n19356_), .ZN(new_n19760_));
  XOR2_X1    g19568(.A1(new_n19760_), .A2(new_n19371_), .Z(new_n19761_));
  OAI21_X1   g19569(.A1(new_n19331_), .A2(new_n19333_), .B(new_n19336_), .ZN(new_n19762_));
  NOR2_X1    g19570(.A1(new_n19653_), .A2(new_n19762_), .ZN(new_n19763_));
  XOR2_X1    g19571(.A1(new_n19763_), .A2(new_n19136_), .Z(new_n19764_));
  INV_X1     g19572(.I(new_n19764_), .ZN(new_n19765_));
  NAND3_X1   g19573(.A1(\asqrt[2] ), .A2(new_n19350_), .A3(new_n19332_), .ZN(new_n19766_));
  XOR2_X1    g19574(.A1(new_n19766_), .A2(new_n19140_), .Z(new_n19767_));
  INV_X1     g19575(.I(new_n19767_), .ZN(new_n19768_));
  OAI21_X1   g19576(.A1(new_n19345_), .A2(new_n19346_), .B(new_n19349_), .ZN(new_n19769_));
  NOR2_X1    g19577(.A1(new_n19653_), .A2(new_n19769_), .ZN(new_n19770_));
  XOR2_X1    g19578(.A1(new_n19770_), .A2(new_n19142_), .Z(new_n19771_));
  NAND3_X1   g19579(.A1(\asqrt[2] ), .A2(new_n19309_), .A3(new_n19328_), .ZN(new_n19772_));
  XOR2_X1    g19580(.A1(new_n19772_), .A2(new_n19343_), .Z(new_n19773_));
  OAI21_X1   g19581(.A1(new_n19303_), .A2(new_n19305_), .B(new_n19308_), .ZN(new_n19774_));
  NOR2_X1    g19582(.A1(new_n19653_), .A2(new_n19774_), .ZN(new_n19775_));
  XOR2_X1    g19583(.A1(new_n19775_), .A2(new_n19148_), .Z(new_n19776_));
  INV_X1     g19584(.I(new_n19776_), .ZN(new_n19777_));
  NAND3_X1   g19585(.A1(\asqrt[2] ), .A2(new_n19322_), .A3(new_n19304_), .ZN(new_n19778_));
  XOR2_X1    g19586(.A1(new_n19778_), .A2(new_n19152_), .Z(new_n19779_));
  INV_X1     g19587(.I(new_n19779_), .ZN(new_n19780_));
  OAI21_X1   g19588(.A1(new_n19317_), .A2(new_n19318_), .B(new_n19321_), .ZN(new_n19781_));
  NOR2_X1    g19589(.A1(new_n19653_), .A2(new_n19781_), .ZN(new_n19782_));
  XOR2_X1    g19590(.A1(new_n19782_), .A2(new_n19154_), .Z(new_n19783_));
  NAND3_X1   g19591(.A1(\asqrt[2] ), .A2(new_n19281_), .A3(new_n19300_), .ZN(new_n19784_));
  XOR2_X1    g19592(.A1(new_n19784_), .A2(new_n19315_), .Z(new_n19785_));
  OAI21_X1   g19593(.A1(new_n19275_), .A2(new_n19277_), .B(new_n19280_), .ZN(new_n19786_));
  NOR2_X1    g19594(.A1(new_n19653_), .A2(new_n19786_), .ZN(new_n19787_));
  XOR2_X1    g19595(.A1(new_n19787_), .A2(new_n19160_), .Z(new_n19788_));
  INV_X1     g19596(.I(new_n19788_), .ZN(new_n19789_));
  NAND3_X1   g19597(.A1(\asqrt[2] ), .A2(new_n19294_), .A3(new_n19276_), .ZN(new_n19790_));
  XOR2_X1    g19598(.A1(new_n19790_), .A2(new_n19164_), .Z(new_n19791_));
  INV_X1     g19599(.I(new_n19791_), .ZN(new_n19792_));
  OAI21_X1   g19600(.A1(new_n19289_), .A2(new_n19290_), .B(new_n19293_), .ZN(new_n19793_));
  NOR2_X1    g19601(.A1(new_n19653_), .A2(new_n19793_), .ZN(new_n19794_));
  XOR2_X1    g19602(.A1(new_n19794_), .A2(new_n19166_), .Z(new_n19795_));
  NAND3_X1   g19603(.A1(\asqrt[2] ), .A2(new_n19253_), .A3(new_n19272_), .ZN(new_n19796_));
  XOR2_X1    g19604(.A1(new_n19796_), .A2(new_n19287_), .Z(new_n19797_));
  AOI21_X1   g19605(.A1(new_n19267_), .A2(new_n19269_), .B(new_n19271_), .ZN(new_n19798_));
  NAND2_X1   g19606(.A1(\asqrt[2] ), .A2(new_n19798_), .ZN(new_n19799_));
  XOR2_X1    g19607(.A1(new_n19799_), .A2(new_n19258_), .Z(new_n19800_));
  INV_X1     g19608(.I(new_n19800_), .ZN(new_n19801_));
  NAND3_X1   g19609(.A1(\asqrt[2] ), .A2(new_n19266_), .A3(new_n19248_), .ZN(new_n19802_));
  XOR2_X1    g19610(.A1(new_n19802_), .A2(new_n19182_), .Z(new_n19803_));
  INV_X1     g19611(.I(new_n19803_), .ZN(new_n19804_));
  OAI21_X1   g19612(.A1(new_n19261_), .A2(new_n19262_), .B(new_n19265_), .ZN(new_n19805_));
  NOR2_X1    g19613(.A1(new_n19653_), .A2(new_n19805_), .ZN(new_n19806_));
  XOR2_X1    g19614(.A1(new_n19806_), .A2(new_n19185_), .Z(new_n19807_));
  NAND3_X1   g19615(.A1(\asqrt[2] ), .A2(new_n19225_), .A3(new_n19244_), .ZN(new_n19808_));
  XOR2_X1    g19616(.A1(new_n19808_), .A2(new_n19259_), .Z(new_n19809_));
  OAI21_X1   g19617(.A1(new_n19220_), .A2(new_n19221_), .B(new_n19224_), .ZN(new_n19810_));
  NOR2_X1    g19618(.A1(new_n19653_), .A2(new_n19810_), .ZN(new_n19811_));
  XOR2_X1    g19619(.A1(new_n19811_), .A2(new_n19191_), .Z(new_n19812_));
  INV_X1     g19620(.I(new_n19812_), .ZN(new_n19813_));
  NAND2_X1   g19621(.A1(new_n19216_), .A2(new_n17242_), .ZN(new_n19814_));
  NAND3_X1   g19622(.A1(\asqrt[2] ), .A2(new_n19814_), .A3(new_n19242_), .ZN(new_n19815_));
  XOR2_X1    g19623(.A1(new_n19815_), .A2(new_n19219_), .Z(new_n19816_));
  INV_X1     g19624(.I(new_n19816_), .ZN(new_n19817_));
  NOR3_X1    g19625(.A1(new_n19653_), .A2(new_n19236_), .A3(new_n19215_), .ZN(new_n19818_));
  XOR2_X1    g19626(.A1(new_n19818_), .A2(new_n19200_), .Z(new_n19819_));
  NAND4_X1   g19627(.A1(new_n19636_), .A2(\asqrt[3] ), .A3(new_n19626_), .A4(new_n19638_), .ZN(new_n19820_));
  INV_X1     g19628(.I(new_n19820_), .ZN(new_n19821_));
  NOR3_X1    g19629(.A1(new_n19653_), .A2(\a[4] ), .A3(\a[5] ), .ZN(new_n19822_));
  OAI21_X1   g19630(.A1(new_n19822_), .A2(new_n19821_), .B(new_n19196_), .ZN(new_n19823_));
  INV_X1     g19631(.I(\a[4] ), .ZN(new_n19824_));
  INV_X1     g19632(.I(\a[5] ), .ZN(new_n19825_));
  NAND3_X1   g19633(.A1(\asqrt[2] ), .A2(new_n19824_), .A3(new_n19825_), .ZN(new_n19826_));
  NAND3_X1   g19634(.A1(new_n19826_), .A2(\a[6] ), .A3(new_n19820_), .ZN(new_n19827_));
  NAND2_X1   g19635(.A1(new_n19823_), .A2(new_n19827_), .ZN(new_n19828_));
  NOR2_X1    g19636(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n19829_));
  NAND2_X1   g19637(.A1(new_n19829_), .A2(new_n19824_), .ZN(new_n19830_));
  NOR3_X1    g19638(.A1(new_n19637_), .A2(new_n19629_), .A3(new_n19647_), .ZN(new_n19831_));
  OAI21_X1   g19639(.A1(new_n19831_), .A2(\asqrt[63] ), .B(new_n19638_), .ZN(new_n19832_));
  OAI21_X1   g19640(.A1(new_n19832_), .A2(new_n19625_), .B(\a[4] ), .ZN(new_n19833_));
  AOI21_X1   g19641(.A1(new_n19833_), .A2(new_n19830_), .B(new_n19173_), .ZN(new_n19834_));
  AOI21_X1   g19642(.A1(\asqrt[2] ), .A2(new_n19824_), .B(new_n19825_), .ZN(new_n19835_));
  NOR2_X1    g19643(.A1(new_n19835_), .A2(new_n19822_), .ZN(new_n19836_));
  NAND3_X1   g19644(.A1(new_n19833_), .A2(new_n19173_), .A3(new_n19830_), .ZN(new_n19837_));
  AOI21_X1   g19645(.A1(new_n19836_), .A2(new_n19837_), .B(new_n19834_), .ZN(new_n19838_));
  AOI21_X1   g19646(.A1(new_n18424_), .A2(new_n19838_), .B(new_n19828_), .ZN(new_n19839_));
  NOR2_X1    g19647(.A1(new_n19838_), .A2(new_n18424_), .ZN(new_n19840_));
  NOR3_X1    g19648(.A1(new_n19839_), .A2(\asqrt[5] ), .A3(new_n19840_), .ZN(new_n19841_));
  NOR2_X1    g19649(.A1(new_n19232_), .A2(new_n19193_), .ZN(new_n19842_));
  NOR3_X1    g19650(.A1(new_n19653_), .A2(new_n19209_), .A3(new_n19234_), .ZN(new_n19843_));
  XOR2_X1    g19651(.A1(new_n19843_), .A2(new_n19842_), .Z(new_n19844_));
  INV_X1     g19652(.I(new_n19844_), .ZN(new_n19845_));
  OAI21_X1   g19653(.A1(new_n19839_), .A2(new_n19840_), .B(\asqrt[5] ), .ZN(new_n19846_));
  OAI21_X1   g19654(.A1(new_n19841_), .A2(new_n19845_), .B(new_n19846_), .ZN(new_n19847_));
  OAI21_X1   g19655(.A1(new_n19847_), .A2(\asqrt[6] ), .B(new_n19819_), .ZN(new_n19848_));
  AOI21_X1   g19656(.A1(new_n19847_), .A2(\asqrt[6] ), .B(\asqrt[7] ), .ZN(new_n19849_));
  AOI21_X1   g19657(.A1(new_n19849_), .A2(new_n19848_), .B(new_n19817_), .ZN(new_n19850_));
  NAND2_X1   g19658(.A1(new_n19847_), .A2(\asqrt[6] ), .ZN(new_n19851_));
  AOI21_X1   g19659(.A1(new_n19848_), .A2(new_n19851_), .B(new_n16649_), .ZN(new_n19852_));
  NOR2_X1    g19660(.A1(new_n19850_), .A2(new_n19852_), .ZN(new_n19853_));
  AOI21_X1   g19661(.A1(new_n19853_), .A2(new_n16093_), .B(new_n19813_), .ZN(new_n19854_));
  OAI21_X1   g19662(.A1(new_n19850_), .A2(new_n19852_), .B(\asqrt[8] ), .ZN(new_n19855_));
  NAND2_X1   g19663(.A1(new_n19855_), .A2(new_n15518_), .ZN(new_n19856_));
  OAI21_X1   g19664(.A1(new_n19854_), .A2(new_n19856_), .B(new_n19809_), .ZN(new_n19857_));
  INV_X1     g19665(.I(new_n19855_), .ZN(new_n19858_));
  OAI21_X1   g19666(.A1(new_n19854_), .A2(new_n19858_), .B(\asqrt[9] ), .ZN(new_n19859_));
  NAND3_X1   g19667(.A1(new_n19857_), .A2(new_n19859_), .A3(new_n14985_), .ZN(new_n19860_));
  NAND2_X1   g19668(.A1(new_n19860_), .A2(new_n19807_), .ZN(new_n19861_));
  NAND2_X1   g19669(.A1(new_n19857_), .A2(new_n19859_), .ZN(new_n19862_));
  AOI21_X1   g19670(.A1(new_n19862_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n19863_));
  AOI21_X1   g19671(.A1(new_n19863_), .A2(new_n19861_), .B(new_n19804_), .ZN(new_n19864_));
  INV_X1     g19672(.I(new_n19809_), .ZN(new_n19865_));
  INV_X1     g19673(.I(new_n19819_), .ZN(new_n19866_));
  INV_X1     g19674(.I(new_n19828_), .ZN(new_n19867_));
  INV_X1     g19675(.I(new_n19834_), .ZN(new_n19868_));
  NAND2_X1   g19676(.A1(new_n19836_), .A2(new_n19837_), .ZN(new_n19869_));
  NAND3_X1   g19677(.A1(new_n19869_), .A2(new_n18424_), .A3(new_n19868_), .ZN(new_n19870_));
  NAND2_X1   g19678(.A1(new_n19870_), .A2(new_n19867_), .ZN(new_n19871_));
  OR2_X2     g19679(.A1(new_n19838_), .A2(new_n18424_), .Z(new_n19872_));
  NAND3_X1   g19680(.A1(new_n19871_), .A2(new_n19872_), .A3(new_n17816_), .ZN(new_n19873_));
  AOI21_X1   g19681(.A1(new_n19871_), .A2(new_n19872_), .B(new_n17816_), .ZN(new_n19874_));
  AOI21_X1   g19682(.A1(new_n19873_), .A2(new_n19844_), .B(new_n19874_), .ZN(new_n19875_));
  AOI21_X1   g19683(.A1(new_n19875_), .A2(new_n17242_), .B(new_n19866_), .ZN(new_n19876_));
  OAI21_X1   g19684(.A1(new_n19875_), .A2(new_n17242_), .B(new_n16649_), .ZN(new_n19877_));
  OAI21_X1   g19685(.A1(new_n19876_), .A2(new_n19877_), .B(new_n19816_), .ZN(new_n19878_));
  NOR2_X1    g19686(.A1(new_n19875_), .A2(new_n17242_), .ZN(new_n19879_));
  OAI21_X1   g19687(.A1(new_n19876_), .A2(new_n19879_), .B(\asqrt[7] ), .ZN(new_n19880_));
  NAND3_X1   g19688(.A1(new_n19878_), .A2(new_n19880_), .A3(new_n16093_), .ZN(new_n19881_));
  NAND2_X1   g19689(.A1(new_n19881_), .A2(new_n19812_), .ZN(new_n19882_));
  NAND2_X1   g19690(.A1(new_n19878_), .A2(new_n19880_), .ZN(new_n19883_));
  AOI21_X1   g19691(.A1(new_n19883_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n19884_));
  AOI21_X1   g19692(.A1(new_n19884_), .A2(new_n19882_), .B(new_n19865_), .ZN(new_n19885_));
  AOI21_X1   g19693(.A1(new_n19882_), .A2(new_n19855_), .B(new_n15518_), .ZN(new_n19886_));
  OAI21_X1   g19694(.A1(new_n19885_), .A2(new_n19886_), .B(\asqrt[10] ), .ZN(new_n19887_));
  AOI21_X1   g19695(.A1(new_n19861_), .A2(new_n19887_), .B(new_n14430_), .ZN(new_n19888_));
  NOR2_X1    g19696(.A1(new_n19864_), .A2(new_n19888_), .ZN(new_n19889_));
  AOI21_X1   g19697(.A1(new_n19889_), .A2(new_n13917_), .B(new_n19801_), .ZN(new_n19890_));
  OAI21_X1   g19698(.A1(new_n19864_), .A2(new_n19888_), .B(\asqrt[12] ), .ZN(new_n19891_));
  NAND2_X1   g19699(.A1(new_n19891_), .A2(new_n13382_), .ZN(new_n19892_));
  OAI21_X1   g19700(.A1(new_n19890_), .A2(new_n19892_), .B(new_n19797_), .ZN(new_n19893_));
  INV_X1     g19701(.I(new_n19891_), .ZN(new_n19894_));
  OAI21_X1   g19702(.A1(new_n19890_), .A2(new_n19894_), .B(\asqrt[13] ), .ZN(new_n19895_));
  NAND3_X1   g19703(.A1(new_n19893_), .A2(new_n19895_), .A3(new_n12889_), .ZN(new_n19896_));
  NAND2_X1   g19704(.A1(new_n19896_), .A2(new_n19795_), .ZN(new_n19897_));
  NAND2_X1   g19705(.A1(new_n19893_), .A2(new_n19895_), .ZN(new_n19898_));
  AOI21_X1   g19706(.A1(new_n19898_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n19899_));
  AOI21_X1   g19707(.A1(new_n19899_), .A2(new_n19897_), .B(new_n19792_), .ZN(new_n19900_));
  INV_X1     g19708(.I(new_n19797_), .ZN(new_n19901_));
  INV_X1     g19709(.I(new_n19807_), .ZN(new_n19902_));
  NOR2_X1    g19710(.A1(new_n19885_), .A2(new_n19886_), .ZN(new_n19903_));
  AOI21_X1   g19711(.A1(new_n19903_), .A2(new_n14985_), .B(new_n19902_), .ZN(new_n19904_));
  NAND2_X1   g19712(.A1(new_n19887_), .A2(new_n14430_), .ZN(new_n19905_));
  OAI21_X1   g19713(.A1(new_n19904_), .A2(new_n19905_), .B(new_n19803_), .ZN(new_n19906_));
  INV_X1     g19714(.I(new_n19887_), .ZN(new_n19907_));
  OAI21_X1   g19715(.A1(new_n19904_), .A2(new_n19907_), .B(\asqrt[11] ), .ZN(new_n19908_));
  NAND3_X1   g19716(.A1(new_n19906_), .A2(new_n19908_), .A3(new_n13917_), .ZN(new_n19909_));
  NAND2_X1   g19717(.A1(new_n19909_), .A2(new_n19800_), .ZN(new_n19910_));
  NAND2_X1   g19718(.A1(new_n19906_), .A2(new_n19908_), .ZN(new_n19911_));
  AOI21_X1   g19719(.A1(new_n19911_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n19912_));
  AOI21_X1   g19720(.A1(new_n19912_), .A2(new_n19910_), .B(new_n19901_), .ZN(new_n19913_));
  AOI21_X1   g19721(.A1(new_n19910_), .A2(new_n19891_), .B(new_n13382_), .ZN(new_n19914_));
  OAI21_X1   g19722(.A1(new_n19913_), .A2(new_n19914_), .B(\asqrt[14] ), .ZN(new_n19915_));
  AOI21_X1   g19723(.A1(new_n19897_), .A2(new_n19915_), .B(new_n12374_), .ZN(new_n19916_));
  NOR2_X1    g19724(.A1(new_n19900_), .A2(new_n19916_), .ZN(new_n19917_));
  AOI21_X1   g19725(.A1(new_n19917_), .A2(new_n11901_), .B(new_n19789_), .ZN(new_n19918_));
  OAI21_X1   g19726(.A1(new_n19900_), .A2(new_n19916_), .B(\asqrt[16] ), .ZN(new_n19919_));
  NAND2_X1   g19727(.A1(new_n19919_), .A2(new_n11406_), .ZN(new_n19920_));
  OAI21_X1   g19728(.A1(new_n19918_), .A2(new_n19920_), .B(new_n19785_), .ZN(new_n19921_));
  INV_X1     g19729(.I(new_n19919_), .ZN(new_n19922_));
  OAI21_X1   g19730(.A1(new_n19918_), .A2(new_n19922_), .B(\asqrt[17] ), .ZN(new_n19923_));
  NAND3_X1   g19731(.A1(new_n19921_), .A2(new_n19923_), .A3(new_n10953_), .ZN(new_n19924_));
  NAND2_X1   g19732(.A1(new_n19924_), .A2(new_n19783_), .ZN(new_n19925_));
  NAND2_X1   g19733(.A1(new_n19921_), .A2(new_n19923_), .ZN(new_n19926_));
  AOI21_X1   g19734(.A1(new_n19926_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n19927_));
  AOI21_X1   g19735(.A1(new_n19927_), .A2(new_n19925_), .B(new_n19780_), .ZN(new_n19928_));
  INV_X1     g19736(.I(new_n19785_), .ZN(new_n19929_));
  INV_X1     g19737(.I(new_n19795_), .ZN(new_n19930_));
  NOR2_X1    g19738(.A1(new_n19913_), .A2(new_n19914_), .ZN(new_n19931_));
  AOI21_X1   g19739(.A1(new_n19931_), .A2(new_n12889_), .B(new_n19930_), .ZN(new_n19932_));
  NAND2_X1   g19740(.A1(new_n19915_), .A2(new_n12374_), .ZN(new_n19933_));
  OAI21_X1   g19741(.A1(new_n19932_), .A2(new_n19933_), .B(new_n19791_), .ZN(new_n19934_));
  INV_X1     g19742(.I(new_n19915_), .ZN(new_n19935_));
  OAI21_X1   g19743(.A1(new_n19932_), .A2(new_n19935_), .B(\asqrt[15] ), .ZN(new_n19936_));
  NAND3_X1   g19744(.A1(new_n19934_), .A2(new_n19936_), .A3(new_n11901_), .ZN(new_n19937_));
  NAND2_X1   g19745(.A1(new_n19937_), .A2(new_n19788_), .ZN(new_n19938_));
  NAND2_X1   g19746(.A1(new_n19934_), .A2(new_n19936_), .ZN(new_n19939_));
  AOI21_X1   g19747(.A1(new_n19939_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n19940_));
  AOI21_X1   g19748(.A1(new_n19940_), .A2(new_n19938_), .B(new_n19929_), .ZN(new_n19941_));
  AOI21_X1   g19749(.A1(new_n19938_), .A2(new_n19919_), .B(new_n11406_), .ZN(new_n19942_));
  OAI21_X1   g19750(.A1(new_n19941_), .A2(new_n19942_), .B(\asqrt[18] ), .ZN(new_n19943_));
  AOI21_X1   g19751(.A1(new_n19925_), .A2(new_n19943_), .B(new_n10478_), .ZN(new_n19944_));
  NOR2_X1    g19752(.A1(new_n19928_), .A2(new_n19944_), .ZN(new_n19945_));
  AOI21_X1   g19753(.A1(new_n19945_), .A2(new_n10045_), .B(new_n19777_), .ZN(new_n19946_));
  OAI21_X1   g19754(.A1(new_n19928_), .A2(new_n19944_), .B(\asqrt[20] ), .ZN(new_n19947_));
  NAND2_X1   g19755(.A1(new_n19947_), .A2(new_n9590_), .ZN(new_n19948_));
  OAI21_X1   g19756(.A1(new_n19946_), .A2(new_n19948_), .B(new_n19773_), .ZN(new_n19949_));
  INV_X1     g19757(.I(new_n19947_), .ZN(new_n19950_));
  OAI21_X1   g19758(.A1(new_n19946_), .A2(new_n19950_), .B(\asqrt[21] ), .ZN(new_n19951_));
  NAND3_X1   g19759(.A1(new_n19949_), .A2(new_n19951_), .A3(new_n9177_), .ZN(new_n19952_));
  NAND2_X1   g19760(.A1(new_n19952_), .A2(new_n19771_), .ZN(new_n19953_));
  NAND2_X1   g19761(.A1(new_n19949_), .A2(new_n19951_), .ZN(new_n19954_));
  AOI21_X1   g19762(.A1(new_n19954_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n19955_));
  AOI21_X1   g19763(.A1(new_n19955_), .A2(new_n19953_), .B(new_n19768_), .ZN(new_n19956_));
  INV_X1     g19764(.I(new_n19773_), .ZN(new_n19957_));
  INV_X1     g19765(.I(new_n19783_), .ZN(new_n19958_));
  NOR2_X1    g19766(.A1(new_n19941_), .A2(new_n19942_), .ZN(new_n19959_));
  AOI21_X1   g19767(.A1(new_n19959_), .A2(new_n10953_), .B(new_n19958_), .ZN(new_n19960_));
  NAND2_X1   g19768(.A1(new_n19943_), .A2(new_n10478_), .ZN(new_n19961_));
  OAI21_X1   g19769(.A1(new_n19960_), .A2(new_n19961_), .B(new_n19779_), .ZN(new_n19962_));
  INV_X1     g19770(.I(new_n19943_), .ZN(new_n19963_));
  OAI21_X1   g19771(.A1(new_n19960_), .A2(new_n19963_), .B(\asqrt[19] ), .ZN(new_n19964_));
  NAND3_X1   g19772(.A1(new_n19962_), .A2(new_n19964_), .A3(new_n10045_), .ZN(new_n19965_));
  NAND2_X1   g19773(.A1(new_n19965_), .A2(new_n19776_), .ZN(new_n19966_));
  NAND2_X1   g19774(.A1(new_n19962_), .A2(new_n19964_), .ZN(new_n19967_));
  AOI21_X1   g19775(.A1(new_n19967_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n19968_));
  AOI21_X1   g19776(.A1(new_n19968_), .A2(new_n19966_), .B(new_n19957_), .ZN(new_n19969_));
  AOI21_X1   g19777(.A1(new_n19966_), .A2(new_n19947_), .B(new_n9590_), .ZN(new_n19970_));
  OAI21_X1   g19778(.A1(new_n19969_), .A2(new_n19970_), .B(\asqrt[22] ), .ZN(new_n19971_));
  AOI21_X1   g19779(.A1(new_n19953_), .A2(new_n19971_), .B(new_n8742_), .ZN(new_n19972_));
  NOR2_X1    g19780(.A1(new_n19956_), .A2(new_n19972_), .ZN(new_n19973_));
  AOI21_X1   g19781(.A1(new_n19973_), .A2(new_n8349_), .B(new_n19765_), .ZN(new_n19974_));
  OAI21_X1   g19782(.A1(new_n19956_), .A2(new_n19972_), .B(\asqrt[24] ), .ZN(new_n19975_));
  NAND2_X1   g19783(.A1(new_n19975_), .A2(new_n7934_), .ZN(new_n19976_));
  OAI21_X1   g19784(.A1(new_n19974_), .A2(new_n19976_), .B(new_n19761_), .ZN(new_n19977_));
  INV_X1     g19785(.I(new_n19975_), .ZN(new_n19978_));
  OAI21_X1   g19786(.A1(new_n19974_), .A2(new_n19978_), .B(\asqrt[25] ), .ZN(new_n19979_));
  NAND3_X1   g19787(.A1(new_n19977_), .A2(new_n19979_), .A3(new_n7561_), .ZN(new_n19980_));
  NAND2_X1   g19788(.A1(new_n19980_), .A2(new_n19759_), .ZN(new_n19981_));
  NAND2_X1   g19789(.A1(new_n19977_), .A2(new_n19979_), .ZN(new_n19982_));
  AOI21_X1   g19790(.A1(new_n19982_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n19983_));
  AOI21_X1   g19791(.A1(new_n19983_), .A2(new_n19981_), .B(new_n19756_), .ZN(new_n19984_));
  INV_X1     g19792(.I(new_n19761_), .ZN(new_n19985_));
  INV_X1     g19793(.I(new_n19771_), .ZN(new_n19986_));
  NOR2_X1    g19794(.A1(new_n19969_), .A2(new_n19970_), .ZN(new_n19987_));
  AOI21_X1   g19795(.A1(new_n19987_), .A2(new_n9177_), .B(new_n19986_), .ZN(new_n19988_));
  NAND2_X1   g19796(.A1(new_n19971_), .A2(new_n8742_), .ZN(new_n19989_));
  OAI21_X1   g19797(.A1(new_n19988_), .A2(new_n19989_), .B(new_n19767_), .ZN(new_n19990_));
  INV_X1     g19798(.I(new_n19971_), .ZN(new_n19991_));
  OAI21_X1   g19799(.A1(new_n19988_), .A2(new_n19991_), .B(\asqrt[23] ), .ZN(new_n19992_));
  NAND3_X1   g19800(.A1(new_n19990_), .A2(new_n19992_), .A3(new_n8349_), .ZN(new_n19993_));
  NAND2_X1   g19801(.A1(new_n19993_), .A2(new_n19764_), .ZN(new_n19994_));
  NAND2_X1   g19802(.A1(new_n19990_), .A2(new_n19992_), .ZN(new_n19995_));
  AOI21_X1   g19803(.A1(new_n19995_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n19996_));
  AOI21_X1   g19804(.A1(new_n19996_), .A2(new_n19994_), .B(new_n19985_), .ZN(new_n19997_));
  AOI21_X1   g19805(.A1(new_n19994_), .A2(new_n19975_), .B(new_n7934_), .ZN(new_n19998_));
  OAI21_X1   g19806(.A1(new_n19997_), .A2(new_n19998_), .B(\asqrt[26] ), .ZN(new_n19999_));
  AOI21_X1   g19807(.A1(new_n19981_), .A2(new_n19999_), .B(new_n7166_), .ZN(new_n20000_));
  NOR2_X1    g19808(.A1(new_n19984_), .A2(new_n20000_), .ZN(new_n20001_));
  AOI21_X1   g19809(.A1(new_n20001_), .A2(new_n6813_), .B(new_n19753_), .ZN(new_n20002_));
  OAI21_X1   g19810(.A1(new_n19984_), .A2(new_n20000_), .B(\asqrt[28] ), .ZN(new_n20003_));
  NAND2_X1   g19811(.A1(new_n20003_), .A2(new_n6454_), .ZN(new_n20004_));
  OAI21_X1   g19812(.A1(new_n20002_), .A2(new_n20004_), .B(new_n19749_), .ZN(new_n20005_));
  INV_X1     g19813(.I(new_n20003_), .ZN(new_n20006_));
  OAI21_X1   g19814(.A1(new_n20002_), .A2(new_n20006_), .B(\asqrt[29] ), .ZN(new_n20007_));
  NAND3_X1   g19815(.A1(new_n20005_), .A2(new_n20007_), .A3(new_n6106_), .ZN(new_n20008_));
  NAND2_X1   g19816(.A1(new_n20008_), .A2(new_n19747_), .ZN(new_n20009_));
  NAND2_X1   g19817(.A1(new_n20005_), .A2(new_n20007_), .ZN(new_n20010_));
  AOI21_X1   g19818(.A1(new_n20010_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n20011_));
  AOI21_X1   g19819(.A1(new_n20011_), .A2(new_n20009_), .B(new_n19744_), .ZN(new_n20012_));
  INV_X1     g19820(.I(new_n19749_), .ZN(new_n20013_));
  INV_X1     g19821(.I(new_n19759_), .ZN(new_n20014_));
  NOR2_X1    g19822(.A1(new_n19997_), .A2(new_n19998_), .ZN(new_n20015_));
  AOI21_X1   g19823(.A1(new_n20015_), .A2(new_n7561_), .B(new_n20014_), .ZN(new_n20016_));
  NAND2_X1   g19824(.A1(new_n19999_), .A2(new_n7166_), .ZN(new_n20017_));
  OAI21_X1   g19825(.A1(new_n20016_), .A2(new_n20017_), .B(new_n19755_), .ZN(new_n20018_));
  INV_X1     g19826(.I(new_n19999_), .ZN(new_n20019_));
  OAI21_X1   g19827(.A1(new_n20016_), .A2(new_n20019_), .B(\asqrt[27] ), .ZN(new_n20020_));
  NAND3_X1   g19828(.A1(new_n20018_), .A2(new_n20020_), .A3(new_n6813_), .ZN(new_n20021_));
  NAND2_X1   g19829(.A1(new_n20021_), .A2(new_n19752_), .ZN(new_n20022_));
  NAND2_X1   g19830(.A1(new_n20018_), .A2(new_n20020_), .ZN(new_n20023_));
  AOI21_X1   g19831(.A1(new_n20023_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n20024_));
  AOI21_X1   g19832(.A1(new_n20024_), .A2(new_n20022_), .B(new_n20013_), .ZN(new_n20025_));
  AOI21_X1   g19833(.A1(new_n20022_), .A2(new_n20003_), .B(new_n6454_), .ZN(new_n20026_));
  OAI21_X1   g19834(.A1(new_n20025_), .A2(new_n20026_), .B(\asqrt[30] ), .ZN(new_n20027_));
  AOI21_X1   g19835(.A1(new_n20009_), .A2(new_n20027_), .B(new_n5750_), .ZN(new_n20028_));
  NOR2_X1    g19836(.A1(new_n20012_), .A2(new_n20028_), .ZN(new_n20029_));
  AOI21_X1   g19837(.A1(new_n20029_), .A2(new_n5435_), .B(new_n19741_), .ZN(new_n20030_));
  OAI21_X1   g19838(.A1(new_n20012_), .A2(new_n20028_), .B(\asqrt[32] ), .ZN(new_n20031_));
  NAND2_X1   g19839(.A1(new_n20031_), .A2(new_n5110_), .ZN(new_n20032_));
  OAI21_X1   g19840(.A1(new_n20030_), .A2(new_n20032_), .B(new_n19737_), .ZN(new_n20033_));
  INV_X1     g19841(.I(new_n20031_), .ZN(new_n20034_));
  OAI21_X1   g19842(.A1(new_n20030_), .A2(new_n20034_), .B(\asqrt[33] ), .ZN(new_n20035_));
  NAND3_X1   g19843(.A1(new_n20033_), .A2(new_n20035_), .A3(new_n4810_), .ZN(new_n20036_));
  NAND2_X1   g19844(.A1(new_n20036_), .A2(new_n19735_), .ZN(new_n20037_));
  NAND2_X1   g19845(.A1(new_n20033_), .A2(new_n20035_), .ZN(new_n20038_));
  AOI21_X1   g19846(.A1(new_n20038_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n20039_));
  AOI21_X1   g19847(.A1(new_n20039_), .A2(new_n20037_), .B(new_n19732_), .ZN(new_n20040_));
  INV_X1     g19848(.I(new_n19737_), .ZN(new_n20041_));
  INV_X1     g19849(.I(new_n19747_), .ZN(new_n20042_));
  NOR2_X1    g19850(.A1(new_n20025_), .A2(new_n20026_), .ZN(new_n20043_));
  AOI21_X1   g19851(.A1(new_n20043_), .A2(new_n6106_), .B(new_n20042_), .ZN(new_n20044_));
  NAND2_X1   g19852(.A1(new_n20027_), .A2(new_n5750_), .ZN(new_n20045_));
  OAI21_X1   g19853(.A1(new_n20044_), .A2(new_n20045_), .B(new_n19743_), .ZN(new_n20046_));
  INV_X1     g19854(.I(new_n20027_), .ZN(new_n20047_));
  OAI21_X1   g19855(.A1(new_n20044_), .A2(new_n20047_), .B(\asqrt[31] ), .ZN(new_n20048_));
  NAND3_X1   g19856(.A1(new_n20046_), .A2(new_n20048_), .A3(new_n5435_), .ZN(new_n20049_));
  NAND2_X1   g19857(.A1(new_n20049_), .A2(new_n19740_), .ZN(new_n20050_));
  NAND2_X1   g19858(.A1(new_n20046_), .A2(new_n20048_), .ZN(new_n20051_));
  AOI21_X1   g19859(.A1(new_n20051_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n20052_));
  AOI21_X1   g19860(.A1(new_n20052_), .A2(new_n20050_), .B(new_n20041_), .ZN(new_n20053_));
  AOI21_X1   g19861(.A1(new_n20050_), .A2(new_n20031_), .B(new_n5110_), .ZN(new_n20054_));
  OAI21_X1   g19862(.A1(new_n20053_), .A2(new_n20054_), .B(\asqrt[34] ), .ZN(new_n20055_));
  AOI21_X1   g19863(.A1(new_n20037_), .A2(new_n20055_), .B(new_n4510_), .ZN(new_n20056_));
  NOR2_X1    g19864(.A1(new_n20040_), .A2(new_n20056_), .ZN(new_n20057_));
  AOI21_X1   g19865(.A1(new_n20057_), .A2(new_n4224_), .B(new_n19729_), .ZN(new_n20058_));
  OAI21_X1   g19866(.A1(new_n20040_), .A2(new_n20056_), .B(\asqrt[36] ), .ZN(new_n20059_));
  NAND2_X1   g19867(.A1(new_n20059_), .A2(new_n3928_), .ZN(new_n20060_));
  OAI21_X1   g19868(.A1(new_n20058_), .A2(new_n20060_), .B(new_n19725_), .ZN(new_n20061_));
  INV_X1     g19869(.I(new_n20059_), .ZN(new_n20062_));
  OAI21_X1   g19870(.A1(new_n20058_), .A2(new_n20062_), .B(\asqrt[37] ), .ZN(new_n20063_));
  NAND3_X1   g19871(.A1(new_n20061_), .A2(new_n20063_), .A3(new_n3675_), .ZN(new_n20064_));
  NAND2_X1   g19872(.A1(new_n20064_), .A2(new_n19723_), .ZN(new_n20065_));
  NAND2_X1   g19873(.A1(new_n20061_), .A2(new_n20063_), .ZN(new_n20066_));
  AOI21_X1   g19874(.A1(new_n20066_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n20067_));
  AOI21_X1   g19875(.A1(new_n20067_), .A2(new_n20065_), .B(new_n19720_), .ZN(new_n20068_));
  INV_X1     g19876(.I(new_n19725_), .ZN(new_n20069_));
  INV_X1     g19877(.I(new_n19735_), .ZN(new_n20070_));
  NOR2_X1    g19878(.A1(new_n20053_), .A2(new_n20054_), .ZN(new_n20071_));
  AOI21_X1   g19879(.A1(new_n20071_), .A2(new_n4810_), .B(new_n20070_), .ZN(new_n20072_));
  NAND2_X1   g19880(.A1(new_n20055_), .A2(new_n4510_), .ZN(new_n20073_));
  OAI21_X1   g19881(.A1(new_n20072_), .A2(new_n20073_), .B(new_n19731_), .ZN(new_n20074_));
  INV_X1     g19882(.I(new_n20055_), .ZN(new_n20075_));
  OAI21_X1   g19883(.A1(new_n20072_), .A2(new_n20075_), .B(\asqrt[35] ), .ZN(new_n20076_));
  NAND3_X1   g19884(.A1(new_n20074_), .A2(new_n20076_), .A3(new_n4224_), .ZN(new_n20077_));
  NAND2_X1   g19885(.A1(new_n20077_), .A2(new_n19728_), .ZN(new_n20078_));
  NAND2_X1   g19886(.A1(new_n20074_), .A2(new_n20076_), .ZN(new_n20079_));
  AOI21_X1   g19887(.A1(new_n20079_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n20080_));
  AOI21_X1   g19888(.A1(new_n20080_), .A2(new_n20078_), .B(new_n20069_), .ZN(new_n20081_));
  AOI21_X1   g19889(.A1(new_n20078_), .A2(new_n20059_), .B(new_n3928_), .ZN(new_n20082_));
  OAI21_X1   g19890(.A1(new_n20081_), .A2(new_n20082_), .B(\asqrt[38] ), .ZN(new_n20083_));
  AOI21_X1   g19891(.A1(new_n20065_), .A2(new_n20083_), .B(new_n3400_), .ZN(new_n20084_));
  NOR2_X1    g19892(.A1(new_n20068_), .A2(new_n20084_), .ZN(new_n20085_));
  AOI21_X1   g19893(.A1(new_n20085_), .A2(new_n3167_), .B(new_n19717_), .ZN(new_n20086_));
  OAI21_X1   g19894(.A1(new_n20068_), .A2(new_n20084_), .B(\asqrt[40] ), .ZN(new_n20087_));
  NAND2_X1   g19895(.A1(new_n20087_), .A2(new_n2912_), .ZN(new_n20088_));
  OAI21_X1   g19896(.A1(new_n20086_), .A2(new_n20088_), .B(new_n19713_), .ZN(new_n20089_));
  INV_X1     g19897(.I(new_n20087_), .ZN(new_n20090_));
  OAI21_X1   g19898(.A1(new_n20086_), .A2(new_n20090_), .B(\asqrt[41] ), .ZN(new_n20091_));
  NAND3_X1   g19899(.A1(new_n20089_), .A2(new_n20091_), .A3(new_n2699_), .ZN(new_n20092_));
  NAND2_X1   g19900(.A1(new_n20092_), .A2(new_n19711_), .ZN(new_n20093_));
  NAND2_X1   g19901(.A1(new_n20089_), .A2(new_n20091_), .ZN(new_n20094_));
  AOI21_X1   g19902(.A1(new_n20094_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n20095_));
  AOI21_X1   g19903(.A1(new_n20095_), .A2(new_n20093_), .B(new_n19708_), .ZN(new_n20096_));
  INV_X1     g19904(.I(new_n19713_), .ZN(new_n20097_));
  INV_X1     g19905(.I(new_n19723_), .ZN(new_n20098_));
  NOR2_X1    g19906(.A1(new_n20081_), .A2(new_n20082_), .ZN(new_n20099_));
  AOI21_X1   g19907(.A1(new_n20099_), .A2(new_n3675_), .B(new_n20098_), .ZN(new_n20100_));
  NAND2_X1   g19908(.A1(new_n20083_), .A2(new_n3400_), .ZN(new_n20101_));
  OAI21_X1   g19909(.A1(new_n20100_), .A2(new_n20101_), .B(new_n19719_), .ZN(new_n20102_));
  INV_X1     g19910(.I(new_n20083_), .ZN(new_n20103_));
  OAI21_X1   g19911(.A1(new_n20100_), .A2(new_n20103_), .B(\asqrt[39] ), .ZN(new_n20104_));
  NAND3_X1   g19912(.A1(new_n20102_), .A2(new_n20104_), .A3(new_n3167_), .ZN(new_n20105_));
  NAND2_X1   g19913(.A1(new_n20105_), .A2(new_n19716_), .ZN(new_n20106_));
  NAND2_X1   g19914(.A1(new_n20102_), .A2(new_n20104_), .ZN(new_n20107_));
  AOI21_X1   g19915(.A1(new_n20107_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n20108_));
  AOI21_X1   g19916(.A1(new_n20108_), .A2(new_n20106_), .B(new_n20097_), .ZN(new_n20109_));
  AOI21_X1   g19917(.A1(new_n20106_), .A2(new_n20087_), .B(new_n2912_), .ZN(new_n20110_));
  OAI21_X1   g19918(.A1(new_n20109_), .A2(new_n20110_), .B(\asqrt[42] ), .ZN(new_n20111_));
  AOI21_X1   g19919(.A1(new_n20093_), .A2(new_n20111_), .B(new_n2464_), .ZN(new_n20112_));
  NOR2_X1    g19920(.A1(new_n20096_), .A2(new_n20112_), .ZN(new_n20113_));
  AOI21_X1   g19921(.A1(new_n20113_), .A2(new_n2271_), .B(new_n19705_), .ZN(new_n20114_));
  OAI21_X1   g19922(.A1(new_n20096_), .A2(new_n20112_), .B(\asqrt[44] ), .ZN(new_n20115_));
  NAND2_X1   g19923(.A1(new_n20115_), .A2(new_n2072_), .ZN(new_n20116_));
  OAI21_X1   g19924(.A1(new_n20114_), .A2(new_n20116_), .B(new_n19701_), .ZN(new_n20117_));
  INV_X1     g19925(.I(new_n20115_), .ZN(new_n20118_));
  OAI21_X1   g19926(.A1(new_n20114_), .A2(new_n20118_), .B(\asqrt[45] ), .ZN(new_n20119_));
  NAND3_X1   g19927(.A1(new_n20117_), .A2(new_n20119_), .A3(new_n1884_), .ZN(new_n20120_));
  NAND2_X1   g19928(.A1(new_n20120_), .A2(new_n19699_), .ZN(new_n20121_));
  NAND2_X1   g19929(.A1(new_n20117_), .A2(new_n20119_), .ZN(new_n20122_));
  AOI21_X1   g19930(.A1(new_n20122_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n20123_));
  AOI21_X1   g19931(.A1(new_n20123_), .A2(new_n20121_), .B(new_n19696_), .ZN(new_n20124_));
  INV_X1     g19932(.I(new_n19701_), .ZN(new_n20125_));
  INV_X1     g19933(.I(new_n19711_), .ZN(new_n20126_));
  NOR2_X1    g19934(.A1(new_n20109_), .A2(new_n20110_), .ZN(new_n20127_));
  AOI21_X1   g19935(.A1(new_n20127_), .A2(new_n2699_), .B(new_n20126_), .ZN(new_n20128_));
  NAND2_X1   g19936(.A1(new_n20111_), .A2(new_n2464_), .ZN(new_n20129_));
  OAI21_X1   g19937(.A1(new_n20128_), .A2(new_n20129_), .B(new_n19707_), .ZN(new_n20130_));
  INV_X1     g19938(.I(new_n20111_), .ZN(new_n20131_));
  OAI21_X1   g19939(.A1(new_n20128_), .A2(new_n20131_), .B(\asqrt[43] ), .ZN(new_n20132_));
  NAND3_X1   g19940(.A1(new_n20130_), .A2(new_n20132_), .A3(new_n2271_), .ZN(new_n20133_));
  NAND2_X1   g19941(.A1(new_n20133_), .A2(new_n19704_), .ZN(new_n20134_));
  NAND2_X1   g19942(.A1(new_n20130_), .A2(new_n20132_), .ZN(new_n20135_));
  AOI21_X1   g19943(.A1(new_n20135_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n20136_));
  AOI21_X1   g19944(.A1(new_n20136_), .A2(new_n20134_), .B(new_n20125_), .ZN(new_n20137_));
  AOI21_X1   g19945(.A1(new_n20134_), .A2(new_n20115_), .B(new_n2072_), .ZN(new_n20138_));
  OAI21_X1   g19946(.A1(new_n20137_), .A2(new_n20138_), .B(\asqrt[46] ), .ZN(new_n20139_));
  AOI21_X1   g19947(.A1(new_n20121_), .A2(new_n20139_), .B(new_n1688_), .ZN(new_n20140_));
  NOR2_X1    g19948(.A1(new_n20124_), .A2(new_n20140_), .ZN(new_n20141_));
  AOI21_X1   g19949(.A1(new_n20141_), .A2(new_n1533_), .B(new_n19693_), .ZN(new_n20142_));
  OAI21_X1   g19950(.A1(new_n20124_), .A2(new_n20140_), .B(\asqrt[48] ), .ZN(new_n20143_));
  NAND2_X1   g19951(.A1(new_n20143_), .A2(new_n1368_), .ZN(new_n20144_));
  OAI21_X1   g19952(.A1(new_n20142_), .A2(new_n20144_), .B(new_n19689_), .ZN(new_n20145_));
  INV_X1     g19953(.I(new_n20143_), .ZN(new_n20146_));
  OAI21_X1   g19954(.A1(new_n20142_), .A2(new_n20146_), .B(\asqrt[49] ), .ZN(new_n20147_));
  NAND3_X1   g19955(.A1(new_n20145_), .A2(new_n20147_), .A3(new_n1228_), .ZN(new_n20148_));
  NAND2_X1   g19956(.A1(new_n20148_), .A2(new_n19687_), .ZN(new_n20149_));
  NAND2_X1   g19957(.A1(new_n20145_), .A2(new_n20147_), .ZN(new_n20150_));
  AOI21_X1   g19958(.A1(new_n20150_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n20151_));
  AOI21_X1   g19959(.A1(new_n20151_), .A2(new_n20149_), .B(new_n19684_), .ZN(new_n20152_));
  INV_X1     g19960(.I(new_n19689_), .ZN(new_n20153_));
  INV_X1     g19961(.I(new_n19699_), .ZN(new_n20154_));
  NOR2_X1    g19962(.A1(new_n20137_), .A2(new_n20138_), .ZN(new_n20155_));
  AOI21_X1   g19963(.A1(new_n20155_), .A2(new_n1884_), .B(new_n20154_), .ZN(new_n20156_));
  NAND2_X1   g19964(.A1(new_n20139_), .A2(new_n1688_), .ZN(new_n20157_));
  OAI21_X1   g19965(.A1(new_n20156_), .A2(new_n20157_), .B(new_n19695_), .ZN(new_n20158_));
  INV_X1     g19966(.I(new_n20139_), .ZN(new_n20159_));
  OAI21_X1   g19967(.A1(new_n20156_), .A2(new_n20159_), .B(\asqrt[47] ), .ZN(new_n20160_));
  NAND3_X1   g19968(.A1(new_n20158_), .A2(new_n20160_), .A3(new_n1533_), .ZN(new_n20161_));
  NAND2_X1   g19969(.A1(new_n20161_), .A2(new_n19692_), .ZN(new_n20162_));
  NAND2_X1   g19970(.A1(new_n20158_), .A2(new_n20160_), .ZN(new_n20163_));
  AOI21_X1   g19971(.A1(new_n20163_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n20164_));
  AOI21_X1   g19972(.A1(new_n20164_), .A2(new_n20162_), .B(new_n20153_), .ZN(new_n20165_));
  AOI21_X1   g19973(.A1(new_n20162_), .A2(new_n20143_), .B(new_n1368_), .ZN(new_n20166_));
  OAI21_X1   g19974(.A1(new_n20165_), .A2(new_n20166_), .B(\asqrt[50] ), .ZN(new_n20167_));
  AOI21_X1   g19975(.A1(new_n20149_), .A2(new_n20167_), .B(new_n1088_), .ZN(new_n20168_));
  NOR2_X1    g19976(.A1(new_n20152_), .A2(new_n20168_), .ZN(new_n20169_));
  AOI21_X1   g19977(.A1(new_n20169_), .A2(new_n962_), .B(new_n19681_), .ZN(new_n20170_));
  OAI21_X1   g19978(.A1(new_n20152_), .A2(new_n20168_), .B(\asqrt[52] ), .ZN(new_n20171_));
  NAND2_X1   g19979(.A1(new_n20171_), .A2(new_n842_), .ZN(new_n20172_));
  OAI21_X1   g19980(.A1(new_n20170_), .A2(new_n20172_), .B(new_n19677_), .ZN(new_n20173_));
  INV_X1     g19981(.I(new_n20171_), .ZN(new_n20174_));
  OAI21_X1   g19982(.A1(new_n20170_), .A2(new_n20174_), .B(\asqrt[53] ), .ZN(new_n20175_));
  NAND3_X1   g19983(.A1(new_n20173_), .A2(new_n20175_), .A3(new_n720_), .ZN(new_n20176_));
  NAND2_X1   g19984(.A1(new_n20176_), .A2(new_n19675_), .ZN(new_n20177_));
  NAND2_X1   g19985(.A1(new_n20173_), .A2(new_n20175_), .ZN(new_n20178_));
  AOI21_X1   g19986(.A1(new_n20178_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n20179_));
  AOI21_X1   g19987(.A1(new_n20179_), .A2(new_n20177_), .B(new_n19672_), .ZN(new_n20180_));
  INV_X1     g19988(.I(new_n19677_), .ZN(new_n20181_));
  INV_X1     g19989(.I(new_n19687_), .ZN(new_n20182_));
  NOR2_X1    g19990(.A1(new_n20165_), .A2(new_n20166_), .ZN(new_n20183_));
  AOI21_X1   g19991(.A1(new_n20183_), .A2(new_n1228_), .B(new_n20182_), .ZN(new_n20184_));
  NAND2_X1   g19992(.A1(new_n20167_), .A2(new_n1088_), .ZN(new_n20185_));
  OAI21_X1   g19993(.A1(new_n20184_), .A2(new_n20185_), .B(new_n19683_), .ZN(new_n20186_));
  INV_X1     g19994(.I(new_n20167_), .ZN(new_n20187_));
  OAI21_X1   g19995(.A1(new_n20184_), .A2(new_n20187_), .B(\asqrt[51] ), .ZN(new_n20188_));
  NAND3_X1   g19996(.A1(new_n20186_), .A2(new_n20188_), .A3(new_n962_), .ZN(new_n20189_));
  NAND2_X1   g19997(.A1(new_n20189_), .A2(new_n19680_), .ZN(new_n20190_));
  NAND2_X1   g19998(.A1(new_n20186_), .A2(new_n20188_), .ZN(new_n20191_));
  AOI21_X1   g19999(.A1(new_n20191_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n20192_));
  AOI21_X1   g20000(.A1(new_n20192_), .A2(new_n20190_), .B(new_n20181_), .ZN(new_n20193_));
  AOI21_X1   g20001(.A1(new_n20190_), .A2(new_n20171_), .B(new_n842_), .ZN(new_n20194_));
  OAI21_X1   g20002(.A1(new_n20193_), .A2(new_n20194_), .B(\asqrt[54] ), .ZN(new_n20195_));
  AOI21_X1   g20003(.A1(new_n20177_), .A2(new_n20195_), .B(new_n630_), .ZN(new_n20196_));
  NOR2_X1    g20004(.A1(new_n20180_), .A2(new_n20196_), .ZN(new_n20197_));
  AOI21_X1   g20005(.A1(new_n20197_), .A2(new_n545_), .B(new_n19669_), .ZN(new_n20198_));
  OAI21_X1   g20006(.A1(new_n20180_), .A2(new_n20196_), .B(\asqrt[56] ), .ZN(new_n20199_));
  NAND2_X1   g20007(.A1(new_n20199_), .A2(new_n450_), .ZN(new_n20200_));
  OAI21_X1   g20008(.A1(new_n20198_), .A2(new_n20200_), .B(new_n19665_), .ZN(new_n20201_));
  INV_X1     g20009(.I(new_n20199_), .ZN(new_n20202_));
  OAI21_X1   g20010(.A1(new_n20198_), .A2(new_n20202_), .B(\asqrt[57] ), .ZN(new_n20203_));
  NAND3_X1   g20011(.A1(new_n20201_), .A2(new_n20203_), .A3(new_n403_), .ZN(new_n20204_));
  NAND2_X1   g20012(.A1(new_n20204_), .A2(new_n19663_), .ZN(new_n20205_));
  NAND2_X1   g20013(.A1(new_n20201_), .A2(new_n20203_), .ZN(new_n20206_));
  AOI21_X1   g20014(.A1(new_n20206_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n20207_));
  AOI21_X1   g20015(.A1(new_n20207_), .A2(new_n20205_), .B(new_n19660_), .ZN(new_n20208_));
  INV_X1     g20016(.I(new_n19665_), .ZN(new_n20209_));
  INV_X1     g20017(.I(new_n19675_), .ZN(new_n20210_));
  NOR2_X1    g20018(.A1(new_n20193_), .A2(new_n20194_), .ZN(new_n20211_));
  AOI21_X1   g20019(.A1(new_n20211_), .A2(new_n720_), .B(new_n20210_), .ZN(new_n20212_));
  NAND2_X1   g20020(.A1(new_n20195_), .A2(new_n630_), .ZN(new_n20213_));
  OAI21_X1   g20021(.A1(new_n20212_), .A2(new_n20213_), .B(new_n19671_), .ZN(new_n20214_));
  INV_X1     g20022(.I(new_n20195_), .ZN(new_n20215_));
  OAI21_X1   g20023(.A1(new_n20212_), .A2(new_n20215_), .B(\asqrt[55] ), .ZN(new_n20216_));
  NAND3_X1   g20024(.A1(new_n20214_), .A2(new_n20216_), .A3(new_n545_), .ZN(new_n20217_));
  NAND2_X1   g20025(.A1(new_n20217_), .A2(new_n19668_), .ZN(new_n20218_));
  NAND2_X1   g20026(.A1(new_n20214_), .A2(new_n20216_), .ZN(new_n20219_));
  AOI21_X1   g20027(.A1(new_n20219_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n20220_));
  AOI21_X1   g20028(.A1(new_n20220_), .A2(new_n20218_), .B(new_n20209_), .ZN(new_n20221_));
  AOI21_X1   g20029(.A1(new_n20218_), .A2(new_n20199_), .B(new_n450_), .ZN(new_n20222_));
  OAI21_X1   g20030(.A1(new_n20221_), .A2(new_n20222_), .B(\asqrt[58] ), .ZN(new_n20223_));
  AOI21_X1   g20031(.A1(new_n20205_), .A2(new_n20223_), .B(new_n339_), .ZN(new_n20224_));
  NOR2_X1    g20032(.A1(new_n20208_), .A2(new_n20224_), .ZN(new_n20225_));
  AOI21_X1   g20033(.A1(new_n20225_), .A2(new_n288_), .B(new_n19657_), .ZN(new_n20226_));
  OAI21_X1   g20034(.A1(new_n20208_), .A2(new_n20224_), .B(\asqrt[60] ), .ZN(new_n20227_));
  NAND2_X1   g20035(.A1(new_n20227_), .A2(new_n242_), .ZN(new_n20228_));
  OAI21_X1   g20036(.A1(new_n20226_), .A2(new_n20228_), .B(new_n19646_), .ZN(new_n20229_));
  INV_X1     g20037(.I(new_n20227_), .ZN(new_n20230_));
  OAI21_X1   g20038(.A1(new_n20226_), .A2(new_n20230_), .B(\asqrt[61] ), .ZN(new_n20231_));
  NAND3_X1   g20039(.A1(new_n20229_), .A2(new_n20231_), .A3(new_n234_), .ZN(new_n20232_));
  AOI21_X1   g20040(.A1(new_n20229_), .A2(new_n20231_), .B(new_n234_), .ZN(new_n20233_));
  AOI21_X1   g20041(.A1(new_n19644_), .A2(new_n20232_), .B(new_n20233_), .ZN(new_n20234_));
  NOR2_X1    g20042(.A1(new_n20234_), .A2(new_n19641_), .ZN(new_n20235_));
  INV_X1     g20043(.I(new_n19641_), .ZN(new_n20236_));
  INV_X1     g20044(.I(new_n20234_), .ZN(new_n20237_));
  NAND2_X1   g20045(.A1(new_n19651_), .A2(new_n19629_), .ZN(new_n20238_));
  NOR2_X1    g20046(.A1(new_n19653_), .A2(new_n19629_), .ZN(new_n20239_));
  NAND2_X1   g20047(.A1(new_n20239_), .A2(new_n19637_), .ZN(new_n20240_));
  AOI21_X1   g20048(.A1(new_n20240_), .A2(new_n20238_), .B(new_n193_), .ZN(new_n20241_));
  AOI21_X1   g20049(.A1(new_n20234_), .A2(new_n20236_), .B(new_n20241_), .ZN(new_n20242_));
  AOI21_X1   g20050(.A1(new_n20239_), .A2(new_n19651_), .B(new_n19652_), .ZN(new_n20243_));
  INV_X1     g20051(.I(new_n20243_), .ZN(new_n20244_));
  NOR3_X1    g20052(.A1(new_n20234_), .A2(new_n20236_), .A3(new_n20244_), .ZN(new_n20245_));
  OAI21_X1   g20053(.A1(\asqrt[63] ), .A2(new_n20245_), .B(new_n20242_), .ZN(\asqrt[1] ));
  INV_X1     g20054(.I(\asqrt[1] ), .ZN(new_n20247_));
  NOR3_X1    g20055(.A1(new_n20247_), .A2(new_n20236_), .A3(new_n20237_), .ZN(new_n20248_));
  OAI21_X1   g20056(.A1(new_n20248_), .A2(new_n20235_), .B(\asqrt[63] ), .ZN(new_n20249_));
  INV_X1     g20057(.I(new_n20232_), .ZN(new_n20250_));
  NOR3_X1    g20058(.A1(new_n20247_), .A2(new_n20250_), .A3(new_n20233_), .ZN(new_n20251_));
  XOR2_X1    g20059(.A1(new_n20251_), .A2(new_n19644_), .Z(new_n20252_));
  INV_X1     g20060(.I(new_n20252_), .ZN(new_n20253_));
  INV_X1     g20061(.I(new_n19646_), .ZN(new_n20254_));
  INV_X1     g20062(.I(new_n19663_), .ZN(new_n20255_));
  NOR2_X1    g20063(.A1(new_n20221_), .A2(new_n20222_), .ZN(new_n20256_));
  AOI21_X1   g20064(.A1(new_n20256_), .A2(new_n403_), .B(new_n20255_), .ZN(new_n20257_));
  NAND2_X1   g20065(.A1(new_n20223_), .A2(new_n339_), .ZN(new_n20258_));
  OAI21_X1   g20066(.A1(new_n20257_), .A2(new_n20258_), .B(new_n19659_), .ZN(new_n20259_));
  INV_X1     g20067(.I(new_n20223_), .ZN(new_n20260_));
  OAI21_X1   g20068(.A1(new_n20257_), .A2(new_n20260_), .B(\asqrt[59] ), .ZN(new_n20261_));
  NAND3_X1   g20069(.A1(new_n20259_), .A2(new_n20261_), .A3(new_n288_), .ZN(new_n20262_));
  NAND2_X1   g20070(.A1(new_n20262_), .A2(new_n19656_), .ZN(new_n20263_));
  NAND2_X1   g20071(.A1(new_n20259_), .A2(new_n20261_), .ZN(new_n20264_));
  AOI21_X1   g20072(.A1(new_n20264_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n20265_));
  AOI21_X1   g20073(.A1(new_n20263_), .A2(new_n20227_), .B(new_n242_), .ZN(new_n20266_));
  AOI21_X1   g20074(.A1(new_n20263_), .A2(new_n20265_), .B(new_n20266_), .ZN(new_n20267_));
  NAND2_X1   g20075(.A1(\asqrt[1] ), .A2(new_n20267_), .ZN(new_n20268_));
  XOR2_X1    g20076(.A1(new_n20268_), .A2(new_n20254_), .Z(new_n20269_));
  INV_X1     g20077(.I(new_n20269_), .ZN(new_n20270_));
  NAND3_X1   g20078(.A1(\asqrt[1] ), .A2(new_n20262_), .A3(new_n20227_), .ZN(new_n20271_));
  XOR2_X1    g20079(.A1(new_n20271_), .A2(new_n19657_), .Z(new_n20272_));
  OAI21_X1   g20080(.A1(new_n20257_), .A2(new_n20258_), .B(new_n20261_), .ZN(new_n20273_));
  NOR2_X1    g20081(.A1(new_n20247_), .A2(new_n20273_), .ZN(new_n20274_));
  XOR2_X1    g20082(.A1(new_n20274_), .A2(new_n19659_), .Z(new_n20275_));
  NAND3_X1   g20083(.A1(\asqrt[1] ), .A2(new_n20204_), .A3(new_n20223_), .ZN(new_n20276_));
  XOR2_X1    g20084(.A1(new_n20276_), .A2(new_n20255_), .Z(new_n20277_));
  INV_X1     g20085(.I(new_n20277_), .ZN(new_n20278_));
  OAI21_X1   g20086(.A1(new_n20198_), .A2(new_n20200_), .B(new_n20203_), .ZN(new_n20279_));
  NOR2_X1    g20087(.A1(new_n20247_), .A2(new_n20279_), .ZN(new_n20280_));
  XOR2_X1    g20088(.A1(new_n20280_), .A2(new_n19665_), .Z(new_n20281_));
  INV_X1     g20089(.I(new_n20281_), .ZN(new_n20282_));
  NAND3_X1   g20090(.A1(\asqrt[1] ), .A2(new_n20217_), .A3(new_n20199_), .ZN(new_n20283_));
  XOR2_X1    g20091(.A1(new_n20283_), .A2(new_n19669_), .Z(new_n20284_));
  OAI21_X1   g20092(.A1(new_n20212_), .A2(new_n20213_), .B(new_n20216_), .ZN(new_n20285_));
  NOR2_X1    g20093(.A1(new_n20247_), .A2(new_n20285_), .ZN(new_n20286_));
  XOR2_X1    g20094(.A1(new_n20286_), .A2(new_n19671_), .Z(new_n20287_));
  NAND3_X1   g20095(.A1(\asqrt[1] ), .A2(new_n20176_), .A3(new_n20195_), .ZN(new_n20288_));
  XOR2_X1    g20096(.A1(new_n20288_), .A2(new_n20210_), .Z(new_n20289_));
  INV_X1     g20097(.I(new_n20289_), .ZN(new_n20290_));
  OAI21_X1   g20098(.A1(new_n20170_), .A2(new_n20172_), .B(new_n20175_), .ZN(new_n20291_));
  NOR2_X1    g20099(.A1(new_n20247_), .A2(new_n20291_), .ZN(new_n20292_));
  XOR2_X1    g20100(.A1(new_n20292_), .A2(new_n19677_), .Z(new_n20293_));
  INV_X1     g20101(.I(new_n20293_), .ZN(new_n20294_));
  NAND3_X1   g20102(.A1(\asqrt[1] ), .A2(new_n20189_), .A3(new_n20171_), .ZN(new_n20295_));
  XOR2_X1    g20103(.A1(new_n20295_), .A2(new_n19681_), .Z(new_n20296_));
  OAI21_X1   g20104(.A1(new_n20184_), .A2(new_n20185_), .B(new_n20188_), .ZN(new_n20297_));
  NOR2_X1    g20105(.A1(new_n20247_), .A2(new_n20297_), .ZN(new_n20298_));
  XOR2_X1    g20106(.A1(new_n20298_), .A2(new_n19683_), .Z(new_n20299_));
  NAND3_X1   g20107(.A1(\asqrt[1] ), .A2(new_n20148_), .A3(new_n20167_), .ZN(new_n20300_));
  XOR2_X1    g20108(.A1(new_n20300_), .A2(new_n20182_), .Z(new_n20301_));
  INV_X1     g20109(.I(new_n20301_), .ZN(new_n20302_));
  OAI21_X1   g20110(.A1(new_n20142_), .A2(new_n20144_), .B(new_n20147_), .ZN(new_n20303_));
  NOR2_X1    g20111(.A1(new_n20247_), .A2(new_n20303_), .ZN(new_n20304_));
  XOR2_X1    g20112(.A1(new_n20304_), .A2(new_n19689_), .Z(new_n20305_));
  INV_X1     g20113(.I(new_n20305_), .ZN(new_n20306_));
  NAND3_X1   g20114(.A1(\asqrt[1] ), .A2(new_n20161_), .A3(new_n20143_), .ZN(new_n20307_));
  XOR2_X1    g20115(.A1(new_n20307_), .A2(new_n19693_), .Z(new_n20308_));
  OAI21_X1   g20116(.A1(new_n20156_), .A2(new_n20157_), .B(new_n20160_), .ZN(new_n20309_));
  NOR2_X1    g20117(.A1(new_n20247_), .A2(new_n20309_), .ZN(new_n20310_));
  XOR2_X1    g20118(.A1(new_n20310_), .A2(new_n19695_), .Z(new_n20311_));
  NAND3_X1   g20119(.A1(\asqrt[1] ), .A2(new_n20120_), .A3(new_n20139_), .ZN(new_n20312_));
  XOR2_X1    g20120(.A1(new_n20312_), .A2(new_n20154_), .Z(new_n20313_));
  INV_X1     g20121(.I(new_n20313_), .ZN(new_n20314_));
  OAI21_X1   g20122(.A1(new_n20114_), .A2(new_n20116_), .B(new_n20119_), .ZN(new_n20315_));
  NOR2_X1    g20123(.A1(new_n20247_), .A2(new_n20315_), .ZN(new_n20316_));
  XOR2_X1    g20124(.A1(new_n20316_), .A2(new_n19701_), .Z(new_n20317_));
  INV_X1     g20125(.I(new_n20317_), .ZN(new_n20318_));
  NAND3_X1   g20126(.A1(\asqrt[1] ), .A2(new_n20133_), .A3(new_n20115_), .ZN(new_n20319_));
  XOR2_X1    g20127(.A1(new_n20319_), .A2(new_n19705_), .Z(new_n20320_));
  OAI21_X1   g20128(.A1(new_n20128_), .A2(new_n20129_), .B(new_n20132_), .ZN(new_n20321_));
  NOR2_X1    g20129(.A1(new_n20247_), .A2(new_n20321_), .ZN(new_n20322_));
  XOR2_X1    g20130(.A1(new_n20322_), .A2(new_n19707_), .Z(new_n20323_));
  NAND3_X1   g20131(.A1(\asqrt[1] ), .A2(new_n20092_), .A3(new_n20111_), .ZN(new_n20324_));
  XOR2_X1    g20132(.A1(new_n20324_), .A2(new_n20126_), .Z(new_n20325_));
  INV_X1     g20133(.I(new_n20325_), .ZN(new_n20326_));
  OAI21_X1   g20134(.A1(new_n20086_), .A2(new_n20088_), .B(new_n20091_), .ZN(new_n20327_));
  NOR2_X1    g20135(.A1(new_n20247_), .A2(new_n20327_), .ZN(new_n20328_));
  XOR2_X1    g20136(.A1(new_n20328_), .A2(new_n19713_), .Z(new_n20329_));
  INV_X1     g20137(.I(new_n20329_), .ZN(new_n20330_));
  NAND3_X1   g20138(.A1(\asqrt[1] ), .A2(new_n20105_), .A3(new_n20087_), .ZN(new_n20331_));
  XOR2_X1    g20139(.A1(new_n20331_), .A2(new_n19717_), .Z(new_n20332_));
  OAI21_X1   g20140(.A1(new_n20100_), .A2(new_n20101_), .B(new_n20104_), .ZN(new_n20333_));
  NOR2_X1    g20141(.A1(new_n20247_), .A2(new_n20333_), .ZN(new_n20334_));
  XOR2_X1    g20142(.A1(new_n20334_), .A2(new_n19719_), .Z(new_n20335_));
  NAND3_X1   g20143(.A1(\asqrt[1] ), .A2(new_n20064_), .A3(new_n20083_), .ZN(new_n20336_));
  XOR2_X1    g20144(.A1(new_n20336_), .A2(new_n20098_), .Z(new_n20337_));
  INV_X1     g20145(.I(new_n20337_), .ZN(new_n20338_));
  OAI21_X1   g20146(.A1(new_n20058_), .A2(new_n20060_), .B(new_n20063_), .ZN(new_n20339_));
  NOR2_X1    g20147(.A1(new_n20247_), .A2(new_n20339_), .ZN(new_n20340_));
  XOR2_X1    g20148(.A1(new_n20340_), .A2(new_n19725_), .Z(new_n20341_));
  INV_X1     g20149(.I(new_n20341_), .ZN(new_n20342_));
  NAND3_X1   g20150(.A1(\asqrt[1] ), .A2(new_n20077_), .A3(new_n20059_), .ZN(new_n20343_));
  XOR2_X1    g20151(.A1(new_n20343_), .A2(new_n19729_), .Z(new_n20344_));
  OAI21_X1   g20152(.A1(new_n20072_), .A2(new_n20073_), .B(new_n20076_), .ZN(new_n20345_));
  NOR2_X1    g20153(.A1(new_n20247_), .A2(new_n20345_), .ZN(new_n20346_));
  XOR2_X1    g20154(.A1(new_n20346_), .A2(new_n19731_), .Z(new_n20347_));
  NAND3_X1   g20155(.A1(\asqrt[1] ), .A2(new_n20036_), .A3(new_n20055_), .ZN(new_n20348_));
  XOR2_X1    g20156(.A1(new_n20348_), .A2(new_n20070_), .Z(new_n20349_));
  INV_X1     g20157(.I(new_n20349_), .ZN(new_n20350_));
  OAI21_X1   g20158(.A1(new_n20030_), .A2(new_n20032_), .B(new_n20035_), .ZN(new_n20351_));
  NOR2_X1    g20159(.A1(new_n20247_), .A2(new_n20351_), .ZN(new_n20352_));
  XOR2_X1    g20160(.A1(new_n20352_), .A2(new_n19737_), .Z(new_n20353_));
  INV_X1     g20161(.I(new_n20353_), .ZN(new_n20354_));
  NAND3_X1   g20162(.A1(\asqrt[1] ), .A2(new_n20049_), .A3(new_n20031_), .ZN(new_n20355_));
  XOR2_X1    g20163(.A1(new_n20355_), .A2(new_n19741_), .Z(new_n20356_));
  OAI21_X1   g20164(.A1(new_n20044_), .A2(new_n20045_), .B(new_n20048_), .ZN(new_n20357_));
  NOR2_X1    g20165(.A1(new_n20247_), .A2(new_n20357_), .ZN(new_n20358_));
  XOR2_X1    g20166(.A1(new_n20358_), .A2(new_n19743_), .Z(new_n20359_));
  NAND3_X1   g20167(.A1(\asqrt[1] ), .A2(new_n20008_), .A3(new_n20027_), .ZN(new_n20360_));
  XOR2_X1    g20168(.A1(new_n20360_), .A2(new_n20042_), .Z(new_n20361_));
  INV_X1     g20169(.I(new_n20361_), .ZN(new_n20362_));
  OAI21_X1   g20170(.A1(new_n20002_), .A2(new_n20004_), .B(new_n20007_), .ZN(new_n20363_));
  NOR2_X1    g20171(.A1(new_n20247_), .A2(new_n20363_), .ZN(new_n20364_));
  XOR2_X1    g20172(.A1(new_n20364_), .A2(new_n19749_), .Z(new_n20365_));
  INV_X1     g20173(.I(new_n20365_), .ZN(new_n20366_));
  NAND3_X1   g20174(.A1(\asqrt[1] ), .A2(new_n20021_), .A3(new_n20003_), .ZN(new_n20367_));
  XOR2_X1    g20175(.A1(new_n20367_), .A2(new_n19753_), .Z(new_n20368_));
  OAI21_X1   g20176(.A1(new_n20016_), .A2(new_n20017_), .B(new_n20020_), .ZN(new_n20369_));
  NOR2_X1    g20177(.A1(new_n20247_), .A2(new_n20369_), .ZN(new_n20370_));
  XOR2_X1    g20178(.A1(new_n20370_), .A2(new_n19755_), .Z(new_n20371_));
  NAND3_X1   g20179(.A1(\asqrt[1] ), .A2(new_n19980_), .A3(new_n19999_), .ZN(new_n20372_));
  XOR2_X1    g20180(.A1(new_n20372_), .A2(new_n20014_), .Z(new_n20373_));
  INV_X1     g20181(.I(new_n20373_), .ZN(new_n20374_));
  OAI21_X1   g20182(.A1(new_n19974_), .A2(new_n19976_), .B(new_n19979_), .ZN(new_n20375_));
  NOR2_X1    g20183(.A1(new_n20247_), .A2(new_n20375_), .ZN(new_n20376_));
  XOR2_X1    g20184(.A1(new_n20376_), .A2(new_n19761_), .Z(new_n20377_));
  INV_X1     g20185(.I(new_n20377_), .ZN(new_n20378_));
  NAND3_X1   g20186(.A1(\asqrt[1] ), .A2(new_n19993_), .A3(new_n19975_), .ZN(new_n20379_));
  XOR2_X1    g20187(.A1(new_n20379_), .A2(new_n19765_), .Z(new_n20380_));
  OAI21_X1   g20188(.A1(new_n19988_), .A2(new_n19989_), .B(new_n19992_), .ZN(new_n20381_));
  NOR2_X1    g20189(.A1(new_n20247_), .A2(new_n20381_), .ZN(new_n20382_));
  XOR2_X1    g20190(.A1(new_n20382_), .A2(new_n19767_), .Z(new_n20383_));
  NAND3_X1   g20191(.A1(\asqrt[1] ), .A2(new_n19952_), .A3(new_n19971_), .ZN(new_n20384_));
  XOR2_X1    g20192(.A1(new_n20384_), .A2(new_n19986_), .Z(new_n20385_));
  INV_X1     g20193(.I(new_n20385_), .ZN(new_n20386_));
  OAI21_X1   g20194(.A1(new_n19946_), .A2(new_n19948_), .B(new_n19951_), .ZN(new_n20387_));
  NOR2_X1    g20195(.A1(new_n20247_), .A2(new_n20387_), .ZN(new_n20388_));
  XOR2_X1    g20196(.A1(new_n20388_), .A2(new_n19773_), .Z(new_n20389_));
  INV_X1     g20197(.I(new_n20389_), .ZN(new_n20390_));
  NAND3_X1   g20198(.A1(\asqrt[1] ), .A2(new_n19965_), .A3(new_n19947_), .ZN(new_n20391_));
  XOR2_X1    g20199(.A1(new_n20391_), .A2(new_n19777_), .Z(new_n20392_));
  OAI21_X1   g20200(.A1(new_n19960_), .A2(new_n19961_), .B(new_n19964_), .ZN(new_n20393_));
  NOR2_X1    g20201(.A1(new_n20247_), .A2(new_n20393_), .ZN(new_n20394_));
  XOR2_X1    g20202(.A1(new_n20394_), .A2(new_n19779_), .Z(new_n20395_));
  NAND3_X1   g20203(.A1(\asqrt[1] ), .A2(new_n19924_), .A3(new_n19943_), .ZN(new_n20396_));
  XOR2_X1    g20204(.A1(new_n20396_), .A2(new_n19958_), .Z(new_n20397_));
  INV_X1     g20205(.I(new_n20397_), .ZN(new_n20398_));
  OAI21_X1   g20206(.A1(new_n19918_), .A2(new_n19920_), .B(new_n19923_), .ZN(new_n20399_));
  NOR2_X1    g20207(.A1(new_n20247_), .A2(new_n20399_), .ZN(new_n20400_));
  XOR2_X1    g20208(.A1(new_n20400_), .A2(new_n19785_), .Z(new_n20401_));
  INV_X1     g20209(.I(new_n20401_), .ZN(new_n20402_));
  NAND3_X1   g20210(.A1(\asqrt[1] ), .A2(new_n19937_), .A3(new_n19919_), .ZN(new_n20403_));
  XOR2_X1    g20211(.A1(new_n20403_), .A2(new_n19789_), .Z(new_n20404_));
  OAI21_X1   g20212(.A1(new_n19932_), .A2(new_n19933_), .B(new_n19936_), .ZN(new_n20405_));
  NOR2_X1    g20213(.A1(new_n20247_), .A2(new_n20405_), .ZN(new_n20406_));
  XOR2_X1    g20214(.A1(new_n20406_), .A2(new_n19791_), .Z(new_n20407_));
  NAND3_X1   g20215(.A1(\asqrt[1] ), .A2(new_n19896_), .A3(new_n19915_), .ZN(new_n20408_));
  XOR2_X1    g20216(.A1(new_n20408_), .A2(new_n19930_), .Z(new_n20409_));
  INV_X1     g20217(.I(new_n20409_), .ZN(new_n20410_));
  OAI21_X1   g20218(.A1(new_n19890_), .A2(new_n19892_), .B(new_n19895_), .ZN(new_n20411_));
  NOR2_X1    g20219(.A1(new_n20247_), .A2(new_n20411_), .ZN(new_n20412_));
  XOR2_X1    g20220(.A1(new_n20412_), .A2(new_n19797_), .Z(new_n20413_));
  INV_X1     g20221(.I(new_n20413_), .ZN(new_n20414_));
  NAND3_X1   g20222(.A1(\asqrt[1] ), .A2(new_n19909_), .A3(new_n19891_), .ZN(new_n20415_));
  XOR2_X1    g20223(.A1(new_n20415_), .A2(new_n19801_), .Z(new_n20416_));
  OAI21_X1   g20224(.A1(new_n19904_), .A2(new_n19905_), .B(new_n19908_), .ZN(new_n20417_));
  NOR2_X1    g20225(.A1(new_n20247_), .A2(new_n20417_), .ZN(new_n20418_));
  XOR2_X1    g20226(.A1(new_n20418_), .A2(new_n19803_), .Z(new_n20419_));
  NAND3_X1   g20227(.A1(\asqrt[1] ), .A2(new_n19860_), .A3(new_n19887_), .ZN(new_n20420_));
  XOR2_X1    g20228(.A1(new_n20420_), .A2(new_n19902_), .Z(new_n20421_));
  INV_X1     g20229(.I(new_n20421_), .ZN(new_n20422_));
  OAI21_X1   g20230(.A1(new_n19854_), .A2(new_n19856_), .B(new_n19859_), .ZN(new_n20423_));
  NOR2_X1    g20231(.A1(new_n20247_), .A2(new_n20423_), .ZN(new_n20424_));
  XOR2_X1    g20232(.A1(new_n20424_), .A2(new_n19809_), .Z(new_n20425_));
  INV_X1     g20233(.I(new_n20425_), .ZN(new_n20426_));
  NAND3_X1   g20234(.A1(\asqrt[1] ), .A2(new_n19881_), .A3(new_n19855_), .ZN(new_n20427_));
  XOR2_X1    g20235(.A1(new_n20427_), .A2(new_n19813_), .Z(new_n20428_));
  OAI21_X1   g20236(.A1(new_n19876_), .A2(new_n19877_), .B(new_n19880_), .ZN(new_n20429_));
  NOR2_X1    g20237(.A1(new_n20247_), .A2(new_n20429_), .ZN(new_n20430_));
  XOR2_X1    g20238(.A1(new_n20430_), .A2(new_n19816_), .Z(new_n20431_));
  NAND2_X1   g20239(.A1(new_n19875_), .A2(new_n17242_), .ZN(new_n20432_));
  NAND3_X1   g20240(.A1(\asqrt[1] ), .A2(new_n20432_), .A3(new_n19851_), .ZN(new_n20433_));
  XOR2_X1    g20241(.A1(new_n20433_), .A2(new_n19866_), .Z(new_n20434_));
  INV_X1     g20242(.I(new_n20434_), .ZN(new_n20435_));
  NAND3_X1   g20243(.A1(\asqrt[1] ), .A2(new_n19873_), .A3(new_n19846_), .ZN(new_n20436_));
  XOR2_X1    g20244(.A1(new_n20436_), .A2(new_n19845_), .Z(new_n20437_));
  INV_X1     g20245(.I(new_n20437_), .ZN(new_n20438_));
  NAND3_X1   g20246(.A1(\asqrt[1] ), .A2(new_n19870_), .A3(new_n19872_), .ZN(new_n20439_));
  XOR2_X1    g20247(.A1(new_n20439_), .A2(new_n19828_), .Z(new_n20440_));
  NOR2_X1    g20248(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n20441_));
  NOR2_X1    g20249(.A1(new_n20441_), .A2(\a[2] ), .ZN(new_n20442_));
  AOI21_X1   g20250(.A1(new_n20247_), .A2(\a[2] ), .B(new_n20442_), .ZN(new_n20443_));
  INV_X1     g20251(.I(new_n19829_), .ZN(new_n20444_));
  INV_X1     g20252(.I(new_n19644_), .ZN(new_n20445_));
  AOI21_X1   g20253(.A1(new_n20265_), .A2(new_n20263_), .B(new_n20254_), .ZN(new_n20446_));
  NOR2_X1    g20254(.A1(new_n20446_), .A2(new_n20266_), .ZN(new_n20447_));
  AOI21_X1   g20255(.A1(new_n20447_), .A2(new_n234_), .B(new_n20445_), .ZN(new_n20448_));
  OAI21_X1   g20256(.A1(new_n20448_), .A2(new_n20233_), .B(new_n20243_), .ZN(new_n20449_));
  OAI21_X1   g20257(.A1(new_n20449_), .A2(new_n20236_), .B(new_n193_), .ZN(new_n20450_));
  AOI21_X1   g20258(.A1(new_n20450_), .A2(new_n20242_), .B(new_n20444_), .ZN(new_n20451_));
  INV_X1     g20259(.I(\a[2] ), .ZN(new_n20452_));
  INV_X1     g20260(.I(\a[3] ), .ZN(new_n20453_));
  AOI21_X1   g20261(.A1(\asqrt[1] ), .A2(new_n20452_), .B(new_n20453_), .ZN(new_n20454_));
  OAI21_X1   g20262(.A1(new_n20454_), .A2(new_n20451_), .B(new_n19653_), .ZN(new_n20455_));
  NOR3_X1    g20263(.A1(new_n20454_), .A2(new_n19653_), .A3(new_n20451_), .ZN(new_n20456_));
  AOI21_X1   g20264(.A1(new_n20443_), .A2(new_n20455_), .B(new_n20456_), .ZN(new_n20457_));
  NAND2_X1   g20265(.A1(new_n20457_), .A2(new_n19173_), .ZN(new_n20458_));
  NOR2_X1    g20266(.A1(\asqrt[1] ), .A2(new_n19653_), .ZN(new_n20459_));
  OAI21_X1   g20267(.A1(new_n20459_), .A2(new_n20451_), .B(new_n19824_), .ZN(new_n20460_));
  NAND2_X1   g20268(.A1(\asqrt[1] ), .A2(new_n19829_), .ZN(new_n20461_));
  NAND3_X1   g20269(.A1(new_n20450_), .A2(\asqrt[2] ), .A3(new_n20242_), .ZN(new_n20462_));
  NAND3_X1   g20270(.A1(new_n20461_), .A2(new_n20462_), .A3(\a[4] ), .ZN(new_n20463_));
  NAND2_X1   g20271(.A1(new_n20460_), .A2(new_n20463_), .ZN(new_n20464_));
  OAI21_X1   g20272(.A1(new_n20457_), .A2(new_n19173_), .B(new_n20464_), .ZN(new_n20465_));
  AND3_X2    g20273(.A1(\asqrt[1] ), .A2(new_n19868_), .A3(new_n19837_), .Z(new_n20466_));
  XOR2_X1    g20274(.A1(new_n20466_), .A2(new_n19836_), .Z(new_n20467_));
  AOI21_X1   g20275(.A1(new_n20465_), .A2(new_n20458_), .B(new_n20467_), .ZN(new_n20468_));
  INV_X1     g20276(.I(new_n20468_), .ZN(new_n20469_));
  NAND3_X1   g20277(.A1(new_n20465_), .A2(new_n20458_), .A3(new_n20467_), .ZN(new_n20470_));
  NAND2_X1   g20278(.A1(new_n20470_), .A2(new_n18424_), .ZN(new_n20471_));
  AOI21_X1   g20279(.A1(new_n20471_), .A2(new_n20469_), .B(new_n20440_), .ZN(new_n20472_));
  AOI21_X1   g20280(.A1(new_n18424_), .A2(new_n20470_), .B(new_n20468_), .ZN(new_n20473_));
  AOI21_X1   g20281(.A1(new_n20473_), .A2(new_n20440_), .B(\asqrt[5] ), .ZN(new_n20474_));
  OAI21_X1   g20282(.A1(new_n20474_), .A2(new_n20472_), .B(new_n20438_), .ZN(new_n20475_));
  NOR3_X1    g20283(.A1(new_n20474_), .A2(new_n20438_), .A3(new_n20472_), .ZN(new_n20476_));
  OAI21_X1   g20284(.A1(\asqrt[6] ), .A2(new_n20476_), .B(new_n20475_), .ZN(new_n20477_));
  NAND2_X1   g20285(.A1(new_n20477_), .A2(new_n20435_), .ZN(new_n20478_));
  OAI21_X1   g20286(.A1(new_n20477_), .A2(new_n20435_), .B(new_n16649_), .ZN(new_n20479_));
  AOI21_X1   g20287(.A1(new_n20479_), .A2(new_n20478_), .B(new_n20431_), .ZN(new_n20480_));
  INV_X1     g20288(.I(new_n20480_), .ZN(new_n20481_));
  NAND3_X1   g20289(.A1(new_n20479_), .A2(new_n20478_), .A3(new_n20431_), .ZN(new_n20482_));
  NAND2_X1   g20290(.A1(new_n20482_), .A2(new_n16093_), .ZN(new_n20483_));
  AOI21_X1   g20291(.A1(new_n20483_), .A2(new_n20481_), .B(new_n20428_), .ZN(new_n20484_));
  AOI21_X1   g20292(.A1(new_n16093_), .A2(new_n20482_), .B(new_n20480_), .ZN(new_n20485_));
  AOI21_X1   g20293(.A1(new_n20485_), .A2(new_n20428_), .B(\asqrt[9] ), .ZN(new_n20486_));
  OAI21_X1   g20294(.A1(new_n20486_), .A2(new_n20484_), .B(new_n20426_), .ZN(new_n20487_));
  NOR3_X1    g20295(.A1(new_n20486_), .A2(new_n20426_), .A3(new_n20484_), .ZN(new_n20488_));
  OAI21_X1   g20296(.A1(\asqrt[10] ), .A2(new_n20488_), .B(new_n20487_), .ZN(new_n20489_));
  NAND2_X1   g20297(.A1(new_n20489_), .A2(new_n20422_), .ZN(new_n20490_));
  OAI21_X1   g20298(.A1(new_n20489_), .A2(new_n20422_), .B(new_n14430_), .ZN(new_n20491_));
  AOI21_X1   g20299(.A1(new_n20491_), .A2(new_n20490_), .B(new_n20419_), .ZN(new_n20492_));
  INV_X1     g20300(.I(new_n20492_), .ZN(new_n20493_));
  NAND3_X1   g20301(.A1(new_n20491_), .A2(new_n20490_), .A3(new_n20419_), .ZN(new_n20494_));
  NAND2_X1   g20302(.A1(new_n20494_), .A2(new_n13917_), .ZN(new_n20495_));
  AOI21_X1   g20303(.A1(new_n20495_), .A2(new_n20493_), .B(new_n20416_), .ZN(new_n20496_));
  AOI21_X1   g20304(.A1(new_n13917_), .A2(new_n20494_), .B(new_n20492_), .ZN(new_n20497_));
  AOI21_X1   g20305(.A1(new_n20497_), .A2(new_n20416_), .B(\asqrt[13] ), .ZN(new_n20498_));
  OAI21_X1   g20306(.A1(new_n20498_), .A2(new_n20496_), .B(new_n20414_), .ZN(new_n20499_));
  NOR3_X1    g20307(.A1(new_n20498_), .A2(new_n20414_), .A3(new_n20496_), .ZN(new_n20500_));
  OAI21_X1   g20308(.A1(\asqrt[14] ), .A2(new_n20500_), .B(new_n20499_), .ZN(new_n20501_));
  NAND2_X1   g20309(.A1(new_n20501_), .A2(new_n20410_), .ZN(new_n20502_));
  OAI21_X1   g20310(.A1(new_n20501_), .A2(new_n20410_), .B(new_n12374_), .ZN(new_n20503_));
  AOI21_X1   g20311(.A1(new_n20503_), .A2(new_n20502_), .B(new_n20407_), .ZN(new_n20504_));
  INV_X1     g20312(.I(new_n20504_), .ZN(new_n20505_));
  NAND3_X1   g20313(.A1(new_n20503_), .A2(new_n20502_), .A3(new_n20407_), .ZN(new_n20506_));
  NAND2_X1   g20314(.A1(new_n20506_), .A2(new_n11901_), .ZN(new_n20507_));
  AOI21_X1   g20315(.A1(new_n20507_), .A2(new_n20505_), .B(new_n20404_), .ZN(new_n20508_));
  AOI21_X1   g20316(.A1(new_n11901_), .A2(new_n20506_), .B(new_n20504_), .ZN(new_n20509_));
  AOI21_X1   g20317(.A1(new_n20509_), .A2(new_n20404_), .B(\asqrt[17] ), .ZN(new_n20510_));
  OAI21_X1   g20318(.A1(new_n20510_), .A2(new_n20508_), .B(new_n20402_), .ZN(new_n20511_));
  NOR3_X1    g20319(.A1(new_n20510_), .A2(new_n20402_), .A3(new_n20508_), .ZN(new_n20512_));
  OAI21_X1   g20320(.A1(\asqrt[18] ), .A2(new_n20512_), .B(new_n20511_), .ZN(new_n20513_));
  NAND2_X1   g20321(.A1(new_n20513_), .A2(new_n20398_), .ZN(new_n20514_));
  OAI21_X1   g20322(.A1(new_n20513_), .A2(new_n20398_), .B(new_n10478_), .ZN(new_n20515_));
  AOI21_X1   g20323(.A1(new_n20515_), .A2(new_n20514_), .B(new_n20395_), .ZN(new_n20516_));
  INV_X1     g20324(.I(new_n20516_), .ZN(new_n20517_));
  NAND3_X1   g20325(.A1(new_n20515_), .A2(new_n20514_), .A3(new_n20395_), .ZN(new_n20518_));
  NAND2_X1   g20326(.A1(new_n20518_), .A2(new_n10045_), .ZN(new_n20519_));
  AOI21_X1   g20327(.A1(new_n20519_), .A2(new_n20517_), .B(new_n20392_), .ZN(new_n20520_));
  AOI21_X1   g20328(.A1(new_n10045_), .A2(new_n20518_), .B(new_n20516_), .ZN(new_n20521_));
  AOI21_X1   g20329(.A1(new_n20521_), .A2(new_n20392_), .B(\asqrt[21] ), .ZN(new_n20522_));
  OAI21_X1   g20330(.A1(new_n20522_), .A2(new_n20520_), .B(new_n20390_), .ZN(new_n20523_));
  NOR3_X1    g20331(.A1(new_n20522_), .A2(new_n20390_), .A3(new_n20520_), .ZN(new_n20524_));
  OAI21_X1   g20332(.A1(\asqrt[22] ), .A2(new_n20524_), .B(new_n20523_), .ZN(new_n20525_));
  NAND2_X1   g20333(.A1(new_n20525_), .A2(new_n20386_), .ZN(new_n20526_));
  OAI21_X1   g20334(.A1(new_n20525_), .A2(new_n20386_), .B(new_n8742_), .ZN(new_n20527_));
  AOI21_X1   g20335(.A1(new_n20527_), .A2(new_n20526_), .B(new_n20383_), .ZN(new_n20528_));
  INV_X1     g20336(.I(new_n20528_), .ZN(new_n20529_));
  NAND3_X1   g20337(.A1(new_n20527_), .A2(new_n20526_), .A3(new_n20383_), .ZN(new_n20530_));
  NAND2_X1   g20338(.A1(new_n20530_), .A2(new_n8349_), .ZN(new_n20531_));
  AOI21_X1   g20339(.A1(new_n20531_), .A2(new_n20529_), .B(new_n20380_), .ZN(new_n20532_));
  AOI21_X1   g20340(.A1(new_n8349_), .A2(new_n20530_), .B(new_n20528_), .ZN(new_n20533_));
  AOI21_X1   g20341(.A1(new_n20533_), .A2(new_n20380_), .B(\asqrt[25] ), .ZN(new_n20534_));
  OAI21_X1   g20342(.A1(new_n20534_), .A2(new_n20532_), .B(new_n20378_), .ZN(new_n20535_));
  NOR3_X1    g20343(.A1(new_n20534_), .A2(new_n20378_), .A3(new_n20532_), .ZN(new_n20536_));
  OAI21_X1   g20344(.A1(\asqrt[26] ), .A2(new_n20536_), .B(new_n20535_), .ZN(new_n20537_));
  NAND2_X1   g20345(.A1(new_n20537_), .A2(new_n20374_), .ZN(new_n20538_));
  OAI21_X1   g20346(.A1(new_n20537_), .A2(new_n20374_), .B(new_n7166_), .ZN(new_n20539_));
  AOI21_X1   g20347(.A1(new_n20539_), .A2(new_n20538_), .B(new_n20371_), .ZN(new_n20540_));
  INV_X1     g20348(.I(new_n20540_), .ZN(new_n20541_));
  NAND3_X1   g20349(.A1(new_n20539_), .A2(new_n20538_), .A3(new_n20371_), .ZN(new_n20542_));
  NAND2_X1   g20350(.A1(new_n20542_), .A2(new_n6813_), .ZN(new_n20543_));
  AOI21_X1   g20351(.A1(new_n20543_), .A2(new_n20541_), .B(new_n20368_), .ZN(new_n20544_));
  AOI21_X1   g20352(.A1(new_n6813_), .A2(new_n20542_), .B(new_n20540_), .ZN(new_n20545_));
  AOI21_X1   g20353(.A1(new_n20545_), .A2(new_n20368_), .B(\asqrt[29] ), .ZN(new_n20546_));
  OAI21_X1   g20354(.A1(new_n20546_), .A2(new_n20544_), .B(new_n20366_), .ZN(new_n20547_));
  NOR3_X1    g20355(.A1(new_n20546_), .A2(new_n20366_), .A3(new_n20544_), .ZN(new_n20548_));
  OAI21_X1   g20356(.A1(\asqrt[30] ), .A2(new_n20548_), .B(new_n20547_), .ZN(new_n20549_));
  NAND2_X1   g20357(.A1(new_n20549_), .A2(new_n20362_), .ZN(new_n20550_));
  OAI21_X1   g20358(.A1(new_n20549_), .A2(new_n20362_), .B(new_n5750_), .ZN(new_n20551_));
  AOI21_X1   g20359(.A1(new_n20551_), .A2(new_n20550_), .B(new_n20359_), .ZN(new_n20552_));
  INV_X1     g20360(.I(new_n20552_), .ZN(new_n20553_));
  NAND3_X1   g20361(.A1(new_n20551_), .A2(new_n20550_), .A3(new_n20359_), .ZN(new_n20554_));
  NAND2_X1   g20362(.A1(new_n20554_), .A2(new_n5435_), .ZN(new_n20555_));
  AOI21_X1   g20363(.A1(new_n20555_), .A2(new_n20553_), .B(new_n20356_), .ZN(new_n20556_));
  AOI21_X1   g20364(.A1(new_n5435_), .A2(new_n20554_), .B(new_n20552_), .ZN(new_n20557_));
  AOI21_X1   g20365(.A1(new_n20557_), .A2(new_n20356_), .B(\asqrt[33] ), .ZN(new_n20558_));
  OAI21_X1   g20366(.A1(new_n20558_), .A2(new_n20556_), .B(new_n20354_), .ZN(new_n20559_));
  NOR3_X1    g20367(.A1(new_n20558_), .A2(new_n20354_), .A3(new_n20556_), .ZN(new_n20560_));
  OAI21_X1   g20368(.A1(\asqrt[34] ), .A2(new_n20560_), .B(new_n20559_), .ZN(new_n20561_));
  NAND2_X1   g20369(.A1(new_n20561_), .A2(new_n20350_), .ZN(new_n20562_));
  OAI21_X1   g20370(.A1(new_n20561_), .A2(new_n20350_), .B(new_n4510_), .ZN(new_n20563_));
  AOI21_X1   g20371(.A1(new_n20563_), .A2(new_n20562_), .B(new_n20347_), .ZN(new_n20564_));
  INV_X1     g20372(.I(new_n20564_), .ZN(new_n20565_));
  NAND3_X1   g20373(.A1(new_n20563_), .A2(new_n20562_), .A3(new_n20347_), .ZN(new_n20566_));
  NAND2_X1   g20374(.A1(new_n20566_), .A2(new_n4224_), .ZN(new_n20567_));
  AOI21_X1   g20375(.A1(new_n20567_), .A2(new_n20565_), .B(new_n20344_), .ZN(new_n20568_));
  AOI21_X1   g20376(.A1(new_n4224_), .A2(new_n20566_), .B(new_n20564_), .ZN(new_n20569_));
  AOI21_X1   g20377(.A1(new_n20569_), .A2(new_n20344_), .B(\asqrt[37] ), .ZN(new_n20570_));
  OAI21_X1   g20378(.A1(new_n20570_), .A2(new_n20568_), .B(new_n20342_), .ZN(new_n20571_));
  NOR3_X1    g20379(.A1(new_n20570_), .A2(new_n20342_), .A3(new_n20568_), .ZN(new_n20572_));
  OAI21_X1   g20380(.A1(\asqrt[38] ), .A2(new_n20572_), .B(new_n20571_), .ZN(new_n20573_));
  NAND2_X1   g20381(.A1(new_n20573_), .A2(new_n20338_), .ZN(new_n20574_));
  OAI21_X1   g20382(.A1(new_n20573_), .A2(new_n20338_), .B(new_n3400_), .ZN(new_n20575_));
  AOI21_X1   g20383(.A1(new_n20575_), .A2(new_n20574_), .B(new_n20335_), .ZN(new_n20576_));
  INV_X1     g20384(.I(new_n20576_), .ZN(new_n20577_));
  NAND3_X1   g20385(.A1(new_n20575_), .A2(new_n20574_), .A3(new_n20335_), .ZN(new_n20578_));
  NAND2_X1   g20386(.A1(new_n20578_), .A2(new_n3167_), .ZN(new_n20579_));
  AOI21_X1   g20387(.A1(new_n20579_), .A2(new_n20577_), .B(new_n20332_), .ZN(new_n20580_));
  AOI21_X1   g20388(.A1(new_n3167_), .A2(new_n20578_), .B(new_n20576_), .ZN(new_n20581_));
  AOI21_X1   g20389(.A1(new_n20581_), .A2(new_n20332_), .B(\asqrt[41] ), .ZN(new_n20582_));
  OAI21_X1   g20390(.A1(new_n20582_), .A2(new_n20580_), .B(new_n20330_), .ZN(new_n20583_));
  NOR3_X1    g20391(.A1(new_n20582_), .A2(new_n20330_), .A3(new_n20580_), .ZN(new_n20584_));
  OAI21_X1   g20392(.A1(\asqrt[42] ), .A2(new_n20584_), .B(new_n20583_), .ZN(new_n20585_));
  NAND2_X1   g20393(.A1(new_n20585_), .A2(new_n20326_), .ZN(new_n20586_));
  OAI21_X1   g20394(.A1(new_n20585_), .A2(new_n20326_), .B(new_n2464_), .ZN(new_n20587_));
  AOI21_X1   g20395(.A1(new_n20587_), .A2(new_n20586_), .B(new_n20323_), .ZN(new_n20588_));
  INV_X1     g20396(.I(new_n20588_), .ZN(new_n20589_));
  NAND3_X1   g20397(.A1(new_n20587_), .A2(new_n20586_), .A3(new_n20323_), .ZN(new_n20590_));
  NAND2_X1   g20398(.A1(new_n20590_), .A2(new_n2271_), .ZN(new_n20591_));
  AOI21_X1   g20399(.A1(new_n20591_), .A2(new_n20589_), .B(new_n20320_), .ZN(new_n20592_));
  AOI21_X1   g20400(.A1(new_n2271_), .A2(new_n20590_), .B(new_n20588_), .ZN(new_n20593_));
  AOI21_X1   g20401(.A1(new_n20593_), .A2(new_n20320_), .B(\asqrt[45] ), .ZN(new_n20594_));
  OAI21_X1   g20402(.A1(new_n20594_), .A2(new_n20592_), .B(new_n20318_), .ZN(new_n20595_));
  NOR3_X1    g20403(.A1(new_n20594_), .A2(new_n20318_), .A3(new_n20592_), .ZN(new_n20596_));
  OAI21_X1   g20404(.A1(\asqrt[46] ), .A2(new_n20596_), .B(new_n20595_), .ZN(new_n20597_));
  NAND2_X1   g20405(.A1(new_n20597_), .A2(new_n20314_), .ZN(new_n20598_));
  OAI21_X1   g20406(.A1(new_n20597_), .A2(new_n20314_), .B(new_n1688_), .ZN(new_n20599_));
  AOI21_X1   g20407(.A1(new_n20599_), .A2(new_n20598_), .B(new_n20311_), .ZN(new_n20600_));
  INV_X1     g20408(.I(new_n20600_), .ZN(new_n20601_));
  NAND3_X1   g20409(.A1(new_n20599_), .A2(new_n20598_), .A3(new_n20311_), .ZN(new_n20602_));
  NAND2_X1   g20410(.A1(new_n20602_), .A2(new_n1533_), .ZN(new_n20603_));
  AOI21_X1   g20411(.A1(new_n20603_), .A2(new_n20601_), .B(new_n20308_), .ZN(new_n20604_));
  AOI21_X1   g20412(.A1(new_n1533_), .A2(new_n20602_), .B(new_n20600_), .ZN(new_n20605_));
  AOI21_X1   g20413(.A1(new_n20605_), .A2(new_n20308_), .B(\asqrt[49] ), .ZN(new_n20606_));
  OAI21_X1   g20414(.A1(new_n20606_), .A2(new_n20604_), .B(new_n20306_), .ZN(new_n20607_));
  NOR3_X1    g20415(.A1(new_n20606_), .A2(new_n20306_), .A3(new_n20604_), .ZN(new_n20608_));
  OAI21_X1   g20416(.A1(\asqrt[50] ), .A2(new_n20608_), .B(new_n20607_), .ZN(new_n20609_));
  NAND2_X1   g20417(.A1(new_n20609_), .A2(new_n20302_), .ZN(new_n20610_));
  OAI21_X1   g20418(.A1(new_n20609_), .A2(new_n20302_), .B(new_n1088_), .ZN(new_n20611_));
  AOI21_X1   g20419(.A1(new_n20611_), .A2(new_n20610_), .B(new_n20299_), .ZN(new_n20612_));
  INV_X1     g20420(.I(new_n20612_), .ZN(new_n20613_));
  NAND3_X1   g20421(.A1(new_n20611_), .A2(new_n20610_), .A3(new_n20299_), .ZN(new_n20614_));
  NAND2_X1   g20422(.A1(new_n20614_), .A2(new_n962_), .ZN(new_n20615_));
  AOI21_X1   g20423(.A1(new_n20615_), .A2(new_n20613_), .B(new_n20296_), .ZN(new_n20616_));
  AOI21_X1   g20424(.A1(new_n962_), .A2(new_n20614_), .B(new_n20612_), .ZN(new_n20617_));
  AOI21_X1   g20425(.A1(new_n20617_), .A2(new_n20296_), .B(\asqrt[53] ), .ZN(new_n20618_));
  OAI21_X1   g20426(.A1(new_n20618_), .A2(new_n20616_), .B(new_n20294_), .ZN(new_n20619_));
  NOR3_X1    g20427(.A1(new_n20618_), .A2(new_n20294_), .A3(new_n20616_), .ZN(new_n20620_));
  OAI21_X1   g20428(.A1(\asqrt[54] ), .A2(new_n20620_), .B(new_n20619_), .ZN(new_n20621_));
  NAND2_X1   g20429(.A1(new_n20621_), .A2(new_n20290_), .ZN(new_n20622_));
  OAI21_X1   g20430(.A1(new_n20621_), .A2(new_n20290_), .B(new_n630_), .ZN(new_n20623_));
  AOI21_X1   g20431(.A1(new_n20623_), .A2(new_n20622_), .B(new_n20287_), .ZN(new_n20624_));
  INV_X1     g20432(.I(new_n20624_), .ZN(new_n20625_));
  NAND3_X1   g20433(.A1(new_n20623_), .A2(new_n20622_), .A3(new_n20287_), .ZN(new_n20626_));
  NAND2_X1   g20434(.A1(new_n20626_), .A2(new_n545_), .ZN(new_n20627_));
  AOI21_X1   g20435(.A1(new_n20627_), .A2(new_n20625_), .B(new_n20284_), .ZN(new_n20628_));
  AOI21_X1   g20436(.A1(new_n545_), .A2(new_n20626_), .B(new_n20624_), .ZN(new_n20629_));
  AOI21_X1   g20437(.A1(new_n20629_), .A2(new_n20284_), .B(\asqrt[57] ), .ZN(new_n20630_));
  OAI21_X1   g20438(.A1(new_n20630_), .A2(new_n20628_), .B(new_n20282_), .ZN(new_n20631_));
  NOR3_X1    g20439(.A1(new_n20630_), .A2(new_n20282_), .A3(new_n20628_), .ZN(new_n20632_));
  OAI21_X1   g20440(.A1(\asqrt[58] ), .A2(new_n20632_), .B(new_n20631_), .ZN(new_n20633_));
  NAND2_X1   g20441(.A1(new_n20633_), .A2(new_n20278_), .ZN(new_n20634_));
  OAI21_X1   g20442(.A1(new_n20633_), .A2(new_n20278_), .B(new_n339_), .ZN(new_n20635_));
  AOI21_X1   g20443(.A1(new_n20635_), .A2(new_n20634_), .B(new_n20275_), .ZN(new_n20636_));
  INV_X1     g20444(.I(new_n20636_), .ZN(new_n20637_));
  NAND3_X1   g20445(.A1(new_n20635_), .A2(new_n20634_), .A3(new_n20275_), .ZN(new_n20638_));
  NAND2_X1   g20446(.A1(new_n20638_), .A2(new_n288_), .ZN(new_n20639_));
  AOI21_X1   g20447(.A1(new_n20639_), .A2(new_n20637_), .B(new_n20272_), .ZN(new_n20640_));
  AOI21_X1   g20448(.A1(new_n288_), .A2(new_n20638_), .B(new_n20636_), .ZN(new_n20641_));
  AOI21_X1   g20449(.A1(new_n20641_), .A2(new_n20272_), .B(\asqrt[61] ), .ZN(new_n20642_));
  OAI21_X1   g20450(.A1(new_n20642_), .A2(new_n20640_), .B(new_n20270_), .ZN(new_n20643_));
  INV_X1     g20451(.I(new_n20643_), .ZN(new_n20644_));
  NOR3_X1    g20452(.A1(new_n20642_), .A2(new_n20270_), .A3(new_n20640_), .ZN(new_n20645_));
  NOR2_X1    g20453(.A1(new_n20645_), .A2(\asqrt[62] ), .ZN(new_n20646_));
  OAI21_X1   g20454(.A1(new_n20646_), .A2(new_n20644_), .B(new_n20253_), .ZN(new_n20647_));
  OAI21_X1   g20455(.A1(\asqrt[62] ), .A2(new_n20645_), .B(new_n20643_), .ZN(new_n20648_));
  NAND2_X1   g20456(.A1(new_n20234_), .A2(new_n20236_), .ZN(new_n20649_));
  NAND3_X1   g20457(.A1(\asqrt[1] ), .A2(new_n19641_), .A3(new_n20237_), .ZN(new_n20650_));
  NAND3_X1   g20458(.A1(new_n20252_), .A2(new_n20649_), .A3(new_n20650_), .ZN(new_n20651_));
  OAI21_X1   g20459(.A1(new_n20648_), .A2(new_n20651_), .B(new_n193_), .ZN(new_n20652_));
  NAND3_X1   g20460(.A1(new_n20652_), .A2(new_n20249_), .A3(new_n20647_), .ZN(\asqrt[0] ));
endmodule


