// Benchmark "multiplier" written by ABC on Tue Sep  5 18:12:39 2023

module multiplier ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257_, new_n258_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_,
    new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_,
    new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_,
    new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_,
    new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_,
    new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_,
    new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_,
    new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_,
    new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_,
    new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_,
    new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_,
    new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_,
    new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_,
    new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_,
    new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_,
    new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_,
    new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_,
    new_n3257_, new_n3258_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_,
    new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_,
    new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_,
    new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_,
    new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_,
    new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_,
    new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_,
    new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_,
    new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_,
    new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_,
    new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_,
    new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_,
    new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_,
    new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_,
    new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_,
    new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_,
    new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_,
    new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_,
    new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_,
    new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_,
    new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_,
    new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_,
    new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_,
    new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_,
    new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_,
    new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_,
    new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_,
    new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_,
    new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_,
    new_n4163_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_,
    new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_,
    new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_,
    new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_,
    new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_,
    new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_,
    new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_,
    new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_,
    new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_,
    new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_,
    new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_,
    new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_,
    new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_,
    new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_,
    new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_,
    new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_,
    new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_,
    new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_,
    new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_,
    new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_,
    new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_,
    new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_,
    new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_,
    new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_,
    new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_,
    new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_,
    new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_,
    new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_,
    new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_,
    new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_,
    new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_,
    new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_,
    new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_,
    new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_,
    new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_,
    new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_,
    new_n5189_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5756_,
    new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_,
    new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_,
    new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_,
    new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_,
    new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_,
    new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_,
    new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_,
    new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_,
    new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_,
    new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_,
    new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_,
    new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_,
    new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_,
    new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_,
    new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6229_, new_n6230_, new_n6231_, new_n6232_,
    new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_,
    new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_,
    new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_,
    new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_,
    new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_,
    new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_,
    new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_,
    new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_,
    new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_,
    new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_,
    new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_,
    new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_,
    new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_,
    new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_,
    new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_,
    new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_,
    new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_,
    new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_,
    new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_,
    new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_,
    new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_,
    new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_,
    new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_,
    new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8286_,
    new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_,
    new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_,
    new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_,
    new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_,
    new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_,
    new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_,
    new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_,
    new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_,
    new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_,
    new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_,
    new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_,
    new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_,
    new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_,
    new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_,
    new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_,
    new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_,
    new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_,
    new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_,
    new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_,
    new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8578_, new_n8579_, new_n8580_, new_n8581_,
    new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8954_,
    new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_,
    new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_,
    new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_,
    new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_,
    new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_,
    new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_,
    new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_,
    new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_,
    new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_,
    new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_,
    new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_,
    new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_,
    new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_,
    new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_,
    new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_,
    new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_,
    new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_,
    new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_,
    new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_,
    new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_,
    new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_,
    new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_,
    new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_,
    new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_,
    new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_,
    new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_,
    new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_,
    new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_,
    new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_,
    new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_,
    new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_,
    new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_,
    new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_,
    new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_,
    new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_,
    new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_,
    new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_,
    new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_,
    new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_,
    new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_,
    new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_,
    new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_,
    new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_,
    new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_,
    new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_,
    new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_,
    new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_,
    new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_,
    new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_,
    new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_,
    new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_,
    new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_,
    new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_,
    new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_,
    new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_,
    new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_,
    new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_,
    new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_,
    new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_,
    new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_,
    new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_,
    new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_,
    new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_,
    new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_,
    new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_,
    new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_,
    new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_,
    new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_,
    new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_,
    new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_,
    new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_,
    new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_,
    new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_,
    new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_,
    new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_,
    new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_,
    new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_,
    new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_,
    new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_,
    new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_,
    new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_,
    new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_,
    new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_,
    new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_,
    new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_,
    new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_,
    new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_,
    new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_,
    new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_,
    new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_,
    new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_,
    new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_,
    new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_,
    new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_,
    new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_,
    new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_,
    new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_,
    new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_,
    new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_,
    new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_,
    new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_,
    new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_,
    new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_,
    new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_,
    new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_,
    new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_,
    new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_,
    new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_,
    new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_,
    new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_,
    new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_,
    new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_,
    new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_,
    new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_,
    new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_,
    new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_,
    new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_,
    new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_,
    new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_,
    new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_,
    new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_,
    new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_,
    new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_,
    new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_,
    new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_,
    new_n9989_, new_n9990_, new_n9991_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10397_, new_n10398_, new_n10399_, new_n10400_, new_n10401_,
    new_n10402_, new_n10403_, new_n10404_, new_n10405_, new_n10406_,
    new_n10407_, new_n10408_, new_n10409_, new_n10410_, new_n10411_,
    new_n10412_, new_n10413_, new_n10414_, new_n10415_, new_n10416_,
    new_n10417_, new_n10418_, new_n10419_, new_n10420_, new_n10421_,
    new_n10422_, new_n10423_, new_n10424_, new_n10425_, new_n10426_,
    new_n10427_, new_n10428_, new_n10429_, new_n10430_, new_n10431_,
    new_n10432_, new_n10433_, new_n10434_, new_n10435_, new_n10436_,
    new_n10437_, new_n10438_, new_n10439_, new_n10440_, new_n10441_,
    new_n10442_, new_n10443_, new_n10444_, new_n10445_, new_n10446_,
    new_n10447_, new_n10448_, new_n10449_, new_n10450_, new_n10451_,
    new_n10452_, new_n10453_, new_n10454_, new_n10455_, new_n10456_,
    new_n10457_, new_n10458_, new_n10459_, new_n10460_, new_n10461_,
    new_n10462_, new_n10463_, new_n10464_, new_n10465_, new_n10466_,
    new_n10467_, new_n10468_, new_n10469_, new_n10470_, new_n10471_,
    new_n10472_, new_n10473_, new_n10474_, new_n10475_, new_n10476_,
    new_n10477_, new_n10478_, new_n10479_, new_n10480_, new_n10481_,
    new_n10482_, new_n10483_, new_n10484_, new_n10485_, new_n10486_,
    new_n10487_, new_n10488_, new_n10489_, new_n10490_, new_n10491_,
    new_n10492_, new_n10493_, new_n10494_, new_n10495_, new_n10496_,
    new_n10497_, new_n10498_, new_n10499_, new_n10500_, new_n10501_,
    new_n10502_, new_n10503_, new_n10504_, new_n10505_, new_n10506_,
    new_n10507_, new_n10508_, new_n10509_, new_n10510_, new_n10511_,
    new_n10512_, new_n10513_, new_n10514_, new_n10515_, new_n10516_,
    new_n10517_, new_n10518_, new_n10519_, new_n10520_, new_n10521_,
    new_n10522_, new_n10523_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10530_, new_n10531_,
    new_n10532_, new_n10533_, new_n10534_, new_n10535_, new_n10536_,
    new_n10537_, new_n10538_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10590_, new_n10591_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10615_, new_n10616_,
    new_n10617_, new_n10618_, new_n10619_, new_n10620_, new_n10621_,
    new_n10622_, new_n10623_, new_n10624_, new_n10625_, new_n10626_,
    new_n10627_, new_n10628_, new_n10629_, new_n10630_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10701_,
    new_n10702_, new_n10703_, new_n10704_, new_n10705_, new_n10706_,
    new_n10707_, new_n10708_, new_n10709_, new_n10710_, new_n10711_,
    new_n10712_, new_n10713_, new_n10714_, new_n10715_, new_n10716_,
    new_n10717_, new_n10718_, new_n10719_, new_n10720_, new_n10721_,
    new_n10722_, new_n10723_, new_n10724_, new_n10725_, new_n10726_,
    new_n10727_, new_n10728_, new_n10729_, new_n10730_, new_n10731_,
    new_n10732_, new_n10733_, new_n10734_, new_n10735_, new_n10736_,
    new_n10737_, new_n10738_, new_n10739_, new_n10740_, new_n10741_,
    new_n10742_, new_n10743_, new_n10744_, new_n10745_, new_n10746_,
    new_n10747_, new_n10748_, new_n10749_, new_n10750_, new_n10751_,
    new_n10752_, new_n10753_, new_n10754_, new_n10755_, new_n10756_,
    new_n10757_, new_n10758_, new_n10759_, new_n10760_, new_n10761_,
    new_n10762_, new_n10763_, new_n10764_, new_n10765_, new_n10766_,
    new_n10767_, new_n10768_, new_n10769_, new_n10770_, new_n10771_,
    new_n10772_, new_n10773_, new_n10774_, new_n10775_, new_n10776_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10785_, new_n10786_,
    new_n10787_, new_n10788_, new_n10789_, new_n10790_, new_n10791_,
    new_n10792_, new_n10793_, new_n10794_, new_n10795_, new_n10796_,
    new_n10797_, new_n10798_, new_n10799_, new_n10800_, new_n10801_,
    new_n10802_, new_n10803_, new_n10804_, new_n10805_, new_n10806_,
    new_n10807_, new_n10808_, new_n10809_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10863_, new_n10864_, new_n10865_, new_n10866_, new_n10867_,
    new_n10868_, new_n10869_, new_n10870_, new_n10871_, new_n10872_,
    new_n10873_, new_n10874_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10880_, new_n10881_, new_n10882_,
    new_n10883_, new_n10884_, new_n10885_, new_n10886_, new_n10887_,
    new_n10888_, new_n10889_, new_n10890_, new_n10891_, new_n10892_,
    new_n10893_, new_n10894_, new_n10895_, new_n10896_, new_n10897_,
    new_n10898_, new_n10899_, new_n10900_, new_n10901_, new_n10902_,
    new_n10903_, new_n10904_, new_n10905_, new_n10906_, new_n10907_,
    new_n10908_, new_n10909_, new_n10910_, new_n10911_, new_n10912_,
    new_n10913_, new_n10914_, new_n10915_, new_n10916_, new_n10917_,
    new_n10918_, new_n10919_, new_n10920_, new_n10921_, new_n10922_,
    new_n10923_, new_n10924_, new_n10925_, new_n10926_, new_n10927_,
    new_n10928_, new_n10929_, new_n10930_, new_n10931_, new_n10932_,
    new_n10933_, new_n10934_, new_n10935_, new_n10936_, new_n10937_,
    new_n10938_, new_n10939_, new_n10940_, new_n10941_, new_n10942_,
    new_n10943_, new_n10944_, new_n10945_, new_n10946_, new_n10947_,
    new_n10948_, new_n10949_, new_n10950_, new_n10951_, new_n10952_,
    new_n10953_, new_n10954_, new_n10955_, new_n10956_, new_n10957_,
    new_n10958_, new_n10959_, new_n10960_, new_n10961_, new_n10962_,
    new_n10963_, new_n10964_, new_n10965_, new_n10966_, new_n10967_,
    new_n10968_, new_n10969_, new_n10970_, new_n10971_, new_n10972_,
    new_n10973_, new_n10974_, new_n10975_, new_n10976_, new_n10977_,
    new_n10978_, new_n10979_, new_n10980_, new_n10981_, new_n10982_,
    new_n10983_, new_n10984_, new_n10985_, new_n10986_, new_n10987_,
    new_n10988_, new_n10989_, new_n10990_, new_n10991_, new_n10992_,
    new_n10993_, new_n10994_, new_n10995_, new_n10996_, new_n10997_,
    new_n10998_, new_n10999_, new_n11000_, new_n11001_, new_n11002_,
    new_n11003_, new_n11004_, new_n11005_, new_n11006_, new_n11007_,
    new_n11008_, new_n11009_, new_n11010_, new_n11011_, new_n11012_,
    new_n11013_, new_n11014_, new_n11015_, new_n11016_, new_n11017_,
    new_n11018_, new_n11019_, new_n11020_, new_n11021_, new_n11022_,
    new_n11023_, new_n11024_, new_n11025_, new_n11026_, new_n11027_,
    new_n11028_, new_n11029_, new_n11030_, new_n11031_, new_n11032_,
    new_n11033_, new_n11034_, new_n11035_, new_n11036_, new_n11037_,
    new_n11038_, new_n11039_, new_n11040_, new_n11041_, new_n11042_,
    new_n11043_, new_n11044_, new_n11045_, new_n11046_, new_n11047_,
    new_n11048_, new_n11049_, new_n11050_, new_n11051_, new_n11052_,
    new_n11053_, new_n11054_, new_n11055_, new_n11056_, new_n11057_,
    new_n11058_, new_n11059_, new_n11060_, new_n11061_, new_n11062_,
    new_n11063_, new_n11064_, new_n11065_, new_n11066_, new_n11067_,
    new_n11068_, new_n11069_, new_n11070_, new_n11071_, new_n11072_,
    new_n11073_, new_n11074_, new_n11075_, new_n11076_, new_n11077_,
    new_n11078_, new_n11079_, new_n11080_, new_n11081_, new_n11082_,
    new_n11083_, new_n11084_, new_n11085_, new_n11086_, new_n11087_,
    new_n11088_, new_n11089_, new_n11090_, new_n11091_, new_n11092_,
    new_n11093_, new_n11094_, new_n11095_, new_n11096_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11101_, new_n11102_,
    new_n11103_, new_n11104_, new_n11105_, new_n11106_, new_n11107_,
    new_n11108_, new_n11109_, new_n11110_, new_n11111_, new_n11112_,
    new_n11113_, new_n11114_, new_n11115_, new_n11116_, new_n11117_,
    new_n11118_, new_n11119_, new_n11120_, new_n11121_, new_n11122_,
    new_n11123_, new_n11124_, new_n11125_, new_n11126_, new_n11127_,
    new_n11128_, new_n11129_, new_n11130_, new_n11131_, new_n11132_,
    new_n11133_, new_n11134_, new_n11135_, new_n11136_, new_n11137_,
    new_n11138_, new_n11139_, new_n11140_, new_n11141_, new_n11142_,
    new_n11143_, new_n11144_, new_n11145_, new_n11146_, new_n11147_,
    new_n11148_, new_n11149_, new_n11150_, new_n11151_, new_n11152_,
    new_n11153_, new_n11154_, new_n11155_, new_n11156_, new_n11157_,
    new_n11158_, new_n11159_, new_n11160_, new_n11161_, new_n11162_,
    new_n11163_, new_n11164_, new_n11165_, new_n11166_, new_n11167_,
    new_n11168_, new_n11169_, new_n11170_, new_n11171_, new_n11172_,
    new_n11173_, new_n11174_, new_n11175_, new_n11176_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11206_, new_n11207_, new_n11208_,
    new_n11209_, new_n11210_, new_n11211_, new_n11212_, new_n11213_,
    new_n11214_, new_n11215_, new_n11216_, new_n11217_, new_n11218_,
    new_n11219_, new_n11220_, new_n11221_, new_n11222_, new_n11223_,
    new_n11224_, new_n11225_, new_n11226_, new_n11227_, new_n11228_,
    new_n11229_, new_n11230_, new_n11231_, new_n11232_, new_n11233_,
    new_n11234_, new_n11235_, new_n11236_, new_n11237_, new_n11238_,
    new_n11239_, new_n11240_, new_n11241_, new_n11242_, new_n11243_,
    new_n11244_, new_n11245_, new_n11246_, new_n11247_, new_n11248_,
    new_n11249_, new_n11250_, new_n11251_, new_n11252_, new_n11253_,
    new_n11254_, new_n11255_, new_n11256_, new_n11257_, new_n11258_,
    new_n11259_, new_n11260_, new_n11261_, new_n11262_, new_n11263_,
    new_n11264_, new_n11265_, new_n11266_, new_n11267_, new_n11268_,
    new_n11269_, new_n11270_, new_n11271_, new_n11272_, new_n11273_,
    new_n11274_, new_n11275_, new_n11276_, new_n11277_, new_n11278_,
    new_n11279_, new_n11280_, new_n11281_, new_n11282_, new_n11283_,
    new_n11284_, new_n11285_, new_n11286_, new_n11287_, new_n11288_,
    new_n11289_, new_n11290_, new_n11291_, new_n11292_, new_n11293_,
    new_n11294_, new_n11295_, new_n11296_, new_n11297_, new_n11298_,
    new_n11299_, new_n11300_, new_n11301_, new_n11302_, new_n11303_,
    new_n11304_, new_n11305_, new_n11306_, new_n11307_, new_n11308_,
    new_n11309_, new_n11310_, new_n11311_, new_n11312_, new_n11313_,
    new_n11314_, new_n11315_, new_n11316_, new_n11317_, new_n11318_,
    new_n11319_, new_n11320_, new_n11321_, new_n11322_, new_n11323_,
    new_n11324_, new_n11325_, new_n11326_, new_n11327_, new_n11328_,
    new_n11329_, new_n11330_, new_n11331_, new_n11332_, new_n11333_,
    new_n11334_, new_n11335_, new_n11336_, new_n11337_, new_n11338_,
    new_n11339_, new_n11340_, new_n11341_, new_n11342_, new_n11343_,
    new_n11344_, new_n11345_, new_n11346_, new_n11347_, new_n11348_,
    new_n11349_, new_n11350_, new_n11351_, new_n11352_, new_n11353_,
    new_n11354_, new_n11355_, new_n11356_, new_n11357_, new_n11358_,
    new_n11359_, new_n11360_, new_n11361_, new_n11362_, new_n11363_,
    new_n11364_, new_n11365_, new_n11366_, new_n11367_, new_n11368_,
    new_n11369_, new_n11370_, new_n11371_, new_n11372_, new_n11373_,
    new_n11374_, new_n11375_, new_n11376_, new_n11377_, new_n11378_,
    new_n11379_, new_n11380_, new_n11381_, new_n11382_, new_n11383_,
    new_n11384_, new_n11385_, new_n11386_, new_n11387_, new_n11388_,
    new_n11389_, new_n11390_, new_n11391_, new_n11392_, new_n11393_,
    new_n11394_, new_n11395_, new_n11396_, new_n11397_, new_n11398_,
    new_n11399_, new_n11400_, new_n11401_, new_n11402_, new_n11403_,
    new_n11404_, new_n11405_, new_n11406_, new_n11407_, new_n11408_,
    new_n11409_, new_n11410_, new_n11411_, new_n11412_, new_n11413_,
    new_n11414_, new_n11415_, new_n11416_, new_n11417_, new_n11418_,
    new_n11419_, new_n11420_, new_n11421_, new_n11422_, new_n11423_,
    new_n11424_, new_n11425_, new_n11426_, new_n11427_, new_n11428_,
    new_n11429_, new_n11430_, new_n11431_, new_n11432_, new_n11433_,
    new_n11434_, new_n11435_, new_n11436_, new_n11437_, new_n11438_,
    new_n11439_, new_n11440_, new_n11441_, new_n11442_, new_n11443_,
    new_n11444_, new_n11445_, new_n11446_, new_n11447_, new_n11448_,
    new_n11449_, new_n11450_, new_n11451_, new_n11452_, new_n11453_,
    new_n11454_, new_n11455_, new_n11456_, new_n11457_, new_n11458_,
    new_n11459_, new_n11460_, new_n11461_, new_n11462_, new_n11463_,
    new_n11464_, new_n11465_, new_n11466_, new_n11467_, new_n11468_,
    new_n11469_, new_n11470_, new_n11471_, new_n11472_, new_n11473_,
    new_n11474_, new_n11475_, new_n11476_, new_n11477_, new_n11478_,
    new_n11479_, new_n11480_, new_n11481_, new_n11482_, new_n11483_,
    new_n11484_, new_n11485_, new_n11486_, new_n11487_, new_n11488_,
    new_n11489_, new_n11490_, new_n11491_, new_n11492_, new_n11493_,
    new_n11494_, new_n11495_, new_n11496_, new_n11497_, new_n11498_,
    new_n11499_, new_n11500_, new_n11501_, new_n11502_, new_n11503_,
    new_n11504_, new_n11505_, new_n11506_, new_n11507_, new_n11508_,
    new_n11509_, new_n11510_, new_n11511_, new_n11512_, new_n11513_,
    new_n11514_, new_n11515_, new_n11516_, new_n11517_, new_n11518_,
    new_n11519_, new_n11520_, new_n11521_, new_n11522_, new_n11523_,
    new_n11524_, new_n11525_, new_n11526_, new_n11527_, new_n11528_,
    new_n11529_, new_n11530_, new_n11531_, new_n11532_, new_n11533_,
    new_n11534_, new_n11535_, new_n11536_, new_n11537_, new_n11538_,
    new_n11539_, new_n11540_, new_n11541_, new_n11542_, new_n11543_,
    new_n11544_, new_n11545_, new_n11546_, new_n11547_, new_n11548_,
    new_n11549_, new_n11550_, new_n11551_, new_n11552_, new_n11553_,
    new_n11554_, new_n11555_, new_n11556_, new_n11557_, new_n11558_,
    new_n11559_, new_n11560_, new_n11561_, new_n11562_, new_n11563_,
    new_n11564_, new_n11565_, new_n11566_, new_n11567_, new_n11568_,
    new_n11569_, new_n11570_, new_n11571_, new_n11572_, new_n11573_,
    new_n11574_, new_n11575_, new_n11576_, new_n11577_, new_n11578_,
    new_n11579_, new_n11580_, new_n11581_, new_n11582_, new_n11583_,
    new_n11585_, new_n11586_, new_n11587_, new_n11588_, new_n11589_,
    new_n11590_, new_n11591_, new_n11592_, new_n11593_, new_n11594_,
    new_n11595_, new_n11596_, new_n11597_, new_n11598_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11606_, new_n11607_, new_n11608_, new_n11609_,
    new_n11610_, new_n11611_, new_n11612_, new_n11613_, new_n11614_,
    new_n11615_, new_n11616_, new_n11617_, new_n11618_, new_n11619_,
    new_n11620_, new_n11621_, new_n11622_, new_n11623_, new_n11624_,
    new_n11625_, new_n11626_, new_n11627_, new_n11628_, new_n11629_,
    new_n11630_, new_n11631_, new_n11632_, new_n11633_, new_n11634_,
    new_n11635_, new_n11636_, new_n11637_, new_n11638_, new_n11639_,
    new_n11640_, new_n11641_, new_n11642_, new_n11643_, new_n11644_,
    new_n11645_, new_n11646_, new_n11647_, new_n11648_, new_n11649_,
    new_n11650_, new_n11651_, new_n11652_, new_n11653_, new_n11654_,
    new_n11655_, new_n11656_, new_n11657_, new_n11658_, new_n11659_,
    new_n11660_, new_n11661_, new_n11662_, new_n11663_, new_n11664_,
    new_n11665_, new_n11666_, new_n11667_, new_n11668_, new_n11669_,
    new_n11670_, new_n11671_, new_n11672_, new_n11673_, new_n11674_,
    new_n11675_, new_n11676_, new_n11677_, new_n11678_, new_n11679_,
    new_n11680_, new_n11681_, new_n11682_, new_n11683_, new_n11684_,
    new_n11685_, new_n11686_, new_n11687_, new_n11688_, new_n11689_,
    new_n11690_, new_n11691_, new_n11692_, new_n11693_, new_n11694_,
    new_n11695_, new_n11696_, new_n11697_, new_n11698_, new_n11699_,
    new_n11700_, new_n11701_, new_n11702_, new_n11703_, new_n11704_,
    new_n11705_, new_n11706_, new_n11707_, new_n11708_, new_n11709_,
    new_n11710_, new_n11711_, new_n11712_, new_n11713_, new_n11714_,
    new_n11715_, new_n11716_, new_n11717_, new_n11718_, new_n11719_,
    new_n11720_, new_n11721_, new_n11722_, new_n11723_, new_n11724_,
    new_n11725_, new_n11726_, new_n11727_, new_n11728_, new_n11729_,
    new_n11730_, new_n11731_, new_n11732_, new_n11733_, new_n11734_,
    new_n11735_, new_n11736_, new_n11737_, new_n11738_, new_n11739_,
    new_n11740_, new_n11741_, new_n11742_, new_n11743_, new_n11744_,
    new_n11745_, new_n11746_, new_n11747_, new_n11748_, new_n11749_,
    new_n11750_, new_n11751_, new_n11752_, new_n11753_, new_n11754_,
    new_n11755_, new_n11756_, new_n11757_, new_n11758_, new_n11759_,
    new_n11760_, new_n11761_, new_n11762_, new_n11763_, new_n11764_,
    new_n11765_, new_n11766_, new_n11767_, new_n11768_, new_n11769_,
    new_n11770_, new_n11771_, new_n11772_, new_n11773_, new_n11774_,
    new_n11775_, new_n11776_, new_n11777_, new_n11778_, new_n11779_,
    new_n11780_, new_n11781_, new_n11782_, new_n11783_, new_n11784_,
    new_n11785_, new_n11786_, new_n11787_, new_n11788_, new_n11789_,
    new_n11790_, new_n11791_, new_n11792_, new_n11793_, new_n11794_,
    new_n11795_, new_n11796_, new_n11797_, new_n11798_, new_n11799_,
    new_n11800_, new_n11801_, new_n11802_, new_n11803_, new_n11804_,
    new_n11805_, new_n11806_, new_n11807_, new_n11808_, new_n11809_,
    new_n11810_, new_n11811_, new_n11812_, new_n11813_, new_n11814_,
    new_n11815_, new_n11816_, new_n11817_, new_n11818_, new_n11819_,
    new_n11820_, new_n11821_, new_n11822_, new_n11823_, new_n11824_,
    new_n11825_, new_n11826_, new_n11827_, new_n11828_, new_n11829_,
    new_n11830_, new_n11831_, new_n11832_, new_n11833_, new_n11834_,
    new_n11835_, new_n11836_, new_n11837_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11850_, new_n11851_, new_n11852_, new_n11853_, new_n11854_,
    new_n11855_, new_n11856_, new_n11857_, new_n11858_, new_n11859_,
    new_n11860_, new_n11861_, new_n11862_, new_n11863_, new_n11864_,
    new_n11865_, new_n11866_, new_n11867_, new_n11868_, new_n11869_,
    new_n11870_, new_n11871_, new_n11872_, new_n11873_, new_n11874_,
    new_n11875_, new_n11876_, new_n11877_, new_n11878_, new_n11879_,
    new_n11880_, new_n11881_, new_n11882_, new_n11883_, new_n11884_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11891_, new_n11892_, new_n11893_, new_n11894_,
    new_n11895_, new_n11896_, new_n11897_, new_n11898_, new_n11899_,
    new_n11900_, new_n11901_, new_n11902_, new_n11903_, new_n11904_,
    new_n11905_, new_n11906_, new_n11907_, new_n11908_, new_n11909_,
    new_n11910_, new_n11911_, new_n11912_, new_n11913_, new_n11914_,
    new_n11915_, new_n11916_, new_n11917_, new_n11918_, new_n11919_,
    new_n11920_, new_n11921_, new_n11922_, new_n11923_, new_n11924_,
    new_n11925_, new_n11926_, new_n11927_, new_n11928_, new_n11929_,
    new_n11930_, new_n11931_, new_n11932_, new_n11933_, new_n11934_,
    new_n11935_, new_n11936_, new_n11937_, new_n11938_, new_n11939_,
    new_n11940_, new_n11941_, new_n11942_, new_n11943_, new_n11944_,
    new_n11945_, new_n11946_, new_n11947_, new_n11948_, new_n11949_,
    new_n11950_, new_n11951_, new_n11952_, new_n11953_, new_n11954_,
    new_n11955_, new_n11956_, new_n11957_, new_n11958_, new_n11959_,
    new_n11960_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11965_, new_n11966_, new_n11967_, new_n11968_, new_n11969_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12147_, new_n12148_, new_n12149_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12338_, new_n12339_, new_n12340_, new_n12341_,
    new_n12342_, new_n12343_, new_n12344_, new_n12345_, new_n12346_,
    new_n12347_, new_n12348_, new_n12349_, new_n12350_, new_n12351_,
    new_n12352_, new_n12353_, new_n12354_, new_n12355_, new_n12356_,
    new_n12357_, new_n12358_, new_n12359_, new_n12360_, new_n12361_,
    new_n12362_, new_n12363_, new_n12364_, new_n12365_, new_n12366_,
    new_n12367_, new_n12368_, new_n12369_, new_n12370_, new_n12371_,
    new_n12372_, new_n12373_, new_n12374_, new_n12375_, new_n12376_,
    new_n12377_, new_n12378_, new_n12379_, new_n12380_, new_n12381_,
    new_n12382_, new_n12383_, new_n12384_, new_n12385_, new_n12386_,
    new_n12387_, new_n12388_, new_n12389_, new_n12390_, new_n12391_,
    new_n12392_, new_n12393_, new_n12394_, new_n12395_, new_n12396_,
    new_n12397_, new_n12398_, new_n12399_, new_n12400_, new_n12401_,
    new_n12402_, new_n12403_, new_n12404_, new_n12405_, new_n12406_,
    new_n12407_, new_n12408_, new_n12409_, new_n12410_, new_n12411_,
    new_n12412_, new_n12413_, new_n12414_, new_n12415_, new_n12416_,
    new_n12417_, new_n12418_, new_n12419_, new_n12420_, new_n12421_,
    new_n12422_, new_n12423_, new_n12424_, new_n12425_, new_n12426_,
    new_n12427_, new_n12428_, new_n12429_, new_n12430_, new_n12431_,
    new_n12432_, new_n12433_, new_n12434_, new_n12435_, new_n12436_,
    new_n12437_, new_n12438_, new_n12439_, new_n12440_, new_n12441_,
    new_n12442_, new_n12443_, new_n12444_, new_n12445_, new_n12446_,
    new_n12447_, new_n12448_, new_n12449_, new_n12450_, new_n12451_,
    new_n12452_, new_n12453_, new_n12454_, new_n12455_, new_n12456_,
    new_n12457_, new_n12458_, new_n12459_, new_n12460_, new_n12461_,
    new_n12462_, new_n12463_, new_n12464_, new_n12465_, new_n12466_,
    new_n12467_, new_n12468_, new_n12469_, new_n12470_, new_n12471_,
    new_n12472_, new_n12473_, new_n12474_, new_n12475_, new_n12476_,
    new_n12477_, new_n12478_, new_n12479_, new_n12480_, new_n12481_,
    new_n12482_, new_n12483_, new_n12484_, new_n12485_, new_n12486_,
    new_n12487_, new_n12488_, new_n12489_, new_n12490_, new_n12491_,
    new_n12492_, new_n12493_, new_n12494_, new_n12495_, new_n12496_,
    new_n12497_, new_n12498_, new_n12499_, new_n12500_, new_n12501_,
    new_n12502_, new_n12503_, new_n12504_, new_n12505_, new_n12506_,
    new_n12507_, new_n12508_, new_n12509_, new_n12510_, new_n12511_,
    new_n12512_, new_n12513_, new_n12514_, new_n12515_, new_n12516_,
    new_n12517_, new_n12518_, new_n12519_, new_n12520_, new_n12521_,
    new_n12522_, new_n12523_, new_n12524_, new_n12525_, new_n12526_,
    new_n12527_, new_n12528_, new_n12529_, new_n12530_, new_n12531_,
    new_n12532_, new_n12533_, new_n12534_, new_n12535_, new_n12536_,
    new_n12537_, new_n12538_, new_n12539_, new_n12540_, new_n12541_,
    new_n12542_, new_n12543_, new_n12544_, new_n12545_, new_n12546_,
    new_n12547_, new_n12548_, new_n12549_, new_n12550_, new_n12551_,
    new_n12552_, new_n12553_, new_n12554_, new_n12555_, new_n12556_,
    new_n12557_, new_n12558_, new_n12559_, new_n12560_, new_n12561_,
    new_n12562_, new_n12563_, new_n12564_, new_n12565_, new_n12566_,
    new_n12567_, new_n12568_, new_n12569_, new_n12570_, new_n12571_,
    new_n12572_, new_n12573_, new_n12574_, new_n12575_, new_n12576_,
    new_n12577_, new_n12578_, new_n12579_, new_n12580_, new_n12581_,
    new_n12582_, new_n12583_, new_n12584_, new_n12585_, new_n12586_,
    new_n12587_, new_n12588_, new_n12589_, new_n12590_, new_n12591_,
    new_n12592_, new_n12593_, new_n12594_, new_n12595_, new_n12596_,
    new_n12597_, new_n12598_, new_n12599_, new_n12600_, new_n12601_,
    new_n12602_, new_n12603_, new_n12604_, new_n12605_, new_n12606_,
    new_n12607_, new_n12608_, new_n12609_, new_n12610_, new_n12611_,
    new_n12612_, new_n12613_, new_n12614_, new_n12615_, new_n12616_,
    new_n12617_, new_n12618_, new_n12619_, new_n12620_, new_n12621_,
    new_n12622_, new_n12623_, new_n12624_, new_n12625_, new_n12626_,
    new_n12627_, new_n12628_, new_n12629_, new_n12630_, new_n12631_,
    new_n12632_, new_n12633_, new_n12634_, new_n12635_, new_n12636_,
    new_n12637_, new_n12638_, new_n12639_, new_n12640_, new_n12641_,
    new_n12642_, new_n12643_, new_n12644_, new_n12645_, new_n12646_,
    new_n12647_, new_n12648_, new_n12649_, new_n12650_, new_n12651_,
    new_n12652_, new_n12653_, new_n12654_, new_n12655_, new_n12656_,
    new_n12657_, new_n12658_, new_n12659_, new_n12660_, new_n12661_,
    new_n12662_, new_n12663_, new_n12664_, new_n12665_, new_n12666_,
    new_n12667_, new_n12668_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12766_, new_n12767_,
    new_n12768_, new_n12769_, new_n12770_, new_n12771_, new_n12772_,
    new_n12773_, new_n12774_, new_n12775_, new_n12776_, new_n12777_,
    new_n12778_, new_n12779_, new_n12780_, new_n12781_, new_n12782_,
    new_n12783_, new_n12784_, new_n12785_, new_n12786_, new_n12787_,
    new_n12788_, new_n12789_, new_n12790_, new_n12791_, new_n12792_,
    new_n12793_, new_n12794_, new_n12795_, new_n12796_, new_n12797_,
    new_n12798_, new_n12799_, new_n12800_, new_n12801_, new_n12802_,
    new_n12803_, new_n12804_, new_n12805_, new_n12806_, new_n12807_,
    new_n12808_, new_n12809_, new_n12810_, new_n12811_, new_n12812_,
    new_n12813_, new_n12814_, new_n12815_, new_n12816_, new_n12817_,
    new_n12818_, new_n12819_, new_n12820_, new_n12821_, new_n12822_,
    new_n12823_, new_n12824_, new_n12825_, new_n12826_, new_n12827_,
    new_n12828_, new_n12829_, new_n12830_, new_n12831_, new_n12832_,
    new_n12833_, new_n12834_, new_n12835_, new_n12836_, new_n12837_,
    new_n12838_, new_n12839_, new_n12840_, new_n12841_, new_n12842_,
    new_n12843_, new_n12844_, new_n12845_, new_n12846_, new_n12847_,
    new_n12848_, new_n12849_, new_n12850_, new_n12851_, new_n12852_,
    new_n12853_, new_n12854_, new_n12855_, new_n12856_, new_n12857_,
    new_n12858_, new_n12859_, new_n12860_, new_n12861_, new_n12862_,
    new_n12863_, new_n12864_, new_n12865_, new_n12866_, new_n12867_,
    new_n12868_, new_n12869_, new_n12870_, new_n12871_, new_n12872_,
    new_n12873_, new_n12874_, new_n12875_, new_n12876_, new_n12877_,
    new_n12878_, new_n12879_, new_n12880_, new_n12881_, new_n12882_,
    new_n12883_, new_n12884_, new_n12885_, new_n12886_, new_n12887_,
    new_n12888_, new_n12889_, new_n12890_, new_n12891_, new_n12892_,
    new_n12893_, new_n12894_, new_n12895_, new_n12896_, new_n12897_,
    new_n12898_, new_n12899_, new_n12900_, new_n12901_, new_n12902_,
    new_n12903_, new_n12904_, new_n12905_, new_n12906_, new_n12907_,
    new_n12908_, new_n12909_, new_n12910_, new_n12911_, new_n12912_,
    new_n12913_, new_n12914_, new_n12915_, new_n12916_, new_n12917_,
    new_n12918_, new_n12919_, new_n12920_, new_n12921_, new_n12922_,
    new_n12923_, new_n12924_, new_n12925_, new_n12926_, new_n12927_,
    new_n12928_, new_n12929_, new_n12930_, new_n12931_, new_n12932_,
    new_n12933_, new_n12934_, new_n12935_, new_n12936_, new_n12937_,
    new_n12938_, new_n12939_, new_n12940_, new_n12941_, new_n12942_,
    new_n12943_, new_n12944_, new_n12945_, new_n12946_, new_n12947_,
    new_n12948_, new_n12949_, new_n12950_, new_n12951_, new_n12952_,
    new_n12953_, new_n12954_, new_n12955_, new_n12956_, new_n12957_,
    new_n12958_, new_n12959_, new_n12960_, new_n12961_, new_n12962_,
    new_n12963_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12993_, new_n12994_, new_n12995_, new_n12996_, new_n12997_,
    new_n12998_, new_n12999_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13006_, new_n13007_, new_n13008_,
    new_n13009_, new_n13010_, new_n13011_, new_n13012_, new_n13013_,
    new_n13014_, new_n13015_, new_n13016_, new_n13017_, new_n13018_,
    new_n13019_, new_n13020_, new_n13021_, new_n13022_, new_n13023_,
    new_n13024_, new_n13025_, new_n13026_, new_n13027_, new_n13028_,
    new_n13029_, new_n13030_, new_n13031_, new_n13032_, new_n13033_,
    new_n13034_, new_n13035_, new_n13036_, new_n13037_, new_n13038_,
    new_n13039_, new_n13040_, new_n13041_, new_n13042_, new_n13043_,
    new_n13044_, new_n13045_, new_n13046_, new_n13047_, new_n13048_,
    new_n13049_, new_n13050_, new_n13051_, new_n13052_, new_n13053_,
    new_n13054_, new_n13055_, new_n13056_, new_n13057_, new_n13058_,
    new_n13059_, new_n13060_, new_n13061_, new_n13062_, new_n13063_,
    new_n13064_, new_n13065_, new_n13066_, new_n13067_, new_n13068_,
    new_n13069_, new_n13070_, new_n13071_, new_n13072_, new_n13073_,
    new_n13074_, new_n13075_, new_n13076_, new_n13077_, new_n13078_,
    new_n13079_, new_n13080_, new_n13081_, new_n13082_, new_n13083_,
    new_n13084_, new_n13085_, new_n13086_, new_n13087_, new_n13088_,
    new_n13089_, new_n13090_, new_n13091_, new_n13092_, new_n13093_,
    new_n13094_, new_n13095_, new_n13096_, new_n13097_, new_n13098_,
    new_n13099_, new_n13100_, new_n13101_, new_n13102_, new_n13103_,
    new_n13104_, new_n13105_, new_n13106_, new_n13107_, new_n13108_,
    new_n13109_, new_n13110_, new_n13111_, new_n13112_, new_n13113_,
    new_n13114_, new_n13115_, new_n13116_, new_n13117_, new_n13118_,
    new_n13119_, new_n13120_, new_n13121_, new_n13122_, new_n13123_,
    new_n13124_, new_n13125_, new_n13126_, new_n13127_, new_n13128_,
    new_n13129_, new_n13130_, new_n13131_, new_n13132_, new_n13133_,
    new_n13134_, new_n13135_, new_n13136_, new_n13137_, new_n13138_,
    new_n13139_, new_n13140_, new_n13141_, new_n13142_, new_n13143_,
    new_n13144_, new_n13145_, new_n13146_, new_n13147_, new_n13148_,
    new_n13149_, new_n13150_, new_n13151_, new_n13152_, new_n13153_,
    new_n13154_, new_n13155_, new_n13156_, new_n13157_, new_n13158_,
    new_n13159_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13165_, new_n13166_, new_n13167_, new_n13168_,
    new_n13169_, new_n13170_, new_n13171_, new_n13172_, new_n13173_,
    new_n13174_, new_n13175_, new_n13176_, new_n13177_, new_n13178_,
    new_n13179_, new_n13180_, new_n13181_, new_n13182_, new_n13183_,
    new_n13184_, new_n13185_, new_n13186_, new_n13187_, new_n13188_,
    new_n13189_, new_n13190_, new_n13191_, new_n13192_, new_n13193_,
    new_n13194_, new_n13195_, new_n13196_, new_n13197_, new_n13198_,
    new_n13199_, new_n13200_, new_n13201_, new_n13202_, new_n13203_,
    new_n13204_, new_n13205_, new_n13206_, new_n13207_, new_n13208_,
    new_n13209_, new_n13210_, new_n13211_, new_n13212_, new_n13213_,
    new_n13214_, new_n13215_, new_n13216_, new_n13217_, new_n13218_,
    new_n13219_, new_n13220_, new_n13221_, new_n13222_, new_n13223_,
    new_n13224_, new_n13225_, new_n13226_, new_n13227_, new_n13228_,
    new_n13229_, new_n13230_, new_n13231_, new_n13232_, new_n13233_,
    new_n13234_, new_n13235_, new_n13236_, new_n13237_, new_n13238_,
    new_n13239_, new_n13240_, new_n13241_, new_n13242_, new_n13243_,
    new_n13244_, new_n13245_, new_n13246_, new_n13247_, new_n13248_,
    new_n13249_, new_n13250_, new_n13251_, new_n13252_, new_n13253_,
    new_n13254_, new_n13255_, new_n13256_, new_n13257_, new_n13258_,
    new_n13259_, new_n13260_, new_n13261_, new_n13262_, new_n13263_,
    new_n13264_, new_n13265_, new_n13266_, new_n13267_, new_n13268_,
    new_n13269_, new_n13270_, new_n13271_, new_n13272_, new_n13273_,
    new_n13274_, new_n13275_, new_n13276_, new_n13277_, new_n13278_,
    new_n13279_, new_n13280_, new_n13281_, new_n13282_, new_n13283_,
    new_n13284_, new_n13285_, new_n13286_, new_n13287_, new_n13288_,
    new_n13289_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13334_,
    new_n13335_, new_n13336_, new_n13337_, new_n13338_, new_n13339_,
    new_n13340_, new_n13341_, new_n13342_, new_n13343_, new_n13344_,
    new_n13345_, new_n13346_, new_n13347_, new_n13348_, new_n13349_,
    new_n13350_, new_n13351_, new_n13352_, new_n13353_, new_n13354_,
    new_n13355_, new_n13356_, new_n13357_, new_n13358_, new_n13359_,
    new_n13360_, new_n13361_, new_n13362_, new_n13363_, new_n13364_,
    new_n13365_, new_n13366_, new_n13367_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13375_, new_n13376_, new_n13377_, new_n13378_, new_n13379_,
    new_n13380_, new_n13381_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13407_, new_n13408_, new_n13409_,
    new_n13410_, new_n13411_, new_n13412_, new_n13413_, new_n13414_,
    new_n13415_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13438_, new_n13439_,
    new_n13440_, new_n13441_, new_n13442_, new_n13443_, new_n13444_,
    new_n13445_, new_n13446_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13452_, new_n13453_, new_n13454_,
    new_n13455_, new_n13456_, new_n13457_, new_n13458_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13464_,
    new_n13465_, new_n13466_, new_n13467_, new_n13468_, new_n13469_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13511_, new_n13512_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13539_,
    new_n13540_, new_n13541_, new_n13542_, new_n13543_, new_n13544_,
    new_n13545_, new_n13546_, new_n13547_, new_n13548_, new_n13549_,
    new_n13550_, new_n13551_, new_n13552_, new_n13553_, new_n13554_,
    new_n13555_, new_n13556_, new_n13557_, new_n13558_, new_n13559_,
    new_n13560_, new_n13561_, new_n13562_, new_n13563_, new_n13564_,
    new_n13565_, new_n13566_, new_n13567_, new_n13568_, new_n13569_,
    new_n13570_, new_n13571_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13591_, new_n13592_, new_n13593_, new_n13594_,
    new_n13595_, new_n13596_, new_n13597_, new_n13598_, new_n13599_,
    new_n13600_, new_n13601_, new_n13602_, new_n13603_, new_n13604_,
    new_n13605_, new_n13606_, new_n13607_, new_n13608_, new_n13609_,
    new_n13610_, new_n13611_, new_n13612_, new_n13613_, new_n13614_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13660_, new_n13661_, new_n13662_, new_n13663_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14536_, new_n14537_, new_n14538_,
    new_n14539_, new_n14540_, new_n14541_, new_n14542_, new_n14543_,
    new_n14544_, new_n14545_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14606_, new_n14607_, new_n14608_,
    new_n14609_, new_n14610_, new_n14611_, new_n14612_, new_n14613_,
    new_n14614_, new_n14615_, new_n14616_, new_n14617_, new_n14618_,
    new_n14619_, new_n14620_, new_n14621_, new_n14622_, new_n14623_,
    new_n14624_, new_n14625_, new_n14626_, new_n14627_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14633_,
    new_n14634_, new_n14635_, new_n14636_, new_n14637_, new_n14638_,
    new_n14639_, new_n14640_, new_n14641_, new_n14642_, new_n14643_,
    new_n14644_, new_n14645_, new_n14646_, new_n14647_, new_n14648_,
    new_n14649_, new_n14650_, new_n14651_, new_n14652_, new_n14653_,
    new_n14654_, new_n14655_, new_n14656_, new_n14657_, new_n14658_,
    new_n14659_, new_n14660_, new_n14661_, new_n14662_, new_n14663_,
    new_n14664_, new_n14665_, new_n14666_, new_n14667_, new_n14668_,
    new_n14669_, new_n14670_, new_n14671_, new_n14672_, new_n14673_,
    new_n14674_, new_n14675_, new_n14676_, new_n14677_, new_n14678_,
    new_n14679_, new_n14680_, new_n14681_, new_n14682_, new_n14683_,
    new_n14684_, new_n14685_, new_n14686_, new_n14687_, new_n14688_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14693_,
    new_n14694_, new_n14695_, new_n14696_, new_n14697_, new_n14698_,
    new_n14699_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14705_, new_n14706_, new_n14707_, new_n14708_,
    new_n14709_, new_n14710_, new_n14711_, new_n14712_, new_n14713_,
    new_n14714_, new_n14715_, new_n14716_, new_n14717_, new_n14718_,
    new_n14719_, new_n14720_, new_n14721_, new_n14722_, new_n14723_,
    new_n14724_, new_n14725_, new_n14726_, new_n14727_, new_n14728_,
    new_n14729_, new_n14730_, new_n14731_, new_n14732_, new_n14733_,
    new_n14734_, new_n14735_, new_n14736_, new_n14737_, new_n14738_,
    new_n14739_, new_n14740_, new_n14741_, new_n14742_, new_n14743_,
    new_n14744_, new_n14745_, new_n14746_, new_n14747_, new_n14748_,
    new_n14749_, new_n14750_, new_n14751_, new_n14752_, new_n14753_,
    new_n14754_, new_n14755_, new_n14756_, new_n14757_, new_n14758_,
    new_n14759_, new_n14760_, new_n14761_, new_n14762_, new_n14763_,
    new_n14764_, new_n14765_, new_n14766_, new_n14767_, new_n14768_,
    new_n14769_, new_n14770_, new_n14771_, new_n14772_, new_n14773_,
    new_n14774_, new_n14775_, new_n14776_, new_n14777_, new_n14778_,
    new_n14779_, new_n14780_, new_n14781_, new_n14782_, new_n14783_,
    new_n14785_, new_n14786_, new_n14787_, new_n14788_, new_n14789_,
    new_n14790_, new_n14791_, new_n14792_, new_n14793_, new_n14794_,
    new_n14795_, new_n14796_, new_n14797_, new_n14798_, new_n14799_,
    new_n14800_, new_n14801_, new_n14802_, new_n14803_, new_n14804_,
    new_n14805_, new_n14806_, new_n14807_, new_n14808_, new_n14809_,
    new_n14810_, new_n14811_, new_n14812_, new_n14813_, new_n14814_,
    new_n14815_, new_n14816_, new_n14817_, new_n14818_, new_n14819_,
    new_n14820_, new_n14821_, new_n14822_, new_n14823_, new_n14824_,
    new_n14825_, new_n14826_, new_n14827_, new_n14828_, new_n14829_,
    new_n14830_, new_n14831_, new_n14832_, new_n14833_, new_n14834_,
    new_n14835_, new_n14836_, new_n14837_, new_n14838_, new_n14839_,
    new_n14840_, new_n14841_, new_n14842_, new_n14843_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14908_, new_n14909_,
    new_n14910_, new_n14911_, new_n14912_, new_n14913_, new_n14914_,
    new_n14915_, new_n14916_, new_n14917_, new_n14918_, new_n14919_,
    new_n14920_, new_n14921_, new_n14922_, new_n14923_, new_n14924_,
    new_n14925_, new_n14926_, new_n14927_, new_n14928_, new_n14929_,
    new_n14930_, new_n14931_, new_n14932_, new_n14933_, new_n14934_,
    new_n14935_, new_n14936_, new_n14937_, new_n14938_, new_n14939_,
    new_n14940_, new_n14941_, new_n14942_, new_n14943_, new_n14944_,
    new_n14945_, new_n14946_, new_n14947_, new_n14948_, new_n14949_,
    new_n14950_, new_n14951_, new_n14952_, new_n14953_, new_n14954_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14963_, new_n14964_,
    new_n14965_, new_n14966_, new_n14967_, new_n14968_, new_n14969_,
    new_n14970_, new_n14971_, new_n14972_, new_n14973_, new_n14974_,
    new_n14975_, new_n14976_, new_n14977_, new_n14978_, new_n14979_,
    new_n14980_, new_n14981_, new_n14982_, new_n14983_, new_n14984_,
    new_n14985_, new_n14986_, new_n14987_, new_n14988_, new_n14989_,
    new_n14990_, new_n14991_, new_n14992_, new_n14993_, new_n14994_,
    new_n14995_, new_n14996_, new_n14997_, new_n14998_, new_n14999_,
    new_n15000_, new_n15001_, new_n15002_, new_n15003_, new_n15004_,
    new_n15005_, new_n15006_, new_n15007_, new_n15008_, new_n15009_,
    new_n15010_, new_n15011_, new_n15012_, new_n15013_, new_n15014_,
    new_n15015_, new_n15016_, new_n15017_, new_n15018_, new_n15019_,
    new_n15020_, new_n15021_, new_n15022_, new_n15023_, new_n15024_,
    new_n15025_, new_n15026_, new_n15027_, new_n15028_, new_n15029_,
    new_n15030_, new_n15031_, new_n15032_, new_n15033_, new_n15034_,
    new_n15035_, new_n15036_, new_n15037_, new_n15038_, new_n15039_,
    new_n15040_, new_n15041_, new_n15042_, new_n15043_, new_n15044_,
    new_n15045_, new_n15046_, new_n15047_, new_n15048_, new_n15049_,
    new_n15050_, new_n15051_, new_n15052_, new_n15053_, new_n15054_,
    new_n15055_, new_n15056_, new_n15057_, new_n15058_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15328_, new_n15329_, new_n15330_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15366_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15374_, new_n15375_, new_n15376_,
    new_n15377_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15422_, new_n15423_, new_n15424_, new_n15425_, new_n15426_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15433_, new_n15434_, new_n15435_, new_n15436_,
    new_n15437_, new_n15438_, new_n15439_, new_n15440_, new_n15441_,
    new_n15442_, new_n15443_, new_n15444_, new_n15445_, new_n15446_,
    new_n15447_, new_n15448_, new_n15449_, new_n15450_, new_n15451_,
    new_n15452_, new_n15453_, new_n15454_, new_n15455_, new_n15456_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15464_, new_n15465_, new_n15466_,
    new_n15467_, new_n15468_, new_n15469_, new_n15470_, new_n15471_,
    new_n15472_, new_n15473_, new_n15474_, new_n15475_, new_n15476_,
    new_n15477_, new_n15478_, new_n15479_, new_n15480_, new_n15481_,
    new_n15482_, new_n15483_, new_n15484_, new_n15485_, new_n15486_,
    new_n15487_, new_n15488_, new_n15489_, new_n15490_, new_n15491_,
    new_n15492_, new_n15493_, new_n15494_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15542_, new_n15543_, new_n15544_, new_n15545_, new_n15546_,
    new_n15547_, new_n15548_, new_n15549_, new_n15550_, new_n15551_,
    new_n15552_, new_n15553_, new_n15554_, new_n15555_, new_n15556_,
    new_n15557_, new_n15558_, new_n15559_, new_n15560_, new_n15561_,
    new_n15562_, new_n15563_, new_n15564_, new_n15565_, new_n15566_,
    new_n15567_, new_n15568_, new_n15569_, new_n15571_, new_n15572_,
    new_n15573_, new_n15574_, new_n15575_, new_n15576_, new_n15577_,
    new_n15578_, new_n15579_, new_n15580_, new_n15581_, new_n15582_,
    new_n15583_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15590_, new_n15591_, new_n15592_,
    new_n15593_, new_n15594_, new_n15595_, new_n15596_, new_n15597_,
    new_n15598_, new_n15599_, new_n15600_, new_n15601_, new_n15602_,
    new_n15603_, new_n15604_, new_n15605_, new_n15606_, new_n15607_,
    new_n15608_, new_n15609_, new_n15610_, new_n15611_, new_n15612_,
    new_n15613_, new_n15614_, new_n15615_, new_n15616_, new_n15617_,
    new_n15618_, new_n15619_, new_n15620_, new_n15621_, new_n15622_,
    new_n15623_, new_n15624_, new_n15625_, new_n15626_, new_n15627_,
    new_n15628_, new_n15629_, new_n15630_, new_n15631_, new_n15632_,
    new_n15633_, new_n15634_, new_n15635_, new_n15636_, new_n15637_,
    new_n15638_, new_n15639_, new_n15640_, new_n15641_, new_n15642_,
    new_n15643_, new_n15644_, new_n15645_, new_n15646_, new_n15647_,
    new_n15648_, new_n15649_, new_n15650_, new_n15651_, new_n15652_,
    new_n15653_, new_n15654_, new_n15655_, new_n15656_, new_n15657_,
    new_n15658_, new_n15659_, new_n15660_, new_n15661_, new_n15662_,
    new_n15663_, new_n15664_, new_n15665_, new_n15666_, new_n15667_,
    new_n15668_, new_n15669_, new_n15670_, new_n15671_, new_n15672_,
    new_n15673_, new_n15674_, new_n15675_, new_n15676_, new_n15677_,
    new_n15678_, new_n15679_, new_n15680_, new_n15681_, new_n15682_,
    new_n15683_, new_n15684_, new_n15685_, new_n15686_, new_n15687_,
    new_n15688_, new_n15689_, new_n15690_, new_n15691_, new_n15692_,
    new_n15693_, new_n15694_, new_n15695_, new_n15696_, new_n15697_,
    new_n15698_, new_n15699_, new_n15700_, new_n15701_, new_n15702_,
    new_n15703_, new_n15704_, new_n15705_, new_n15706_, new_n15707_,
    new_n15708_, new_n15709_, new_n15710_, new_n15711_, new_n15712_,
    new_n15713_, new_n15714_, new_n15715_, new_n15716_, new_n15717_,
    new_n15718_, new_n15719_, new_n15720_, new_n15721_, new_n15722_,
    new_n15723_, new_n15724_, new_n15725_, new_n15726_, new_n15727_,
    new_n15728_, new_n15729_, new_n15730_, new_n15731_, new_n15732_,
    new_n15733_, new_n15734_, new_n15735_, new_n15736_, new_n15737_,
    new_n15738_, new_n15739_, new_n15740_, new_n15741_, new_n15742_,
    new_n15743_, new_n15744_, new_n15745_, new_n15746_, new_n15747_,
    new_n15748_, new_n15749_, new_n15750_, new_n15751_, new_n15752_,
    new_n15753_, new_n15754_, new_n15755_, new_n15756_, new_n15757_,
    new_n15758_, new_n15759_, new_n15760_, new_n15761_, new_n15762_,
    new_n15763_, new_n15764_, new_n15765_, new_n15766_, new_n15767_,
    new_n15768_, new_n15769_, new_n15770_, new_n15771_, new_n15772_,
    new_n15773_, new_n15774_, new_n15775_, new_n15776_, new_n15777_,
    new_n15778_, new_n15779_, new_n15780_, new_n15781_, new_n15782_,
    new_n15784_, new_n15785_, new_n15786_, new_n15787_, new_n15788_,
    new_n15789_, new_n15790_, new_n15791_, new_n15792_, new_n15793_,
    new_n15794_, new_n15795_, new_n15796_, new_n15797_, new_n15798_,
    new_n15799_, new_n15800_, new_n15801_, new_n15802_, new_n15803_,
    new_n15804_, new_n15805_, new_n15806_, new_n15807_, new_n15808_,
    new_n15809_, new_n15810_, new_n15811_, new_n15812_, new_n15813_,
    new_n15814_, new_n15815_, new_n15816_, new_n15817_, new_n15818_,
    new_n15819_, new_n15820_, new_n15821_, new_n15822_, new_n15823_,
    new_n15824_, new_n15825_, new_n15826_, new_n15827_, new_n15828_,
    new_n15829_, new_n15830_, new_n15831_, new_n15832_, new_n15833_,
    new_n15834_, new_n15835_, new_n15836_, new_n15837_, new_n15838_,
    new_n15839_, new_n15840_, new_n15841_, new_n15842_, new_n15843_,
    new_n15844_, new_n15845_, new_n15846_, new_n15847_, new_n15848_,
    new_n15849_, new_n15850_, new_n15851_, new_n15852_, new_n15853_,
    new_n15854_, new_n15855_, new_n15856_, new_n15857_, new_n15858_,
    new_n15859_, new_n15860_, new_n15861_, new_n15862_, new_n15863_,
    new_n15864_, new_n15865_, new_n15866_, new_n15867_, new_n15868_,
    new_n15869_, new_n15870_, new_n15871_, new_n15872_, new_n15873_,
    new_n15874_, new_n15875_, new_n15876_, new_n15877_, new_n15878_,
    new_n15879_, new_n15880_, new_n15881_, new_n15882_, new_n15883_,
    new_n15884_, new_n15885_, new_n15886_, new_n15887_, new_n15888_,
    new_n15889_, new_n15890_, new_n15891_, new_n15892_, new_n15893_,
    new_n15894_, new_n15895_, new_n15896_, new_n15897_, new_n15898_,
    new_n15899_, new_n15900_, new_n15901_, new_n15902_, new_n15903_,
    new_n15904_, new_n15905_, new_n15906_, new_n15907_, new_n15908_,
    new_n15909_, new_n15910_, new_n15911_, new_n15912_, new_n15913_,
    new_n15914_, new_n15915_, new_n15916_, new_n15917_, new_n15918_,
    new_n15919_, new_n15920_, new_n15921_, new_n15922_, new_n15923_,
    new_n15924_, new_n15925_, new_n15926_, new_n15927_, new_n15928_,
    new_n15929_, new_n15930_, new_n15931_, new_n15932_, new_n15933_,
    new_n15934_, new_n15935_, new_n15936_, new_n15937_, new_n15938_,
    new_n15939_, new_n15940_, new_n15941_, new_n15942_, new_n15943_,
    new_n15944_, new_n15945_, new_n15946_, new_n15947_, new_n15948_,
    new_n15949_, new_n15950_, new_n15951_, new_n15952_, new_n15953_,
    new_n15954_, new_n15955_, new_n15956_, new_n15957_, new_n15958_,
    new_n15959_, new_n15960_, new_n15961_, new_n15962_, new_n15963_,
    new_n15964_, new_n15965_, new_n15966_, new_n15967_, new_n15968_,
    new_n15969_, new_n15970_, new_n15971_, new_n15972_, new_n15973_,
    new_n15974_, new_n15975_, new_n15976_, new_n15977_, new_n15978_,
    new_n15979_, new_n15980_, new_n15981_, new_n15982_, new_n15983_,
    new_n15984_, new_n15985_, new_n15986_, new_n15987_, new_n15988_,
    new_n15989_, new_n15990_, new_n15991_, new_n15992_, new_n15993_,
    new_n15994_, new_n15995_, new_n15996_, new_n15997_, new_n15998_,
    new_n15999_, new_n16000_, new_n16001_, new_n16002_, new_n16003_,
    new_n16004_, new_n16005_, new_n16006_, new_n16007_, new_n16008_,
    new_n16009_, new_n16010_, new_n16011_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16067_, new_n16068_, new_n16069_,
    new_n16070_, new_n16071_, new_n16072_, new_n16073_, new_n16074_,
    new_n16075_, new_n16076_, new_n16077_, new_n16078_, new_n16079_,
    new_n16080_, new_n16081_, new_n16082_, new_n16083_, new_n16084_,
    new_n16085_, new_n16086_, new_n16087_, new_n16088_, new_n16089_,
    new_n16090_, new_n16091_, new_n16092_, new_n16093_, new_n16094_,
    new_n16095_, new_n16096_, new_n16097_, new_n16098_, new_n16099_,
    new_n16100_, new_n16101_, new_n16102_, new_n16103_, new_n16104_,
    new_n16105_, new_n16106_, new_n16107_, new_n16108_, new_n16109_,
    new_n16110_, new_n16111_, new_n16112_, new_n16113_, new_n16114_,
    new_n16115_, new_n16116_, new_n16117_, new_n16118_, new_n16119_,
    new_n16120_, new_n16121_, new_n16122_, new_n16123_, new_n16124_,
    new_n16125_, new_n16126_, new_n16127_, new_n16128_, new_n16129_,
    new_n16130_, new_n16131_, new_n16132_, new_n16133_, new_n16134_,
    new_n16135_, new_n16136_, new_n16137_, new_n16138_, new_n16139_,
    new_n16140_, new_n16141_, new_n16142_, new_n16143_, new_n16144_,
    new_n16145_, new_n16146_, new_n16147_, new_n16148_, new_n16149_,
    new_n16150_, new_n16151_, new_n16152_, new_n16153_, new_n16154_,
    new_n16155_, new_n16156_, new_n16157_, new_n16158_, new_n16159_,
    new_n16160_, new_n16161_, new_n16162_, new_n16163_, new_n16164_,
    new_n16165_, new_n16166_, new_n16167_, new_n16168_, new_n16169_,
    new_n16170_, new_n16171_, new_n16172_, new_n16173_, new_n16174_,
    new_n16175_, new_n16176_, new_n16177_, new_n16178_, new_n16179_,
    new_n16180_, new_n16181_, new_n16182_, new_n16183_, new_n16184_,
    new_n16185_, new_n16186_, new_n16187_, new_n16188_, new_n16189_,
    new_n16190_, new_n16191_, new_n16192_, new_n16193_, new_n16194_,
    new_n16195_, new_n16196_, new_n16197_, new_n16198_, new_n16199_,
    new_n16200_, new_n16201_, new_n16202_, new_n16203_, new_n16204_,
    new_n16205_, new_n16206_, new_n16207_, new_n16208_, new_n16209_,
    new_n16210_, new_n16211_, new_n16212_, new_n16213_, new_n16214_,
    new_n16215_, new_n16216_, new_n16217_, new_n16218_, new_n16219_,
    new_n16220_, new_n16221_, new_n16222_, new_n16223_, new_n16224_,
    new_n16225_, new_n16226_, new_n16227_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16349_, new_n16350_,
    new_n16351_, new_n16352_, new_n16353_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16361_, new_n16362_, new_n16363_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16612_, new_n16613_, new_n16614_, new_n16615_, new_n16616_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16634_, new_n16635_, new_n16636_,
    new_n16637_, new_n16638_, new_n16639_, new_n16640_, new_n16641_,
    new_n16642_, new_n16643_, new_n16644_, new_n16645_, new_n16646_,
    new_n16647_, new_n16648_, new_n16649_, new_n16651_, new_n16652_,
    new_n16653_, new_n16654_, new_n16655_, new_n16656_, new_n16657_,
    new_n16658_, new_n16659_, new_n16660_, new_n16661_, new_n16662_,
    new_n16663_, new_n16664_, new_n16665_, new_n16666_, new_n16667_,
    new_n16668_, new_n16669_, new_n16670_, new_n16671_, new_n16672_,
    new_n16673_, new_n16674_, new_n16675_, new_n16676_, new_n16677_,
    new_n16678_, new_n16679_, new_n16680_, new_n16681_, new_n16682_,
    new_n16683_, new_n16684_, new_n16685_, new_n16686_, new_n16687_,
    new_n16688_, new_n16689_, new_n16690_, new_n16691_, new_n16692_,
    new_n16693_, new_n16694_, new_n16695_, new_n16696_, new_n16697_,
    new_n16698_, new_n16699_, new_n16700_, new_n16701_, new_n16702_,
    new_n16703_, new_n16704_, new_n16705_, new_n16706_, new_n16707_,
    new_n16708_, new_n16709_, new_n16710_, new_n16711_, new_n16712_,
    new_n16713_, new_n16714_, new_n16715_, new_n16716_, new_n16717_,
    new_n16718_, new_n16719_, new_n16720_, new_n16721_, new_n16722_,
    new_n16723_, new_n16724_, new_n16725_, new_n16726_, new_n16727_,
    new_n16728_, new_n16729_, new_n16730_, new_n16731_, new_n16732_,
    new_n16733_, new_n16734_, new_n16735_, new_n16736_, new_n16737_,
    new_n16738_, new_n16739_, new_n16740_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16749_, new_n16750_, new_n16751_, new_n16752_,
    new_n16753_, new_n16754_, new_n16755_, new_n16756_, new_n16757_,
    new_n16758_, new_n16759_, new_n16760_, new_n16761_, new_n16762_,
    new_n16763_, new_n16764_, new_n16765_, new_n16766_, new_n16767_,
    new_n16768_, new_n16769_, new_n16770_, new_n16771_, new_n16772_,
    new_n16773_, new_n16774_, new_n16775_, new_n16776_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16781_, new_n16782_,
    new_n16783_, new_n16784_, new_n16785_, new_n16786_, new_n16787_,
    new_n16788_, new_n16789_, new_n16790_, new_n16791_, new_n16792_,
    new_n16793_, new_n16794_, new_n16795_, new_n16796_, new_n16797_,
    new_n16798_, new_n16799_, new_n16800_, new_n16801_, new_n16802_,
    new_n16803_, new_n16804_, new_n16805_, new_n16806_, new_n16807_,
    new_n16808_, new_n16809_, new_n16810_, new_n16811_, new_n16812_,
    new_n16813_, new_n16814_, new_n16815_, new_n16816_, new_n16817_,
    new_n16818_, new_n16819_, new_n16820_, new_n16821_, new_n16822_,
    new_n16823_, new_n16824_, new_n16825_, new_n16826_, new_n16827_,
    new_n16828_, new_n16829_, new_n16830_, new_n16831_, new_n16832_,
    new_n16833_, new_n16834_, new_n16835_, new_n16836_, new_n16837_,
    new_n16838_, new_n16839_, new_n16840_, new_n16841_, new_n16842_,
    new_n16843_, new_n16844_, new_n16845_, new_n16846_, new_n16847_,
    new_n16848_, new_n16849_, new_n16850_, new_n16851_, new_n16852_,
    new_n16853_, new_n16855_, new_n16856_, new_n16857_, new_n16858_,
    new_n16859_, new_n16860_, new_n16861_, new_n16862_, new_n16863_,
    new_n16864_, new_n16865_, new_n16866_, new_n16867_, new_n16868_,
    new_n16869_, new_n16870_, new_n16871_, new_n16872_, new_n16873_,
    new_n16874_, new_n16875_, new_n16876_, new_n16877_, new_n16878_,
    new_n16879_, new_n16880_, new_n16881_, new_n16882_, new_n16883_,
    new_n16884_, new_n16885_, new_n16886_, new_n16887_, new_n16888_,
    new_n16889_, new_n16890_, new_n16891_, new_n16892_, new_n16893_,
    new_n16894_, new_n16895_, new_n16896_, new_n16897_, new_n16898_,
    new_n16899_, new_n16900_, new_n16901_, new_n16902_, new_n16903_,
    new_n16904_, new_n16905_, new_n16906_, new_n16907_, new_n16908_,
    new_n16909_, new_n16910_, new_n16911_, new_n16912_, new_n16913_,
    new_n16914_, new_n16915_, new_n16916_, new_n16917_, new_n16918_,
    new_n16919_, new_n16920_, new_n16921_, new_n16922_, new_n16923_,
    new_n16924_, new_n16925_, new_n16926_, new_n16927_, new_n16928_,
    new_n16929_, new_n16930_, new_n16931_, new_n16932_, new_n16933_,
    new_n16934_, new_n16935_, new_n16936_, new_n16937_, new_n16938_,
    new_n16939_, new_n16940_, new_n16941_, new_n16942_, new_n16943_,
    new_n16944_, new_n16945_, new_n16946_, new_n16947_, new_n16948_,
    new_n16949_, new_n16950_, new_n16951_, new_n16952_, new_n16953_,
    new_n16954_, new_n16955_, new_n16956_, new_n16957_, new_n16958_,
    new_n16959_, new_n16960_, new_n16961_, new_n16962_, new_n16963_,
    new_n16964_, new_n16965_, new_n16966_, new_n16967_, new_n16968_,
    new_n16969_, new_n16970_, new_n16971_, new_n16972_, new_n16973_,
    new_n16974_, new_n16975_, new_n16976_, new_n16977_, new_n16978_,
    new_n16979_, new_n16980_, new_n16981_, new_n16982_, new_n16983_,
    new_n16984_, new_n16985_, new_n16986_, new_n16987_, new_n16988_,
    new_n16989_, new_n16990_, new_n16991_, new_n16992_, new_n16993_,
    new_n16994_, new_n16995_, new_n16996_, new_n16997_, new_n16998_,
    new_n16999_, new_n17000_, new_n17001_, new_n17002_, new_n17003_,
    new_n17004_, new_n17005_, new_n17006_, new_n17007_, new_n17008_,
    new_n17009_, new_n17010_, new_n17011_, new_n17012_, new_n17013_,
    new_n17014_, new_n17015_, new_n17016_, new_n17017_, new_n17018_,
    new_n17019_, new_n17020_, new_n17021_, new_n17022_, new_n17023_,
    new_n17024_, new_n17025_, new_n17026_, new_n17027_, new_n17028_,
    new_n17029_, new_n17030_, new_n17031_, new_n17032_, new_n17033_,
    new_n17034_, new_n17035_, new_n17036_, new_n17037_, new_n17038_,
    new_n17039_, new_n17040_, new_n17041_, new_n17042_, new_n17043_,
    new_n17044_, new_n17045_, new_n17046_, new_n17047_, new_n17048_,
    new_n17049_, new_n17050_, new_n17051_, new_n17052_, new_n17054_,
    new_n17055_, new_n17056_, new_n17057_, new_n17058_, new_n17059_,
    new_n17060_, new_n17061_, new_n17062_, new_n17063_, new_n17064_,
    new_n17065_, new_n17066_, new_n17067_, new_n17068_, new_n17069_,
    new_n17070_, new_n17071_, new_n17072_, new_n17073_, new_n17074_,
    new_n17075_, new_n17076_, new_n17077_, new_n17078_, new_n17079_,
    new_n17080_, new_n17081_, new_n17082_, new_n17083_, new_n17084_,
    new_n17085_, new_n17086_, new_n17087_, new_n17088_, new_n17089_,
    new_n17090_, new_n17091_, new_n17092_, new_n17093_, new_n17094_,
    new_n17095_, new_n17096_, new_n17097_, new_n17098_, new_n17099_,
    new_n17100_, new_n17101_, new_n17102_, new_n17103_, new_n17104_,
    new_n17105_, new_n17106_, new_n17107_, new_n17108_, new_n17109_,
    new_n17110_, new_n17111_, new_n17112_, new_n17113_, new_n17114_,
    new_n17115_, new_n17116_, new_n17117_, new_n17118_, new_n17119_,
    new_n17120_, new_n17121_, new_n17122_, new_n17123_, new_n17124_,
    new_n17125_, new_n17126_, new_n17127_, new_n17128_, new_n17129_,
    new_n17130_, new_n17131_, new_n17132_, new_n17133_, new_n17134_,
    new_n17135_, new_n17136_, new_n17137_, new_n17138_, new_n17139_,
    new_n17140_, new_n17141_, new_n17142_, new_n17143_, new_n17144_,
    new_n17145_, new_n17146_, new_n17147_, new_n17148_, new_n17149_,
    new_n17150_, new_n17151_, new_n17152_, new_n17153_, new_n17154_,
    new_n17155_, new_n17156_, new_n17157_, new_n17158_, new_n17159_,
    new_n17160_, new_n17161_, new_n17162_, new_n17163_, new_n17164_,
    new_n17165_, new_n17166_, new_n17167_, new_n17168_, new_n17169_,
    new_n17170_, new_n17171_, new_n17172_, new_n17173_, new_n17174_,
    new_n17175_, new_n17176_, new_n17177_, new_n17178_, new_n17179_,
    new_n17180_, new_n17181_, new_n17182_, new_n17183_, new_n17184_,
    new_n17185_, new_n17186_, new_n17187_, new_n17188_, new_n17189_,
    new_n17190_, new_n17191_, new_n17192_, new_n17193_, new_n17194_,
    new_n17195_, new_n17196_, new_n17197_, new_n17198_, new_n17199_,
    new_n17200_, new_n17201_, new_n17202_, new_n17203_, new_n17204_,
    new_n17205_, new_n17206_, new_n17207_, new_n17208_, new_n17209_,
    new_n17210_, new_n17211_, new_n17212_, new_n17213_, new_n17214_,
    new_n17215_, new_n17216_, new_n17217_, new_n17218_, new_n17219_,
    new_n17220_, new_n17221_, new_n17222_, new_n17223_, new_n17224_,
    new_n17225_, new_n17226_, new_n17227_, new_n17228_, new_n17229_,
    new_n17230_, new_n17231_, new_n17232_, new_n17233_, new_n17234_,
    new_n17235_, new_n17236_, new_n17237_, new_n17238_, new_n17239_,
    new_n17240_, new_n17241_, new_n17242_, new_n17243_, new_n17244_,
    new_n17245_, new_n17246_, new_n17247_, new_n17248_, new_n17249_,
    new_n17250_, new_n17251_, new_n17252_, new_n17253_, new_n17254_,
    new_n17255_, new_n17256_, new_n17257_, new_n17258_, new_n17259_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17283_, new_n17284_, new_n17285_,
    new_n17286_, new_n17287_, new_n17288_, new_n17289_, new_n17290_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17345_,
    new_n17346_, new_n17347_, new_n17348_, new_n17349_, new_n17350_,
    new_n17351_, new_n17352_, new_n17353_, new_n17354_, new_n17355_,
    new_n17356_, new_n17357_, new_n17358_, new_n17359_, new_n17360_,
    new_n17361_, new_n17362_, new_n17363_, new_n17364_, new_n17365_,
    new_n17366_, new_n17367_, new_n17368_, new_n17369_, new_n17370_,
    new_n17371_, new_n17372_, new_n17373_, new_n17374_, new_n17375_,
    new_n17376_, new_n17377_, new_n17378_, new_n17379_, new_n17380_,
    new_n17381_, new_n17382_, new_n17383_, new_n17384_, new_n17385_,
    new_n17386_, new_n17387_, new_n17388_, new_n17389_, new_n17390_,
    new_n17391_, new_n17392_, new_n17393_, new_n17394_, new_n17395_,
    new_n17396_, new_n17397_, new_n17398_, new_n17399_, new_n17400_,
    new_n17401_, new_n17402_, new_n17403_, new_n17404_, new_n17405_,
    new_n17406_, new_n17407_, new_n17408_, new_n17409_, new_n17410_,
    new_n17411_, new_n17412_, new_n17413_, new_n17414_, new_n17415_,
    new_n17416_, new_n17417_, new_n17418_, new_n17419_, new_n17420_,
    new_n17421_, new_n17422_, new_n17423_, new_n17424_, new_n17425_,
    new_n17426_, new_n17427_, new_n17428_, new_n17429_, new_n17430_,
    new_n17431_, new_n17432_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17438_, new_n17439_, new_n17440_,
    new_n17441_, new_n17442_, new_n17443_, new_n17444_, new_n17445_,
    new_n17446_, new_n17447_, new_n17448_, new_n17449_, new_n17450_,
    new_n17451_, new_n17453_, new_n17454_, new_n17455_, new_n17456_,
    new_n17457_, new_n17458_, new_n17459_, new_n17460_, new_n17461_,
    new_n17462_, new_n17463_, new_n17464_, new_n17465_, new_n17466_,
    new_n17467_, new_n17468_, new_n17469_, new_n17470_, new_n17471_,
    new_n17472_, new_n17473_, new_n17474_, new_n17475_, new_n17476_,
    new_n17477_, new_n17478_, new_n17479_, new_n17480_, new_n17481_,
    new_n17482_, new_n17483_, new_n17484_, new_n17485_, new_n17486_,
    new_n17487_, new_n17488_, new_n17489_, new_n17490_, new_n17491_,
    new_n17492_, new_n17493_, new_n17494_, new_n17495_, new_n17496_,
    new_n17497_, new_n17498_, new_n17499_, new_n17500_, new_n17501_,
    new_n17502_, new_n17503_, new_n17504_, new_n17505_, new_n17506_,
    new_n17507_, new_n17508_, new_n17509_, new_n17510_, new_n17511_,
    new_n17512_, new_n17513_, new_n17514_, new_n17515_, new_n17516_,
    new_n17517_, new_n17518_, new_n17519_, new_n17520_, new_n17521_,
    new_n17522_, new_n17523_, new_n17524_, new_n17525_, new_n17526_,
    new_n17527_, new_n17528_, new_n17529_, new_n17530_, new_n17531_,
    new_n17532_, new_n17533_, new_n17534_, new_n17535_, new_n17536_,
    new_n17537_, new_n17538_, new_n17539_, new_n17540_, new_n17541_,
    new_n17542_, new_n17543_, new_n17544_, new_n17545_, new_n17546_,
    new_n17547_, new_n17548_, new_n17549_, new_n17550_, new_n17551_,
    new_n17552_, new_n17553_, new_n17554_, new_n17555_, new_n17556_,
    new_n17557_, new_n17558_, new_n17559_, new_n17560_, new_n17561_,
    new_n17562_, new_n17563_, new_n17564_, new_n17565_, new_n17566_,
    new_n17567_, new_n17568_, new_n17569_, new_n17570_, new_n17571_,
    new_n17572_, new_n17573_, new_n17574_, new_n17575_, new_n17576_,
    new_n17577_, new_n17578_, new_n17579_, new_n17580_, new_n17581_,
    new_n17582_, new_n17583_, new_n17584_, new_n17585_, new_n17586_,
    new_n17587_, new_n17588_, new_n17589_, new_n17590_, new_n17591_,
    new_n17592_, new_n17593_, new_n17594_, new_n17595_, new_n17596_,
    new_n17597_, new_n17598_, new_n17599_, new_n17600_, new_n17601_,
    new_n17602_, new_n17603_, new_n17604_, new_n17605_, new_n17606_,
    new_n17607_, new_n17608_, new_n17609_, new_n17610_, new_n17611_,
    new_n17612_, new_n17613_, new_n17614_, new_n17615_, new_n17616_,
    new_n17617_, new_n17618_, new_n17619_, new_n17620_, new_n17621_,
    new_n17622_, new_n17623_, new_n17624_, new_n17625_, new_n17626_,
    new_n17627_, new_n17628_, new_n17629_, new_n17630_, new_n17631_,
    new_n17632_, new_n17633_, new_n17634_, new_n17635_, new_n17636_,
    new_n17637_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17653_, new_n17654_, new_n17655_, new_n17656_, new_n17657_,
    new_n17658_, new_n17659_, new_n17660_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17680_, new_n17681_, new_n17682_,
    new_n17683_, new_n17684_, new_n17685_, new_n17686_, new_n17687_,
    new_n17688_, new_n17689_, new_n17690_, new_n17691_, new_n17692_,
    new_n17693_, new_n17694_, new_n17695_, new_n17696_, new_n17697_,
    new_n17698_, new_n17699_, new_n17700_, new_n17701_, new_n17702_,
    new_n17703_, new_n17704_, new_n17705_, new_n17706_, new_n17707_,
    new_n17708_, new_n17709_, new_n17710_, new_n17711_, new_n17712_,
    new_n17713_, new_n17714_, new_n17715_, new_n17716_, new_n17717_,
    new_n17718_, new_n17719_, new_n17720_, new_n17721_, new_n17722_,
    new_n17723_, new_n17724_, new_n17725_, new_n17726_, new_n17727_,
    new_n17728_, new_n17729_, new_n17730_, new_n17731_, new_n17732_,
    new_n17733_, new_n17734_, new_n17735_, new_n17736_, new_n17737_,
    new_n17738_, new_n17739_, new_n17740_, new_n17741_, new_n17742_,
    new_n17743_, new_n17744_, new_n17745_, new_n17746_, new_n17747_,
    new_n17748_, new_n17749_, new_n17750_, new_n17751_, new_n17752_,
    new_n17753_, new_n17754_, new_n17755_, new_n17756_, new_n17757_,
    new_n17758_, new_n17759_, new_n17760_, new_n17761_, new_n17762_,
    new_n17763_, new_n17764_, new_n17765_, new_n17766_, new_n17767_,
    new_n17768_, new_n17769_, new_n17770_, new_n17771_, new_n17772_,
    new_n17773_, new_n17774_, new_n17775_, new_n17776_, new_n17777_,
    new_n17778_, new_n17779_, new_n17780_, new_n17781_, new_n17782_,
    new_n17783_, new_n17784_, new_n17785_, new_n17786_, new_n17787_,
    new_n17788_, new_n17789_, new_n17790_, new_n17791_, new_n17792_,
    new_n17793_, new_n17794_, new_n17795_, new_n17796_, new_n17797_,
    new_n17798_, new_n17799_, new_n17800_, new_n17801_, new_n17802_,
    new_n17803_, new_n17804_, new_n17805_, new_n17806_, new_n17807_,
    new_n17808_, new_n17809_, new_n17810_, new_n17811_, new_n17812_,
    new_n17813_, new_n17814_, new_n17816_, new_n17817_, new_n17818_,
    new_n17819_, new_n17820_, new_n17821_, new_n17822_, new_n17823_,
    new_n17824_, new_n17825_, new_n17826_, new_n17827_, new_n17828_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17834_, new_n17835_, new_n17836_, new_n17837_, new_n17838_,
    new_n17839_, new_n17840_, new_n17841_, new_n17842_, new_n17843_,
    new_n17844_, new_n17845_, new_n17846_, new_n17847_, new_n17848_,
    new_n17849_, new_n17850_, new_n17851_, new_n17852_, new_n17853_,
    new_n17854_, new_n17855_, new_n17856_, new_n17857_, new_n17858_,
    new_n17859_, new_n17860_, new_n17861_, new_n17862_, new_n17863_,
    new_n17864_, new_n17865_, new_n17866_, new_n17867_, new_n17868_,
    new_n17869_, new_n17870_, new_n17871_, new_n17872_, new_n17873_,
    new_n17874_, new_n17875_, new_n17876_, new_n17877_, new_n17878_,
    new_n17879_, new_n17880_, new_n17881_, new_n17882_, new_n17883_,
    new_n17884_, new_n17885_, new_n17886_, new_n17887_, new_n17888_,
    new_n17889_, new_n17890_, new_n17891_, new_n17892_, new_n17893_,
    new_n17894_, new_n17895_, new_n17896_, new_n17897_, new_n17898_,
    new_n17899_, new_n17900_, new_n17901_, new_n17902_, new_n17903_,
    new_n17904_, new_n17905_, new_n17906_, new_n17907_, new_n17908_,
    new_n17909_, new_n17910_, new_n17911_, new_n17912_, new_n17913_,
    new_n17914_, new_n17915_, new_n17916_, new_n17917_, new_n17918_,
    new_n17919_, new_n17920_, new_n17921_, new_n17922_, new_n17923_,
    new_n17924_, new_n17925_, new_n17926_, new_n17927_, new_n17928_,
    new_n17929_, new_n17930_, new_n17931_, new_n17932_, new_n17933_,
    new_n17934_, new_n17935_, new_n17936_, new_n17937_, new_n17938_,
    new_n17939_, new_n17940_, new_n17941_, new_n17942_, new_n17943_,
    new_n17944_, new_n17945_, new_n17946_, new_n17947_, new_n17948_,
    new_n17949_, new_n17950_, new_n17951_, new_n17952_, new_n17953_,
    new_n17954_, new_n17955_, new_n17956_, new_n17957_, new_n17958_,
    new_n17959_, new_n17960_, new_n17961_, new_n17962_, new_n17963_,
    new_n17964_, new_n17965_, new_n17966_, new_n17967_, new_n17968_,
    new_n17969_, new_n17970_, new_n17971_, new_n17972_, new_n17973_,
    new_n17974_, new_n17975_, new_n17976_, new_n17977_, new_n17978_,
    new_n17979_, new_n17980_, new_n17981_, new_n17982_, new_n17983_,
    new_n17984_, new_n17985_, new_n17986_, new_n17987_, new_n17988_,
    new_n17989_, new_n17990_, new_n17991_, new_n17992_, new_n17994_,
    new_n17995_, new_n17996_, new_n17997_, new_n17998_, new_n17999_,
    new_n18000_, new_n18001_, new_n18002_, new_n18003_, new_n18004_,
    new_n18005_, new_n18006_, new_n18007_, new_n18008_, new_n18009_,
    new_n18010_, new_n18011_, new_n18012_, new_n18013_, new_n18014_,
    new_n18015_, new_n18016_, new_n18017_, new_n18018_, new_n18019_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18025_, new_n18026_, new_n18027_, new_n18028_, new_n18029_,
    new_n18030_, new_n18031_, new_n18032_, new_n18033_, new_n18034_,
    new_n18035_, new_n18036_, new_n18037_, new_n18038_, new_n18039_,
    new_n18040_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18108_, new_n18109_,
    new_n18110_, new_n18111_, new_n18112_, new_n18113_, new_n18114_,
    new_n18115_, new_n18116_, new_n18117_, new_n18118_, new_n18119_,
    new_n18120_, new_n18121_, new_n18122_, new_n18123_, new_n18124_,
    new_n18125_, new_n18126_, new_n18127_, new_n18128_, new_n18129_,
    new_n18130_, new_n18131_, new_n18132_, new_n18133_, new_n18134_,
    new_n18135_, new_n18136_, new_n18137_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18170_,
    new_n18171_, new_n18172_, new_n18173_, new_n18174_, new_n18175_,
    new_n18176_, new_n18177_, new_n18178_, new_n18179_, new_n18180_,
    new_n18181_, new_n18182_, new_n18183_, new_n18184_, new_n18185_,
    new_n18186_, new_n18187_, new_n18188_, new_n18189_, new_n18190_,
    new_n18191_, new_n18192_, new_n18193_, new_n18194_, new_n18195_,
    new_n18196_, new_n18197_, new_n18198_, new_n18199_, new_n18200_,
    new_n18201_, new_n18202_, new_n18203_, new_n18204_, new_n18205_,
    new_n18206_, new_n18207_, new_n18208_, new_n18209_, new_n18210_,
    new_n18211_, new_n18212_, new_n18213_, new_n18214_, new_n18215_,
    new_n18216_, new_n18217_, new_n18218_, new_n18219_, new_n18220_,
    new_n18221_, new_n18222_, new_n18223_, new_n18224_, new_n18225_,
    new_n18226_, new_n18227_, new_n18228_, new_n18229_, new_n18230_,
    new_n18231_, new_n18232_, new_n18233_, new_n18234_, new_n18235_,
    new_n18236_, new_n18237_, new_n18238_, new_n18239_, new_n18240_,
    new_n18241_, new_n18242_, new_n18243_, new_n18244_, new_n18245_,
    new_n18246_, new_n18247_, new_n18248_, new_n18249_, new_n18250_,
    new_n18251_, new_n18252_, new_n18253_, new_n18254_, new_n18255_,
    new_n18256_, new_n18257_, new_n18258_, new_n18259_, new_n18260_,
    new_n18261_, new_n18262_, new_n18263_, new_n18264_, new_n18265_,
    new_n18266_, new_n18267_, new_n18268_, new_n18269_, new_n18270_,
    new_n18271_, new_n18272_, new_n18273_, new_n18274_, new_n18275_,
    new_n18276_, new_n18277_, new_n18278_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18339_, new_n18340_, new_n18341_,
    new_n18342_, new_n18343_, new_n18344_, new_n18345_, new_n18346_,
    new_n18347_, new_n18348_, new_n18349_, new_n18350_, new_n18351_,
    new_n18352_, new_n18353_, new_n18354_, new_n18355_, new_n18356_,
    new_n18357_, new_n18358_, new_n18359_, new_n18360_, new_n18361_,
    new_n18362_, new_n18363_, new_n18364_, new_n18365_, new_n18366_,
    new_n18367_, new_n18368_, new_n18369_, new_n18370_, new_n18371_,
    new_n18372_, new_n18373_, new_n18374_, new_n18375_, new_n18376_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18393_, new_n18394_, new_n18395_, new_n18396_,
    new_n18397_, new_n18398_, new_n18399_, new_n18400_, new_n18401_,
    new_n18402_, new_n18403_, new_n18404_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18409_, new_n18410_, new_n18411_,
    new_n18412_, new_n18413_, new_n18414_, new_n18415_, new_n18416_,
    new_n18417_, new_n18418_, new_n18419_, new_n18420_, new_n18421_,
    new_n18422_, new_n18423_, new_n18424_, new_n18425_, new_n18426_,
    new_n18427_, new_n18428_, new_n18429_, new_n18430_, new_n18431_,
    new_n18432_, new_n18433_, new_n18434_, new_n18435_, new_n18436_,
    new_n18437_, new_n18438_, new_n18439_, new_n18440_, new_n18441_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18501_, new_n18502_,
    new_n18503_, new_n18504_, new_n18505_, new_n18506_, new_n18507_,
    new_n18508_, new_n18509_, new_n18510_, new_n18511_, new_n18512_,
    new_n18513_, new_n18514_, new_n18515_, new_n18516_, new_n18517_,
    new_n18518_, new_n18519_, new_n18520_, new_n18521_, new_n18522_,
    new_n18523_, new_n18524_, new_n18525_, new_n18526_, new_n18527_,
    new_n18528_, new_n18529_, new_n18530_, new_n18531_, new_n18532_,
    new_n18533_, new_n18534_, new_n18535_, new_n18536_, new_n18537_,
    new_n18538_, new_n18539_, new_n18540_, new_n18541_, new_n18542_,
    new_n18543_, new_n18544_, new_n18545_, new_n18546_, new_n18547_,
    new_n18548_, new_n18549_, new_n18550_, new_n18551_, new_n18552_,
    new_n18553_, new_n18554_, new_n18555_, new_n18556_, new_n18557_,
    new_n18558_, new_n18559_, new_n18560_, new_n18561_, new_n18562_,
    new_n18563_, new_n18564_, new_n18565_, new_n18566_, new_n18567_,
    new_n18568_, new_n18569_, new_n18570_, new_n18571_, new_n18572_,
    new_n18573_, new_n18574_, new_n18575_, new_n18576_, new_n18577_,
    new_n18578_, new_n18579_, new_n18580_, new_n18581_, new_n18582_,
    new_n18583_, new_n18584_, new_n18585_, new_n18586_, new_n18587_,
    new_n18588_, new_n18589_, new_n18590_, new_n18591_, new_n18592_,
    new_n18593_, new_n18594_, new_n18595_, new_n18596_, new_n18597_,
    new_n18598_, new_n18599_, new_n18600_, new_n18601_, new_n18602_,
    new_n18603_, new_n18604_, new_n18605_, new_n18606_, new_n18607_,
    new_n18608_, new_n18609_, new_n18610_, new_n18611_, new_n18612_,
    new_n18613_, new_n18614_, new_n18615_, new_n18616_, new_n18617_,
    new_n18618_, new_n18619_, new_n18620_, new_n18621_, new_n18622_,
    new_n18623_, new_n18624_, new_n18625_, new_n18626_, new_n18627_,
    new_n18628_, new_n18629_, new_n18630_, new_n18631_, new_n18632_,
    new_n18633_, new_n18634_, new_n18635_, new_n18636_, new_n18637_,
    new_n18638_, new_n18639_, new_n18640_, new_n18641_, new_n18642_,
    new_n18643_, new_n18645_, new_n18646_, new_n18647_, new_n18648_,
    new_n18649_, new_n18650_, new_n18651_, new_n18652_, new_n18653_,
    new_n18654_, new_n18655_, new_n18656_, new_n18657_, new_n18658_,
    new_n18659_, new_n18660_, new_n18661_, new_n18662_, new_n18663_,
    new_n18664_, new_n18665_, new_n18666_, new_n18667_, new_n18668_,
    new_n18669_, new_n18670_, new_n18671_, new_n18672_, new_n18673_,
    new_n18674_, new_n18675_, new_n18676_, new_n18677_, new_n18678_,
    new_n18679_, new_n18680_, new_n18681_, new_n18682_, new_n18683_,
    new_n18684_, new_n18685_, new_n18686_, new_n18687_, new_n18688_,
    new_n18689_, new_n18690_, new_n18691_, new_n18692_, new_n18693_,
    new_n18694_, new_n18695_, new_n18696_, new_n18697_, new_n18698_,
    new_n18699_, new_n18700_, new_n18701_, new_n18702_, new_n18703_,
    new_n18704_, new_n18705_, new_n18706_, new_n18707_, new_n18708_,
    new_n18709_, new_n18710_, new_n18711_, new_n18712_, new_n18713_,
    new_n18714_, new_n18715_, new_n18716_, new_n18717_, new_n18718_,
    new_n18719_, new_n18720_, new_n18721_, new_n18722_, new_n18723_,
    new_n18724_, new_n18725_, new_n18726_, new_n18727_, new_n18728_,
    new_n18729_, new_n18730_, new_n18731_, new_n18732_, new_n18733_,
    new_n18734_, new_n18735_, new_n18736_, new_n18737_, new_n18738_,
    new_n18739_, new_n18740_, new_n18741_, new_n18742_, new_n18743_,
    new_n18744_, new_n18745_, new_n18746_, new_n18747_, new_n18748_,
    new_n18749_, new_n18750_, new_n18751_, new_n18752_, new_n18753_,
    new_n18754_, new_n18755_, new_n18756_, new_n18757_, new_n18758_,
    new_n18759_, new_n18760_, new_n18761_, new_n18762_, new_n18763_,
    new_n18764_, new_n18765_, new_n18766_, new_n18767_, new_n18768_,
    new_n18769_, new_n18770_, new_n18771_, new_n18772_, new_n18773_,
    new_n18774_, new_n18775_, new_n18776_, new_n18777_, new_n18778_,
    new_n18779_, new_n18780_, new_n18781_, new_n18782_, new_n18783_,
    new_n18784_, new_n18785_, new_n18786_, new_n18787_, new_n18788_,
    new_n18789_, new_n18790_, new_n18791_, new_n18792_, new_n18793_,
    new_n18794_, new_n18795_, new_n18796_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19090_, new_n19091_,
    new_n19092_, new_n19093_, new_n19094_, new_n19095_, new_n19096_,
    new_n19097_, new_n19098_, new_n19099_, new_n19100_, new_n19101_,
    new_n19102_, new_n19103_, new_n19104_, new_n19105_, new_n19106_,
    new_n19107_, new_n19108_, new_n19109_, new_n19110_, new_n19111_,
    new_n19112_, new_n19113_, new_n19114_, new_n19115_, new_n19116_,
    new_n19117_, new_n19118_, new_n19119_, new_n19120_, new_n19121_,
    new_n19122_, new_n19123_, new_n19124_, new_n19125_, new_n19126_,
    new_n19127_, new_n19128_, new_n19129_, new_n19130_, new_n19131_,
    new_n19132_, new_n19133_, new_n19134_, new_n19135_, new_n19136_,
    new_n19137_, new_n19138_, new_n19139_, new_n19140_, new_n19141_,
    new_n19142_, new_n19143_, new_n19144_, new_n19145_, new_n19146_,
    new_n19147_, new_n19148_, new_n19149_, new_n19150_, new_n19151_,
    new_n19152_, new_n19153_, new_n19154_, new_n19155_, new_n19156_,
    new_n19157_, new_n19158_, new_n19159_, new_n19160_, new_n19161_,
    new_n19162_, new_n19163_, new_n19164_, new_n19165_, new_n19166_,
    new_n19167_, new_n19168_, new_n19169_, new_n19170_, new_n19171_,
    new_n19172_, new_n19173_, new_n19174_, new_n19175_, new_n19176_,
    new_n19177_, new_n19178_, new_n19179_, new_n19180_, new_n19181_,
    new_n19182_, new_n19183_, new_n19184_, new_n19185_, new_n19186_,
    new_n19187_, new_n19188_, new_n19189_, new_n19190_, new_n19191_,
    new_n19192_, new_n19193_, new_n19194_, new_n19195_, new_n19196_,
    new_n19197_, new_n19198_, new_n19199_, new_n19200_, new_n19201_,
    new_n19202_, new_n19203_, new_n19204_, new_n19205_, new_n19206_,
    new_n19207_, new_n19208_, new_n19209_, new_n19210_, new_n19211_,
    new_n19212_, new_n19213_, new_n19214_, new_n19215_, new_n19216_,
    new_n19217_, new_n19218_, new_n19219_, new_n19220_, new_n19221_,
    new_n19222_, new_n19223_, new_n19224_, new_n19225_, new_n19226_,
    new_n19228_, new_n19229_, new_n19230_, new_n19231_, new_n19232_,
    new_n19233_, new_n19234_, new_n19235_, new_n19236_, new_n19237_,
    new_n19238_, new_n19239_, new_n19240_, new_n19241_, new_n19242_,
    new_n19243_, new_n19244_, new_n19245_, new_n19246_, new_n19247_,
    new_n19248_, new_n19249_, new_n19250_, new_n19251_, new_n19252_,
    new_n19253_, new_n19254_, new_n19255_, new_n19256_, new_n19257_,
    new_n19258_, new_n19259_, new_n19260_, new_n19261_, new_n19262_,
    new_n19263_, new_n19264_, new_n19265_, new_n19266_, new_n19267_,
    new_n19268_, new_n19269_, new_n19270_, new_n19271_, new_n19272_,
    new_n19273_, new_n19274_, new_n19275_, new_n19276_, new_n19277_,
    new_n19278_, new_n19279_, new_n19280_, new_n19281_, new_n19282_,
    new_n19283_, new_n19284_, new_n19285_, new_n19286_, new_n19287_,
    new_n19288_, new_n19289_, new_n19290_, new_n19291_, new_n19292_,
    new_n19293_, new_n19294_, new_n19295_, new_n19296_, new_n19297_,
    new_n19298_, new_n19299_, new_n19300_, new_n19301_, new_n19302_,
    new_n19303_, new_n19304_, new_n19305_, new_n19306_, new_n19307_,
    new_n19308_, new_n19309_, new_n19310_, new_n19311_, new_n19312_,
    new_n19313_, new_n19314_, new_n19315_, new_n19316_, new_n19317_,
    new_n19318_, new_n19319_, new_n19320_, new_n19321_, new_n19322_,
    new_n19323_, new_n19324_, new_n19325_, new_n19326_, new_n19327_,
    new_n19328_, new_n19329_, new_n19330_, new_n19331_, new_n19332_,
    new_n19333_, new_n19334_, new_n19335_, new_n19336_, new_n19337_,
    new_n19338_, new_n19339_, new_n19340_, new_n19341_, new_n19342_,
    new_n19343_, new_n19344_, new_n19345_, new_n19346_, new_n19347_,
    new_n19348_, new_n19349_, new_n19350_, new_n19351_, new_n19352_,
    new_n19353_, new_n19354_, new_n19355_, new_n19356_, new_n19357_,
    new_n19358_, new_n19359_, new_n19360_, new_n19361_, new_n19362_,
    new_n19363_, new_n19364_, new_n19365_, new_n19367_, new_n19368_,
    new_n19369_, new_n19370_, new_n19371_, new_n19372_, new_n19373_,
    new_n19374_, new_n19375_, new_n19376_, new_n19377_, new_n19378_,
    new_n19379_, new_n19380_, new_n19381_, new_n19382_, new_n19383_,
    new_n19384_, new_n19385_, new_n19386_, new_n19387_, new_n19388_,
    new_n19389_, new_n19390_, new_n19391_, new_n19392_, new_n19393_,
    new_n19394_, new_n19395_, new_n19396_, new_n19397_, new_n19398_,
    new_n19399_, new_n19400_, new_n19401_, new_n19402_, new_n19403_,
    new_n19404_, new_n19405_, new_n19406_, new_n19407_, new_n19408_,
    new_n19409_, new_n19410_, new_n19411_, new_n19412_, new_n19413_,
    new_n19414_, new_n19415_, new_n19416_, new_n19417_, new_n19418_,
    new_n19419_, new_n19420_, new_n19421_, new_n19422_, new_n19423_,
    new_n19424_, new_n19425_, new_n19426_, new_n19427_, new_n19428_,
    new_n19429_, new_n19430_, new_n19431_, new_n19432_, new_n19433_,
    new_n19434_, new_n19435_, new_n19436_, new_n19437_, new_n19438_,
    new_n19439_, new_n19440_, new_n19441_, new_n19442_, new_n19443_,
    new_n19444_, new_n19445_, new_n19446_, new_n19447_, new_n19448_,
    new_n19449_, new_n19450_, new_n19451_, new_n19452_, new_n19453_,
    new_n19454_, new_n19455_, new_n19456_, new_n19457_, new_n19458_,
    new_n19459_, new_n19460_, new_n19461_, new_n19462_, new_n19463_,
    new_n19464_, new_n19465_, new_n19466_, new_n19467_, new_n19468_,
    new_n19469_, new_n19470_, new_n19471_, new_n19472_, new_n19473_,
    new_n19474_, new_n19475_, new_n19476_, new_n19477_, new_n19478_,
    new_n19479_, new_n19480_, new_n19481_, new_n19482_, new_n19483_,
    new_n19484_, new_n19485_, new_n19486_, new_n19487_, new_n19488_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19531_, new_n19532_, new_n19533_, new_n19534_,
    new_n19535_, new_n19536_, new_n19537_, new_n19538_, new_n19539_,
    new_n19540_, new_n19541_, new_n19542_, new_n19543_, new_n19544_,
    new_n19545_, new_n19546_, new_n19547_, new_n19548_, new_n19549_,
    new_n19550_, new_n19551_, new_n19552_, new_n19553_, new_n19554_,
    new_n19555_, new_n19556_, new_n19557_, new_n19558_, new_n19559_,
    new_n19560_, new_n19561_, new_n19562_, new_n19563_, new_n19564_,
    new_n19565_, new_n19566_, new_n19567_, new_n19568_, new_n19569_,
    new_n19570_, new_n19571_, new_n19572_, new_n19573_, new_n19574_,
    new_n19575_, new_n19576_, new_n19577_, new_n19578_, new_n19579_,
    new_n19580_, new_n19581_, new_n19582_, new_n19583_, new_n19584_,
    new_n19585_, new_n19586_, new_n19587_, new_n19588_, new_n19589_,
    new_n19590_, new_n19591_, new_n19592_, new_n19593_, new_n19594_,
    new_n19595_, new_n19596_, new_n19597_, new_n19598_, new_n19599_,
    new_n19600_, new_n19601_, new_n19602_, new_n19603_, new_n19604_,
    new_n19605_, new_n19606_, new_n19607_, new_n19608_, new_n19609_,
    new_n19610_, new_n19611_, new_n19612_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19841_, new_n19842_,
    new_n19843_, new_n19844_, new_n19845_, new_n19846_, new_n19847_,
    new_n19848_, new_n19849_, new_n19850_, new_n19851_, new_n19852_,
    new_n19853_, new_n19854_, new_n19855_, new_n19856_, new_n19857_,
    new_n19858_, new_n19859_, new_n19860_, new_n19861_, new_n19862_,
    new_n19863_, new_n19864_, new_n19865_, new_n19866_, new_n19867_,
    new_n19868_, new_n19869_, new_n19870_, new_n19871_, new_n19872_,
    new_n19873_, new_n19874_, new_n19875_, new_n19876_, new_n19877_,
    new_n19878_, new_n19879_, new_n19880_, new_n19881_, new_n19882_,
    new_n19883_, new_n19884_, new_n19885_, new_n19886_, new_n19887_,
    new_n19888_, new_n19889_, new_n19890_, new_n19891_, new_n19892_,
    new_n19893_, new_n19894_, new_n19895_, new_n19896_, new_n19897_,
    new_n19898_, new_n19899_, new_n19900_, new_n19901_, new_n19902_,
    new_n19903_, new_n19904_, new_n19905_, new_n19906_, new_n19907_,
    new_n19908_, new_n19909_, new_n19910_, new_n19911_, new_n19912_,
    new_n19913_, new_n19914_, new_n19915_, new_n19916_, new_n19917_,
    new_n19918_, new_n19919_, new_n19920_, new_n19921_, new_n19922_,
    new_n19923_, new_n19924_, new_n19925_, new_n19926_, new_n19927_,
    new_n19928_, new_n19929_, new_n19930_, new_n19931_, new_n19932_,
    new_n19933_, new_n19934_, new_n19935_, new_n19936_, new_n19937_,
    new_n19938_, new_n19939_, new_n19940_, new_n19941_, new_n19942_,
    new_n19943_, new_n19944_, new_n19945_, new_n19946_, new_n19947_,
    new_n19948_, new_n19950_, new_n19951_, new_n19952_, new_n19953_,
    new_n19954_, new_n19955_, new_n19956_, new_n19957_, new_n19958_,
    new_n19959_, new_n19960_, new_n19961_, new_n19962_, new_n19963_,
    new_n19964_, new_n19965_, new_n19966_, new_n19967_, new_n19968_,
    new_n19969_, new_n19970_, new_n19971_, new_n19972_, new_n19973_,
    new_n19974_, new_n19975_, new_n19976_, new_n19977_, new_n19978_,
    new_n19979_, new_n19980_, new_n19981_, new_n19982_, new_n19983_,
    new_n19984_, new_n19985_, new_n19986_, new_n19987_, new_n19988_,
    new_n19989_, new_n19990_, new_n19991_, new_n19992_, new_n19993_,
    new_n19994_, new_n19995_, new_n19996_, new_n19997_, new_n19998_,
    new_n19999_, new_n20000_, new_n20001_, new_n20002_, new_n20003_,
    new_n20004_, new_n20005_, new_n20006_, new_n20007_, new_n20008_,
    new_n20009_, new_n20010_, new_n20011_, new_n20012_, new_n20013_,
    new_n20014_, new_n20015_, new_n20016_, new_n20017_, new_n20018_,
    new_n20019_, new_n20020_, new_n20021_, new_n20022_, new_n20023_,
    new_n20024_, new_n20025_, new_n20026_, new_n20027_, new_n20028_,
    new_n20029_, new_n20030_, new_n20031_, new_n20032_, new_n20033_,
    new_n20034_, new_n20035_, new_n20036_, new_n20037_, new_n20038_,
    new_n20039_, new_n20040_, new_n20041_, new_n20042_, new_n20043_,
    new_n20044_, new_n20045_, new_n20046_, new_n20047_, new_n20048_,
    new_n20049_, new_n20050_, new_n20051_, new_n20052_, new_n20053_,
    new_n20054_, new_n20056_, new_n20057_, new_n20058_, new_n20059_,
    new_n20060_, new_n20061_, new_n20062_, new_n20063_, new_n20064_,
    new_n20065_, new_n20066_, new_n20067_, new_n20068_, new_n20069_,
    new_n20070_, new_n20071_, new_n20072_, new_n20073_, new_n20074_,
    new_n20075_, new_n20076_, new_n20077_, new_n20078_, new_n20079_,
    new_n20080_, new_n20081_, new_n20082_, new_n20083_, new_n20084_,
    new_n20085_, new_n20086_, new_n20087_, new_n20088_, new_n20089_,
    new_n20090_, new_n20091_, new_n20092_, new_n20093_, new_n20094_,
    new_n20095_, new_n20096_, new_n20097_, new_n20098_, new_n20099_,
    new_n20100_, new_n20101_, new_n20102_, new_n20103_, new_n20104_,
    new_n20105_, new_n20106_, new_n20107_, new_n20108_, new_n20109_,
    new_n20110_, new_n20111_, new_n20112_, new_n20113_, new_n20114_,
    new_n20115_, new_n20116_, new_n20117_, new_n20118_, new_n20119_,
    new_n20120_, new_n20121_, new_n20122_, new_n20123_, new_n20124_,
    new_n20125_, new_n20126_, new_n20127_, new_n20128_, new_n20129_,
    new_n20130_, new_n20131_, new_n20132_, new_n20133_, new_n20134_,
    new_n20135_, new_n20136_, new_n20137_, new_n20138_, new_n20139_,
    new_n20140_, new_n20141_, new_n20142_, new_n20143_, new_n20144_,
    new_n20145_, new_n20146_, new_n20148_, new_n20149_, new_n20150_,
    new_n20151_, new_n20152_, new_n20153_, new_n20154_, new_n20155_,
    new_n20156_, new_n20157_, new_n20158_, new_n20159_, new_n20160_,
    new_n20161_, new_n20162_, new_n20163_, new_n20164_, new_n20165_,
    new_n20166_, new_n20167_, new_n20168_, new_n20169_, new_n20170_,
    new_n20171_, new_n20172_, new_n20173_, new_n20174_, new_n20175_,
    new_n20176_, new_n20177_, new_n20178_, new_n20179_, new_n20180_,
    new_n20181_, new_n20182_, new_n20183_, new_n20184_, new_n20185_,
    new_n20186_, new_n20187_, new_n20188_, new_n20189_, new_n20190_,
    new_n20191_, new_n20192_, new_n20193_, new_n20194_, new_n20195_,
    new_n20196_, new_n20197_, new_n20198_, new_n20199_, new_n20200_,
    new_n20201_, new_n20202_, new_n20203_, new_n20204_, new_n20205_,
    new_n20206_, new_n20207_, new_n20208_, new_n20209_, new_n20210_,
    new_n20211_, new_n20212_, new_n20213_, new_n20214_, new_n20215_,
    new_n20216_, new_n20217_, new_n20218_, new_n20219_, new_n20220_,
    new_n20221_, new_n20222_, new_n20223_, new_n20224_, new_n20225_,
    new_n20226_, new_n20227_, new_n20228_, new_n20229_, new_n20230_,
    new_n20231_, new_n20232_, new_n20233_, new_n20234_, new_n20235_,
    new_n20236_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20296_,
    new_n20297_, new_n20298_, new_n20299_, new_n20300_, new_n20301_,
    new_n20302_, new_n20303_, new_n20304_, new_n20305_, new_n20306_,
    new_n20307_, new_n20308_, new_n20309_, new_n20310_, new_n20311_,
    new_n20312_, new_n20313_, new_n20314_, new_n20315_, new_n20316_,
    new_n20317_, new_n20318_, new_n20319_, new_n20320_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20376_, new_n20377_,
    new_n20378_, new_n20379_, new_n20380_, new_n20381_, new_n20382_,
    new_n20383_, new_n20384_, new_n20385_, new_n20386_, new_n20387_,
    new_n20388_, new_n20389_, new_n20390_, new_n20391_, new_n20392_,
    new_n20393_, new_n20394_, new_n20395_, new_n20396_, new_n20397_,
    new_n20398_, new_n20399_, new_n20401_, new_n20402_, new_n20403_,
    new_n20404_, new_n20405_, new_n20406_, new_n20407_, new_n20408_,
    new_n20409_, new_n20410_, new_n20411_, new_n20412_, new_n20413_,
    new_n20414_, new_n20415_, new_n20416_, new_n20417_, new_n20418_,
    new_n20419_, new_n20420_, new_n20421_, new_n20422_, new_n20423_,
    new_n20424_, new_n20425_, new_n20426_, new_n20427_, new_n20428_,
    new_n20429_, new_n20430_, new_n20431_, new_n20432_, new_n20433_,
    new_n20434_, new_n20435_, new_n20436_, new_n20437_, new_n20438_,
    new_n20439_, new_n20440_, new_n20441_, new_n20442_, new_n20443_,
    new_n20444_, new_n20445_, new_n20446_, new_n20447_, new_n20448_,
    new_n20449_, new_n20450_, new_n20451_, new_n20452_, new_n20453_,
    new_n20454_, new_n20455_, new_n20456_, new_n20457_, new_n20458_,
    new_n20459_, new_n20460_, new_n20461_, new_n20462_, new_n20463_,
    new_n20464_, new_n20465_, new_n20466_, new_n20467_, new_n20468_,
    new_n20469_, new_n20470_, new_n20471_, new_n20472_, new_n20473_,
    new_n20474_, new_n20475_, new_n20476_, new_n20477_, new_n20478_,
    new_n20479_, new_n20480_, new_n20482_, new_n20483_, new_n20484_,
    new_n20485_, new_n20486_, new_n20487_, new_n20488_, new_n20489_,
    new_n20490_, new_n20491_, new_n20492_, new_n20493_, new_n20494_,
    new_n20495_, new_n20496_, new_n20497_, new_n20498_, new_n20499_,
    new_n20500_, new_n20501_, new_n20502_, new_n20503_, new_n20504_,
    new_n20505_, new_n20506_, new_n20507_, new_n20508_, new_n20509_,
    new_n20510_, new_n20511_, new_n20512_, new_n20513_, new_n20514_,
    new_n20515_, new_n20516_, new_n20517_, new_n20518_, new_n20519_,
    new_n20520_, new_n20521_, new_n20522_, new_n20523_, new_n20524_,
    new_n20525_, new_n20526_, new_n20527_, new_n20528_, new_n20529_,
    new_n20530_, new_n20531_, new_n20532_, new_n20533_, new_n20534_,
    new_n20535_, new_n20536_, new_n20537_, new_n20538_, new_n20539_,
    new_n20540_, new_n20541_, new_n20542_, new_n20543_, new_n20544_,
    new_n20545_, new_n20546_, new_n20547_, new_n20548_, new_n20549_,
    new_n20550_, new_n20551_, new_n20552_, new_n20553_, new_n20554_,
    new_n20555_, new_n20556_, new_n20557_, new_n20558_, new_n20559_,
    new_n20561_, new_n20562_, new_n20563_, new_n20564_, new_n20565_,
    new_n20566_, new_n20567_, new_n20568_, new_n20569_, new_n20570_,
    new_n20571_, new_n20572_, new_n20573_, new_n20574_, new_n20575_,
    new_n20576_, new_n20577_, new_n20578_, new_n20579_, new_n20580_,
    new_n20581_, new_n20582_, new_n20583_, new_n20584_, new_n20585_,
    new_n20586_, new_n20587_, new_n20588_, new_n20589_, new_n20590_,
    new_n20591_, new_n20592_, new_n20593_, new_n20594_, new_n20595_,
    new_n20596_, new_n20597_, new_n20598_, new_n20599_, new_n20600_,
    new_n20601_, new_n20602_, new_n20603_, new_n20604_, new_n20605_,
    new_n20606_, new_n20607_, new_n20608_, new_n20609_, new_n20610_,
    new_n20611_, new_n20612_, new_n20613_, new_n20614_, new_n20615_,
    new_n20616_, new_n20617_, new_n20618_, new_n20619_, new_n20620_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20677_, new_n20678_, new_n20679_, new_n20680_, new_n20681_,
    new_n20682_, new_n20683_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20713_, new_n20714_, new_n20715_, new_n20716_, new_n20717_,
    new_n20718_, new_n20719_, new_n20720_, new_n20721_, new_n20722_,
    new_n20723_, new_n20724_, new_n20725_, new_n20726_, new_n20727_,
    new_n20728_, new_n20729_, new_n20730_, new_n20731_, new_n20732_,
    new_n20733_, new_n20734_, new_n20735_, new_n20736_, new_n20737_,
    new_n20738_, new_n20739_, new_n20740_, new_n20741_, new_n20743_,
    new_n20744_, new_n20745_, new_n20746_, new_n20747_, new_n20748_,
    new_n20749_, new_n20750_, new_n20751_, new_n20752_, new_n20753_,
    new_n20754_, new_n20755_, new_n20756_, new_n20757_, new_n20758_,
    new_n20759_, new_n20760_, new_n20761_, new_n20762_, new_n20763_,
    new_n20764_, new_n20765_, new_n20766_, new_n20767_, new_n20768_,
    new_n20769_, new_n20770_, new_n20771_, new_n20772_, new_n20773_,
    new_n20774_, new_n20775_, new_n20776_, new_n20777_, new_n20778_,
    new_n20779_, new_n20780_, new_n20781_, new_n20782_, new_n20783_,
    new_n20784_, new_n20785_, new_n20786_, new_n20787_, new_n20788_,
    new_n20789_, new_n20790_, new_n20792_, new_n20793_, new_n20794_,
    new_n20795_, new_n20796_, new_n20797_, new_n20798_, new_n20799_,
    new_n20800_, new_n20801_, new_n20802_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20836_, new_n20837_, new_n20838_, new_n20839_,
    new_n20841_, new_n20842_, new_n20843_, new_n20844_, new_n20845_,
    new_n20846_, new_n20847_, new_n20848_, new_n20849_, new_n20850_,
    new_n20851_, new_n20852_, new_n20853_, new_n20854_, new_n20855_,
    new_n20856_, new_n20857_, new_n20858_, new_n20859_, new_n20860_,
    new_n20861_, new_n20862_, new_n20863_, new_n20864_, new_n20865_,
    new_n20866_, new_n20867_, new_n20868_, new_n20869_, new_n20870_,
    new_n20871_, new_n20872_, new_n20873_, new_n20874_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20889_, new_n20890_, new_n20891_,
    new_n20892_, new_n20893_, new_n20894_, new_n20895_, new_n20896_,
    new_n20897_, new_n20898_, new_n20899_, new_n20900_, new_n20901_,
    new_n20902_, new_n20903_, new_n20904_, new_n20905_, new_n20906_,
    new_n20907_, new_n20908_, new_n20909_, new_n20910_, new_n20911_,
    new_n20912_, new_n20913_, new_n20914_, new_n20915_, new_n20916_,
    new_n20917_, new_n20918_, new_n20919_, new_n20920_, new_n20921_,
    new_n20922_, new_n20923_, new_n20925_, new_n20926_, new_n20927_,
    new_n20928_, new_n20929_, new_n20930_, new_n20931_, new_n20932_,
    new_n20933_, new_n20934_, new_n20935_, new_n20936_, new_n20937_,
    new_n20938_, new_n20939_, new_n20940_, new_n20941_, new_n20942_,
    new_n20943_, new_n20944_, new_n20945_, new_n20946_, new_n20947_,
    new_n20948_, new_n20949_, new_n20950_, new_n20951_, new_n20952_,
    new_n20953_, new_n20954_, new_n20955_, new_n20956_, new_n20957_,
    new_n20959_, new_n20960_, new_n20961_, new_n20962_, new_n20963_,
    new_n20964_, new_n20965_, new_n20966_, new_n20967_, new_n20968_,
    new_n20969_, new_n20970_, new_n20971_, new_n20972_, new_n20973_,
    new_n20974_, new_n20975_, new_n20976_, new_n20977_, new_n20978_,
    new_n20979_, new_n20980_, new_n20981_, new_n20982_, new_n20983_,
    new_n20984_, new_n20985_, new_n20986_, new_n20987_, new_n20988_,
    new_n20990_, new_n20991_, new_n20992_, new_n20993_, new_n20994_,
    new_n20995_, new_n20996_, new_n20997_, new_n20998_, new_n20999_,
    new_n21000_, new_n21001_, new_n21002_, new_n21003_, new_n21004_,
    new_n21005_, new_n21006_, new_n21007_, new_n21008_, new_n21009_,
    new_n21011_, new_n21012_, new_n21013_, new_n21014_, new_n21015_,
    new_n21016_, new_n21017_, new_n21018_, new_n21019_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21029_, new_n21030_, new_n21031_,
    new_n21032_, new_n21033_, new_n21034_, new_n21035_, new_n21036_,
    new_n21037_, new_n21038_, new_n21039_, new_n21040_, new_n21041_,
    new_n21042_, new_n21043_, new_n21044_, new_n21045_, new_n21046_,
    new_n21047_, new_n21048_, new_n21049_, new_n21050_, new_n21051_,
    new_n21052_, new_n21053_;
  INV_X1     g00000(.I(\a[0] ), .ZN(new_n257_));
  INV_X1     g00001(.I(\b[0] ), .ZN(new_n258_));
  NOR2_X1    g00002(.A1(new_n257_), .A2(new_n258_), .ZN(\f[0] ));
  XOR2_X1    g00003(.A1(\b[0] ), .A2(\b[1] ), .Z(new_n260_));
  INV_X1     g00004(.I(new_n260_), .ZN(new_n261_));
  XNOR2_X1   g00005(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n262_));
  NOR2_X1    g00006(.A1(new_n262_), .A2(new_n257_), .ZN(new_n263_));
  INV_X1     g00007(.I(new_n263_), .ZN(new_n264_));
  INV_X1     g00008(.I(\a[1] ), .ZN(new_n265_));
  NOR2_X1    g00009(.A1(new_n265_), .A2(\a[0] ), .ZN(new_n266_));
  INV_X1     g00010(.I(\b[1] ), .ZN(new_n267_));
  NOR2_X1    g00011(.A1(new_n257_), .A2(new_n267_), .ZN(new_n268_));
  AOI22_X1   g00012(.A1(new_n262_), .A2(new_n268_), .B1(\b[0] ), .B2(new_n266_), .ZN(new_n269_));
  OAI21_X1   g00013(.A1(new_n264_), .A2(new_n261_), .B(new_n269_), .ZN(new_n270_));
  INV_X1     g00014(.I(\a[2] ), .ZN(new_n271_));
  INV_X1     g00015(.I(\f[0] ), .ZN(new_n272_));
  NOR2_X1    g00016(.A1(new_n272_), .A2(new_n271_), .ZN(new_n273_));
  XOR2_X1    g00017(.A1(new_n270_), .A2(new_n273_), .Z(\f[1] ));
  NAND3_X1   g00018(.A1(new_n270_), .A2(\a[2] ), .A3(new_n272_), .ZN(new_n275_));
  NAND2_X1   g00019(.A1(new_n258_), .A2(\b[1] ), .ZN(new_n276_));
  NOR2_X1    g00020(.A1(new_n267_), .A2(\b[2] ), .ZN(new_n277_));
  AOI22_X1   g00021(.A1(new_n258_), .A2(new_n277_), .B1(new_n276_), .B2(\b[2] ), .ZN(new_n278_));
  NOR3_X1    g00022(.A1(new_n271_), .A2(\a[0] ), .A3(\a[1] ), .ZN(new_n279_));
  INV_X1     g00023(.I(new_n279_), .ZN(new_n280_));
  OAI22_X1   g00024(.A1(new_n264_), .A2(new_n278_), .B1(new_n258_), .B2(new_n280_), .ZN(new_n281_));
  XOR2_X1    g00025(.A1(\a[1] ), .A2(\a[2] ), .Z(new_n282_));
  NOR2_X1    g00026(.A1(new_n282_), .A2(new_n257_), .ZN(new_n283_));
  AOI22_X1   g00027(.A1(new_n283_), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n266_), .ZN(new_n284_));
  NAND2_X1   g00028(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1    g00029(.A1(new_n285_), .A2(\a[2] ), .Z(new_n286_));
  XNOR2_X1   g00030(.A1(new_n286_), .A2(new_n275_), .ZN(\f[2] ));
  NAND4_X1   g00031(.A1(new_n286_), .A2(\a[2] ), .A3(new_n272_), .A4(new_n270_), .ZN(new_n288_));
  NAND2_X1   g00032(.A1(new_n267_), .A2(\b[3] ), .ZN(new_n289_));
  INV_X1     g00033(.I(\b[3] ), .ZN(new_n290_));
  NAND2_X1   g00034(.A1(new_n290_), .A2(\b[1] ), .ZN(new_n291_));
  INV_X1     g00035(.I(\b[2] ), .ZN(new_n292_));
  OAI21_X1   g00036(.A1(\b[0] ), .A2(new_n267_), .B(new_n292_), .ZN(new_n293_));
  NAND3_X1   g00037(.A1(new_n293_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n294_));
  XOR2_X1    g00038(.A1(\b[1] ), .A2(\b[3] ), .Z(new_n295_));
  AOI21_X1   g00039(.A1(new_n258_), .A2(\b[1] ), .B(\b[2] ), .ZN(new_n296_));
  NAND2_X1   g00040(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1   g00041(.A1(new_n297_), .A2(new_n294_), .ZN(new_n298_));
  AOI21_X1   g00042(.A1(\b[2] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n299_));
  NAND3_X1   g00043(.A1(new_n262_), .A2(\a[0] ), .A3(\b[3] ), .ZN(new_n300_));
  NAND2_X1   g00044(.A1(new_n279_), .A2(\b[1] ), .ZN(new_n301_));
  NAND4_X1   g00045(.A1(new_n299_), .A2(new_n298_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  XOR2_X1    g00046(.A1(new_n302_), .A2(\a[2] ), .Z(new_n303_));
  XNOR2_X1   g00047(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n304_));
  NOR2_X1    g00048(.A1(new_n304_), .A2(new_n258_), .ZN(new_n305_));
  XOR2_X1    g00049(.A1(new_n303_), .A2(new_n305_), .Z(new_n306_));
  XOR2_X1    g00050(.A1(new_n306_), .A2(new_n288_), .Z(\f[3] ));
  INV_X1     g00051(.I(\a[5] ), .ZN(new_n308_));
  NOR2_X1    g00052(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1   g00053(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n310_));
  NOR2_X1    g00054(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1     g00055(.I(new_n311_), .ZN(new_n312_));
  NOR2_X1    g00056(.A1(new_n312_), .A2(new_n261_), .ZN(new_n313_));
  INV_X1     g00057(.I(new_n304_), .ZN(new_n314_));
  NOR2_X1    g00058(.A1(new_n314_), .A2(new_n310_), .ZN(new_n315_));
  INV_X1     g00059(.I(\a[4] ), .ZN(new_n316_));
  NOR3_X1    g00060(.A1(new_n316_), .A2(\a[2] ), .A3(\a[3] ), .ZN(new_n317_));
  NAND3_X1   g00061(.A1(new_n316_), .A2(\a[2] ), .A3(\a[3] ), .ZN(new_n318_));
  INV_X1     g00062(.I(new_n318_), .ZN(new_n319_));
  NOR2_X1    g00063(.A1(new_n319_), .A2(new_n317_), .ZN(new_n320_));
  INV_X1     g00064(.I(new_n320_), .ZN(new_n321_));
  AOI22_X1   g00065(.A1(\b[1] ), .A2(new_n315_), .B1(new_n321_), .B2(\b[0] ), .ZN(new_n322_));
  NOR2_X1    g00066(.A1(new_n322_), .A2(new_n313_), .ZN(new_n323_));
  NOR2_X1    g00067(.A1(new_n323_), .A2(new_n308_), .ZN(new_n324_));
  NOR3_X1    g00068(.A1(new_n322_), .A2(\a[5] ), .A3(new_n313_), .ZN(new_n325_));
  NOR2_X1    g00069(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1   g00070(.A1(\b[1] ), .A2(\b[2] ), .ZN(new_n327_));
  AOI21_X1   g00071(.A1(\b[0] ), .A2(\b[1] ), .B(\b[2] ), .ZN(new_n328_));
  INV_X1     g00072(.I(new_n328_), .ZN(new_n329_));
  OAI21_X1   g00073(.A1(new_n327_), .A2(\b[3] ), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1   g00074(.A1(\b[3] ), .A2(\b[4] ), .ZN(new_n331_));
  XNOR2_X1   g00075(.A1(\b[3] ), .A2(\b[4] ), .ZN(new_n332_));
  NAND2_X1   g00076(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1   g00077(.A1(new_n330_), .A2(new_n331_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1   g00078(.A1(new_n283_), .A2(\b[4] ), .ZN(new_n335_));
  NAND2_X1   g00079(.A1(new_n279_), .A2(\b[2] ), .ZN(new_n336_));
  AOI21_X1   g00080(.A1(\b[3] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n337_));
  NAND4_X1   g00081(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .A4(new_n336_), .ZN(new_n338_));
  XOR2_X1    g00082(.A1(new_n326_), .A2(new_n338_), .Z(new_n339_));
  XOR2_X1    g00083(.A1(new_n339_), .A2(new_n271_), .Z(new_n340_));
  XOR2_X1    g00084(.A1(new_n340_), .A2(new_n309_), .Z(new_n341_));
  NAND2_X1   g00085(.A1(new_n306_), .A2(new_n286_), .ZN(new_n342_));
  NAND2_X1   g00086(.A1(new_n342_), .A2(new_n275_), .ZN(new_n343_));
  NAND2_X1   g00087(.A1(new_n303_), .A2(new_n305_), .ZN(new_n344_));
  XNOR2_X1   g00088(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1    g00089(.A1(new_n345_), .A2(new_n341_), .Z(\f[4] ));
  INV_X1     g00090(.I(\b[5] ), .ZN(new_n347_));
  INV_X1     g00091(.I(new_n331_), .ZN(new_n348_));
  AND2_X2    g00092(.A1(new_n330_), .A2(\b[3] ), .Z(new_n349_));
  NOR2_X1    g00093(.A1(new_n330_), .A2(\b[3] ), .ZN(new_n350_));
  OAI21_X1   g00094(.A1(new_n349_), .A2(new_n350_), .B(new_n348_), .ZN(new_n351_));
  XOR2_X1    g00095(.A1(new_n351_), .A2(new_n347_), .Z(new_n352_));
  AOI21_X1   g00096(.A1(\b[4] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n353_));
  NAND3_X1   g00097(.A1(new_n262_), .A2(\a[0] ), .A3(\b[5] ), .ZN(new_n354_));
  NAND2_X1   g00098(.A1(new_n279_), .A2(\b[3] ), .ZN(new_n355_));
  NAND4_X1   g00099(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  XOR2_X1    g00100(.A1(new_n356_), .A2(\a[2] ), .Z(new_n357_));
  NAND2_X1   g00101(.A1(new_n323_), .A2(new_n309_), .ZN(new_n358_));
  XNOR2_X1   g00102(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n359_));
  XNOR2_X1   g00103(.A1(\a[2] ), .A2(\a[4] ), .ZN(new_n360_));
  NAND2_X1   g00104(.A1(new_n304_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1   g00105(.A1(new_n361_), .A2(new_n359_), .ZN(new_n362_));
  NOR2_X1    g00106(.A1(new_n320_), .A2(new_n267_), .ZN(new_n363_));
  INV_X1     g00107(.I(new_n315_), .ZN(new_n364_));
  NOR2_X1    g00108(.A1(new_n364_), .A2(new_n292_), .ZN(new_n365_));
  NOR4_X1    g00109(.A1(new_n365_), .A2(new_n278_), .A3(new_n312_), .A4(new_n363_), .ZN(new_n366_));
  OAI21_X1   g00110(.A1(new_n258_), .A2(new_n362_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1    g00111(.A1(new_n367_), .A2(new_n358_), .Z(new_n368_));
  XOR2_X1    g00112(.A1(new_n368_), .A2(\a[5] ), .Z(new_n369_));
  XOR2_X1    g00113(.A1(new_n369_), .A2(new_n357_), .Z(new_n370_));
  NAND2_X1   g00114(.A1(new_n345_), .A2(new_n341_), .ZN(new_n371_));
  XNOR2_X1   g00115(.A1(new_n326_), .A2(new_n309_), .ZN(new_n372_));
  XOR2_X1    g00116(.A1(new_n338_), .A2(new_n271_), .Z(new_n373_));
  NOR2_X1    g00117(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1   g00118(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1    g00119(.A1(new_n375_), .A2(new_n370_), .Z(\f[5] ));
  NOR2_X1    g00120(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n377_));
  INV_X1     g00121(.I(\a[6] ), .ZN(new_n378_));
  NOR2_X1    g00122(.A1(new_n308_), .A2(new_n378_), .ZN(new_n379_));
  NOR3_X1    g00123(.A1(new_n379_), .A2(new_n258_), .A3(new_n377_), .ZN(new_n380_));
  INV_X1     g00124(.I(new_n380_), .ZN(new_n381_));
  XOR2_X1    g00125(.A1(new_n367_), .A2(\a[5] ), .Z(new_n382_));
  NOR2_X1    g00126(.A1(new_n382_), .A2(new_n358_), .ZN(new_n383_));
  XOR2_X1    g00127(.A1(new_n383_), .A2(new_n381_), .Z(new_n384_));
  OAI22_X1   g00128(.A1(new_n364_), .A2(new_n290_), .B1(new_n292_), .B2(new_n320_), .ZN(new_n385_));
  OAI21_X1   g00129(.A1(new_n267_), .A2(new_n362_), .B(new_n385_), .ZN(new_n386_));
  NAND3_X1   g00130(.A1(new_n386_), .A2(new_n298_), .A3(new_n311_), .ZN(new_n387_));
  XOR2_X1    g00131(.A1(new_n387_), .A2(\a[5] ), .Z(new_n388_));
  NOR2_X1    g00132(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1     g00133(.I(new_n389_), .ZN(new_n390_));
  NAND2_X1   g00134(.A1(new_n384_), .A2(new_n388_), .ZN(new_n391_));
  NAND2_X1   g00135(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1     g00136(.I(\b[4] ), .ZN(new_n393_));
  OAI21_X1   g00137(.A1(new_n290_), .A2(new_n347_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1   g00138(.A1(new_n330_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1   g00139(.A1(new_n290_), .A2(new_n347_), .B(new_n393_), .ZN(new_n396_));
  INV_X1     g00140(.I(new_n396_), .ZN(new_n397_));
  NAND2_X1   g00141(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  XOR2_X1    g00142(.A1(\b[5] ), .A2(\b[6] ), .Z(new_n399_));
  NAND2_X1   g00143(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1    g00144(.A1(\b[5] ), .A2(\b[6] ), .Z(new_n401_));
  OAI21_X1   g00145(.A1(new_n398_), .A2(new_n401_), .B(new_n400_), .ZN(new_n402_));
  INV_X1     g00146(.I(\b[6] ), .ZN(new_n403_));
  INV_X1     g00147(.I(new_n266_), .ZN(new_n404_));
  INV_X1     g00148(.I(new_n283_), .ZN(new_n405_));
  OAI22_X1   g00149(.A1(new_n405_), .A2(new_n403_), .B1(new_n347_), .B2(new_n404_), .ZN(new_n406_));
  NAND2_X1   g00150(.A1(new_n279_), .A2(\b[4] ), .ZN(new_n407_));
  AOI21_X1   g00151(.A1(new_n406_), .A2(new_n407_), .B(new_n264_), .ZN(new_n408_));
  NAND2_X1   g00152(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1    g00153(.A1(new_n409_), .A2(\a[2] ), .Z(new_n410_));
  INV_X1     g00154(.I(new_n410_), .ZN(new_n411_));
  AND2_X2    g00155(.A1(new_n375_), .A2(new_n370_), .Z(new_n412_));
  XOR2_X1    g00156(.A1(new_n382_), .A2(new_n358_), .Z(new_n413_));
  NAND2_X1   g00157(.A1(new_n413_), .A2(new_n357_), .ZN(new_n414_));
  NAND2_X1   g00158(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1    g00159(.A1(new_n415_), .A2(new_n411_), .Z(new_n416_));
  XOR2_X1    g00160(.A1(new_n416_), .A2(new_n392_), .Z(\f[6] ));
  NAND2_X1   g00161(.A1(new_n392_), .A2(new_n410_), .ZN(new_n418_));
  XOR2_X1    g00162(.A1(new_n392_), .A2(new_n411_), .Z(new_n419_));
  NAND3_X1   g00163(.A1(new_n412_), .A2(new_n419_), .A3(new_n414_), .ZN(new_n420_));
  NAND2_X1   g00164(.A1(new_n420_), .A2(new_n418_), .ZN(new_n421_));
  OAI21_X1   g00165(.A1(new_n383_), .A2(new_n388_), .B(new_n381_), .ZN(new_n422_));
  NOR2_X1    g00166(.A1(new_n330_), .A2(new_n331_), .ZN(new_n423_));
  AOI21_X1   g00167(.A1(new_n330_), .A2(new_n332_), .B(new_n423_), .ZN(new_n424_));
  NOR2_X1    g00168(.A1(new_n362_), .A2(new_n292_), .ZN(new_n425_));
  NOR2_X1    g00169(.A1(new_n320_), .A2(new_n290_), .ZN(new_n426_));
  OAI21_X1   g00170(.A1(new_n364_), .A2(new_n393_), .B(new_n311_), .ZN(new_n427_));
  NOR4_X1    g00171(.A1(new_n427_), .A2(new_n424_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n428_));
  INV_X1     g00172(.I(\a[8] ), .ZN(new_n429_));
  NOR3_X1    g00173(.A1(new_n308_), .A2(new_n378_), .A3(\a[7] ), .ZN(new_n430_));
  AOI21_X1   g00174(.A1(\a[7] ), .A2(new_n377_), .B(new_n430_), .ZN(new_n431_));
  NOR2_X1    g00175(.A1(new_n431_), .A2(new_n258_), .ZN(new_n432_));
  XNOR2_X1   g00176(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n433_));
  INV_X1     g00177(.I(new_n433_), .ZN(new_n434_));
  XNOR2_X1   g00178(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n435_));
  NOR2_X1    g00179(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1     g00180(.I(new_n436_), .ZN(new_n437_));
  NOR2_X1    g00181(.A1(new_n437_), .A2(new_n267_), .ZN(new_n438_));
  NOR2_X1    g00182(.A1(new_n433_), .A2(new_n435_), .ZN(new_n439_));
  INV_X1     g00183(.I(new_n439_), .ZN(new_n440_));
  NOR4_X1    g00184(.A1(new_n438_), .A2(new_n261_), .A3(new_n432_), .A4(new_n440_), .ZN(new_n441_));
  XOR2_X1    g00185(.A1(new_n441_), .A2(\a[8] ), .Z(new_n442_));
  OAI21_X1   g00186(.A1(new_n429_), .A2(new_n380_), .B(new_n442_), .ZN(new_n443_));
  NOR3_X1    g00187(.A1(new_n442_), .A2(new_n429_), .A3(new_n380_), .ZN(new_n444_));
  INV_X1     g00188(.I(new_n444_), .ZN(new_n445_));
  NAND2_X1   g00189(.A1(new_n445_), .A2(new_n443_), .ZN(new_n446_));
  XOR2_X1    g00190(.A1(new_n446_), .A2(new_n308_), .Z(new_n447_));
  XOR2_X1    g00191(.A1(new_n447_), .A2(new_n428_), .Z(new_n448_));
  XOR2_X1    g00192(.A1(new_n448_), .A2(new_n422_), .Z(new_n449_));
  INV_X1     g00193(.I(\b[7] ), .ZN(new_n450_));
  AOI21_X1   g00194(.A1(new_n330_), .A2(new_n394_), .B(new_n396_), .ZN(new_n451_));
  XOR2_X1    g00195(.A1(new_n451_), .A2(new_n347_), .Z(new_n452_));
  NAND2_X1   g00196(.A1(new_n452_), .A2(new_n399_), .ZN(new_n453_));
  XOR2_X1    g00197(.A1(new_n453_), .A2(new_n450_), .Z(new_n454_));
  OAI22_X1   g00198(.A1(new_n405_), .A2(new_n450_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n455_));
  NAND2_X1   g00199(.A1(new_n279_), .A2(\b[5] ), .ZN(new_n456_));
  AOI21_X1   g00200(.A1(new_n455_), .A2(new_n456_), .B(new_n264_), .ZN(new_n457_));
  NAND2_X1   g00201(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1    g00202(.A1(new_n458_), .A2(\a[2] ), .Z(new_n459_));
  INV_X1     g00203(.I(new_n459_), .ZN(new_n460_));
  XOR2_X1    g00204(.A1(new_n449_), .A2(new_n460_), .Z(new_n461_));
  NAND2_X1   g00205(.A1(new_n449_), .A2(new_n460_), .ZN(new_n462_));
  NOR2_X1    g00206(.A1(new_n449_), .A2(new_n460_), .ZN(new_n463_));
  INV_X1     g00207(.I(new_n463_), .ZN(new_n464_));
  NAND2_X1   g00208(.A1(new_n464_), .A2(new_n462_), .ZN(new_n465_));
  MUX2_X1    g00209(.I0(new_n465_), .I1(new_n461_), .S(new_n421_), .Z(\f[7] ));
  OAI22_X1   g00210(.A1(new_n364_), .A2(new_n347_), .B1(new_n393_), .B2(new_n320_), .ZN(new_n467_));
  OAI21_X1   g00211(.A1(new_n290_), .A2(new_n362_), .B(new_n467_), .ZN(new_n468_));
  AOI21_X1   g00212(.A1(new_n352_), .A2(new_n311_), .B(new_n468_), .ZN(new_n469_));
  NOR2_X1    g00213(.A1(new_n440_), .A2(new_n278_), .ZN(new_n470_));
  XNOR2_X1   g00214(.A1(\a[5] ), .A2(\a[7] ), .ZN(new_n471_));
  NAND2_X1   g00215(.A1(new_n433_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1   g00216(.A1(\a[5] ), .A2(\a[8] ), .ZN(new_n473_));
  NAND2_X1   g00217(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI22_X1   g00218(.A1(new_n437_), .A2(new_n292_), .B1(new_n267_), .B2(new_n431_), .ZN(new_n475_));
  NOR4_X1    g00219(.A1(new_n475_), .A2(new_n258_), .A3(new_n470_), .A4(new_n474_), .ZN(new_n476_));
  XOR2_X1    g00220(.A1(new_n476_), .A2(new_n429_), .Z(new_n477_));
  INV_X1     g00221(.I(new_n477_), .ZN(new_n478_));
  NAND2_X1   g00222(.A1(new_n445_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1    g00223(.A1(new_n445_), .A2(new_n478_), .ZN(new_n480_));
  INV_X1     g00224(.I(new_n480_), .ZN(new_n481_));
  NAND2_X1   g00225(.A1(new_n481_), .A2(new_n479_), .ZN(new_n482_));
  XOR2_X1    g00226(.A1(new_n482_), .A2(new_n308_), .Z(new_n483_));
  XOR2_X1    g00227(.A1(new_n483_), .A2(new_n469_), .Z(new_n484_));
  AOI21_X1   g00228(.A1(\b[5] ), .A2(\b[7] ), .B(\b[6] ), .ZN(new_n485_));
  NOR2_X1    g00229(.A1(new_n398_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1   g00230(.A1(new_n347_), .A2(new_n450_), .B(new_n403_), .ZN(new_n487_));
  NOR2_X1    g00231(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1   g00232(.A1(\b[7] ), .A2(\b[8] ), .ZN(new_n489_));
  NOR2_X1    g00233(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X2     g00234(.A1(new_n486_), .A2(new_n487_), .Z(new_n491_));
  XOR2_X1    g00235(.A1(\b[7] ), .A2(\b[8] ), .Z(new_n492_));
  NOR2_X1    g00236(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OR2_X2     g00237(.A1(new_n493_), .A2(new_n490_), .Z(new_n494_));
  INV_X1     g00238(.I(\b[8] ), .ZN(new_n495_));
  OAI22_X1   g00239(.A1(new_n405_), .A2(new_n495_), .B1(new_n450_), .B2(new_n404_), .ZN(new_n496_));
  NAND2_X1   g00240(.A1(new_n279_), .A2(\b[6] ), .ZN(new_n497_));
  AOI21_X1   g00241(.A1(new_n496_), .A2(new_n497_), .B(new_n264_), .ZN(new_n498_));
  NAND2_X1   g00242(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1    g00243(.A1(new_n499_), .A2(\a[2] ), .Z(new_n500_));
  NAND2_X1   g00244(.A1(new_n448_), .A2(new_n390_), .ZN(new_n501_));
  NOR2_X1    g00245(.A1(new_n383_), .A2(new_n380_), .ZN(new_n502_));
  NAND2_X1   g00246(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1    g00247(.A1(new_n428_), .A2(new_n308_), .Z(new_n504_));
  NAND4_X1   g00248(.A1(new_n503_), .A2(new_n443_), .A3(new_n445_), .A4(new_n504_), .ZN(new_n505_));
  XNOR2_X1   g00249(.A1(new_n505_), .A2(new_n500_), .ZN(new_n506_));
  XOR2_X1    g00250(.A1(new_n506_), .A2(new_n484_), .Z(new_n507_));
  OAI21_X1   g00251(.A1(new_n421_), .A2(new_n449_), .B(new_n460_), .ZN(new_n508_));
  XOR2_X1    g00252(.A1(new_n507_), .A2(new_n508_), .Z(\f[8] ));
  INV_X1     g00253(.I(\b[9] ), .ZN(new_n510_));
  INV_X1     g00254(.I(new_n489_), .ZN(new_n511_));
  XOR2_X1    g00255(.A1(new_n488_), .A2(new_n450_), .Z(new_n512_));
  NAND3_X1   g00256(.A1(new_n512_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n513_));
  NOR2_X1    g00257(.A1(new_n491_), .A2(new_n450_), .ZN(new_n514_));
  NOR2_X1    g00258(.A1(new_n488_), .A2(\b[7] ), .ZN(new_n515_));
  OAI21_X1   g00259(.A1(new_n514_), .A2(new_n515_), .B(new_n511_), .ZN(new_n516_));
  NAND2_X1   g00260(.A1(new_n516_), .A2(\b[9] ), .ZN(new_n517_));
  NAND2_X1   g00261(.A1(new_n517_), .A2(new_n513_), .ZN(new_n518_));
  NOR2_X1    g00262(.A1(new_n405_), .A2(new_n510_), .ZN(new_n519_));
  NOR2_X1    g00263(.A1(new_n280_), .A2(new_n450_), .ZN(new_n520_));
  NOR2_X1    g00264(.A1(new_n404_), .A2(new_n495_), .ZN(new_n521_));
  NOR4_X1    g00265(.A1(new_n519_), .A2(new_n264_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  NAND2_X1   g00266(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1     g00267(.I(new_n402_), .ZN(new_n524_));
  AOI22_X1   g00268(.A1(\b[6] ), .A2(new_n315_), .B1(new_n321_), .B2(\b[5] ), .ZN(new_n525_));
  NOR2_X1    g00269(.A1(new_n362_), .A2(new_n393_), .ZN(new_n526_));
  OAI21_X1   g00270(.A1(new_n525_), .A2(new_n526_), .B(new_n311_), .ZN(new_n527_));
  NOR2_X1    g00271(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1    g00272(.A1(new_n528_), .A2(new_n308_), .Z(new_n529_));
  XNOR2_X1   g00273(.A1(\a[8] ), .A2(\a[9] ), .ZN(new_n530_));
  NOR2_X1    g00274(.A1(new_n530_), .A2(new_n258_), .ZN(new_n531_));
  OAI22_X1   g00275(.A1(new_n437_), .A2(new_n290_), .B1(new_n292_), .B2(new_n431_), .ZN(new_n532_));
  OAI21_X1   g00276(.A1(new_n267_), .A2(new_n474_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1   g00277(.A1(new_n533_), .A2(new_n298_), .A3(new_n439_), .ZN(new_n534_));
  NOR2_X1    g00278(.A1(new_n534_), .A2(\a[8] ), .ZN(new_n535_));
  NAND2_X1   g00279(.A1(new_n534_), .A2(\a[8] ), .ZN(new_n536_));
  INV_X1     g00280(.I(new_n536_), .ZN(new_n537_));
  NOR2_X1    g00281(.A1(new_n537_), .A2(new_n535_), .ZN(new_n538_));
  INV_X1     g00282(.I(new_n538_), .ZN(new_n539_));
  XOR2_X1    g00283(.A1(new_n480_), .A2(new_n539_), .Z(new_n540_));
  XOR2_X1    g00284(.A1(new_n540_), .A2(new_n531_), .Z(new_n541_));
  XOR2_X1    g00285(.A1(new_n541_), .A2(new_n529_), .Z(new_n542_));
  XOR2_X1    g00286(.A1(new_n542_), .A2(\a[2] ), .Z(new_n543_));
  XNOR2_X1   g00287(.A1(new_n543_), .A2(new_n523_), .ZN(new_n544_));
  NAND3_X1   g00288(.A1(new_n420_), .A2(new_n463_), .A3(new_n418_), .ZN(new_n545_));
  NAND3_X1   g00289(.A1(new_n507_), .A2(new_n464_), .A3(new_n545_), .ZN(new_n546_));
  OR2_X2     g00290(.A1(new_n505_), .A2(new_n484_), .Z(new_n547_));
  NAND2_X1   g00291(.A1(new_n505_), .A2(new_n484_), .ZN(new_n548_));
  NAND3_X1   g00292(.A1(new_n547_), .A2(new_n500_), .A3(new_n548_), .ZN(new_n549_));
  NOR2_X1    g00293(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1   g00294(.A1(new_n544_), .A2(new_n500_), .A3(new_n547_), .A4(new_n548_), .ZN(new_n551_));
  OAI22_X1   g00295(.A1(new_n550_), .A2(new_n544_), .B1(new_n546_), .B2(new_n551_), .ZN(\f[9] ));
  INV_X1     g00296(.I(new_n542_), .ZN(new_n553_));
  XOR2_X1    g00297(.A1(new_n523_), .A2(\a[2] ), .Z(new_n554_));
  NOR2_X1    g00298(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1     g00299(.I(new_n555_), .ZN(new_n556_));
  OAI21_X1   g00300(.A1(new_n546_), .A2(new_n549_), .B(new_n544_), .ZN(new_n557_));
  AND2_X2    g00301(.A1(new_n557_), .A2(new_n556_), .Z(new_n558_));
  XOR2_X1    g00302(.A1(new_n538_), .A2(new_n531_), .Z(new_n559_));
  AOI21_X1   g00303(.A1(new_n559_), .A2(new_n477_), .B(new_n444_), .ZN(new_n560_));
  INV_X1     g00304(.I(new_n531_), .ZN(new_n561_));
  NOR2_X1    g00305(.A1(new_n539_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1     g00306(.I(new_n562_), .ZN(new_n563_));
  NOR2_X1    g00307(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1   g00308(.A1(new_n560_), .A2(new_n563_), .ZN(new_n565_));
  INV_X1     g00309(.I(new_n565_), .ZN(new_n566_));
  NOR2_X1    g00310(.A1(new_n566_), .A2(new_n564_), .ZN(new_n567_));
  INV_X1     g00311(.I(new_n567_), .ZN(new_n568_));
  OAI22_X1   g00312(.A1(new_n437_), .A2(new_n393_), .B1(new_n290_), .B2(new_n431_), .ZN(new_n569_));
  OAI21_X1   g00313(.A1(new_n292_), .A2(new_n474_), .B(new_n569_), .ZN(new_n570_));
  AOI21_X1   g00314(.A1(new_n334_), .A2(new_n439_), .B(new_n570_), .ZN(new_n571_));
  INV_X1     g00315(.I(\a[11] ), .ZN(new_n572_));
  INV_X1     g00316(.I(\a[10] ), .ZN(new_n573_));
  NOR3_X1    g00317(.A1(new_n573_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n574_));
  NAND3_X1   g00318(.A1(new_n573_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n575_));
  INV_X1     g00319(.I(new_n575_), .ZN(new_n576_));
  NOR2_X1    g00320(.A1(new_n576_), .A2(new_n574_), .ZN(new_n577_));
  NOR2_X1    g00321(.A1(new_n577_), .A2(new_n258_), .ZN(new_n578_));
  INV_X1     g00322(.I(new_n530_), .ZN(new_n579_));
  XNOR2_X1   g00323(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n580_));
  NOR2_X1    g00324(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1     g00325(.I(new_n581_), .ZN(new_n582_));
  NOR2_X1    g00326(.A1(new_n582_), .A2(new_n267_), .ZN(new_n583_));
  NOR2_X1    g00327(.A1(new_n530_), .A2(new_n580_), .ZN(new_n584_));
  INV_X1     g00328(.I(new_n584_), .ZN(new_n585_));
  NOR4_X1    g00329(.A1(new_n583_), .A2(new_n261_), .A3(new_n578_), .A4(new_n585_), .ZN(new_n586_));
  XOR2_X1    g00330(.A1(new_n586_), .A2(new_n572_), .Z(new_n587_));
  NOR2_X1    g00331(.A1(new_n531_), .A2(new_n572_), .ZN(new_n588_));
  XNOR2_X1   g00332(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1    g00333(.A1(new_n589_), .A2(\a[8] ), .Z(new_n590_));
  XOR2_X1    g00334(.A1(new_n589_), .A2(new_n429_), .Z(new_n591_));
  MUX2_X1    g00335(.I0(new_n591_), .I1(new_n590_), .S(new_n571_), .Z(new_n592_));
  OAI22_X1   g00336(.A1(new_n364_), .A2(new_n450_), .B1(new_n403_), .B2(new_n320_), .ZN(new_n593_));
  INV_X1     g00337(.I(new_n362_), .ZN(new_n594_));
  NAND2_X1   g00338(.A1(new_n594_), .A2(\b[5] ), .ZN(new_n595_));
  AOI21_X1   g00339(.A1(new_n593_), .A2(new_n595_), .B(new_n312_), .ZN(new_n596_));
  NAND2_X1   g00340(.A1(new_n454_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1    g00341(.A1(new_n597_), .A2(\a[5] ), .Z(new_n598_));
  XOR2_X1    g00342(.A1(new_n592_), .A2(new_n598_), .Z(new_n599_));
  NAND2_X1   g00343(.A1(new_n599_), .A2(new_n568_), .ZN(new_n600_));
  XOR2_X1    g00344(.A1(new_n592_), .A2(new_n598_), .Z(new_n601_));
  OAI21_X1   g00345(.A1(new_n568_), .A2(new_n601_), .B(new_n600_), .ZN(new_n602_));
  OR2_X2     g00346(.A1(new_n559_), .A2(new_n481_), .Z(new_n603_));
  XOR2_X1    g00347(.A1(new_n538_), .A2(new_n531_), .Z(new_n604_));
  NAND2_X1   g00348(.A1(new_n604_), .A2(new_n481_), .ZN(new_n605_));
  NAND3_X1   g00349(.A1(new_n603_), .A2(new_n529_), .A3(new_n605_), .ZN(new_n606_));
  XOR2_X1    g00350(.A1(new_n602_), .A2(new_n606_), .Z(new_n607_));
  AOI21_X1   g00351(.A1(\b[7] ), .A2(\b[9] ), .B(\b[8] ), .ZN(new_n608_));
  AOI21_X1   g00352(.A1(new_n450_), .A2(new_n510_), .B(new_n495_), .ZN(new_n609_));
  INV_X1     g00353(.I(new_n609_), .ZN(new_n610_));
  OAI21_X1   g00354(.A1(new_n491_), .A2(new_n608_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1   g00355(.A1(\b[9] ), .A2(\b[10] ), .ZN(new_n612_));
  INV_X1     g00356(.I(new_n612_), .ZN(new_n613_));
  NAND2_X1   g00357(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1    g00358(.A1(\b[9] ), .A2(\b[10] ), .Z(new_n615_));
  OAI21_X1   g00359(.A1(new_n611_), .A2(new_n615_), .B(new_n614_), .ZN(new_n616_));
  INV_X1     g00360(.I(\b[10] ), .ZN(new_n617_));
  OAI22_X1   g00361(.A1(new_n405_), .A2(new_n617_), .B1(new_n510_), .B2(new_n404_), .ZN(new_n618_));
  NAND2_X1   g00362(.A1(new_n279_), .A2(\b[8] ), .ZN(new_n619_));
  AOI21_X1   g00363(.A1(new_n618_), .A2(new_n619_), .B(new_n264_), .ZN(new_n620_));
  NAND2_X1   g00364(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  XOR2_X1    g00365(.A1(new_n621_), .A2(\a[2] ), .Z(new_n622_));
  INV_X1     g00366(.I(new_n622_), .ZN(new_n623_));
  XOR2_X1    g00367(.A1(new_n607_), .A2(new_n623_), .Z(new_n624_));
  XOR2_X1    g00368(.A1(new_n607_), .A2(new_n623_), .Z(new_n625_));
  NAND2_X1   g00369(.A1(new_n558_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1   g00370(.A1(new_n558_), .A2(new_n624_), .B(new_n626_), .ZN(\f[10] ));
  OAI22_X1   g00371(.A1(new_n437_), .A2(new_n347_), .B1(new_n393_), .B2(new_n431_), .ZN(new_n628_));
  OAI21_X1   g00372(.A1(new_n290_), .A2(new_n474_), .B(new_n628_), .ZN(new_n629_));
  AOI21_X1   g00373(.A1(new_n352_), .A2(new_n439_), .B(new_n629_), .ZN(new_n630_));
  NOR2_X1    g00374(.A1(new_n585_), .A2(new_n278_), .ZN(new_n631_));
  XNOR2_X1   g00375(.A1(\a[8] ), .A2(\a[10] ), .ZN(new_n632_));
  NAND2_X1   g00376(.A1(new_n530_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1   g00377(.A1(\a[8] ), .A2(\a[11] ), .ZN(new_n634_));
  NAND2_X1   g00378(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI22_X1   g00379(.A1(new_n582_), .A2(new_n292_), .B1(new_n267_), .B2(new_n577_), .ZN(new_n636_));
  NOR4_X1    g00380(.A1(new_n636_), .A2(new_n258_), .A3(new_n631_), .A4(new_n635_), .ZN(new_n637_));
  XOR2_X1    g00381(.A1(new_n637_), .A2(new_n572_), .Z(new_n638_));
  AOI21_X1   g00382(.A1(new_n587_), .A2(new_n588_), .B(new_n638_), .ZN(new_n639_));
  NAND2_X1   g00383(.A1(new_n587_), .A2(new_n588_), .ZN(new_n640_));
  INV_X1     g00384(.I(new_n638_), .ZN(new_n641_));
  NOR2_X1    g00385(.A1(new_n641_), .A2(new_n640_), .ZN(new_n642_));
  NOR2_X1    g00386(.A1(new_n642_), .A2(new_n639_), .ZN(new_n643_));
  XOR2_X1    g00387(.A1(new_n643_), .A2(\a[8] ), .Z(new_n644_));
  XOR2_X1    g00388(.A1(new_n644_), .A2(new_n630_), .Z(new_n645_));
  INV_X1     g00389(.I(new_n645_), .ZN(new_n646_));
  XOR2_X1    g00390(.A1(new_n571_), .A2(new_n429_), .Z(new_n647_));
  XOR2_X1    g00391(.A1(new_n567_), .A2(new_n647_), .Z(new_n648_));
  NAND2_X1   g00392(.A1(new_n648_), .A2(new_n589_), .ZN(new_n649_));
  XOR2_X1    g00393(.A1(new_n649_), .A2(new_n646_), .Z(new_n650_));
  NOR2_X1    g00394(.A1(new_n567_), .A2(new_n647_), .ZN(new_n651_));
  XOR2_X1    g00395(.A1(new_n650_), .A2(new_n651_), .Z(new_n652_));
  OAI22_X1   g00396(.A1(new_n364_), .A2(new_n495_), .B1(new_n450_), .B2(new_n320_), .ZN(new_n653_));
  NAND2_X1   g00397(.A1(new_n594_), .A2(\b[6] ), .ZN(new_n654_));
  AOI21_X1   g00398(.A1(new_n653_), .A2(new_n654_), .B(new_n312_), .ZN(new_n655_));
  NAND2_X1   g00399(.A1(new_n494_), .A2(new_n655_), .ZN(new_n656_));
  XOR2_X1    g00400(.A1(new_n656_), .A2(new_n308_), .Z(new_n657_));
  XOR2_X1    g00401(.A1(new_n652_), .A2(new_n657_), .Z(new_n658_));
  INV_X1     g00402(.I(\b[11] ), .ZN(new_n659_));
  XOR2_X1    g00403(.A1(new_n611_), .A2(\b[9] ), .Z(new_n660_));
  AND3_X2    g00404(.A1(new_n660_), .A2(new_n659_), .A3(new_n613_), .Z(new_n661_));
  AOI21_X1   g00405(.A1(new_n660_), .A2(new_n613_), .B(new_n659_), .ZN(new_n662_));
  OR2_X2     g00406(.A1(new_n661_), .A2(new_n662_), .Z(new_n663_));
  OAI22_X1   g00407(.A1(new_n405_), .A2(new_n659_), .B1(new_n617_), .B2(new_n404_), .ZN(new_n664_));
  NAND2_X1   g00408(.A1(new_n279_), .A2(\b[9] ), .ZN(new_n665_));
  AOI21_X1   g00409(.A1(new_n664_), .A2(new_n665_), .B(new_n264_), .ZN(new_n666_));
  NAND2_X1   g00410(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  XOR2_X1    g00411(.A1(new_n667_), .A2(\a[2] ), .Z(new_n668_));
  XNOR2_X1   g00412(.A1(new_n567_), .A2(new_n592_), .ZN(new_n669_));
  NAND2_X1   g00413(.A1(new_n669_), .A2(new_n598_), .ZN(new_n670_));
  NAND2_X1   g00414(.A1(new_n670_), .A2(new_n529_), .ZN(new_n671_));
  NOR2_X1    g00415(.A1(new_n671_), .A2(new_n602_), .ZN(new_n672_));
  XOR2_X1    g00416(.A1(new_n672_), .A2(new_n668_), .Z(new_n673_));
  XOR2_X1    g00417(.A1(new_n658_), .A2(new_n673_), .Z(new_n674_));
  AOI21_X1   g00418(.A1(new_n558_), .A2(new_n607_), .B(new_n622_), .ZN(new_n675_));
  XNOR2_X1   g00419(.A1(new_n674_), .A2(new_n675_), .ZN(\f[11] ));
  INV_X1     g00420(.I(new_n298_), .ZN(new_n677_));
  NOR2_X1    g00421(.A1(new_n635_), .A2(new_n267_), .ZN(new_n678_));
  OAI22_X1   g00422(.A1(new_n582_), .A2(new_n290_), .B1(new_n292_), .B2(new_n577_), .ZN(new_n679_));
  NOR4_X1    g00423(.A1(new_n679_), .A2(new_n677_), .A3(new_n585_), .A4(new_n678_), .ZN(new_n680_));
  XOR2_X1    g00424(.A1(new_n680_), .A2(new_n572_), .Z(new_n681_));
  XNOR2_X1   g00425(.A1(\a[11] ), .A2(\a[12] ), .ZN(new_n682_));
  NOR2_X1    g00426(.A1(new_n682_), .A2(new_n258_), .ZN(new_n683_));
  XOR2_X1    g00427(.A1(new_n681_), .A2(new_n683_), .Z(new_n684_));
  XOR2_X1    g00428(.A1(new_n684_), .A2(new_n642_), .Z(new_n685_));
  INV_X1     g00429(.I(new_n431_), .ZN(new_n686_));
  AOI22_X1   g00430(.A1(new_n436_), .A2(\b[6] ), .B1(new_n686_), .B2(\b[5] ), .ZN(new_n687_));
  NOR2_X1    g00431(.A1(new_n474_), .A2(new_n393_), .ZN(new_n688_));
  OAI21_X1   g00432(.A1(new_n687_), .A2(new_n688_), .B(new_n439_), .ZN(new_n689_));
  NOR2_X1    g00433(.A1(new_n524_), .A2(new_n689_), .ZN(new_n690_));
  XOR2_X1    g00434(.A1(new_n690_), .A2(\a[8] ), .Z(new_n691_));
  INV_X1     g00435(.I(new_n647_), .ZN(new_n692_));
  NOR2_X1    g00436(.A1(new_n692_), .A2(new_n589_), .ZN(new_n693_));
  INV_X1     g00437(.I(new_n693_), .ZN(new_n694_));
  NOR2_X1    g00438(.A1(new_n568_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1   g00439(.A1(new_n630_), .A2(new_n429_), .ZN(new_n696_));
  OR2_X2     g00440(.A1(new_n630_), .A2(new_n429_), .Z(new_n697_));
  NAND4_X1   g00441(.A1(new_n694_), .A2(new_n697_), .A3(new_n696_), .A4(new_n643_), .ZN(new_n698_));
  NOR3_X1    g00442(.A1(new_n695_), .A2(new_n646_), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1    g00443(.A1(new_n699_), .A2(new_n691_), .Z(new_n700_));
  XNOR2_X1   g00444(.A1(new_n700_), .A2(new_n685_), .ZN(new_n701_));
  OAI22_X1   g00445(.A1(new_n364_), .A2(new_n510_), .B1(new_n495_), .B2(new_n320_), .ZN(new_n702_));
  NAND2_X1   g00446(.A1(new_n594_), .A2(\b[7] ), .ZN(new_n703_));
  AOI21_X1   g00447(.A1(new_n702_), .A2(new_n703_), .B(new_n312_), .ZN(new_n704_));
  NAND2_X1   g00448(.A1(new_n518_), .A2(new_n704_), .ZN(new_n705_));
  XOR2_X1    g00449(.A1(new_n705_), .A2(\a[5] ), .Z(new_n706_));
  XOR2_X1    g00450(.A1(new_n701_), .A2(new_n706_), .Z(new_n707_));
  AOI21_X1   g00451(.A1(\b[9] ), .A2(\b[11] ), .B(\b[10] ), .ZN(new_n708_));
  NOR2_X1    g00452(.A1(new_n611_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1   g00453(.A1(new_n510_), .A2(new_n659_), .B(new_n617_), .ZN(new_n710_));
  OR2_X2     g00454(.A1(new_n709_), .A2(new_n710_), .Z(new_n711_));
  XNOR2_X1   g00455(.A1(\b[11] ), .A2(\b[12] ), .ZN(new_n712_));
  INV_X1     g00456(.I(new_n712_), .ZN(new_n713_));
  NAND2_X1   g00457(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1    g00458(.A1(\b[11] ), .A2(\b[12] ), .Z(new_n715_));
  OAI21_X1   g00459(.A1(new_n711_), .A2(new_n715_), .B(new_n714_), .ZN(new_n716_));
  INV_X1     g00460(.I(\b[12] ), .ZN(new_n717_));
  OAI22_X1   g00461(.A1(new_n405_), .A2(new_n717_), .B1(new_n659_), .B2(new_n404_), .ZN(new_n718_));
  NAND2_X1   g00462(.A1(new_n279_), .A2(\b[10] ), .ZN(new_n719_));
  AOI21_X1   g00463(.A1(new_n718_), .A2(new_n719_), .B(new_n264_), .ZN(new_n720_));
  NAND2_X1   g00464(.A1(new_n716_), .A2(new_n720_), .ZN(new_n721_));
  XOR2_X1    g00465(.A1(new_n721_), .A2(\a[2] ), .Z(new_n722_));
  INV_X1     g00466(.I(new_n672_), .ZN(new_n723_));
  NOR2_X1    g00467(.A1(new_n658_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1   g00468(.A1(new_n607_), .A2(new_n622_), .ZN(new_n725_));
  NAND2_X1   g00469(.A1(new_n658_), .A2(new_n723_), .ZN(new_n726_));
  NAND3_X1   g00470(.A1(new_n726_), .A2(new_n725_), .A3(new_n668_), .ZN(new_n727_));
  INV_X1     g00471(.I(new_n558_), .ZN(new_n728_));
  OAI21_X1   g00472(.A1(new_n728_), .A2(new_n725_), .B(new_n674_), .ZN(new_n729_));
  NOR3_X1    g00473(.A1(new_n729_), .A2(new_n724_), .A3(new_n727_), .ZN(new_n730_));
  XOR2_X1    g00474(.A1(new_n730_), .A2(new_n722_), .Z(new_n731_));
  XOR2_X1    g00475(.A1(new_n731_), .A2(new_n707_), .Z(\f[12] ));
  INV_X1     g00476(.I(new_n701_), .ZN(new_n733_));
  NOR2_X1    g00477(.A1(new_n733_), .A2(new_n706_), .ZN(new_n734_));
  NAND2_X1   g00478(.A1(new_n684_), .A2(new_n638_), .ZN(new_n735_));
  NAND2_X1   g00479(.A1(new_n735_), .A2(new_n640_), .ZN(new_n736_));
  INV_X1     g00480(.I(new_n736_), .ZN(new_n737_));
  NAND2_X1   g00481(.A1(new_n681_), .A2(new_n683_), .ZN(new_n738_));
  NOR2_X1    g00482(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1   g00483(.A1(new_n737_), .A2(new_n738_), .ZN(new_n740_));
  INV_X1     g00484(.I(new_n740_), .ZN(new_n741_));
  NOR2_X1    g00485(.A1(new_n741_), .A2(new_n739_), .ZN(new_n742_));
  OAI22_X1   g00486(.A1(new_n582_), .A2(new_n393_), .B1(new_n290_), .B2(new_n577_), .ZN(new_n743_));
  OAI21_X1   g00487(.A1(new_n292_), .A2(new_n635_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1   g00488(.A1(new_n744_), .A2(new_n334_), .A3(new_n584_), .ZN(new_n745_));
  XOR2_X1    g00489(.A1(new_n745_), .A2(\a[11] ), .Z(new_n746_));
  INV_X1     g00490(.I(\a[14] ), .ZN(new_n747_));
  INV_X1     g00491(.I(\a[13] ), .ZN(new_n748_));
  NOR3_X1    g00492(.A1(new_n748_), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n749_));
  NAND3_X1   g00493(.A1(new_n748_), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n750_));
  INV_X1     g00494(.I(new_n750_), .ZN(new_n751_));
  NOR2_X1    g00495(.A1(new_n751_), .A2(new_n749_), .ZN(new_n752_));
  NOR2_X1    g00496(.A1(new_n752_), .A2(new_n258_), .ZN(new_n753_));
  INV_X1     g00497(.I(new_n682_), .ZN(new_n754_));
  XNOR2_X1   g00498(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n755_));
  NOR2_X1    g00499(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1     g00500(.I(new_n756_), .ZN(new_n757_));
  NOR2_X1    g00501(.A1(new_n757_), .A2(new_n267_), .ZN(new_n758_));
  NOR2_X1    g00502(.A1(new_n682_), .A2(new_n755_), .ZN(new_n759_));
  INV_X1     g00503(.I(new_n759_), .ZN(new_n760_));
  NOR4_X1    g00504(.A1(new_n758_), .A2(new_n261_), .A3(new_n753_), .A4(new_n760_), .ZN(new_n761_));
  XOR2_X1    g00505(.A1(new_n761_), .A2(new_n747_), .Z(new_n762_));
  NOR2_X1    g00506(.A1(new_n683_), .A2(new_n747_), .ZN(new_n763_));
  XNOR2_X1   g00507(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  XOR2_X1    g00508(.A1(new_n764_), .A2(new_n746_), .Z(new_n765_));
  NOR2_X1    g00509(.A1(new_n742_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1     g00510(.I(new_n746_), .ZN(new_n767_));
  NOR2_X1    g00511(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1     g00512(.I(new_n768_), .ZN(new_n769_));
  NAND2_X1   g00513(.A1(new_n764_), .A2(new_n767_), .ZN(new_n770_));
  NAND2_X1   g00514(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1   g00515(.A1(new_n742_), .A2(new_n771_), .B(new_n766_), .ZN(new_n772_));
  INV_X1     g00516(.I(new_n772_), .ZN(new_n773_));
  OAI22_X1   g00517(.A1(new_n437_), .A2(new_n450_), .B1(new_n403_), .B2(new_n431_), .ZN(new_n774_));
  INV_X1     g00518(.I(new_n474_), .ZN(new_n775_));
  NAND2_X1   g00519(.A1(new_n775_), .A2(\b[5] ), .ZN(new_n776_));
  AOI21_X1   g00520(.A1(new_n774_), .A2(new_n776_), .B(new_n440_), .ZN(new_n777_));
  NAND2_X1   g00521(.A1(new_n454_), .A2(new_n777_), .ZN(new_n778_));
  XOR2_X1    g00522(.A1(new_n778_), .A2(\a[8] ), .Z(new_n779_));
  NOR2_X1    g00523(.A1(new_n773_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1   g00524(.A1(new_n773_), .A2(new_n779_), .ZN(new_n781_));
  INV_X1     g00525(.I(new_n781_), .ZN(new_n782_));
  OAI22_X1   g00526(.A1(new_n364_), .A2(new_n617_), .B1(new_n510_), .B2(new_n320_), .ZN(new_n783_));
  NAND2_X1   g00527(.A1(new_n594_), .A2(\b[8] ), .ZN(new_n784_));
  AOI21_X1   g00528(.A1(new_n783_), .A2(new_n784_), .B(new_n312_), .ZN(new_n785_));
  NAND2_X1   g00529(.A1(new_n616_), .A2(new_n785_), .ZN(new_n786_));
  XOR2_X1    g00530(.A1(new_n786_), .A2(\a[5] ), .Z(new_n787_));
  NOR3_X1    g00531(.A1(new_n782_), .A2(new_n780_), .A3(new_n787_), .ZN(new_n788_));
  NOR2_X1    g00532(.A1(new_n782_), .A2(new_n780_), .ZN(new_n789_));
  INV_X1     g00533(.I(new_n787_), .ZN(new_n790_));
  NOR2_X1    g00534(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1   g00535(.A1(new_n788_), .A2(new_n791_), .B(new_n734_), .ZN(new_n792_));
  XOR2_X1    g00536(.A1(new_n789_), .A2(new_n787_), .Z(new_n793_));
  OAI21_X1   g00537(.A1(new_n734_), .A2(new_n793_), .B(new_n792_), .ZN(new_n794_));
  INV_X1     g00538(.I(\b[13] ), .ZN(new_n795_));
  NOR2_X1    g00539(.A1(new_n709_), .A2(new_n710_), .ZN(new_n796_));
  XOR2_X1    g00540(.A1(new_n796_), .A2(new_n659_), .Z(new_n797_));
  NAND2_X1   g00541(.A1(new_n797_), .A2(new_n713_), .ZN(new_n798_));
  XOR2_X1    g00542(.A1(new_n798_), .A2(new_n795_), .Z(new_n799_));
  OAI22_X1   g00543(.A1(new_n405_), .A2(new_n795_), .B1(new_n717_), .B2(new_n404_), .ZN(new_n800_));
  NAND2_X1   g00544(.A1(new_n279_), .A2(\b[11] ), .ZN(new_n801_));
  AOI21_X1   g00545(.A1(new_n800_), .A2(new_n801_), .B(new_n264_), .ZN(new_n802_));
  NAND2_X1   g00546(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  XOR2_X1    g00547(.A1(new_n803_), .A2(\a[2] ), .Z(new_n804_));
  XOR2_X1    g00548(.A1(new_n794_), .A2(new_n804_), .Z(\f[13] ));
  INV_X1     g00549(.I(new_n804_), .ZN(new_n806_));
  NAND2_X1   g00550(.A1(new_n794_), .A2(new_n806_), .ZN(new_n807_));
  OAI22_X1   g00551(.A1(new_n582_), .A2(new_n347_), .B1(new_n393_), .B2(new_n577_), .ZN(new_n808_));
  OAI21_X1   g00552(.A1(new_n290_), .A2(new_n635_), .B(new_n808_), .ZN(new_n809_));
  AOI21_X1   g00553(.A1(new_n352_), .A2(new_n584_), .B(new_n809_), .ZN(new_n810_));
  XOR2_X1    g00554(.A1(new_n810_), .A2(new_n572_), .Z(new_n811_));
  OAI22_X1   g00555(.A1(new_n437_), .A2(new_n495_), .B1(new_n450_), .B2(new_n431_), .ZN(new_n812_));
  NAND2_X1   g00556(.A1(new_n775_), .A2(\b[6] ), .ZN(new_n813_));
  AOI21_X1   g00557(.A1(new_n812_), .A2(new_n813_), .B(new_n440_), .ZN(new_n814_));
  NAND2_X1   g00558(.A1(new_n494_), .A2(new_n814_), .ZN(new_n815_));
  XOR2_X1    g00559(.A1(new_n815_), .A2(\a[8] ), .Z(new_n816_));
  OAI21_X1   g00560(.A1(new_n742_), .A2(new_n768_), .B(new_n770_), .ZN(new_n817_));
  NAND2_X1   g00561(.A1(new_n762_), .A2(new_n763_), .ZN(new_n818_));
  NOR2_X1    g00562(.A1(new_n760_), .A2(new_n278_), .ZN(new_n819_));
  XNOR2_X1   g00563(.A1(\a[11] ), .A2(\a[13] ), .ZN(new_n820_));
  NAND2_X1   g00564(.A1(new_n682_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1   g00565(.A1(\a[11] ), .A2(\a[14] ), .ZN(new_n822_));
  NAND2_X1   g00566(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI22_X1   g00567(.A1(new_n757_), .A2(new_n292_), .B1(new_n267_), .B2(new_n752_), .ZN(new_n824_));
  NOR4_X1    g00568(.A1(new_n824_), .A2(new_n258_), .A3(new_n819_), .A4(new_n823_), .ZN(new_n825_));
  XOR2_X1    g00569(.A1(new_n825_), .A2(new_n747_), .Z(new_n826_));
  XOR2_X1    g00570(.A1(new_n818_), .A2(new_n826_), .Z(new_n827_));
  INV_X1     g00571(.I(new_n827_), .ZN(new_n828_));
  XOR2_X1    g00572(.A1(new_n817_), .A2(new_n828_), .Z(new_n829_));
  XOR2_X1    g00573(.A1(new_n829_), .A2(new_n816_), .Z(new_n830_));
  XOR2_X1    g00574(.A1(new_n830_), .A2(new_n811_), .Z(new_n831_));
  XOR2_X1    g00575(.A1(new_n831_), .A2(new_n780_), .Z(new_n832_));
  OAI22_X1   g00576(.A1(new_n364_), .A2(new_n659_), .B1(new_n617_), .B2(new_n320_), .ZN(new_n833_));
  NAND2_X1   g00577(.A1(new_n594_), .A2(\b[9] ), .ZN(new_n834_));
  AOI21_X1   g00578(.A1(new_n833_), .A2(new_n834_), .B(new_n312_), .ZN(new_n835_));
  NAND2_X1   g00579(.A1(new_n663_), .A2(new_n835_), .ZN(new_n836_));
  XOR2_X1    g00580(.A1(new_n836_), .A2(\a[5] ), .Z(new_n837_));
  XOR2_X1    g00581(.A1(new_n832_), .A2(new_n837_), .Z(new_n838_));
  AOI21_X1   g00582(.A1(\b[11] ), .A2(\b[13] ), .B(\b[12] ), .ZN(new_n839_));
  AOI21_X1   g00583(.A1(new_n659_), .A2(new_n795_), .B(new_n717_), .ZN(new_n840_));
  INV_X1     g00584(.I(new_n840_), .ZN(new_n841_));
  OAI21_X1   g00585(.A1(new_n711_), .A2(new_n839_), .B(new_n841_), .ZN(new_n842_));
  XNOR2_X1   g00586(.A1(\b[13] ), .A2(\b[14] ), .ZN(new_n843_));
  INV_X1     g00587(.I(new_n843_), .ZN(new_n844_));
  NAND2_X1   g00588(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  XOR2_X1    g00589(.A1(\b[13] ), .A2(\b[14] ), .Z(new_n846_));
  OAI21_X1   g00590(.A1(new_n842_), .A2(new_n846_), .B(new_n845_), .ZN(new_n847_));
  INV_X1     g00591(.I(\b[14] ), .ZN(new_n848_));
  OAI22_X1   g00592(.A1(new_n405_), .A2(new_n848_), .B1(new_n795_), .B2(new_n404_), .ZN(new_n849_));
  NAND2_X1   g00593(.A1(new_n279_), .A2(\b[12] ), .ZN(new_n850_));
  AOI21_X1   g00594(.A1(new_n849_), .A2(new_n850_), .B(new_n264_), .ZN(new_n851_));
  NAND2_X1   g00595(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  XOR2_X1    g00596(.A1(new_n852_), .A2(\a[2] ), .Z(new_n853_));
  NOR2_X1    g00597(.A1(new_n734_), .A2(new_n791_), .ZN(new_n854_));
  XNOR2_X1   g00598(.A1(new_n854_), .A2(new_n853_), .ZN(new_n855_));
  XOR2_X1    g00599(.A1(new_n838_), .A2(new_n855_), .Z(new_n856_));
  XOR2_X1    g00600(.A1(new_n856_), .A2(new_n807_), .Z(\f[14] ));
  NAND3_X1   g00601(.A1(new_n826_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n858_));
  NOR2_X1    g00602(.A1(new_n823_), .A2(new_n267_), .ZN(new_n859_));
  OAI22_X1   g00603(.A1(new_n757_), .A2(new_n290_), .B1(new_n292_), .B2(new_n752_), .ZN(new_n860_));
  NOR4_X1    g00604(.A1(new_n860_), .A2(new_n677_), .A3(new_n760_), .A4(new_n859_), .ZN(new_n861_));
  XOR2_X1    g00605(.A1(new_n861_), .A2(new_n747_), .Z(new_n862_));
  XNOR2_X1   g00606(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n863_));
  NOR2_X1    g00607(.A1(new_n863_), .A2(new_n258_), .ZN(new_n864_));
  XOR2_X1    g00608(.A1(new_n862_), .A2(new_n864_), .Z(new_n865_));
  XNOR2_X1   g00609(.A1(new_n865_), .A2(new_n858_), .ZN(new_n866_));
  INV_X1     g00610(.I(new_n577_), .ZN(new_n867_));
  AOI22_X1   g00611(.A1(\b[6] ), .A2(new_n581_), .B1(new_n867_), .B2(\b[5] ), .ZN(new_n868_));
  NOR2_X1    g00612(.A1(new_n635_), .A2(new_n393_), .ZN(new_n869_));
  OAI21_X1   g00613(.A1(new_n868_), .A2(new_n869_), .B(new_n584_), .ZN(new_n870_));
  NOR2_X1    g00614(.A1(new_n524_), .A2(new_n870_), .ZN(new_n871_));
  XOR2_X1    g00615(.A1(new_n871_), .A2(new_n572_), .Z(new_n872_));
  NAND2_X1   g00616(.A1(new_n828_), .A2(new_n811_), .ZN(new_n873_));
  XOR2_X1    g00617(.A1(new_n742_), .A2(new_n767_), .Z(new_n874_));
  XOR2_X1    g00618(.A1(new_n818_), .A2(new_n826_), .Z(new_n875_));
  XOR2_X1    g00619(.A1(new_n875_), .A2(new_n572_), .Z(new_n876_));
  NAND2_X1   g00620(.A1(new_n876_), .A2(new_n810_), .ZN(new_n877_));
  OR2_X2     g00621(.A1(new_n876_), .A2(new_n810_), .Z(new_n878_));
  NAND3_X1   g00622(.A1(new_n878_), .A2(new_n767_), .A3(new_n877_), .ZN(new_n879_));
  OAI21_X1   g00623(.A1(new_n879_), .A2(new_n742_), .B(new_n764_), .ZN(new_n880_));
  OAI21_X1   g00624(.A1(new_n874_), .A2(new_n880_), .B(new_n873_), .ZN(new_n881_));
  XOR2_X1    g00625(.A1(new_n881_), .A2(new_n872_), .Z(new_n882_));
  XNOR2_X1   g00626(.A1(new_n882_), .A2(new_n866_), .ZN(new_n883_));
  OAI22_X1   g00627(.A1(new_n437_), .A2(new_n510_), .B1(new_n495_), .B2(new_n431_), .ZN(new_n884_));
  NAND2_X1   g00628(.A1(new_n775_), .A2(\b[7] ), .ZN(new_n885_));
  AOI21_X1   g00629(.A1(new_n884_), .A2(new_n885_), .B(new_n440_), .ZN(new_n886_));
  NAND2_X1   g00630(.A1(new_n518_), .A2(new_n886_), .ZN(new_n887_));
  XOR2_X1    g00631(.A1(new_n887_), .A2(new_n429_), .Z(new_n888_));
  XOR2_X1    g00632(.A1(new_n883_), .A2(new_n888_), .Z(new_n889_));
  XOR2_X1    g00633(.A1(new_n827_), .A2(new_n811_), .Z(new_n890_));
  XOR2_X1    g00634(.A1(new_n817_), .A2(new_n890_), .Z(new_n891_));
  AOI21_X1   g00635(.A1(new_n891_), .A2(new_n816_), .B(new_n780_), .ZN(new_n892_));
  XOR2_X1    g00636(.A1(new_n889_), .A2(new_n892_), .Z(new_n893_));
  INV_X1     g00637(.I(new_n893_), .ZN(new_n894_));
  OAI22_X1   g00638(.A1(new_n364_), .A2(new_n717_), .B1(new_n659_), .B2(new_n320_), .ZN(new_n895_));
  NAND2_X1   g00639(.A1(new_n594_), .A2(\b[10] ), .ZN(new_n896_));
  AOI21_X1   g00640(.A1(new_n895_), .A2(new_n896_), .B(new_n312_), .ZN(new_n897_));
  NAND2_X1   g00641(.A1(new_n716_), .A2(new_n897_), .ZN(new_n898_));
  XOR2_X1    g00642(.A1(new_n898_), .A2(\a[5] ), .Z(new_n899_));
  NOR2_X1    g00643(.A1(new_n894_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1     g00644(.I(new_n900_), .ZN(new_n901_));
  NAND2_X1   g00645(.A1(new_n894_), .A2(new_n899_), .ZN(new_n902_));
  NAND2_X1   g00646(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1     g00647(.I(\b[15] ), .ZN(new_n904_));
  XOR2_X1    g00648(.A1(new_n842_), .A2(\b[13] ), .Z(new_n905_));
  NAND2_X1   g00649(.A1(new_n905_), .A2(new_n844_), .ZN(new_n906_));
  XOR2_X1    g00650(.A1(new_n906_), .A2(new_n904_), .Z(new_n907_));
  OAI22_X1   g00651(.A1(new_n405_), .A2(new_n904_), .B1(new_n848_), .B2(new_n404_), .ZN(new_n908_));
  NAND2_X1   g00652(.A1(new_n279_), .A2(\b[13] ), .ZN(new_n909_));
  AOI21_X1   g00653(.A1(new_n908_), .A2(new_n909_), .B(new_n264_), .ZN(new_n910_));
  NAND2_X1   g00654(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  XOR2_X1    g00655(.A1(new_n911_), .A2(new_n271_), .Z(new_n912_));
  XNOR2_X1   g00656(.A1(new_n838_), .A2(new_n854_), .ZN(new_n913_));
  NAND2_X1   g00657(.A1(new_n913_), .A2(new_n853_), .ZN(new_n914_));
  NAND3_X1   g00658(.A1(new_n914_), .A2(new_n807_), .A3(new_n856_), .ZN(new_n915_));
  XOR2_X1    g00659(.A1(new_n915_), .A2(new_n912_), .Z(new_n916_));
  XOR2_X1    g00660(.A1(new_n916_), .A2(new_n903_), .Z(\f[15] ));
  NAND2_X1   g00661(.A1(new_n865_), .A2(new_n826_), .ZN(new_n918_));
  NAND2_X1   g00662(.A1(new_n918_), .A2(new_n818_), .ZN(new_n919_));
  INV_X1     g00663(.I(new_n919_), .ZN(new_n920_));
  NAND2_X1   g00664(.A1(new_n862_), .A2(new_n864_), .ZN(new_n921_));
  NOR2_X1    g00665(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1   g00666(.A1(new_n920_), .A2(new_n921_), .ZN(new_n923_));
  INV_X1     g00667(.I(new_n923_), .ZN(new_n924_));
  NOR2_X1    g00668(.A1(new_n924_), .A2(new_n922_), .ZN(new_n925_));
  OAI22_X1   g00669(.A1(new_n757_), .A2(new_n393_), .B1(new_n290_), .B2(new_n752_), .ZN(new_n926_));
  OAI21_X1   g00670(.A1(new_n292_), .A2(new_n823_), .B(new_n926_), .ZN(new_n927_));
  NAND3_X1   g00671(.A1(new_n927_), .A2(new_n334_), .A3(new_n759_), .ZN(new_n928_));
  XOR2_X1    g00672(.A1(new_n928_), .A2(\a[14] ), .Z(new_n929_));
  INV_X1     g00673(.I(\a[17] ), .ZN(new_n930_));
  INV_X1     g00674(.I(\a[16] ), .ZN(new_n931_));
  NOR3_X1    g00675(.A1(new_n931_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n932_));
  NAND3_X1   g00676(.A1(new_n931_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n933_));
  INV_X1     g00677(.I(new_n933_), .ZN(new_n934_));
  NOR2_X1    g00678(.A1(new_n934_), .A2(new_n932_), .ZN(new_n935_));
  NOR2_X1    g00679(.A1(new_n935_), .A2(new_n258_), .ZN(new_n936_));
  INV_X1     g00680(.I(new_n863_), .ZN(new_n937_));
  XNOR2_X1   g00681(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n938_));
  NOR2_X1    g00682(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  INV_X1     g00683(.I(new_n939_), .ZN(new_n940_));
  NOR2_X1    g00684(.A1(new_n940_), .A2(new_n267_), .ZN(new_n941_));
  NOR2_X1    g00685(.A1(new_n863_), .A2(new_n938_), .ZN(new_n942_));
  INV_X1     g00686(.I(new_n942_), .ZN(new_n943_));
  NOR4_X1    g00687(.A1(new_n941_), .A2(new_n261_), .A3(new_n936_), .A4(new_n943_), .ZN(new_n944_));
  XOR2_X1    g00688(.A1(new_n944_), .A2(new_n930_), .Z(new_n945_));
  NOR2_X1    g00689(.A1(new_n864_), .A2(new_n930_), .ZN(new_n946_));
  XNOR2_X1   g00690(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  XOR2_X1    g00691(.A1(new_n947_), .A2(new_n929_), .Z(new_n948_));
  NOR2_X1    g00692(.A1(new_n925_), .A2(new_n948_), .ZN(new_n949_));
  INV_X1     g00693(.I(new_n925_), .ZN(new_n950_));
  INV_X1     g00694(.I(new_n929_), .ZN(new_n951_));
  NOR2_X1    g00695(.A1(new_n947_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1     g00696(.I(new_n947_), .ZN(new_n953_));
  NOR2_X1    g00697(.A1(new_n953_), .A2(new_n929_), .ZN(new_n954_));
  NOR2_X1    g00698(.A1(new_n954_), .A2(new_n952_), .ZN(new_n955_));
  NOR2_X1    g00699(.A1(new_n950_), .A2(new_n955_), .ZN(new_n956_));
  NOR2_X1    g00700(.A1(new_n956_), .A2(new_n949_), .ZN(new_n957_));
  INV_X1     g00701(.I(new_n957_), .ZN(new_n958_));
  OAI22_X1   g00702(.A1(new_n582_), .A2(new_n450_), .B1(new_n403_), .B2(new_n577_), .ZN(new_n959_));
  INV_X1     g00703(.I(new_n635_), .ZN(new_n960_));
  NAND2_X1   g00704(.A1(new_n960_), .A2(\b[5] ), .ZN(new_n961_));
  AOI21_X1   g00705(.A1(new_n959_), .A2(new_n961_), .B(new_n585_), .ZN(new_n962_));
  NAND2_X1   g00706(.A1(new_n454_), .A2(new_n962_), .ZN(new_n963_));
  XOR2_X1    g00707(.A1(new_n963_), .A2(\a[11] ), .Z(new_n964_));
  NOR2_X1    g00708(.A1(new_n958_), .A2(new_n964_), .ZN(new_n965_));
  INV_X1     g00709(.I(new_n965_), .ZN(new_n966_));
  NAND2_X1   g00710(.A1(new_n958_), .A2(new_n964_), .ZN(new_n967_));
  NAND2_X1   g00711(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  OAI22_X1   g00712(.A1(new_n437_), .A2(new_n617_), .B1(new_n510_), .B2(new_n431_), .ZN(new_n969_));
  NAND2_X1   g00713(.A1(new_n775_), .A2(\b[8] ), .ZN(new_n970_));
  AOI21_X1   g00714(.A1(new_n969_), .A2(new_n970_), .B(new_n440_), .ZN(new_n971_));
  NAND2_X1   g00715(.A1(new_n616_), .A2(new_n971_), .ZN(new_n972_));
  XOR2_X1    g00716(.A1(new_n972_), .A2(\a[8] ), .Z(new_n973_));
  XNOR2_X1   g00717(.A1(new_n968_), .A2(new_n973_), .ZN(new_n974_));
  OAI22_X1   g00718(.A1(new_n364_), .A2(new_n795_), .B1(new_n717_), .B2(new_n320_), .ZN(new_n975_));
  NAND2_X1   g00719(.A1(new_n594_), .A2(\b[11] ), .ZN(new_n976_));
  AOI21_X1   g00720(.A1(new_n975_), .A2(new_n976_), .B(new_n312_), .ZN(new_n977_));
  NAND2_X1   g00721(.A1(new_n799_), .A2(new_n977_), .ZN(new_n978_));
  XOR2_X1    g00722(.A1(new_n978_), .A2(\a[5] ), .Z(new_n979_));
  XNOR2_X1   g00723(.A1(new_n974_), .A2(new_n979_), .ZN(new_n980_));
  XOR2_X1    g00724(.A1(new_n900_), .A2(new_n980_), .Z(new_n981_));
  AOI21_X1   g00725(.A1(\b[13] ), .A2(\b[15] ), .B(\b[14] ), .ZN(new_n982_));
  NOR2_X1    g00726(.A1(new_n842_), .A2(new_n982_), .ZN(new_n983_));
  AOI21_X1   g00727(.A1(new_n795_), .A2(new_n904_), .B(new_n848_), .ZN(new_n984_));
  NOR2_X1    g00728(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  INV_X1     g00729(.I(new_n985_), .ZN(new_n986_));
  XNOR2_X1   g00730(.A1(\b[15] ), .A2(\b[16] ), .ZN(new_n987_));
  INV_X1     g00731(.I(new_n987_), .ZN(new_n988_));
  NAND2_X1   g00732(.A1(new_n986_), .A2(new_n988_), .ZN(new_n989_));
  XOR2_X1    g00733(.A1(\b[15] ), .A2(\b[16] ), .Z(new_n990_));
  OAI21_X1   g00734(.A1(new_n986_), .A2(new_n990_), .B(new_n989_), .ZN(new_n991_));
  INV_X1     g00735(.I(\b[16] ), .ZN(new_n992_));
  OAI22_X1   g00736(.A1(new_n405_), .A2(new_n992_), .B1(new_n904_), .B2(new_n404_), .ZN(new_n993_));
  NAND2_X1   g00737(.A1(new_n279_), .A2(\b[14] ), .ZN(new_n994_));
  AOI21_X1   g00738(.A1(new_n993_), .A2(new_n994_), .B(new_n264_), .ZN(new_n995_));
  NAND2_X1   g00739(.A1(new_n991_), .A2(new_n995_), .ZN(new_n996_));
  XOR2_X1    g00740(.A1(new_n996_), .A2(\a[2] ), .Z(new_n997_));
  INV_X1     g00741(.I(new_n997_), .ZN(new_n998_));
  NAND2_X1   g00742(.A1(new_n981_), .A2(new_n998_), .ZN(new_n999_));
  NOR2_X1    g00743(.A1(new_n981_), .A2(new_n998_), .ZN(new_n1000_));
  INV_X1     g00744(.I(new_n1000_), .ZN(new_n1001_));
  NAND2_X1   g00745(.A1(new_n1001_), .A2(new_n999_), .ZN(\f[16] ));
  OAI22_X1   g00746(.A1(new_n757_), .A2(new_n347_), .B1(new_n393_), .B2(new_n752_), .ZN(new_n1003_));
  OAI21_X1   g00747(.A1(new_n290_), .A2(new_n823_), .B(new_n1003_), .ZN(new_n1004_));
  AOI21_X1   g00748(.A1(new_n352_), .A2(new_n759_), .B(new_n1004_), .ZN(new_n1005_));
  XOR2_X1    g00749(.A1(new_n1005_), .A2(new_n747_), .Z(new_n1006_));
  INV_X1     g00750(.I(new_n1006_), .ZN(new_n1007_));
  OAI22_X1   g00751(.A1(new_n582_), .A2(new_n495_), .B1(new_n450_), .B2(new_n577_), .ZN(new_n1008_));
  NAND2_X1   g00752(.A1(new_n960_), .A2(\b[6] ), .ZN(new_n1009_));
  AOI21_X1   g00753(.A1(new_n1008_), .A2(new_n1009_), .B(new_n585_), .ZN(new_n1010_));
  NAND2_X1   g00754(.A1(new_n494_), .A2(new_n1010_), .ZN(new_n1011_));
  XOR2_X1    g00755(.A1(new_n1011_), .A2(\a[11] ), .Z(new_n1012_));
  INV_X1     g00756(.I(new_n954_), .ZN(new_n1013_));
  OAI21_X1   g00757(.A1(new_n925_), .A2(new_n952_), .B(new_n1013_), .ZN(new_n1014_));
  NAND2_X1   g00758(.A1(new_n945_), .A2(new_n946_), .ZN(new_n1015_));
  NOR2_X1    g00759(.A1(new_n943_), .A2(new_n278_), .ZN(new_n1016_));
  XNOR2_X1   g00760(.A1(\a[14] ), .A2(\a[16] ), .ZN(new_n1017_));
  NAND2_X1   g00761(.A1(new_n863_), .A2(new_n1017_), .ZN(new_n1018_));
  XNOR2_X1   g00762(.A1(\a[14] ), .A2(\a[17] ), .ZN(new_n1019_));
  NAND2_X1   g00763(.A1(new_n1018_), .A2(new_n1019_), .ZN(new_n1020_));
  OAI22_X1   g00764(.A1(new_n940_), .A2(new_n292_), .B1(new_n267_), .B2(new_n935_), .ZN(new_n1021_));
  NOR4_X1    g00765(.A1(new_n1021_), .A2(new_n258_), .A3(new_n1016_), .A4(new_n1020_), .ZN(new_n1022_));
  XOR2_X1    g00766(.A1(new_n1022_), .A2(new_n930_), .Z(new_n1023_));
  XOR2_X1    g00767(.A1(new_n1015_), .A2(new_n1023_), .Z(new_n1024_));
  INV_X1     g00768(.I(new_n1024_), .ZN(new_n1025_));
  XOR2_X1    g00769(.A1(new_n1014_), .A2(new_n1025_), .Z(new_n1026_));
  XOR2_X1    g00770(.A1(new_n1026_), .A2(new_n1012_), .Z(new_n1027_));
  XOR2_X1    g00771(.A1(new_n1027_), .A2(new_n1007_), .Z(new_n1028_));
  XOR2_X1    g00772(.A1(new_n1028_), .A2(new_n966_), .Z(new_n1029_));
  OAI22_X1   g00773(.A1(new_n437_), .A2(new_n659_), .B1(new_n617_), .B2(new_n431_), .ZN(new_n1030_));
  NAND2_X1   g00774(.A1(new_n775_), .A2(\b[9] ), .ZN(new_n1031_));
  AOI21_X1   g00775(.A1(new_n1030_), .A2(new_n1031_), .B(new_n440_), .ZN(new_n1032_));
  NAND2_X1   g00776(.A1(new_n663_), .A2(new_n1032_), .ZN(new_n1033_));
  XOR2_X1    g00777(.A1(new_n1033_), .A2(\a[8] ), .Z(new_n1034_));
  XOR2_X1    g00778(.A1(new_n1029_), .A2(new_n1034_), .Z(new_n1035_));
  NOR2_X1    g00779(.A1(new_n968_), .A2(new_n973_), .ZN(new_n1036_));
  XOR2_X1    g00780(.A1(new_n1035_), .A2(new_n1036_), .Z(new_n1037_));
  OAI22_X1   g00781(.A1(new_n364_), .A2(new_n848_), .B1(new_n795_), .B2(new_n320_), .ZN(new_n1038_));
  NAND2_X1   g00782(.A1(new_n594_), .A2(\b[12] ), .ZN(new_n1039_));
  AOI21_X1   g00783(.A1(new_n1038_), .A2(new_n1039_), .B(new_n312_), .ZN(new_n1040_));
  NAND2_X1   g00784(.A1(new_n847_), .A2(new_n1040_), .ZN(new_n1041_));
  XOR2_X1    g00785(.A1(new_n1041_), .A2(\a[5] ), .Z(new_n1042_));
  XOR2_X1    g00786(.A1(new_n1037_), .A2(new_n1042_), .Z(new_n1043_));
  INV_X1     g00787(.I(\b[17] ), .ZN(new_n1044_));
  XOR2_X1    g00788(.A1(new_n985_), .A2(new_n904_), .Z(new_n1045_));
  NAND2_X1   g00789(.A1(new_n1045_), .A2(new_n988_), .ZN(new_n1046_));
  XOR2_X1    g00790(.A1(new_n1046_), .A2(new_n1044_), .Z(new_n1047_));
  OAI22_X1   g00791(.A1(new_n405_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n404_), .ZN(new_n1048_));
  NAND2_X1   g00792(.A1(new_n279_), .A2(\b[15] ), .ZN(new_n1049_));
  AOI21_X1   g00793(.A1(new_n1048_), .A2(new_n1049_), .B(new_n264_), .ZN(new_n1050_));
  NAND2_X1   g00794(.A1(new_n1047_), .A2(new_n1050_), .ZN(new_n1051_));
  XOR2_X1    g00795(.A1(new_n1051_), .A2(\a[2] ), .Z(new_n1052_));
  NAND2_X1   g00796(.A1(new_n974_), .A2(new_n979_), .ZN(new_n1053_));
  NAND2_X1   g00797(.A1(new_n901_), .A2(new_n1053_), .ZN(new_n1054_));
  XOR2_X1    g00798(.A1(new_n1054_), .A2(new_n1052_), .Z(new_n1055_));
  XOR2_X1    g00799(.A1(new_n1055_), .A2(new_n1043_), .Z(new_n1056_));
  NAND2_X1   g00800(.A1(new_n981_), .A2(new_n998_), .ZN(new_n1057_));
  XOR2_X1    g00801(.A1(new_n1056_), .A2(new_n1057_), .Z(\f[17] ));
  INV_X1     g00802(.I(new_n752_), .ZN(new_n1059_));
  AOI22_X1   g00803(.A1(\b[6] ), .A2(new_n756_), .B1(new_n1059_), .B2(\b[5] ), .ZN(new_n1060_));
  NOR2_X1    g00804(.A1(new_n823_), .A2(new_n393_), .ZN(new_n1061_));
  OAI21_X1   g00805(.A1(new_n1060_), .A2(new_n1061_), .B(new_n759_), .ZN(new_n1062_));
  NOR2_X1    g00806(.A1(new_n524_), .A2(new_n1062_), .ZN(new_n1063_));
  XOR2_X1    g00807(.A1(new_n1063_), .A2(\a[14] ), .Z(new_n1064_));
  XNOR2_X1   g00808(.A1(\a[17] ), .A2(\a[18] ), .ZN(new_n1065_));
  NOR2_X1    g00809(.A1(new_n1065_), .A2(new_n258_), .ZN(new_n1066_));
  INV_X1     g00810(.I(new_n1023_), .ZN(new_n1067_));
  NOR2_X1    g00811(.A1(new_n1067_), .A2(new_n1015_), .ZN(new_n1068_));
  NOR2_X1    g00812(.A1(new_n1020_), .A2(new_n267_), .ZN(new_n1069_));
  OAI22_X1   g00813(.A1(new_n940_), .A2(new_n290_), .B1(new_n292_), .B2(new_n935_), .ZN(new_n1070_));
  NOR4_X1    g00814(.A1(new_n1070_), .A2(new_n677_), .A3(new_n943_), .A4(new_n1069_), .ZN(new_n1071_));
  XOR2_X1    g00815(.A1(new_n1071_), .A2(new_n930_), .Z(new_n1072_));
  XOR2_X1    g00816(.A1(new_n1068_), .A2(new_n1072_), .Z(new_n1073_));
  XOR2_X1    g00817(.A1(new_n1073_), .A2(new_n1066_), .Z(new_n1074_));
  XOR2_X1    g00818(.A1(new_n1074_), .A2(new_n1064_), .Z(new_n1075_));
  XOR2_X1    g00819(.A1(new_n925_), .A2(new_n929_), .Z(new_n1076_));
  INV_X1     g00820(.I(new_n1015_), .ZN(new_n1077_));
  NOR2_X1    g00821(.A1(new_n1077_), .A2(new_n1023_), .ZN(new_n1078_));
  NOR2_X1    g00822(.A1(new_n1078_), .A2(new_n1068_), .ZN(new_n1079_));
  XOR2_X1    g00823(.A1(new_n1079_), .A2(\a[14] ), .Z(new_n1080_));
  OAI21_X1   g00824(.A1(new_n1080_), .A2(new_n1005_), .B(new_n951_), .ZN(new_n1081_));
  AOI21_X1   g00825(.A1(new_n1005_), .A2(new_n1080_), .B(new_n1081_), .ZN(new_n1082_));
  AOI21_X1   g00826(.A1(new_n950_), .A2(new_n1082_), .B(new_n953_), .ZN(new_n1083_));
  NAND2_X1   g00827(.A1(new_n1076_), .A2(new_n1083_), .ZN(new_n1084_));
  OAI21_X1   g00828(.A1(new_n1007_), .A2(new_n1024_), .B(new_n1084_), .ZN(new_n1085_));
  NAND2_X1   g00829(.A1(new_n1085_), .A2(new_n1075_), .ZN(new_n1086_));
  AOI21_X1   g00830(.A1(new_n1006_), .A2(new_n1025_), .B(new_n1075_), .ZN(new_n1087_));
  NAND2_X1   g00831(.A1(new_n1084_), .A2(new_n1087_), .ZN(new_n1088_));
  NAND2_X1   g00832(.A1(new_n1086_), .A2(new_n1088_), .ZN(new_n1089_));
  OAI22_X1   g00833(.A1(new_n582_), .A2(new_n510_), .B1(new_n495_), .B2(new_n577_), .ZN(new_n1090_));
  NAND2_X1   g00834(.A1(new_n960_), .A2(\b[7] ), .ZN(new_n1091_));
  AOI21_X1   g00835(.A1(new_n1090_), .A2(new_n1091_), .B(new_n585_), .ZN(new_n1092_));
  NAND2_X1   g00836(.A1(new_n518_), .A2(new_n1092_), .ZN(new_n1093_));
  XOR2_X1    g00837(.A1(new_n1093_), .A2(\a[11] ), .Z(new_n1094_));
  XOR2_X1    g00838(.A1(new_n1024_), .A2(new_n1006_), .Z(new_n1095_));
  XOR2_X1    g00839(.A1(new_n1014_), .A2(new_n1095_), .Z(new_n1096_));
  NAND2_X1   g00840(.A1(new_n1096_), .A2(new_n1012_), .ZN(new_n1097_));
  NAND2_X1   g00841(.A1(new_n966_), .A2(new_n1097_), .ZN(new_n1098_));
  XOR2_X1    g00842(.A1(new_n1098_), .A2(new_n1094_), .Z(new_n1099_));
  XOR2_X1    g00843(.A1(new_n1099_), .A2(new_n1089_), .Z(new_n1100_));
  OAI22_X1   g00844(.A1(new_n437_), .A2(new_n717_), .B1(new_n659_), .B2(new_n431_), .ZN(new_n1101_));
  NAND2_X1   g00845(.A1(new_n775_), .A2(\b[10] ), .ZN(new_n1102_));
  AOI21_X1   g00846(.A1(new_n1101_), .A2(new_n1102_), .B(new_n440_), .ZN(new_n1103_));
  NAND2_X1   g00847(.A1(new_n716_), .A2(new_n1103_), .ZN(new_n1104_));
  XOR2_X1    g00848(.A1(new_n1104_), .A2(new_n429_), .Z(new_n1105_));
  AOI21_X1   g00849(.A1(new_n1029_), .A2(new_n1034_), .B(new_n1036_), .ZN(new_n1106_));
  XOR2_X1    g00850(.A1(new_n1106_), .A2(new_n1105_), .Z(new_n1107_));
  XNOR2_X1   g00851(.A1(new_n1107_), .A2(new_n1100_), .ZN(new_n1108_));
  OAI22_X1   g00852(.A1(new_n364_), .A2(new_n904_), .B1(new_n848_), .B2(new_n320_), .ZN(new_n1109_));
  NAND2_X1   g00853(.A1(new_n594_), .A2(\b[13] ), .ZN(new_n1110_));
  AOI21_X1   g00854(.A1(new_n1109_), .A2(new_n1110_), .B(new_n312_), .ZN(new_n1111_));
  NAND2_X1   g00855(.A1(new_n907_), .A2(new_n1111_), .ZN(new_n1112_));
  XOR2_X1    g00856(.A1(new_n1112_), .A2(\a[5] ), .Z(new_n1113_));
  XOR2_X1    g00857(.A1(new_n1108_), .A2(new_n1113_), .Z(new_n1114_));
  AOI21_X1   g00858(.A1(\b[15] ), .A2(\b[17] ), .B(\b[16] ), .ZN(new_n1115_));
  AOI21_X1   g00859(.A1(new_n904_), .A2(new_n1044_), .B(new_n992_), .ZN(new_n1116_));
  INV_X1     g00860(.I(new_n1116_), .ZN(new_n1117_));
  OAI21_X1   g00861(.A1(new_n986_), .A2(new_n1115_), .B(new_n1117_), .ZN(new_n1118_));
  XNOR2_X1   g00862(.A1(\b[17] ), .A2(\b[18] ), .ZN(new_n1119_));
  INV_X1     g00863(.I(new_n1119_), .ZN(new_n1120_));
  NAND2_X1   g00864(.A1(new_n1118_), .A2(new_n1120_), .ZN(new_n1121_));
  XOR2_X1    g00865(.A1(\b[17] ), .A2(\b[18] ), .Z(new_n1122_));
  OAI21_X1   g00866(.A1(new_n1118_), .A2(new_n1122_), .B(new_n1121_), .ZN(new_n1123_));
  INV_X1     g00867(.I(\b[18] ), .ZN(new_n1124_));
  OAI22_X1   g00868(.A1(new_n405_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n404_), .ZN(new_n1125_));
  NAND2_X1   g00869(.A1(new_n279_), .A2(\b[16] ), .ZN(new_n1126_));
  AOI21_X1   g00870(.A1(new_n1125_), .A2(new_n1126_), .B(new_n264_), .ZN(new_n1127_));
  NAND2_X1   g00871(.A1(new_n1123_), .A2(new_n1127_), .ZN(new_n1128_));
  XOR2_X1    g00872(.A1(new_n1128_), .A2(\a[2] ), .Z(new_n1129_));
  XOR2_X1    g00873(.A1(new_n1114_), .A2(new_n1129_), .Z(new_n1130_));
  INV_X1     g00874(.I(new_n1130_), .ZN(new_n1131_));
  NAND2_X1   g00875(.A1(new_n1056_), .A2(new_n1001_), .ZN(new_n1132_));
  XNOR2_X1   g00876(.A1(new_n1043_), .A2(new_n1054_), .ZN(new_n1133_));
  INV_X1     g00877(.I(new_n1133_), .ZN(new_n1134_));
  AOI21_X1   g00878(.A1(new_n1052_), .A2(new_n1134_), .B(new_n1132_), .ZN(new_n1135_));
  XOR2_X1    g00879(.A1(new_n1135_), .A2(new_n1131_), .Z(\f[18] ));
  INV_X1     g00880(.I(new_n1094_), .ZN(new_n1137_));
  XOR2_X1    g00881(.A1(new_n1089_), .A2(new_n1094_), .Z(new_n1138_));
  AOI21_X1   g00882(.A1(new_n1137_), .A2(new_n1098_), .B(new_n1138_), .ZN(new_n1139_));
  INV_X1     g00883(.I(new_n1139_), .ZN(new_n1140_));
  XOR2_X1    g00884(.A1(new_n1072_), .A2(new_n1066_), .Z(new_n1141_));
  NAND2_X1   g00885(.A1(new_n1141_), .A2(new_n1068_), .ZN(new_n1142_));
  NOR2_X1    g00886(.A1(new_n1141_), .A2(new_n1068_), .ZN(new_n1143_));
  NOR2_X1    g00887(.A1(new_n1143_), .A2(new_n1064_), .ZN(new_n1144_));
  NAND3_X1   g00888(.A1(new_n1086_), .A2(new_n1142_), .A3(new_n1144_), .ZN(new_n1145_));
  AOI21_X1   g00889(.A1(new_n1141_), .A2(new_n1023_), .B(new_n1077_), .ZN(new_n1146_));
  NAND2_X1   g00890(.A1(new_n1072_), .A2(new_n1066_), .ZN(new_n1147_));
  NOR2_X1    g00891(.A1(new_n1146_), .A2(new_n1147_), .ZN(new_n1148_));
  NAND2_X1   g00892(.A1(new_n1146_), .A2(new_n1147_), .ZN(new_n1149_));
  INV_X1     g00893(.I(new_n1149_), .ZN(new_n1150_));
  NOR2_X1    g00894(.A1(new_n1150_), .A2(new_n1148_), .ZN(new_n1151_));
  INV_X1     g00895(.I(new_n1151_), .ZN(new_n1152_));
  OAI22_X1   g00896(.A1(new_n940_), .A2(new_n393_), .B1(new_n290_), .B2(new_n935_), .ZN(new_n1153_));
  OAI21_X1   g00897(.A1(new_n292_), .A2(new_n1020_), .B(new_n1153_), .ZN(new_n1154_));
  NAND3_X1   g00898(.A1(new_n1154_), .A2(new_n334_), .A3(new_n942_), .ZN(new_n1155_));
  XOR2_X1    g00899(.A1(new_n1155_), .A2(\a[17] ), .Z(new_n1156_));
  INV_X1     g00900(.I(new_n1156_), .ZN(new_n1157_));
  INV_X1     g00901(.I(\a[20] ), .ZN(new_n1158_));
  INV_X1     g00902(.I(\a[19] ), .ZN(new_n1159_));
  NOR3_X1    g00903(.A1(new_n1159_), .A2(\a[17] ), .A3(\a[18] ), .ZN(new_n1160_));
  NAND3_X1   g00904(.A1(new_n1159_), .A2(\a[17] ), .A3(\a[18] ), .ZN(new_n1161_));
  INV_X1     g00905(.I(new_n1161_), .ZN(new_n1162_));
  NOR2_X1    g00906(.A1(new_n1162_), .A2(new_n1160_), .ZN(new_n1163_));
  NOR2_X1    g00907(.A1(new_n1163_), .A2(new_n258_), .ZN(new_n1164_));
  INV_X1     g00908(.I(new_n1065_), .ZN(new_n1165_));
  XNOR2_X1   g00909(.A1(\a[19] ), .A2(\a[20] ), .ZN(new_n1166_));
  NOR2_X1    g00910(.A1(new_n1165_), .A2(new_n1166_), .ZN(new_n1167_));
  INV_X1     g00911(.I(new_n1167_), .ZN(new_n1168_));
  NOR2_X1    g00912(.A1(new_n1168_), .A2(new_n267_), .ZN(new_n1169_));
  NOR2_X1    g00913(.A1(new_n1065_), .A2(new_n1166_), .ZN(new_n1170_));
  INV_X1     g00914(.I(new_n1170_), .ZN(new_n1171_));
  NOR4_X1    g00915(.A1(new_n1169_), .A2(new_n261_), .A3(new_n1164_), .A4(new_n1171_), .ZN(new_n1172_));
  XOR2_X1    g00916(.A1(new_n1172_), .A2(new_n1158_), .Z(new_n1173_));
  NOR2_X1    g00917(.A1(new_n1066_), .A2(new_n1158_), .ZN(new_n1174_));
  XNOR2_X1   g00918(.A1(new_n1173_), .A2(new_n1174_), .ZN(new_n1175_));
  XOR2_X1    g00919(.A1(new_n1175_), .A2(new_n1157_), .Z(new_n1176_));
  OR2_X2     g00920(.A1(new_n1175_), .A2(new_n1157_), .Z(new_n1177_));
  NAND2_X1   g00921(.A1(new_n1175_), .A2(new_n1157_), .ZN(new_n1178_));
  AOI21_X1   g00922(.A1(new_n1177_), .A2(new_n1178_), .B(new_n1152_), .ZN(new_n1179_));
  AOI21_X1   g00923(.A1(new_n1152_), .A2(new_n1176_), .B(new_n1179_), .ZN(new_n1180_));
  OAI22_X1   g00924(.A1(new_n757_), .A2(new_n450_), .B1(new_n403_), .B2(new_n752_), .ZN(new_n1181_));
  INV_X1     g00925(.I(new_n823_), .ZN(new_n1182_));
  NAND2_X1   g00926(.A1(new_n1182_), .A2(\b[5] ), .ZN(new_n1183_));
  AOI21_X1   g00927(.A1(new_n1181_), .A2(new_n1183_), .B(new_n760_), .ZN(new_n1184_));
  NAND2_X1   g00928(.A1(new_n454_), .A2(new_n1184_), .ZN(new_n1185_));
  XOR2_X1    g00929(.A1(new_n1185_), .A2(\a[14] ), .Z(new_n1186_));
  INV_X1     g00930(.I(new_n1186_), .ZN(new_n1187_));
  XOR2_X1    g00931(.A1(new_n1180_), .A2(new_n1187_), .Z(new_n1188_));
  NAND2_X1   g00932(.A1(new_n1145_), .A2(new_n1188_), .ZN(new_n1189_));
  XOR2_X1    g00933(.A1(new_n1180_), .A2(new_n1187_), .Z(new_n1190_));
  OAI21_X1   g00934(.A1(new_n1145_), .A2(new_n1190_), .B(new_n1189_), .ZN(new_n1191_));
  OAI22_X1   g00935(.A1(new_n582_), .A2(new_n617_), .B1(new_n510_), .B2(new_n577_), .ZN(new_n1192_));
  NAND2_X1   g00936(.A1(new_n960_), .A2(\b[8] ), .ZN(new_n1193_));
  AOI21_X1   g00937(.A1(new_n1192_), .A2(new_n1193_), .B(new_n585_), .ZN(new_n1194_));
  NAND2_X1   g00938(.A1(new_n616_), .A2(new_n1194_), .ZN(new_n1195_));
  XOR2_X1    g00939(.A1(new_n1195_), .A2(\a[11] ), .Z(new_n1196_));
  INV_X1     g00940(.I(new_n1196_), .ZN(new_n1197_));
  XOR2_X1    g00941(.A1(new_n1191_), .A2(new_n1197_), .Z(new_n1198_));
  NOR2_X1    g00942(.A1(new_n1198_), .A2(new_n1140_), .ZN(new_n1199_));
  XOR2_X1    g00943(.A1(new_n1191_), .A2(new_n1196_), .Z(new_n1200_));
  NOR2_X1    g00944(.A1(new_n1200_), .A2(new_n1139_), .ZN(new_n1201_));
  NOR2_X1    g00945(.A1(new_n1199_), .A2(new_n1201_), .ZN(new_n1202_));
  OAI22_X1   g00946(.A1(new_n437_), .A2(new_n795_), .B1(new_n717_), .B2(new_n431_), .ZN(new_n1203_));
  NAND2_X1   g00947(.A1(new_n775_), .A2(\b[11] ), .ZN(new_n1204_));
  AOI21_X1   g00948(.A1(new_n1203_), .A2(new_n1204_), .B(new_n440_), .ZN(new_n1205_));
  NAND2_X1   g00949(.A1(new_n799_), .A2(new_n1205_), .ZN(new_n1206_));
  XOR2_X1    g00950(.A1(new_n1206_), .A2(\a[8] ), .Z(new_n1207_));
  XOR2_X1    g00951(.A1(new_n1202_), .A2(new_n1207_), .Z(new_n1208_));
  OAI22_X1   g00952(.A1(new_n364_), .A2(new_n992_), .B1(new_n904_), .B2(new_n320_), .ZN(new_n1209_));
  NAND2_X1   g00953(.A1(new_n594_), .A2(\b[14] ), .ZN(new_n1210_));
  AOI21_X1   g00954(.A1(new_n1209_), .A2(new_n1210_), .B(new_n312_), .ZN(new_n1211_));
  NAND2_X1   g00955(.A1(new_n991_), .A2(new_n1211_), .ZN(new_n1212_));
  XOR2_X1    g00956(.A1(new_n1212_), .A2(\a[5] ), .Z(new_n1213_));
  NOR2_X1    g00957(.A1(new_n1208_), .A2(new_n1213_), .ZN(new_n1214_));
  NAND2_X1   g00958(.A1(new_n1208_), .A2(new_n1213_), .ZN(new_n1215_));
  INV_X1     g00959(.I(new_n1215_), .ZN(new_n1216_));
  NOR2_X1    g00960(.A1(new_n1216_), .A2(new_n1214_), .ZN(new_n1217_));
  INV_X1     g00961(.I(new_n1113_), .ZN(new_n1218_));
  NAND2_X1   g00962(.A1(new_n1108_), .A2(new_n1218_), .ZN(new_n1219_));
  XNOR2_X1   g00963(.A1(new_n1217_), .A2(new_n1219_), .ZN(new_n1220_));
  INV_X1     g00964(.I(new_n1220_), .ZN(new_n1221_));
  INV_X1     g00965(.I(\b[19] ), .ZN(new_n1222_));
  XOR2_X1    g00966(.A1(new_n1118_), .A2(\b[17] ), .Z(new_n1223_));
  NAND2_X1   g00967(.A1(new_n1223_), .A2(new_n1120_), .ZN(new_n1224_));
  XOR2_X1    g00968(.A1(new_n1224_), .A2(new_n1222_), .Z(new_n1225_));
  NAND2_X1   g00969(.A1(new_n283_), .A2(\b[19] ), .ZN(new_n1226_));
  NAND2_X1   g00970(.A1(new_n279_), .A2(\b[17] ), .ZN(new_n1227_));
  AOI21_X1   g00971(.A1(\b[18] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n1228_));
  NAND4_X1   g00972(.A1(new_n1225_), .A2(new_n1226_), .A3(new_n1227_), .A4(new_n1228_), .ZN(new_n1229_));
  XOR2_X1    g00973(.A1(new_n1229_), .A2(new_n271_), .Z(new_n1230_));
  NOR2_X1    g00974(.A1(new_n1220_), .A2(new_n1230_), .ZN(new_n1231_));
  INV_X1     g00975(.I(new_n1231_), .ZN(new_n1232_));
  XOR2_X1    g00976(.A1(new_n1229_), .A2(\a[2] ), .Z(new_n1233_));
  OAI21_X1   g00977(.A1(new_n1221_), .A2(new_n1233_), .B(new_n1232_), .ZN(new_n1234_));
  NAND2_X1   g00978(.A1(new_n1114_), .A2(new_n1129_), .ZN(new_n1235_));
  OAI21_X1   g00979(.A1(new_n1135_), .A2(new_n1131_), .B(new_n1235_), .ZN(new_n1236_));
  XOR2_X1    g00980(.A1(new_n1236_), .A2(new_n1234_), .Z(\f[19] ));
  OAI22_X1   g00981(.A1(new_n940_), .A2(new_n347_), .B1(new_n393_), .B2(new_n935_), .ZN(new_n1238_));
  OAI21_X1   g00982(.A1(new_n290_), .A2(new_n1020_), .B(new_n1238_), .ZN(new_n1239_));
  AOI21_X1   g00983(.A1(new_n352_), .A2(new_n942_), .B(new_n1239_), .ZN(new_n1240_));
  XOR2_X1    g00984(.A1(new_n1240_), .A2(new_n930_), .Z(new_n1241_));
  INV_X1     g00985(.I(new_n1241_), .ZN(new_n1242_));
  OAI22_X1   g00986(.A1(new_n757_), .A2(new_n495_), .B1(new_n450_), .B2(new_n752_), .ZN(new_n1243_));
  NAND2_X1   g00987(.A1(new_n1182_), .A2(\b[6] ), .ZN(new_n1244_));
  AOI21_X1   g00988(.A1(new_n1243_), .A2(new_n1244_), .B(new_n760_), .ZN(new_n1245_));
  NAND2_X1   g00989(.A1(new_n494_), .A2(new_n1245_), .ZN(new_n1246_));
  XOR2_X1    g00990(.A1(new_n1246_), .A2(\a[14] ), .Z(new_n1247_));
  NAND2_X1   g00991(.A1(new_n1152_), .A2(new_n1177_), .ZN(new_n1248_));
  NAND2_X1   g00992(.A1(new_n1248_), .A2(new_n1178_), .ZN(new_n1249_));
  NAND2_X1   g00993(.A1(new_n1173_), .A2(new_n1174_), .ZN(new_n1250_));
  NOR2_X1    g00994(.A1(new_n1171_), .A2(new_n278_), .ZN(new_n1251_));
  XNOR2_X1   g00995(.A1(\a[17] ), .A2(\a[19] ), .ZN(new_n1252_));
  NAND2_X1   g00996(.A1(new_n1065_), .A2(new_n1252_), .ZN(new_n1253_));
  XNOR2_X1   g00997(.A1(\a[17] ), .A2(\a[20] ), .ZN(new_n1254_));
  NAND2_X1   g00998(.A1(new_n1253_), .A2(new_n1254_), .ZN(new_n1255_));
  OAI22_X1   g00999(.A1(new_n1168_), .A2(new_n292_), .B1(new_n267_), .B2(new_n1163_), .ZN(new_n1256_));
  NOR4_X1    g01000(.A1(new_n1256_), .A2(new_n258_), .A3(new_n1251_), .A4(new_n1255_), .ZN(new_n1257_));
  XOR2_X1    g01001(.A1(new_n1257_), .A2(new_n1158_), .Z(new_n1258_));
  XOR2_X1    g01002(.A1(new_n1250_), .A2(new_n1258_), .Z(new_n1259_));
  INV_X1     g01003(.I(new_n1259_), .ZN(new_n1260_));
  XOR2_X1    g01004(.A1(new_n1249_), .A2(new_n1260_), .Z(new_n1261_));
  XOR2_X1    g01005(.A1(new_n1261_), .A2(new_n1247_), .Z(new_n1262_));
  XOR2_X1    g01006(.A1(new_n1262_), .A2(new_n1242_), .Z(new_n1263_));
  INV_X1     g01007(.I(new_n1263_), .ZN(new_n1264_));
  XOR2_X1    g01008(.A1(new_n1145_), .A2(new_n1187_), .Z(new_n1265_));
  NAND2_X1   g01009(.A1(new_n1265_), .A2(new_n1180_), .ZN(new_n1266_));
  XOR2_X1    g01010(.A1(new_n1266_), .A2(new_n1264_), .Z(new_n1267_));
  NAND2_X1   g01011(.A1(new_n1145_), .A2(new_n1187_), .ZN(new_n1268_));
  XNOR2_X1   g01012(.A1(new_n1267_), .A2(new_n1268_), .ZN(new_n1269_));
  OAI22_X1   g01013(.A1(new_n582_), .A2(new_n659_), .B1(new_n617_), .B2(new_n577_), .ZN(new_n1270_));
  NAND2_X1   g01014(.A1(new_n960_), .A2(\b[9] ), .ZN(new_n1271_));
  AOI21_X1   g01015(.A1(new_n1270_), .A2(new_n1271_), .B(new_n585_), .ZN(new_n1272_));
  NAND2_X1   g01016(.A1(new_n663_), .A2(new_n1272_), .ZN(new_n1273_));
  XOR2_X1    g01017(.A1(new_n1273_), .A2(\a[11] ), .Z(new_n1274_));
  XOR2_X1    g01018(.A1(new_n1269_), .A2(new_n1274_), .Z(new_n1275_));
  XOR2_X1    g01019(.A1(new_n1139_), .A2(new_n1196_), .Z(new_n1276_));
  NOR2_X1    g01020(.A1(new_n1276_), .A2(new_n1191_), .ZN(new_n1277_));
  XOR2_X1    g01021(.A1(new_n1275_), .A2(new_n1277_), .Z(new_n1278_));
  NAND2_X1   g01022(.A1(new_n1139_), .A2(new_n1197_), .ZN(new_n1279_));
  XNOR2_X1   g01023(.A1(new_n1278_), .A2(new_n1279_), .ZN(new_n1280_));
  OAI22_X1   g01024(.A1(new_n437_), .A2(new_n848_), .B1(new_n795_), .B2(new_n431_), .ZN(new_n1281_));
  NAND2_X1   g01025(.A1(new_n775_), .A2(\b[12] ), .ZN(new_n1282_));
  AOI21_X1   g01026(.A1(new_n1281_), .A2(new_n1282_), .B(new_n440_), .ZN(new_n1283_));
  NAND2_X1   g01027(.A1(new_n847_), .A2(new_n1283_), .ZN(new_n1284_));
  XOR2_X1    g01028(.A1(new_n1284_), .A2(\a[8] ), .Z(new_n1285_));
  XNOR2_X1   g01029(.A1(new_n1280_), .A2(new_n1285_), .ZN(new_n1286_));
  INV_X1     g01030(.I(new_n1202_), .ZN(new_n1287_));
  NOR2_X1    g01031(.A1(new_n1287_), .A2(new_n1207_), .ZN(new_n1288_));
  XOR2_X1    g01032(.A1(new_n1286_), .A2(new_n1288_), .Z(new_n1289_));
  OAI22_X1   g01033(.A1(new_n364_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n320_), .ZN(new_n1290_));
  NAND2_X1   g01034(.A1(new_n594_), .A2(\b[15] ), .ZN(new_n1291_));
  AOI21_X1   g01035(.A1(new_n1290_), .A2(new_n1291_), .B(new_n312_), .ZN(new_n1292_));
  NAND2_X1   g01036(.A1(new_n1047_), .A2(new_n1292_), .ZN(new_n1293_));
  XOR2_X1    g01037(.A1(new_n1293_), .A2(new_n308_), .Z(new_n1294_));
  XOR2_X1    g01038(.A1(new_n1289_), .A2(new_n1294_), .Z(new_n1295_));
  AOI21_X1   g01039(.A1(\b[17] ), .A2(\b[19] ), .B(\b[18] ), .ZN(new_n1296_));
  NOR2_X1    g01040(.A1(new_n1118_), .A2(new_n1296_), .ZN(new_n1297_));
  AOI21_X1   g01041(.A1(new_n1044_), .A2(new_n1222_), .B(new_n1124_), .ZN(new_n1298_));
  OR2_X2     g01042(.A1(new_n1297_), .A2(new_n1298_), .Z(new_n1299_));
  XNOR2_X1   g01043(.A1(\b[19] ), .A2(\b[20] ), .ZN(new_n1300_));
  INV_X1     g01044(.I(new_n1300_), .ZN(new_n1301_));
  NAND2_X1   g01045(.A1(new_n1299_), .A2(new_n1301_), .ZN(new_n1302_));
  XOR2_X1    g01046(.A1(\b[19] ), .A2(\b[20] ), .Z(new_n1303_));
  OAI21_X1   g01047(.A1(new_n1299_), .A2(new_n1303_), .B(new_n1302_), .ZN(new_n1304_));
  INV_X1     g01048(.I(\b[20] ), .ZN(new_n1305_));
  OAI22_X1   g01049(.A1(new_n405_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n404_), .ZN(new_n1306_));
  NAND2_X1   g01050(.A1(new_n279_), .A2(\b[18] ), .ZN(new_n1307_));
  AOI21_X1   g01051(.A1(new_n1306_), .A2(new_n1307_), .B(new_n264_), .ZN(new_n1308_));
  NAND2_X1   g01052(.A1(new_n1304_), .A2(new_n1308_), .ZN(new_n1309_));
  XOR2_X1    g01053(.A1(new_n1309_), .A2(\a[2] ), .Z(new_n1310_));
  NOR2_X1    g01054(.A1(new_n1108_), .A2(new_n1218_), .ZN(new_n1311_));
  NOR3_X1    g01055(.A1(new_n1311_), .A2(new_n1216_), .A3(new_n1214_), .ZN(new_n1312_));
  XOR2_X1    g01056(.A1(new_n1312_), .A2(new_n1310_), .Z(new_n1313_));
  XOR2_X1    g01057(.A1(new_n1295_), .A2(new_n1313_), .Z(new_n1314_));
  OAI21_X1   g01058(.A1(new_n1236_), .A2(new_n1234_), .B(new_n1232_), .ZN(new_n1315_));
  XOR2_X1    g01059(.A1(new_n1314_), .A2(new_n1315_), .Z(\f[20] ));
  INV_X1     g01060(.I(new_n935_), .ZN(new_n1317_));
  AOI22_X1   g01061(.A1(\b[6] ), .A2(new_n939_), .B1(new_n1317_), .B2(\b[5] ), .ZN(new_n1318_));
  NOR2_X1    g01062(.A1(new_n1020_), .A2(new_n393_), .ZN(new_n1319_));
  OAI21_X1   g01063(.A1(new_n1318_), .A2(new_n1319_), .B(new_n942_), .ZN(new_n1320_));
  NOR2_X1    g01064(.A1(new_n524_), .A2(new_n1320_), .ZN(new_n1321_));
  XOR2_X1    g01065(.A1(new_n1321_), .A2(\a[17] ), .Z(new_n1322_));
  XNOR2_X1   g01066(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n1323_));
  NOR2_X1    g01067(.A1(new_n1323_), .A2(new_n258_), .ZN(new_n1324_));
  INV_X1     g01068(.I(new_n1258_), .ZN(new_n1325_));
  NOR2_X1    g01069(.A1(new_n1325_), .A2(new_n1250_), .ZN(new_n1326_));
  NOR2_X1    g01070(.A1(new_n1255_), .A2(new_n267_), .ZN(new_n1327_));
  OAI22_X1   g01071(.A1(new_n1168_), .A2(new_n290_), .B1(new_n292_), .B2(new_n1163_), .ZN(new_n1328_));
  NOR4_X1    g01072(.A1(new_n1328_), .A2(new_n677_), .A3(new_n1171_), .A4(new_n1327_), .ZN(new_n1329_));
  XOR2_X1    g01073(.A1(new_n1329_), .A2(new_n1158_), .Z(new_n1330_));
  XOR2_X1    g01074(.A1(new_n1326_), .A2(new_n1330_), .Z(new_n1331_));
  XOR2_X1    g01075(.A1(new_n1331_), .A2(new_n1324_), .Z(new_n1332_));
  XOR2_X1    g01076(.A1(new_n1332_), .A2(new_n1322_), .Z(new_n1333_));
  XOR2_X1    g01077(.A1(new_n1151_), .A2(new_n1156_), .Z(new_n1334_));
  INV_X1     g01078(.I(new_n1250_), .ZN(new_n1335_));
  NOR2_X1    g01079(.A1(new_n1335_), .A2(new_n1258_), .ZN(new_n1336_));
  NOR2_X1    g01080(.A1(new_n1336_), .A2(new_n1326_), .ZN(new_n1337_));
  XOR2_X1    g01081(.A1(new_n1337_), .A2(\a[17] ), .Z(new_n1338_));
  OAI21_X1   g01082(.A1(new_n1338_), .A2(new_n1240_), .B(new_n1157_), .ZN(new_n1339_));
  AOI21_X1   g01083(.A1(new_n1240_), .A2(new_n1338_), .B(new_n1339_), .ZN(new_n1340_));
  NAND2_X1   g01084(.A1(new_n1340_), .A2(new_n1152_), .ZN(new_n1341_));
  NAND3_X1   g01085(.A1(new_n1341_), .A2(new_n1175_), .A3(new_n1334_), .ZN(new_n1342_));
  OAI21_X1   g01086(.A1(new_n1242_), .A2(new_n1259_), .B(new_n1342_), .ZN(new_n1343_));
  NAND2_X1   g01087(.A1(new_n1343_), .A2(new_n1333_), .ZN(new_n1344_));
  AOI21_X1   g01088(.A1(new_n1241_), .A2(new_n1260_), .B(new_n1333_), .ZN(new_n1345_));
  NAND2_X1   g01089(.A1(new_n1345_), .A2(new_n1342_), .ZN(new_n1346_));
  NAND2_X1   g01090(.A1(new_n1344_), .A2(new_n1346_), .ZN(new_n1347_));
  OAI22_X1   g01091(.A1(new_n757_), .A2(new_n510_), .B1(new_n495_), .B2(new_n752_), .ZN(new_n1348_));
  NAND2_X1   g01092(.A1(new_n1182_), .A2(\b[7] ), .ZN(new_n1349_));
  AOI21_X1   g01093(.A1(new_n1348_), .A2(new_n1349_), .B(new_n760_), .ZN(new_n1350_));
  NAND2_X1   g01094(.A1(new_n518_), .A2(new_n1350_), .ZN(new_n1351_));
  XOR2_X1    g01095(.A1(new_n1351_), .A2(\a[14] ), .Z(new_n1352_));
  NOR2_X1    g01096(.A1(new_n1264_), .A2(new_n1268_), .ZN(new_n1353_));
  OR2_X2     g01097(.A1(new_n1266_), .A2(new_n1353_), .Z(new_n1354_));
  XOR2_X1    g01098(.A1(new_n1259_), .A2(new_n1241_), .Z(new_n1355_));
  XOR2_X1    g01099(.A1(new_n1249_), .A2(new_n1355_), .Z(new_n1356_));
  NAND2_X1   g01100(.A1(new_n1356_), .A2(new_n1247_), .ZN(new_n1357_));
  NAND2_X1   g01101(.A1(new_n1354_), .A2(new_n1357_), .ZN(new_n1358_));
  XOR2_X1    g01102(.A1(new_n1358_), .A2(new_n1352_), .Z(new_n1359_));
  XOR2_X1    g01103(.A1(new_n1359_), .A2(new_n1347_), .Z(new_n1360_));
  OAI22_X1   g01104(.A1(new_n582_), .A2(new_n717_), .B1(new_n659_), .B2(new_n577_), .ZN(new_n1361_));
  NAND2_X1   g01105(.A1(new_n960_), .A2(\b[10] ), .ZN(new_n1362_));
  AOI21_X1   g01106(.A1(new_n1361_), .A2(new_n1362_), .B(new_n585_), .ZN(new_n1363_));
  NAND2_X1   g01107(.A1(new_n716_), .A2(new_n1363_), .ZN(new_n1364_));
  XOR2_X1    g01108(.A1(new_n1364_), .A2(\a[11] ), .Z(new_n1365_));
  INV_X1     g01109(.I(new_n1275_), .ZN(new_n1366_));
  OAI21_X1   g01110(.A1(new_n1366_), .A2(new_n1279_), .B(new_n1277_), .ZN(new_n1367_));
  INV_X1     g01111(.I(new_n1269_), .ZN(new_n1368_));
  NAND2_X1   g01112(.A1(new_n1368_), .A2(new_n1274_), .ZN(new_n1369_));
  NAND2_X1   g01113(.A1(new_n1367_), .A2(new_n1369_), .ZN(new_n1370_));
  XOR2_X1    g01114(.A1(new_n1370_), .A2(new_n1365_), .Z(new_n1371_));
  XNOR2_X1   g01115(.A1(new_n1371_), .A2(new_n1360_), .ZN(new_n1372_));
  OAI22_X1   g01116(.A1(new_n437_), .A2(new_n904_), .B1(new_n848_), .B2(new_n431_), .ZN(new_n1373_));
  NAND2_X1   g01117(.A1(new_n775_), .A2(\b[13] ), .ZN(new_n1374_));
  AOI21_X1   g01118(.A1(new_n1373_), .A2(new_n1374_), .B(new_n440_), .ZN(new_n1375_));
  NAND2_X1   g01119(.A1(new_n907_), .A2(new_n1375_), .ZN(new_n1376_));
  XOR2_X1    g01120(.A1(new_n1376_), .A2(\a[8] ), .Z(new_n1377_));
  INV_X1     g01121(.I(new_n1280_), .ZN(new_n1378_));
  AOI22_X1   g01122(.A1(new_n1378_), .A2(new_n1285_), .B1(new_n1287_), .B2(new_n1207_), .ZN(new_n1379_));
  NAND2_X1   g01123(.A1(new_n1379_), .A2(new_n1286_), .ZN(new_n1380_));
  XOR2_X1    g01124(.A1(new_n1380_), .A2(new_n1377_), .Z(new_n1381_));
  XNOR2_X1   g01125(.A1(new_n1381_), .A2(new_n1372_), .ZN(new_n1382_));
  INV_X1     g01126(.I(new_n1382_), .ZN(new_n1383_));
  OAI22_X1   g01127(.A1(new_n364_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n320_), .ZN(new_n1384_));
  NAND2_X1   g01128(.A1(new_n594_), .A2(\b[16] ), .ZN(new_n1385_));
  AOI21_X1   g01129(.A1(new_n1384_), .A2(new_n1385_), .B(new_n312_), .ZN(new_n1386_));
  NAND2_X1   g01130(.A1(new_n1123_), .A2(new_n1386_), .ZN(new_n1387_));
  XOR2_X1    g01131(.A1(new_n1387_), .A2(\a[5] ), .Z(new_n1388_));
  NOR2_X1    g01132(.A1(new_n1383_), .A2(new_n1388_), .ZN(new_n1389_));
  NAND2_X1   g01133(.A1(new_n1383_), .A2(new_n1388_), .ZN(new_n1390_));
  INV_X1     g01134(.I(new_n1390_), .ZN(new_n1391_));
  NOR2_X1    g01135(.A1(new_n1391_), .A2(new_n1389_), .ZN(new_n1392_));
  INV_X1     g01136(.I(\b[21] ), .ZN(new_n1393_));
  XOR2_X1    g01137(.A1(new_n1299_), .A2(\b[19] ), .Z(new_n1394_));
  NAND2_X1   g01138(.A1(new_n1394_), .A2(new_n1301_), .ZN(new_n1395_));
  XOR2_X1    g01139(.A1(new_n1395_), .A2(new_n1393_), .Z(new_n1396_));
  NAND2_X1   g01140(.A1(new_n283_), .A2(\b[21] ), .ZN(new_n1397_));
  NAND2_X1   g01141(.A1(new_n279_), .A2(\b[19] ), .ZN(new_n1398_));
  AOI21_X1   g01142(.A1(\b[20] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n1399_));
  NAND4_X1   g01143(.A1(new_n1396_), .A2(new_n1397_), .A3(new_n1398_), .A4(new_n1399_), .ZN(new_n1400_));
  XOR2_X1    g01144(.A1(new_n1400_), .A2(\a[2] ), .Z(new_n1401_));
  INV_X1     g01145(.I(new_n1401_), .ZN(new_n1402_));
  XOR2_X1    g01146(.A1(new_n1392_), .A2(new_n1402_), .Z(new_n1403_));
  INV_X1     g01147(.I(new_n1312_), .ZN(new_n1404_));
  NOR2_X1    g01148(.A1(new_n1295_), .A2(new_n1404_), .ZN(new_n1405_));
  NAND2_X1   g01149(.A1(new_n1295_), .A2(new_n1404_), .ZN(new_n1406_));
  NAND2_X1   g01150(.A1(new_n1406_), .A2(new_n1310_), .ZN(new_n1407_));
  NOR2_X1    g01151(.A1(new_n1407_), .A2(new_n1405_), .ZN(new_n1408_));
  NAND2_X1   g01152(.A1(new_n1314_), .A2(new_n1315_), .ZN(new_n1409_));
  NOR2_X1    g01153(.A1(new_n1409_), .A2(new_n1408_), .ZN(new_n1410_));
  INV_X1     g01154(.I(new_n1410_), .ZN(new_n1411_));
  XOR2_X1    g01155(.A1(new_n1403_), .A2(new_n1411_), .Z(\f[21] ));
  NOR2_X1    g01156(.A1(new_n1392_), .A2(new_n1402_), .ZN(new_n1413_));
  AOI21_X1   g01157(.A1(new_n1403_), .A2(new_n1411_), .B(new_n1413_), .ZN(new_n1414_));
  NAND2_X1   g01158(.A1(new_n1347_), .A2(new_n1352_), .ZN(new_n1415_));
  XNOR2_X1   g01159(.A1(new_n1347_), .A2(new_n1352_), .ZN(new_n1416_));
  NAND3_X1   g01160(.A1(new_n1354_), .A2(new_n1357_), .A3(new_n1416_), .ZN(new_n1417_));
  XOR2_X1    g01161(.A1(new_n1330_), .A2(new_n1324_), .Z(new_n1418_));
  AND2_X2    g01162(.A1(new_n1418_), .A2(new_n1326_), .Z(new_n1419_));
  NOR2_X1    g01163(.A1(new_n1418_), .A2(new_n1326_), .ZN(new_n1420_));
  NOR3_X1    g01164(.A1(new_n1419_), .A2(new_n1420_), .A3(new_n1322_), .ZN(new_n1421_));
  AOI21_X1   g01165(.A1(new_n1418_), .A2(new_n1258_), .B(new_n1335_), .ZN(new_n1422_));
  NAND2_X1   g01166(.A1(new_n1330_), .A2(new_n1324_), .ZN(new_n1423_));
  NOR2_X1    g01167(.A1(new_n1422_), .A2(new_n1423_), .ZN(new_n1424_));
  NAND2_X1   g01168(.A1(new_n1422_), .A2(new_n1423_), .ZN(new_n1425_));
  INV_X1     g01169(.I(new_n1425_), .ZN(new_n1426_));
  NOR2_X1    g01170(.A1(new_n1426_), .A2(new_n1424_), .ZN(new_n1427_));
  INV_X1     g01171(.I(new_n1427_), .ZN(new_n1428_));
  OAI22_X1   g01172(.A1(new_n1168_), .A2(new_n393_), .B1(new_n290_), .B2(new_n1163_), .ZN(new_n1429_));
  OAI21_X1   g01173(.A1(new_n292_), .A2(new_n1255_), .B(new_n1429_), .ZN(new_n1430_));
  NAND3_X1   g01174(.A1(new_n1430_), .A2(new_n334_), .A3(new_n1170_), .ZN(new_n1431_));
  XOR2_X1    g01175(.A1(new_n1431_), .A2(\a[20] ), .Z(new_n1432_));
  INV_X1     g01176(.I(new_n1432_), .ZN(new_n1433_));
  INV_X1     g01177(.I(\a[23] ), .ZN(new_n1434_));
  INV_X1     g01178(.I(\a[22] ), .ZN(new_n1435_));
  NOR3_X1    g01179(.A1(new_n1435_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n1436_));
  NAND3_X1   g01180(.A1(new_n1435_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n1437_));
  INV_X1     g01181(.I(new_n1437_), .ZN(new_n1438_));
  NOR2_X1    g01182(.A1(new_n1438_), .A2(new_n1436_), .ZN(new_n1439_));
  NOR2_X1    g01183(.A1(new_n1439_), .A2(new_n258_), .ZN(new_n1440_));
  INV_X1     g01184(.I(new_n1323_), .ZN(new_n1441_));
  XNOR2_X1   g01185(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n1442_));
  NOR2_X1    g01186(.A1(new_n1441_), .A2(new_n1442_), .ZN(new_n1443_));
  INV_X1     g01187(.I(new_n1443_), .ZN(new_n1444_));
  NOR2_X1    g01188(.A1(new_n1444_), .A2(new_n267_), .ZN(new_n1445_));
  NOR2_X1    g01189(.A1(new_n1323_), .A2(new_n1442_), .ZN(new_n1446_));
  INV_X1     g01190(.I(new_n1446_), .ZN(new_n1447_));
  NOR4_X1    g01191(.A1(new_n1445_), .A2(new_n261_), .A3(new_n1440_), .A4(new_n1447_), .ZN(new_n1448_));
  XOR2_X1    g01192(.A1(new_n1448_), .A2(new_n1434_), .Z(new_n1449_));
  NOR2_X1    g01193(.A1(new_n1324_), .A2(new_n1434_), .ZN(new_n1450_));
  XNOR2_X1   g01194(.A1(new_n1449_), .A2(new_n1450_), .ZN(new_n1451_));
  XOR2_X1    g01195(.A1(new_n1451_), .A2(new_n1433_), .Z(new_n1452_));
  OR2_X2     g01196(.A1(new_n1451_), .A2(new_n1433_), .Z(new_n1453_));
  NAND2_X1   g01197(.A1(new_n1451_), .A2(new_n1433_), .ZN(new_n1454_));
  AOI21_X1   g01198(.A1(new_n1453_), .A2(new_n1454_), .B(new_n1428_), .ZN(new_n1455_));
  AOI21_X1   g01199(.A1(new_n1428_), .A2(new_n1452_), .B(new_n1455_), .ZN(new_n1456_));
  OAI22_X1   g01200(.A1(new_n940_), .A2(new_n450_), .B1(new_n403_), .B2(new_n935_), .ZN(new_n1457_));
  INV_X1     g01201(.I(new_n1020_), .ZN(new_n1458_));
  NAND2_X1   g01202(.A1(new_n1458_), .A2(\b[5] ), .ZN(new_n1459_));
  AOI21_X1   g01203(.A1(new_n1457_), .A2(new_n1459_), .B(new_n943_), .ZN(new_n1460_));
  NAND2_X1   g01204(.A1(new_n454_), .A2(new_n1460_), .ZN(new_n1461_));
  XOR2_X1    g01205(.A1(new_n1461_), .A2(\a[17] ), .Z(new_n1462_));
  XOR2_X1    g01206(.A1(new_n1456_), .A2(new_n1462_), .Z(new_n1463_));
  AOI21_X1   g01207(.A1(new_n1344_), .A2(new_n1421_), .B(new_n1463_), .ZN(new_n1464_));
  NAND2_X1   g01208(.A1(new_n1344_), .A2(new_n1421_), .ZN(new_n1465_));
  INV_X1     g01209(.I(new_n1462_), .ZN(new_n1466_));
  XOR2_X1    g01210(.A1(new_n1456_), .A2(new_n1466_), .Z(new_n1467_));
  NOR2_X1    g01211(.A1(new_n1465_), .A2(new_n1467_), .ZN(new_n1468_));
  NOR2_X1    g01212(.A1(new_n1468_), .A2(new_n1464_), .ZN(new_n1469_));
  OAI22_X1   g01213(.A1(new_n757_), .A2(new_n617_), .B1(new_n510_), .B2(new_n752_), .ZN(new_n1470_));
  NAND2_X1   g01214(.A1(new_n1182_), .A2(\b[8] ), .ZN(new_n1471_));
  AOI21_X1   g01215(.A1(new_n1470_), .A2(new_n1471_), .B(new_n760_), .ZN(new_n1472_));
  NAND2_X1   g01216(.A1(new_n616_), .A2(new_n1472_), .ZN(new_n1473_));
  XOR2_X1    g01217(.A1(new_n1473_), .A2(\a[14] ), .Z(new_n1474_));
  XOR2_X1    g01218(.A1(new_n1469_), .A2(new_n1474_), .Z(new_n1475_));
  AOI21_X1   g01219(.A1(new_n1417_), .A2(new_n1415_), .B(new_n1475_), .ZN(new_n1476_));
  NAND2_X1   g01220(.A1(new_n1417_), .A2(new_n1415_), .ZN(new_n1477_));
  INV_X1     g01221(.I(new_n1474_), .ZN(new_n1478_));
  XOR2_X1    g01222(.A1(new_n1469_), .A2(new_n1478_), .Z(new_n1479_));
  NOR2_X1    g01223(.A1(new_n1477_), .A2(new_n1479_), .ZN(new_n1480_));
  NOR2_X1    g01224(.A1(new_n1480_), .A2(new_n1476_), .ZN(new_n1481_));
  INV_X1     g01225(.I(new_n1481_), .ZN(new_n1482_));
  OAI22_X1   g01226(.A1(new_n582_), .A2(new_n795_), .B1(new_n717_), .B2(new_n577_), .ZN(new_n1483_));
  NAND2_X1   g01227(.A1(new_n960_), .A2(\b[11] ), .ZN(new_n1484_));
  AOI21_X1   g01228(.A1(new_n1483_), .A2(new_n1484_), .B(new_n585_), .ZN(new_n1485_));
  NAND2_X1   g01229(.A1(new_n799_), .A2(new_n1485_), .ZN(new_n1486_));
  XOR2_X1    g01230(.A1(new_n1486_), .A2(\a[11] ), .Z(new_n1487_));
  NOR2_X1    g01231(.A1(new_n1482_), .A2(new_n1487_), .ZN(new_n1488_));
  INV_X1     g01232(.I(new_n1487_), .ZN(new_n1489_));
  NOR2_X1    g01233(.A1(new_n1481_), .A2(new_n1489_), .ZN(new_n1490_));
  NOR2_X1    g01234(.A1(new_n1488_), .A2(new_n1490_), .ZN(new_n1491_));
  OAI22_X1   g01235(.A1(new_n437_), .A2(new_n992_), .B1(new_n904_), .B2(new_n431_), .ZN(new_n1492_));
  NAND2_X1   g01236(.A1(new_n775_), .A2(\b[14] ), .ZN(new_n1493_));
  AOI21_X1   g01237(.A1(new_n1492_), .A2(new_n1493_), .B(new_n440_), .ZN(new_n1494_));
  NAND2_X1   g01238(.A1(new_n991_), .A2(new_n1494_), .ZN(new_n1495_));
  XOR2_X1    g01239(.A1(new_n1495_), .A2(\a[8] ), .Z(new_n1496_));
  XOR2_X1    g01240(.A1(new_n1491_), .A2(new_n1496_), .Z(new_n1497_));
  OAI22_X1   g01241(.A1(new_n364_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n320_), .ZN(new_n1498_));
  NAND2_X1   g01242(.A1(new_n594_), .A2(\b[17] ), .ZN(new_n1499_));
  AOI21_X1   g01243(.A1(new_n1498_), .A2(new_n1499_), .B(new_n312_), .ZN(new_n1500_));
  NAND2_X1   g01244(.A1(new_n1225_), .A2(new_n1500_), .ZN(new_n1501_));
  XOR2_X1    g01245(.A1(new_n1501_), .A2(\a[5] ), .Z(new_n1502_));
  NOR2_X1    g01246(.A1(new_n1497_), .A2(new_n1502_), .ZN(new_n1503_));
  NAND2_X1   g01247(.A1(new_n1497_), .A2(new_n1502_), .ZN(new_n1504_));
  INV_X1     g01248(.I(new_n1504_), .ZN(new_n1505_));
  NOR2_X1    g01249(.A1(new_n1505_), .A2(new_n1503_), .ZN(new_n1506_));
  NOR2_X1    g01250(.A1(new_n1383_), .A2(new_n1388_), .ZN(new_n1507_));
  XOR2_X1    g01251(.A1(new_n1507_), .A2(new_n1506_), .Z(new_n1508_));
  AOI21_X1   g01252(.A1(\b[19] ), .A2(\b[21] ), .B(\b[20] ), .ZN(new_n1509_));
  AOI21_X1   g01253(.A1(new_n1222_), .A2(new_n1393_), .B(new_n1305_), .ZN(new_n1510_));
  INV_X1     g01254(.I(new_n1510_), .ZN(new_n1511_));
  OAI21_X1   g01255(.A1(new_n1299_), .A2(new_n1509_), .B(new_n1511_), .ZN(new_n1512_));
  XNOR2_X1   g01256(.A1(\b[21] ), .A2(\b[22] ), .ZN(new_n1513_));
  INV_X1     g01257(.I(new_n1513_), .ZN(new_n1514_));
  NAND2_X1   g01258(.A1(new_n1512_), .A2(new_n1514_), .ZN(new_n1515_));
  XOR2_X1    g01259(.A1(\b[21] ), .A2(\b[22] ), .Z(new_n1516_));
  OAI21_X1   g01260(.A1(new_n1512_), .A2(new_n1516_), .B(new_n1515_), .ZN(new_n1517_));
  INV_X1     g01261(.I(\b[22] ), .ZN(new_n1518_));
  OAI22_X1   g01262(.A1(new_n405_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n404_), .ZN(new_n1519_));
  NAND2_X1   g01263(.A1(new_n279_), .A2(\b[20] ), .ZN(new_n1520_));
  AOI21_X1   g01264(.A1(new_n1519_), .A2(new_n1520_), .B(new_n264_), .ZN(new_n1521_));
  NAND2_X1   g01265(.A1(new_n1517_), .A2(new_n1521_), .ZN(new_n1522_));
  XOR2_X1    g01266(.A1(new_n1522_), .A2(\a[2] ), .Z(new_n1523_));
  XOR2_X1    g01267(.A1(new_n1508_), .A2(new_n1523_), .Z(new_n1524_));
  INV_X1     g01268(.I(new_n1508_), .ZN(new_n1525_));
  NOR2_X1    g01269(.A1(new_n1525_), .A2(new_n1523_), .ZN(new_n1526_));
  INV_X1     g01270(.I(new_n1523_), .ZN(new_n1527_));
  NOR2_X1    g01271(.A1(new_n1508_), .A2(new_n1527_), .ZN(new_n1528_));
  OAI21_X1   g01272(.A1(new_n1526_), .A2(new_n1528_), .B(new_n1414_), .ZN(new_n1529_));
  OAI21_X1   g01273(.A1(new_n1414_), .A2(new_n1524_), .B(new_n1529_), .ZN(\f[22] ));
  OAI22_X1   g01274(.A1(new_n1168_), .A2(new_n347_), .B1(new_n393_), .B2(new_n1163_), .ZN(new_n1531_));
  OAI21_X1   g01275(.A1(new_n290_), .A2(new_n1255_), .B(new_n1531_), .ZN(new_n1532_));
  AOI21_X1   g01276(.A1(new_n352_), .A2(new_n1170_), .B(new_n1532_), .ZN(new_n1533_));
  XOR2_X1    g01277(.A1(new_n1533_), .A2(new_n1158_), .Z(new_n1534_));
  INV_X1     g01278(.I(new_n1534_), .ZN(new_n1535_));
  OAI22_X1   g01279(.A1(new_n940_), .A2(new_n495_), .B1(new_n450_), .B2(new_n935_), .ZN(new_n1536_));
  NAND2_X1   g01280(.A1(new_n1458_), .A2(\b[6] ), .ZN(new_n1537_));
  AOI21_X1   g01281(.A1(new_n1536_), .A2(new_n1537_), .B(new_n943_), .ZN(new_n1538_));
  NAND2_X1   g01282(.A1(new_n494_), .A2(new_n1538_), .ZN(new_n1539_));
  XOR2_X1    g01283(.A1(new_n1539_), .A2(\a[17] ), .Z(new_n1540_));
  NAND2_X1   g01284(.A1(new_n1428_), .A2(new_n1453_), .ZN(new_n1541_));
  NAND2_X1   g01285(.A1(new_n1541_), .A2(new_n1454_), .ZN(new_n1542_));
  NAND2_X1   g01286(.A1(new_n1449_), .A2(new_n1450_), .ZN(new_n1543_));
  NOR2_X1    g01287(.A1(new_n1447_), .A2(new_n278_), .ZN(new_n1544_));
  XNOR2_X1   g01288(.A1(\a[20] ), .A2(\a[22] ), .ZN(new_n1545_));
  NAND2_X1   g01289(.A1(new_n1323_), .A2(new_n1545_), .ZN(new_n1546_));
  XNOR2_X1   g01290(.A1(\a[20] ), .A2(\a[23] ), .ZN(new_n1547_));
  NAND2_X1   g01291(.A1(new_n1546_), .A2(new_n1547_), .ZN(new_n1548_));
  OAI22_X1   g01292(.A1(new_n1444_), .A2(new_n292_), .B1(new_n267_), .B2(new_n1439_), .ZN(new_n1549_));
  NOR4_X1    g01293(.A1(new_n1549_), .A2(new_n258_), .A3(new_n1544_), .A4(new_n1548_), .ZN(new_n1550_));
  XOR2_X1    g01294(.A1(new_n1550_), .A2(new_n1434_), .Z(new_n1551_));
  XOR2_X1    g01295(.A1(new_n1543_), .A2(new_n1551_), .Z(new_n1552_));
  INV_X1     g01296(.I(new_n1552_), .ZN(new_n1553_));
  XOR2_X1    g01297(.A1(new_n1542_), .A2(new_n1553_), .Z(new_n1554_));
  XOR2_X1    g01298(.A1(new_n1554_), .A2(new_n1540_), .Z(new_n1555_));
  XOR2_X1    g01299(.A1(new_n1555_), .A2(new_n1535_), .Z(new_n1556_));
  INV_X1     g01300(.I(new_n1556_), .ZN(new_n1557_));
  XOR2_X1    g01301(.A1(new_n1465_), .A2(new_n1466_), .Z(new_n1558_));
  NAND2_X1   g01302(.A1(new_n1558_), .A2(new_n1456_), .ZN(new_n1559_));
  XOR2_X1    g01303(.A1(new_n1559_), .A2(new_n1557_), .Z(new_n1560_));
  NAND2_X1   g01304(.A1(new_n1465_), .A2(new_n1466_), .ZN(new_n1561_));
  XNOR2_X1   g01305(.A1(new_n1560_), .A2(new_n1561_), .ZN(new_n1562_));
  OAI22_X1   g01306(.A1(new_n757_), .A2(new_n659_), .B1(new_n617_), .B2(new_n752_), .ZN(new_n1563_));
  NAND2_X1   g01307(.A1(new_n1182_), .A2(\b[9] ), .ZN(new_n1564_));
  AOI21_X1   g01308(.A1(new_n1563_), .A2(new_n1564_), .B(new_n760_), .ZN(new_n1565_));
  NAND2_X1   g01309(.A1(new_n663_), .A2(new_n1565_), .ZN(new_n1566_));
  XOR2_X1    g01310(.A1(new_n1566_), .A2(\a[14] ), .Z(new_n1567_));
  XOR2_X1    g01311(.A1(new_n1562_), .A2(new_n1567_), .Z(new_n1568_));
  XOR2_X1    g01312(.A1(new_n1477_), .A2(new_n1474_), .Z(new_n1569_));
  NOR3_X1    g01313(.A1(new_n1569_), .A2(new_n1464_), .A3(new_n1468_), .ZN(new_n1570_));
  XOR2_X1    g01314(.A1(new_n1570_), .A2(new_n1568_), .Z(new_n1571_));
  NAND2_X1   g01315(.A1(new_n1477_), .A2(new_n1478_), .ZN(new_n1572_));
  XNOR2_X1   g01316(.A1(new_n1571_), .A2(new_n1572_), .ZN(new_n1573_));
  INV_X1     g01317(.I(new_n1573_), .ZN(new_n1574_));
  OAI22_X1   g01318(.A1(new_n582_), .A2(new_n848_), .B1(new_n795_), .B2(new_n577_), .ZN(new_n1575_));
  NAND2_X1   g01319(.A1(new_n960_), .A2(\b[12] ), .ZN(new_n1576_));
  AOI21_X1   g01320(.A1(new_n1575_), .A2(new_n1576_), .B(new_n585_), .ZN(new_n1577_));
  NAND2_X1   g01321(.A1(new_n847_), .A2(new_n1577_), .ZN(new_n1578_));
  XOR2_X1    g01322(.A1(new_n1578_), .A2(\a[11] ), .Z(new_n1579_));
  NOR2_X1    g01323(.A1(new_n1574_), .A2(new_n1579_), .ZN(new_n1580_));
  NAND2_X1   g01324(.A1(new_n1574_), .A2(new_n1579_), .ZN(new_n1581_));
  INV_X1     g01325(.I(new_n1581_), .ZN(new_n1582_));
  NOR2_X1    g01326(.A1(new_n1582_), .A2(new_n1580_), .ZN(new_n1583_));
  NOR2_X1    g01327(.A1(new_n1482_), .A2(new_n1487_), .ZN(new_n1584_));
  XOR2_X1    g01328(.A1(new_n1583_), .A2(new_n1584_), .Z(new_n1585_));
  OAI22_X1   g01329(.A1(new_n437_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n431_), .ZN(new_n1586_));
  NAND2_X1   g01330(.A1(new_n775_), .A2(\b[15] ), .ZN(new_n1587_));
  AOI21_X1   g01331(.A1(new_n1586_), .A2(new_n1587_), .B(new_n440_), .ZN(new_n1588_));
  NAND2_X1   g01332(.A1(new_n1047_), .A2(new_n1588_), .ZN(new_n1589_));
  XOR2_X1    g01333(.A1(new_n1589_), .A2(\a[8] ), .Z(new_n1590_));
  XNOR2_X1   g01334(.A1(new_n1585_), .A2(new_n1590_), .ZN(new_n1591_));
  INV_X1     g01335(.I(new_n1491_), .ZN(new_n1592_));
  NOR2_X1    g01336(.A1(new_n1592_), .A2(new_n1496_), .ZN(new_n1593_));
  XOR2_X1    g01337(.A1(new_n1591_), .A2(new_n1593_), .Z(new_n1594_));
  OAI22_X1   g01338(.A1(new_n364_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n320_), .ZN(new_n1595_));
  NAND2_X1   g01339(.A1(new_n594_), .A2(\b[18] ), .ZN(new_n1596_));
  AOI21_X1   g01340(.A1(new_n1595_), .A2(new_n1596_), .B(new_n312_), .ZN(new_n1597_));
  NAND2_X1   g01341(.A1(new_n1304_), .A2(new_n1597_), .ZN(new_n1598_));
  XOR2_X1    g01342(.A1(new_n1598_), .A2(\a[5] ), .Z(new_n1599_));
  XOR2_X1    g01343(.A1(new_n1594_), .A2(new_n1599_), .Z(new_n1600_));
  INV_X1     g01344(.I(\b[23] ), .ZN(new_n1601_));
  XOR2_X1    g01345(.A1(new_n1512_), .A2(\b[21] ), .Z(new_n1602_));
  NAND2_X1   g01346(.A1(new_n1602_), .A2(new_n1514_), .ZN(new_n1603_));
  XOR2_X1    g01347(.A1(new_n1603_), .A2(new_n1601_), .Z(new_n1604_));
  NAND2_X1   g01348(.A1(new_n283_), .A2(\b[23] ), .ZN(new_n1605_));
  NAND2_X1   g01349(.A1(new_n279_), .A2(\b[21] ), .ZN(new_n1606_));
  AOI21_X1   g01350(.A1(\b[22] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n1607_));
  NAND4_X1   g01351(.A1(new_n1604_), .A2(new_n1605_), .A3(new_n1606_), .A4(new_n1607_), .ZN(new_n1608_));
  XOR2_X1    g01352(.A1(new_n1608_), .A2(\a[2] ), .Z(new_n1609_));
  NOR3_X1    g01353(.A1(new_n1391_), .A2(new_n1503_), .A3(new_n1505_), .ZN(new_n1610_));
  XOR2_X1    g01354(.A1(new_n1610_), .A2(new_n1609_), .Z(new_n1611_));
  XOR2_X1    g01355(.A1(new_n1611_), .A2(new_n1600_), .Z(new_n1612_));
  AOI21_X1   g01356(.A1(new_n1414_), .A2(new_n1525_), .B(new_n1523_), .ZN(new_n1613_));
  XNOR2_X1   g01357(.A1(new_n1612_), .A2(new_n1613_), .ZN(\f[23] ));
  INV_X1     g01358(.I(new_n1599_), .ZN(new_n1615_));
  INV_X1     g01359(.I(new_n1610_), .ZN(new_n1616_));
  XOR2_X1    g01360(.A1(new_n1594_), .A2(new_n1615_), .Z(new_n1617_));
  AOI21_X1   g01361(.A1(new_n1615_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n1618_));
  INV_X1     g01362(.I(new_n1163_), .ZN(new_n1619_));
  AOI22_X1   g01363(.A1(\b[6] ), .A2(new_n1167_), .B1(new_n1619_), .B2(\b[5] ), .ZN(new_n1620_));
  NOR2_X1    g01364(.A1(new_n1255_), .A2(new_n393_), .ZN(new_n1621_));
  OAI21_X1   g01365(.A1(new_n1620_), .A2(new_n1621_), .B(new_n1170_), .ZN(new_n1622_));
  NOR2_X1    g01366(.A1(new_n524_), .A2(new_n1622_), .ZN(new_n1623_));
  XOR2_X1    g01367(.A1(new_n1623_), .A2(\a[20] ), .Z(new_n1624_));
  XNOR2_X1   g01368(.A1(\a[23] ), .A2(\a[24] ), .ZN(new_n1625_));
  NOR2_X1    g01369(.A1(new_n1625_), .A2(new_n258_), .ZN(new_n1626_));
  INV_X1     g01370(.I(new_n1551_), .ZN(new_n1627_));
  NOR2_X1    g01371(.A1(new_n1627_), .A2(new_n1543_), .ZN(new_n1628_));
  NOR2_X1    g01372(.A1(new_n1548_), .A2(new_n267_), .ZN(new_n1629_));
  OAI22_X1   g01373(.A1(new_n1444_), .A2(new_n290_), .B1(new_n292_), .B2(new_n1439_), .ZN(new_n1630_));
  NOR4_X1    g01374(.A1(new_n1630_), .A2(new_n677_), .A3(new_n1447_), .A4(new_n1629_), .ZN(new_n1631_));
  XOR2_X1    g01375(.A1(new_n1631_), .A2(new_n1434_), .Z(new_n1632_));
  XOR2_X1    g01376(.A1(new_n1628_), .A2(new_n1632_), .Z(new_n1633_));
  XOR2_X1    g01377(.A1(new_n1633_), .A2(new_n1626_), .Z(new_n1634_));
  XOR2_X1    g01378(.A1(new_n1634_), .A2(new_n1624_), .Z(new_n1635_));
  XOR2_X1    g01379(.A1(new_n1427_), .A2(new_n1432_), .Z(new_n1636_));
  INV_X1     g01380(.I(new_n1543_), .ZN(new_n1637_));
  NOR2_X1    g01381(.A1(new_n1637_), .A2(new_n1551_), .ZN(new_n1638_));
  NOR2_X1    g01382(.A1(new_n1638_), .A2(new_n1628_), .ZN(new_n1639_));
  XOR2_X1    g01383(.A1(new_n1639_), .A2(\a[20] ), .Z(new_n1640_));
  OAI21_X1   g01384(.A1(new_n1640_), .A2(new_n1533_), .B(new_n1433_), .ZN(new_n1641_));
  AOI21_X1   g01385(.A1(new_n1533_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n1642_));
  NAND2_X1   g01386(.A1(new_n1642_), .A2(new_n1428_), .ZN(new_n1643_));
  NAND3_X1   g01387(.A1(new_n1643_), .A2(new_n1451_), .A3(new_n1636_), .ZN(new_n1644_));
  OAI21_X1   g01388(.A1(new_n1535_), .A2(new_n1552_), .B(new_n1644_), .ZN(new_n1645_));
  NAND2_X1   g01389(.A1(new_n1645_), .A2(new_n1635_), .ZN(new_n1646_));
  AOI21_X1   g01390(.A1(new_n1534_), .A2(new_n1553_), .B(new_n1635_), .ZN(new_n1647_));
  NAND2_X1   g01391(.A1(new_n1647_), .A2(new_n1644_), .ZN(new_n1648_));
  NAND2_X1   g01392(.A1(new_n1646_), .A2(new_n1648_), .ZN(new_n1649_));
  OAI22_X1   g01393(.A1(new_n940_), .A2(new_n510_), .B1(new_n495_), .B2(new_n935_), .ZN(new_n1650_));
  NAND2_X1   g01394(.A1(new_n1458_), .A2(\b[7] ), .ZN(new_n1651_));
  AOI21_X1   g01395(.A1(new_n1650_), .A2(new_n1651_), .B(new_n943_), .ZN(new_n1652_));
  NAND2_X1   g01396(.A1(new_n518_), .A2(new_n1652_), .ZN(new_n1653_));
  XOR2_X1    g01397(.A1(new_n1653_), .A2(\a[17] ), .Z(new_n1654_));
  NOR2_X1    g01398(.A1(new_n1557_), .A2(new_n1561_), .ZN(new_n1655_));
  OR2_X2     g01399(.A1(new_n1655_), .A2(new_n1559_), .Z(new_n1656_));
  XOR2_X1    g01400(.A1(new_n1552_), .A2(new_n1534_), .Z(new_n1657_));
  XOR2_X1    g01401(.A1(new_n1542_), .A2(new_n1657_), .Z(new_n1658_));
  NAND2_X1   g01402(.A1(new_n1658_), .A2(new_n1540_), .ZN(new_n1659_));
  NAND2_X1   g01403(.A1(new_n1656_), .A2(new_n1659_), .ZN(new_n1660_));
  XOR2_X1    g01404(.A1(new_n1660_), .A2(new_n1654_), .Z(new_n1661_));
  XOR2_X1    g01405(.A1(new_n1661_), .A2(new_n1649_), .Z(new_n1662_));
  OAI22_X1   g01406(.A1(new_n757_), .A2(new_n717_), .B1(new_n659_), .B2(new_n752_), .ZN(new_n1663_));
  NAND2_X1   g01407(.A1(new_n1182_), .A2(\b[10] ), .ZN(new_n1664_));
  AOI21_X1   g01408(.A1(new_n1663_), .A2(new_n1664_), .B(new_n760_), .ZN(new_n1665_));
  NAND2_X1   g01409(.A1(new_n716_), .A2(new_n1665_), .ZN(new_n1666_));
  XOR2_X1    g01410(.A1(new_n1666_), .A2(\a[14] ), .Z(new_n1667_));
  INV_X1     g01411(.I(new_n1568_), .ZN(new_n1668_));
  OAI21_X1   g01412(.A1(new_n1668_), .A2(new_n1572_), .B(new_n1570_), .ZN(new_n1669_));
  INV_X1     g01413(.I(new_n1562_), .ZN(new_n1670_));
  NAND2_X1   g01414(.A1(new_n1670_), .A2(new_n1567_), .ZN(new_n1671_));
  NAND2_X1   g01415(.A1(new_n1669_), .A2(new_n1671_), .ZN(new_n1672_));
  XOR2_X1    g01416(.A1(new_n1672_), .A2(new_n1667_), .Z(new_n1673_));
  XOR2_X1    g01417(.A1(new_n1673_), .A2(new_n1662_), .Z(new_n1674_));
  OAI22_X1   g01418(.A1(new_n582_), .A2(new_n904_), .B1(new_n848_), .B2(new_n577_), .ZN(new_n1675_));
  NAND2_X1   g01419(.A1(new_n960_), .A2(\b[13] ), .ZN(new_n1676_));
  AOI21_X1   g01420(.A1(new_n1675_), .A2(new_n1676_), .B(new_n585_), .ZN(new_n1677_));
  NAND2_X1   g01421(.A1(new_n907_), .A2(new_n1677_), .ZN(new_n1678_));
  XOR2_X1    g01422(.A1(new_n1678_), .A2(new_n572_), .Z(new_n1679_));
  NOR3_X1    g01423(.A1(new_n1582_), .A2(new_n1490_), .A3(new_n1580_), .ZN(new_n1680_));
  XOR2_X1    g01424(.A1(new_n1680_), .A2(new_n1679_), .Z(new_n1681_));
  XOR2_X1    g01425(.A1(new_n1681_), .A2(new_n1674_), .Z(new_n1682_));
  OAI22_X1   g01426(.A1(new_n437_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n431_), .ZN(new_n1683_));
  NAND2_X1   g01427(.A1(new_n775_), .A2(\b[16] ), .ZN(new_n1684_));
  AOI21_X1   g01428(.A1(new_n1683_), .A2(new_n1684_), .B(new_n440_), .ZN(new_n1685_));
  NAND2_X1   g01429(.A1(new_n1123_), .A2(new_n1685_), .ZN(new_n1686_));
  XOR2_X1    g01430(.A1(new_n1686_), .A2(\a[8] ), .Z(new_n1687_));
  INV_X1     g01431(.I(new_n1585_), .ZN(new_n1688_));
  AOI22_X1   g01432(.A1(new_n1688_), .A2(new_n1590_), .B1(new_n1592_), .B2(new_n1496_), .ZN(new_n1689_));
  NAND2_X1   g01433(.A1(new_n1689_), .A2(new_n1591_), .ZN(new_n1690_));
  XOR2_X1    g01434(.A1(new_n1690_), .A2(new_n1687_), .Z(new_n1691_));
  XOR2_X1    g01435(.A1(new_n1691_), .A2(new_n1682_), .Z(new_n1692_));
  OAI22_X1   g01436(.A1(new_n364_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n320_), .ZN(new_n1693_));
  NAND2_X1   g01437(.A1(new_n594_), .A2(\b[19] ), .ZN(new_n1694_));
  AOI21_X1   g01438(.A1(new_n1693_), .A2(new_n1694_), .B(new_n312_), .ZN(new_n1695_));
  NAND2_X1   g01439(.A1(new_n1396_), .A2(new_n1695_), .ZN(new_n1696_));
  XOR2_X1    g01440(.A1(new_n1696_), .A2(\a[5] ), .Z(new_n1697_));
  XNOR2_X1   g01441(.A1(new_n1692_), .A2(new_n1697_), .ZN(new_n1698_));
  AOI21_X1   g01442(.A1(\b[21] ), .A2(\b[23] ), .B(\b[22] ), .ZN(new_n1699_));
  NOR2_X1    g01443(.A1(new_n1512_), .A2(new_n1699_), .ZN(new_n1700_));
  AOI21_X1   g01444(.A1(new_n1393_), .A2(new_n1601_), .B(new_n1518_), .ZN(new_n1701_));
  NOR2_X1    g01445(.A1(new_n1700_), .A2(new_n1701_), .ZN(new_n1702_));
  INV_X1     g01446(.I(new_n1702_), .ZN(new_n1703_));
  XNOR2_X1   g01447(.A1(\b[23] ), .A2(\b[24] ), .ZN(new_n1704_));
  INV_X1     g01448(.I(new_n1704_), .ZN(new_n1705_));
  NAND2_X1   g01449(.A1(new_n1703_), .A2(new_n1705_), .ZN(new_n1706_));
  XOR2_X1    g01450(.A1(\b[23] ), .A2(\b[24] ), .Z(new_n1707_));
  OAI21_X1   g01451(.A1(new_n1703_), .A2(new_n1707_), .B(new_n1706_), .ZN(new_n1708_));
  INV_X1     g01452(.I(\b[24] ), .ZN(new_n1709_));
  OAI22_X1   g01453(.A1(new_n405_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n404_), .ZN(new_n1710_));
  NAND2_X1   g01454(.A1(new_n279_), .A2(\b[22] ), .ZN(new_n1711_));
  AOI21_X1   g01455(.A1(new_n1710_), .A2(new_n1711_), .B(new_n264_), .ZN(new_n1712_));
  NAND2_X1   g01456(.A1(new_n1708_), .A2(new_n1712_), .ZN(new_n1713_));
  XOR2_X1    g01457(.A1(new_n1713_), .A2(\a[2] ), .Z(new_n1714_));
  XOR2_X1    g01458(.A1(new_n1698_), .A2(new_n1714_), .Z(new_n1715_));
  NAND2_X1   g01459(.A1(new_n1715_), .A2(new_n1618_), .ZN(new_n1716_));
  XOR2_X1    g01460(.A1(new_n1698_), .A2(new_n1714_), .Z(new_n1717_));
  OAI21_X1   g01461(.A1(new_n1618_), .A2(new_n1717_), .B(new_n1716_), .ZN(new_n1718_));
  INV_X1     g01462(.I(new_n1528_), .ZN(new_n1719_));
  NAND2_X1   g01463(.A1(new_n1414_), .A2(new_n1528_), .ZN(new_n1720_));
  NAND3_X1   g01464(.A1(new_n1612_), .A2(new_n1719_), .A3(new_n1720_), .ZN(new_n1721_));
  NOR2_X1    g01465(.A1(new_n1600_), .A2(new_n1616_), .ZN(new_n1722_));
  NAND2_X1   g01466(.A1(new_n1600_), .A2(new_n1616_), .ZN(new_n1723_));
  NAND2_X1   g01467(.A1(new_n1723_), .A2(new_n1609_), .ZN(new_n1724_));
  NOR3_X1    g01468(.A1(new_n1721_), .A2(new_n1722_), .A3(new_n1724_), .ZN(new_n1725_));
  XOR2_X1    g01469(.A1(new_n1718_), .A2(new_n1725_), .Z(\f[24] ));
  INV_X1     g01470(.I(new_n1714_), .ZN(new_n1727_));
  INV_X1     g01471(.I(new_n1618_), .ZN(new_n1728_));
  XOR2_X1    g01472(.A1(new_n1698_), .A2(new_n1728_), .Z(new_n1729_));
  OAI22_X1   g01473(.A1(new_n1718_), .A2(new_n1725_), .B1(new_n1727_), .B2(new_n1729_), .ZN(new_n1730_));
  NAND2_X1   g01474(.A1(new_n1649_), .A2(new_n1654_), .ZN(new_n1731_));
  XNOR2_X1   g01475(.A1(new_n1649_), .A2(new_n1654_), .ZN(new_n1732_));
  NAND3_X1   g01476(.A1(new_n1656_), .A2(new_n1659_), .A3(new_n1732_), .ZN(new_n1733_));
  XOR2_X1    g01477(.A1(new_n1632_), .A2(new_n1626_), .Z(new_n1734_));
  AND2_X2    g01478(.A1(new_n1734_), .A2(new_n1628_), .Z(new_n1735_));
  NOR2_X1    g01479(.A1(new_n1734_), .A2(new_n1628_), .ZN(new_n1736_));
  NOR3_X1    g01480(.A1(new_n1735_), .A2(new_n1736_), .A3(new_n1624_), .ZN(new_n1737_));
  AOI21_X1   g01481(.A1(new_n1734_), .A2(new_n1551_), .B(new_n1637_), .ZN(new_n1738_));
  NAND2_X1   g01482(.A1(new_n1632_), .A2(new_n1626_), .ZN(new_n1739_));
  NOR2_X1    g01483(.A1(new_n1738_), .A2(new_n1739_), .ZN(new_n1740_));
  NAND2_X1   g01484(.A1(new_n1738_), .A2(new_n1739_), .ZN(new_n1741_));
  INV_X1     g01485(.I(new_n1741_), .ZN(new_n1742_));
  NOR2_X1    g01486(.A1(new_n1742_), .A2(new_n1740_), .ZN(new_n1743_));
  INV_X1     g01487(.I(new_n1743_), .ZN(new_n1744_));
  OAI22_X1   g01488(.A1(new_n1444_), .A2(new_n393_), .B1(new_n290_), .B2(new_n1439_), .ZN(new_n1745_));
  OAI21_X1   g01489(.A1(new_n292_), .A2(new_n1548_), .B(new_n1745_), .ZN(new_n1746_));
  NAND3_X1   g01490(.A1(new_n1746_), .A2(new_n334_), .A3(new_n1446_), .ZN(new_n1747_));
  XOR2_X1    g01491(.A1(new_n1747_), .A2(\a[23] ), .Z(new_n1748_));
  INV_X1     g01492(.I(new_n1748_), .ZN(new_n1749_));
  INV_X1     g01493(.I(\a[26] ), .ZN(new_n1750_));
  INV_X1     g01494(.I(\a[25] ), .ZN(new_n1751_));
  NOR3_X1    g01495(.A1(new_n1751_), .A2(\a[23] ), .A3(\a[24] ), .ZN(new_n1752_));
  NAND3_X1   g01496(.A1(new_n1751_), .A2(\a[23] ), .A3(\a[24] ), .ZN(new_n1753_));
  INV_X1     g01497(.I(new_n1753_), .ZN(new_n1754_));
  NOR2_X1    g01498(.A1(new_n1754_), .A2(new_n1752_), .ZN(new_n1755_));
  NOR2_X1    g01499(.A1(new_n1755_), .A2(new_n258_), .ZN(new_n1756_));
  INV_X1     g01500(.I(new_n1625_), .ZN(new_n1757_));
  XNOR2_X1   g01501(.A1(\a[25] ), .A2(\a[26] ), .ZN(new_n1758_));
  NOR2_X1    g01502(.A1(new_n1757_), .A2(new_n1758_), .ZN(new_n1759_));
  INV_X1     g01503(.I(new_n1759_), .ZN(new_n1760_));
  NOR2_X1    g01504(.A1(new_n1760_), .A2(new_n267_), .ZN(new_n1761_));
  NOR2_X1    g01505(.A1(new_n1625_), .A2(new_n1758_), .ZN(new_n1762_));
  INV_X1     g01506(.I(new_n1762_), .ZN(new_n1763_));
  NOR4_X1    g01507(.A1(new_n1761_), .A2(new_n261_), .A3(new_n1756_), .A4(new_n1763_), .ZN(new_n1764_));
  XOR2_X1    g01508(.A1(new_n1764_), .A2(new_n1750_), .Z(new_n1765_));
  NOR2_X1    g01509(.A1(new_n1626_), .A2(new_n1750_), .ZN(new_n1766_));
  XNOR2_X1   g01510(.A1(new_n1765_), .A2(new_n1766_), .ZN(new_n1767_));
  XOR2_X1    g01511(.A1(new_n1767_), .A2(new_n1749_), .Z(new_n1768_));
  OR2_X2     g01512(.A1(new_n1767_), .A2(new_n1749_), .Z(new_n1769_));
  NAND2_X1   g01513(.A1(new_n1767_), .A2(new_n1749_), .ZN(new_n1770_));
  AOI21_X1   g01514(.A1(new_n1769_), .A2(new_n1770_), .B(new_n1744_), .ZN(new_n1771_));
  AOI21_X1   g01515(.A1(new_n1744_), .A2(new_n1768_), .B(new_n1771_), .ZN(new_n1772_));
  OAI22_X1   g01516(.A1(new_n1168_), .A2(new_n450_), .B1(new_n403_), .B2(new_n1163_), .ZN(new_n1773_));
  INV_X1     g01517(.I(new_n1255_), .ZN(new_n1774_));
  NAND2_X1   g01518(.A1(new_n1774_), .A2(\b[5] ), .ZN(new_n1775_));
  AOI21_X1   g01519(.A1(new_n1773_), .A2(new_n1775_), .B(new_n1171_), .ZN(new_n1776_));
  NAND2_X1   g01520(.A1(new_n454_), .A2(new_n1776_), .ZN(new_n1777_));
  XOR2_X1    g01521(.A1(new_n1777_), .A2(\a[20] ), .Z(new_n1778_));
  XOR2_X1    g01522(.A1(new_n1772_), .A2(new_n1778_), .Z(new_n1779_));
  AOI21_X1   g01523(.A1(new_n1646_), .A2(new_n1737_), .B(new_n1779_), .ZN(new_n1780_));
  NAND2_X1   g01524(.A1(new_n1646_), .A2(new_n1737_), .ZN(new_n1781_));
  INV_X1     g01525(.I(new_n1778_), .ZN(new_n1782_));
  XOR2_X1    g01526(.A1(new_n1772_), .A2(new_n1782_), .Z(new_n1783_));
  NOR2_X1    g01527(.A1(new_n1781_), .A2(new_n1783_), .ZN(new_n1784_));
  NOR2_X1    g01528(.A1(new_n1784_), .A2(new_n1780_), .ZN(new_n1785_));
  OAI22_X1   g01529(.A1(new_n940_), .A2(new_n617_), .B1(new_n510_), .B2(new_n935_), .ZN(new_n1786_));
  NAND2_X1   g01530(.A1(new_n1458_), .A2(\b[8] ), .ZN(new_n1787_));
  AOI21_X1   g01531(.A1(new_n1786_), .A2(new_n1787_), .B(new_n943_), .ZN(new_n1788_));
  NAND2_X1   g01532(.A1(new_n616_), .A2(new_n1788_), .ZN(new_n1789_));
  XOR2_X1    g01533(.A1(new_n1789_), .A2(\a[17] ), .Z(new_n1790_));
  XOR2_X1    g01534(.A1(new_n1785_), .A2(new_n1790_), .Z(new_n1791_));
  AOI21_X1   g01535(.A1(new_n1733_), .A2(new_n1731_), .B(new_n1791_), .ZN(new_n1792_));
  NAND2_X1   g01536(.A1(new_n1733_), .A2(new_n1731_), .ZN(new_n1793_));
  INV_X1     g01537(.I(new_n1790_), .ZN(new_n1794_));
  XOR2_X1    g01538(.A1(new_n1785_), .A2(new_n1794_), .Z(new_n1795_));
  NOR2_X1    g01539(.A1(new_n1793_), .A2(new_n1795_), .ZN(new_n1796_));
  NOR2_X1    g01540(.A1(new_n1796_), .A2(new_n1792_), .ZN(new_n1797_));
  OAI22_X1   g01541(.A1(new_n757_), .A2(new_n795_), .B1(new_n717_), .B2(new_n752_), .ZN(new_n1798_));
  NAND2_X1   g01542(.A1(new_n1182_), .A2(\b[11] ), .ZN(new_n1799_));
  AOI21_X1   g01543(.A1(new_n1798_), .A2(new_n1799_), .B(new_n760_), .ZN(new_n1800_));
  NAND2_X1   g01544(.A1(new_n799_), .A2(new_n1800_), .ZN(new_n1801_));
  XOR2_X1    g01545(.A1(new_n1801_), .A2(\a[14] ), .Z(new_n1802_));
  XOR2_X1    g01546(.A1(new_n1797_), .A2(new_n1802_), .Z(new_n1803_));
  OAI22_X1   g01547(.A1(new_n582_), .A2(new_n992_), .B1(new_n904_), .B2(new_n577_), .ZN(new_n1804_));
  NAND2_X1   g01548(.A1(new_n960_), .A2(\b[14] ), .ZN(new_n1805_));
  AOI21_X1   g01549(.A1(new_n1804_), .A2(new_n1805_), .B(new_n585_), .ZN(new_n1806_));
  NAND2_X1   g01550(.A1(new_n991_), .A2(new_n1806_), .ZN(new_n1807_));
  XOR2_X1    g01551(.A1(new_n1807_), .A2(\a[11] ), .Z(new_n1808_));
  XOR2_X1    g01552(.A1(new_n1803_), .A2(new_n1808_), .Z(new_n1809_));
  OAI22_X1   g01553(.A1(new_n437_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n431_), .ZN(new_n1810_));
  NAND2_X1   g01554(.A1(new_n775_), .A2(\b[17] ), .ZN(new_n1811_));
  AOI21_X1   g01555(.A1(new_n1810_), .A2(new_n1811_), .B(new_n440_), .ZN(new_n1812_));
  NAND2_X1   g01556(.A1(new_n1225_), .A2(new_n1812_), .ZN(new_n1813_));
  XOR2_X1    g01557(.A1(new_n1813_), .A2(\a[8] ), .Z(new_n1814_));
  INV_X1     g01558(.I(new_n1814_), .ZN(new_n1815_));
  XOR2_X1    g01559(.A1(new_n1809_), .A2(new_n1815_), .Z(new_n1816_));
  OAI22_X1   g01560(.A1(new_n364_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n320_), .ZN(new_n1817_));
  NAND2_X1   g01561(.A1(new_n594_), .A2(\b[20] ), .ZN(new_n1818_));
  AOI21_X1   g01562(.A1(new_n1817_), .A2(new_n1818_), .B(new_n312_), .ZN(new_n1819_));
  NAND2_X1   g01563(.A1(new_n1517_), .A2(new_n1819_), .ZN(new_n1820_));
  XOR2_X1    g01564(.A1(new_n1820_), .A2(\a[5] ), .Z(new_n1821_));
  XNOR2_X1   g01565(.A1(new_n1816_), .A2(new_n1821_), .ZN(new_n1822_));
  AOI21_X1   g01566(.A1(new_n1728_), .A2(new_n1692_), .B(new_n1697_), .ZN(new_n1823_));
  XOR2_X1    g01567(.A1(new_n1823_), .A2(new_n1822_), .Z(new_n1824_));
  INV_X1     g01568(.I(\b[25] ), .ZN(new_n1825_));
  XOR2_X1    g01569(.A1(new_n1702_), .A2(new_n1601_), .Z(new_n1826_));
  NAND2_X1   g01570(.A1(new_n1826_), .A2(new_n1705_), .ZN(new_n1827_));
  XOR2_X1    g01571(.A1(new_n1827_), .A2(new_n1825_), .Z(new_n1828_));
  OAI22_X1   g01572(.A1(new_n405_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n404_), .ZN(new_n1829_));
  NAND2_X1   g01573(.A1(new_n279_), .A2(\b[23] ), .ZN(new_n1830_));
  AOI21_X1   g01574(.A1(new_n1829_), .A2(new_n1830_), .B(new_n264_), .ZN(new_n1831_));
  NAND2_X1   g01575(.A1(new_n1828_), .A2(new_n1831_), .ZN(new_n1832_));
  XOR2_X1    g01576(.A1(new_n1832_), .A2(\a[2] ), .Z(new_n1833_));
  INV_X1     g01577(.I(new_n1833_), .ZN(new_n1834_));
  XOR2_X1    g01578(.A1(new_n1824_), .A2(new_n1834_), .Z(new_n1835_));
  NAND2_X1   g01579(.A1(new_n1730_), .A2(new_n1835_), .ZN(new_n1836_));
  XOR2_X1    g01580(.A1(new_n1824_), .A2(new_n1834_), .Z(new_n1837_));
  OAI21_X1   g01581(.A1(new_n1730_), .A2(new_n1837_), .B(new_n1836_), .ZN(\f[25] ));
  INV_X1     g01582(.I(new_n1797_), .ZN(new_n1839_));
  OAI22_X1   g01583(.A1(new_n1444_), .A2(new_n347_), .B1(new_n393_), .B2(new_n1439_), .ZN(new_n1840_));
  OAI21_X1   g01584(.A1(new_n290_), .A2(new_n1548_), .B(new_n1840_), .ZN(new_n1841_));
  AOI21_X1   g01585(.A1(new_n352_), .A2(new_n1446_), .B(new_n1841_), .ZN(new_n1842_));
  XOR2_X1    g01586(.A1(new_n1842_), .A2(new_n1434_), .Z(new_n1843_));
  INV_X1     g01587(.I(new_n1843_), .ZN(new_n1844_));
  OAI22_X1   g01588(.A1(new_n1168_), .A2(new_n495_), .B1(new_n450_), .B2(new_n1163_), .ZN(new_n1845_));
  NAND2_X1   g01589(.A1(new_n1774_), .A2(\b[6] ), .ZN(new_n1846_));
  AOI21_X1   g01590(.A1(new_n1845_), .A2(new_n1846_), .B(new_n1171_), .ZN(new_n1847_));
  NAND2_X1   g01591(.A1(new_n494_), .A2(new_n1847_), .ZN(new_n1848_));
  XOR2_X1    g01592(.A1(new_n1848_), .A2(\a[20] ), .Z(new_n1849_));
  NAND2_X1   g01593(.A1(new_n1744_), .A2(new_n1769_), .ZN(new_n1850_));
  NAND2_X1   g01594(.A1(new_n1850_), .A2(new_n1770_), .ZN(new_n1851_));
  NAND2_X1   g01595(.A1(new_n1765_), .A2(new_n1766_), .ZN(new_n1852_));
  NOR2_X1    g01596(.A1(new_n1763_), .A2(new_n278_), .ZN(new_n1853_));
  XNOR2_X1   g01597(.A1(\a[23] ), .A2(\a[25] ), .ZN(new_n1854_));
  NAND2_X1   g01598(.A1(new_n1625_), .A2(new_n1854_), .ZN(new_n1855_));
  XNOR2_X1   g01599(.A1(\a[23] ), .A2(\a[26] ), .ZN(new_n1856_));
  NAND2_X1   g01600(.A1(new_n1855_), .A2(new_n1856_), .ZN(new_n1857_));
  OAI22_X1   g01601(.A1(new_n1760_), .A2(new_n292_), .B1(new_n267_), .B2(new_n1755_), .ZN(new_n1858_));
  NOR4_X1    g01602(.A1(new_n1858_), .A2(new_n258_), .A3(new_n1853_), .A4(new_n1857_), .ZN(new_n1859_));
  XOR2_X1    g01603(.A1(new_n1859_), .A2(new_n1750_), .Z(new_n1860_));
  XOR2_X1    g01604(.A1(new_n1852_), .A2(new_n1860_), .Z(new_n1861_));
  INV_X1     g01605(.I(new_n1861_), .ZN(new_n1862_));
  XOR2_X1    g01606(.A1(new_n1851_), .A2(new_n1862_), .Z(new_n1863_));
  XOR2_X1    g01607(.A1(new_n1863_), .A2(new_n1849_), .Z(new_n1864_));
  XOR2_X1    g01608(.A1(new_n1864_), .A2(new_n1844_), .Z(new_n1865_));
  INV_X1     g01609(.I(new_n1865_), .ZN(new_n1866_));
  XOR2_X1    g01610(.A1(new_n1781_), .A2(new_n1782_), .Z(new_n1867_));
  NAND2_X1   g01611(.A1(new_n1867_), .A2(new_n1772_), .ZN(new_n1868_));
  XOR2_X1    g01612(.A1(new_n1868_), .A2(new_n1866_), .Z(new_n1869_));
  NAND2_X1   g01613(.A1(new_n1781_), .A2(new_n1782_), .ZN(new_n1870_));
  XNOR2_X1   g01614(.A1(new_n1869_), .A2(new_n1870_), .ZN(new_n1871_));
  OAI22_X1   g01615(.A1(new_n940_), .A2(new_n659_), .B1(new_n617_), .B2(new_n935_), .ZN(new_n1872_));
  NAND2_X1   g01616(.A1(new_n1458_), .A2(\b[9] ), .ZN(new_n1873_));
  AOI21_X1   g01617(.A1(new_n1872_), .A2(new_n1873_), .B(new_n943_), .ZN(new_n1874_));
  NAND2_X1   g01618(.A1(new_n663_), .A2(new_n1874_), .ZN(new_n1875_));
  XOR2_X1    g01619(.A1(new_n1875_), .A2(\a[17] ), .Z(new_n1876_));
  XOR2_X1    g01620(.A1(new_n1871_), .A2(new_n1876_), .Z(new_n1877_));
  XOR2_X1    g01621(.A1(new_n1793_), .A2(new_n1790_), .Z(new_n1878_));
  NOR3_X1    g01622(.A1(new_n1878_), .A2(new_n1780_), .A3(new_n1784_), .ZN(new_n1879_));
  XOR2_X1    g01623(.A1(new_n1879_), .A2(new_n1877_), .Z(new_n1880_));
  NAND2_X1   g01624(.A1(new_n1793_), .A2(new_n1794_), .ZN(new_n1881_));
  XNOR2_X1   g01625(.A1(new_n1880_), .A2(new_n1881_), .ZN(new_n1882_));
  OAI22_X1   g01626(.A1(new_n757_), .A2(new_n848_), .B1(new_n795_), .B2(new_n752_), .ZN(new_n1883_));
  NAND2_X1   g01627(.A1(new_n1182_), .A2(\b[12] ), .ZN(new_n1884_));
  AOI21_X1   g01628(.A1(new_n1883_), .A2(new_n1884_), .B(new_n760_), .ZN(new_n1885_));
  NAND2_X1   g01629(.A1(new_n847_), .A2(new_n1885_), .ZN(new_n1886_));
  XOR2_X1    g01630(.A1(new_n1886_), .A2(\a[14] ), .Z(new_n1887_));
  XNOR2_X1   g01631(.A1(new_n1882_), .A2(new_n1887_), .ZN(new_n1888_));
  OAI22_X1   g01632(.A1(new_n582_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n577_), .ZN(new_n1889_));
  NAND2_X1   g01633(.A1(new_n960_), .A2(\b[15] ), .ZN(new_n1890_));
  AOI21_X1   g01634(.A1(new_n1889_), .A2(new_n1890_), .B(new_n585_), .ZN(new_n1891_));
  NAND2_X1   g01635(.A1(new_n1047_), .A2(new_n1891_), .ZN(new_n1892_));
  XOR2_X1    g01636(.A1(new_n1892_), .A2(\a[11] ), .Z(new_n1893_));
  INV_X1     g01637(.I(new_n1893_), .ZN(new_n1894_));
  XOR2_X1    g01638(.A1(new_n1888_), .A2(new_n1894_), .Z(new_n1895_));
  NOR3_X1    g01639(.A1(new_n1895_), .A2(new_n1839_), .A3(new_n1802_), .ZN(new_n1896_));
  NOR2_X1    g01640(.A1(new_n1839_), .A2(new_n1802_), .ZN(new_n1897_));
  XOR2_X1    g01641(.A1(new_n1888_), .A2(new_n1893_), .Z(new_n1898_));
  NOR2_X1    g01642(.A1(new_n1898_), .A2(new_n1897_), .ZN(new_n1899_));
  NOR2_X1    g01643(.A1(new_n1896_), .A2(new_n1899_), .ZN(new_n1900_));
  NOR2_X1    g01644(.A1(new_n1803_), .A2(new_n1808_), .ZN(new_n1901_));
  XOR2_X1    g01645(.A1(new_n1900_), .A2(new_n1901_), .Z(new_n1902_));
  OAI22_X1   g01646(.A1(new_n437_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n431_), .ZN(new_n1903_));
  NAND2_X1   g01647(.A1(new_n775_), .A2(\b[18] ), .ZN(new_n1904_));
  AOI21_X1   g01648(.A1(new_n1903_), .A2(new_n1904_), .B(new_n440_), .ZN(new_n1905_));
  NAND2_X1   g01649(.A1(new_n1304_), .A2(new_n1905_), .ZN(new_n1906_));
  XOR2_X1    g01650(.A1(new_n1906_), .A2(\a[8] ), .Z(new_n1907_));
  XNOR2_X1   g01651(.A1(new_n1902_), .A2(new_n1907_), .ZN(new_n1908_));
  NAND2_X1   g01652(.A1(new_n1809_), .A2(new_n1815_), .ZN(new_n1909_));
  XNOR2_X1   g01653(.A1(new_n1908_), .A2(new_n1909_), .ZN(new_n1910_));
  OAI22_X1   g01654(.A1(new_n364_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n320_), .ZN(new_n1911_));
  NAND2_X1   g01655(.A1(new_n594_), .A2(\b[21] ), .ZN(new_n1912_));
  AOI21_X1   g01656(.A1(new_n1911_), .A2(new_n1912_), .B(new_n312_), .ZN(new_n1913_));
  NAND2_X1   g01657(.A1(new_n1604_), .A2(new_n1913_), .ZN(new_n1914_));
  XOR2_X1    g01658(.A1(new_n1914_), .A2(\a[5] ), .Z(new_n1915_));
  XNOR2_X1   g01659(.A1(new_n1910_), .A2(new_n1915_), .ZN(new_n1916_));
  INV_X1     g01660(.I(new_n1916_), .ZN(new_n1917_));
  AOI21_X1   g01661(.A1(\b[23] ), .A2(\b[25] ), .B(\b[24] ), .ZN(new_n1918_));
  AOI21_X1   g01662(.A1(new_n1601_), .A2(new_n1825_), .B(new_n1709_), .ZN(new_n1919_));
  INV_X1     g01663(.I(new_n1919_), .ZN(new_n1920_));
  OAI21_X1   g01664(.A1(new_n1703_), .A2(new_n1918_), .B(new_n1920_), .ZN(new_n1921_));
  XNOR2_X1   g01665(.A1(\b[25] ), .A2(\b[26] ), .ZN(new_n1922_));
  INV_X1     g01666(.I(new_n1922_), .ZN(new_n1923_));
  NAND2_X1   g01667(.A1(new_n1921_), .A2(new_n1923_), .ZN(new_n1924_));
  XOR2_X1    g01668(.A1(\b[25] ), .A2(\b[26] ), .Z(new_n1925_));
  OAI21_X1   g01669(.A1(new_n1921_), .A2(new_n1925_), .B(new_n1924_), .ZN(new_n1926_));
  INV_X1     g01670(.I(\b[26] ), .ZN(new_n1927_));
  OAI22_X1   g01671(.A1(new_n405_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n404_), .ZN(new_n1928_));
  NAND2_X1   g01672(.A1(new_n279_), .A2(\b[24] ), .ZN(new_n1929_));
  AOI21_X1   g01673(.A1(new_n1928_), .A2(new_n1929_), .B(new_n264_), .ZN(new_n1930_));
  NAND2_X1   g01674(.A1(new_n1926_), .A2(new_n1930_), .ZN(new_n1931_));
  XOR2_X1    g01675(.A1(new_n1931_), .A2(new_n271_), .Z(new_n1932_));
  NAND2_X1   g01676(.A1(new_n1692_), .A2(new_n1697_), .ZN(new_n1933_));
  NOR2_X1    g01677(.A1(new_n1933_), .A2(new_n1618_), .ZN(new_n1934_));
  INV_X1     g01678(.I(new_n1816_), .ZN(new_n1935_));
  NAND2_X1   g01679(.A1(new_n1935_), .A2(new_n1821_), .ZN(new_n1936_));
  NAND3_X1   g01680(.A1(new_n1933_), .A2(new_n1936_), .A3(new_n1822_), .ZN(new_n1937_));
  NOR2_X1    g01681(.A1(new_n1937_), .A2(new_n1934_), .ZN(new_n1938_));
  XOR2_X1    g01682(.A1(new_n1938_), .A2(new_n1932_), .Z(new_n1939_));
  XOR2_X1    g01683(.A1(new_n1939_), .A2(new_n1917_), .Z(new_n1940_));
  INV_X1     g01684(.I(new_n1940_), .ZN(new_n1941_));
  XOR2_X1    g01685(.A1(new_n1730_), .A2(new_n1834_), .Z(new_n1942_));
  NAND2_X1   g01686(.A1(new_n1942_), .A2(new_n1824_), .ZN(new_n1943_));
  XOR2_X1    g01687(.A1(new_n1943_), .A2(new_n1941_), .Z(new_n1944_));
  NAND2_X1   g01688(.A1(new_n1730_), .A2(new_n1834_), .ZN(new_n1945_));
  XOR2_X1    g01689(.A1(new_n1944_), .A2(new_n1945_), .Z(\f[26] ));
  INV_X1     g01690(.I(new_n1439_), .ZN(new_n1947_));
  AOI22_X1   g01691(.A1(\b[6] ), .A2(new_n1443_), .B1(new_n1947_), .B2(\b[5] ), .ZN(new_n1948_));
  NOR2_X1    g01692(.A1(new_n1548_), .A2(new_n393_), .ZN(new_n1949_));
  OAI21_X1   g01693(.A1(new_n1948_), .A2(new_n1949_), .B(new_n1446_), .ZN(new_n1950_));
  NOR2_X1    g01694(.A1(new_n524_), .A2(new_n1950_), .ZN(new_n1951_));
  XOR2_X1    g01695(.A1(new_n1951_), .A2(\a[23] ), .Z(new_n1952_));
  XNOR2_X1   g01696(.A1(\a[26] ), .A2(\a[27] ), .ZN(new_n1953_));
  NOR2_X1    g01697(.A1(new_n1953_), .A2(new_n258_), .ZN(new_n1954_));
  INV_X1     g01698(.I(new_n1860_), .ZN(new_n1955_));
  NOR2_X1    g01699(.A1(new_n1955_), .A2(new_n1852_), .ZN(new_n1956_));
  NOR2_X1    g01700(.A1(new_n1857_), .A2(new_n267_), .ZN(new_n1957_));
  OAI22_X1   g01701(.A1(new_n1760_), .A2(new_n290_), .B1(new_n292_), .B2(new_n1755_), .ZN(new_n1958_));
  NOR4_X1    g01702(.A1(new_n1958_), .A2(new_n677_), .A3(new_n1763_), .A4(new_n1957_), .ZN(new_n1959_));
  XOR2_X1    g01703(.A1(new_n1959_), .A2(new_n1750_), .Z(new_n1960_));
  XOR2_X1    g01704(.A1(new_n1956_), .A2(new_n1960_), .Z(new_n1961_));
  XOR2_X1    g01705(.A1(new_n1961_), .A2(new_n1954_), .Z(new_n1962_));
  XOR2_X1    g01706(.A1(new_n1962_), .A2(new_n1952_), .Z(new_n1963_));
  XOR2_X1    g01707(.A1(new_n1743_), .A2(new_n1748_), .Z(new_n1964_));
  INV_X1     g01708(.I(new_n1852_), .ZN(new_n1965_));
  NOR2_X1    g01709(.A1(new_n1965_), .A2(new_n1860_), .ZN(new_n1966_));
  NOR2_X1    g01710(.A1(new_n1966_), .A2(new_n1956_), .ZN(new_n1967_));
  XOR2_X1    g01711(.A1(new_n1967_), .A2(\a[23] ), .Z(new_n1968_));
  OAI21_X1   g01712(.A1(new_n1968_), .A2(new_n1842_), .B(new_n1749_), .ZN(new_n1969_));
  AOI21_X1   g01713(.A1(new_n1842_), .A2(new_n1968_), .B(new_n1969_), .ZN(new_n1970_));
  NAND2_X1   g01714(.A1(new_n1970_), .A2(new_n1744_), .ZN(new_n1971_));
  NAND3_X1   g01715(.A1(new_n1971_), .A2(new_n1767_), .A3(new_n1964_), .ZN(new_n1972_));
  OAI21_X1   g01716(.A1(new_n1844_), .A2(new_n1861_), .B(new_n1972_), .ZN(new_n1973_));
  NAND2_X1   g01717(.A1(new_n1973_), .A2(new_n1963_), .ZN(new_n1974_));
  AOI21_X1   g01718(.A1(new_n1843_), .A2(new_n1862_), .B(new_n1963_), .ZN(new_n1975_));
  NAND2_X1   g01719(.A1(new_n1975_), .A2(new_n1972_), .ZN(new_n1976_));
  NAND2_X1   g01720(.A1(new_n1974_), .A2(new_n1976_), .ZN(new_n1977_));
  OAI22_X1   g01721(.A1(new_n1168_), .A2(new_n510_), .B1(new_n495_), .B2(new_n1163_), .ZN(new_n1978_));
  NAND2_X1   g01722(.A1(new_n1774_), .A2(\b[7] ), .ZN(new_n1979_));
  AOI21_X1   g01723(.A1(new_n1978_), .A2(new_n1979_), .B(new_n1171_), .ZN(new_n1980_));
  NAND2_X1   g01724(.A1(new_n518_), .A2(new_n1980_), .ZN(new_n1981_));
  XOR2_X1    g01725(.A1(new_n1981_), .A2(\a[20] ), .Z(new_n1982_));
  NOR2_X1    g01726(.A1(new_n1866_), .A2(new_n1870_), .ZN(new_n1983_));
  OR2_X2     g01727(.A1(new_n1983_), .A2(new_n1868_), .Z(new_n1984_));
  XOR2_X1    g01728(.A1(new_n1861_), .A2(new_n1843_), .Z(new_n1985_));
  XOR2_X1    g01729(.A1(new_n1851_), .A2(new_n1985_), .Z(new_n1986_));
  NAND2_X1   g01730(.A1(new_n1986_), .A2(new_n1849_), .ZN(new_n1987_));
  NAND2_X1   g01731(.A1(new_n1984_), .A2(new_n1987_), .ZN(new_n1988_));
  XOR2_X1    g01732(.A1(new_n1988_), .A2(new_n1982_), .Z(new_n1989_));
  XOR2_X1    g01733(.A1(new_n1989_), .A2(new_n1977_), .Z(new_n1990_));
  OAI22_X1   g01734(.A1(new_n940_), .A2(new_n717_), .B1(new_n659_), .B2(new_n935_), .ZN(new_n1991_));
  NAND2_X1   g01735(.A1(new_n1458_), .A2(\b[10] ), .ZN(new_n1992_));
  AOI21_X1   g01736(.A1(new_n1991_), .A2(new_n1992_), .B(new_n943_), .ZN(new_n1993_));
  NAND2_X1   g01737(.A1(new_n716_), .A2(new_n1993_), .ZN(new_n1994_));
  XOR2_X1    g01738(.A1(new_n1994_), .A2(\a[17] ), .Z(new_n1995_));
  INV_X1     g01739(.I(new_n1877_), .ZN(new_n1996_));
  OAI21_X1   g01740(.A1(new_n1996_), .A2(new_n1881_), .B(new_n1879_), .ZN(new_n1997_));
  INV_X1     g01741(.I(new_n1871_), .ZN(new_n1998_));
  NAND2_X1   g01742(.A1(new_n1998_), .A2(new_n1876_), .ZN(new_n1999_));
  NAND2_X1   g01743(.A1(new_n1997_), .A2(new_n1999_), .ZN(new_n2000_));
  XOR2_X1    g01744(.A1(new_n2000_), .A2(new_n1995_), .Z(new_n2001_));
  XNOR2_X1   g01745(.A1(new_n2001_), .A2(new_n1990_), .ZN(new_n2002_));
  OAI22_X1   g01746(.A1(new_n757_), .A2(new_n904_), .B1(new_n848_), .B2(new_n752_), .ZN(new_n2003_));
  NAND2_X1   g01747(.A1(new_n1182_), .A2(\b[13] ), .ZN(new_n2004_));
  AOI21_X1   g01748(.A1(new_n2003_), .A2(new_n2004_), .B(new_n760_), .ZN(new_n2005_));
  NAND2_X1   g01749(.A1(new_n907_), .A2(new_n2005_), .ZN(new_n2006_));
  XOR2_X1    g01750(.A1(new_n2006_), .A2(\a[14] ), .Z(new_n2007_));
  INV_X1     g01751(.I(new_n1882_), .ZN(new_n2008_));
  AOI22_X1   g01752(.A1(new_n2008_), .A2(new_n1887_), .B1(new_n1839_), .B2(new_n1802_), .ZN(new_n2009_));
  NAND2_X1   g01753(.A1(new_n2009_), .A2(new_n1888_), .ZN(new_n2010_));
  XOR2_X1    g01754(.A1(new_n2010_), .A2(new_n2007_), .Z(new_n2011_));
  XNOR2_X1   g01755(.A1(new_n2011_), .A2(new_n2002_), .ZN(new_n2012_));
  OAI22_X1   g01756(.A1(new_n582_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n577_), .ZN(new_n2013_));
  NAND2_X1   g01757(.A1(new_n960_), .A2(\b[16] ), .ZN(new_n2014_));
  AOI21_X1   g01758(.A1(new_n2013_), .A2(new_n2014_), .B(new_n585_), .ZN(new_n2015_));
  NAND2_X1   g01759(.A1(new_n1123_), .A2(new_n2015_), .ZN(new_n2016_));
  XOR2_X1    g01760(.A1(new_n2016_), .A2(new_n572_), .Z(new_n2017_));
  XOR2_X1    g01761(.A1(new_n1888_), .A2(new_n1897_), .Z(new_n2018_));
  NOR2_X1    g01762(.A1(new_n2018_), .A2(new_n1894_), .ZN(new_n2019_));
  AOI21_X1   g01763(.A1(new_n1900_), .A2(new_n1901_), .B(new_n2019_), .ZN(new_n2020_));
  XOR2_X1    g01764(.A1(new_n2020_), .A2(new_n2017_), .Z(new_n2021_));
  XNOR2_X1   g01765(.A1(new_n2021_), .A2(new_n2012_), .ZN(new_n2022_));
  OAI22_X1   g01766(.A1(new_n437_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n431_), .ZN(new_n2023_));
  NAND2_X1   g01767(.A1(new_n775_), .A2(\b[19] ), .ZN(new_n2024_));
  AOI21_X1   g01768(.A1(new_n2023_), .A2(new_n2024_), .B(new_n440_), .ZN(new_n2025_));
  NAND2_X1   g01769(.A1(new_n1396_), .A2(new_n2025_), .ZN(new_n2026_));
  XOR2_X1    g01770(.A1(new_n2026_), .A2(\a[8] ), .Z(new_n2027_));
  INV_X1     g01771(.I(new_n1902_), .ZN(new_n2028_));
  NAND2_X1   g01772(.A1(new_n2028_), .A2(new_n1907_), .ZN(new_n2029_));
  NAND3_X1   g01773(.A1(new_n1908_), .A2(new_n2029_), .A3(new_n1909_), .ZN(new_n2030_));
  XOR2_X1    g01774(.A1(new_n2030_), .A2(new_n2027_), .Z(new_n2031_));
  XNOR2_X1   g01775(.A1(new_n2031_), .A2(new_n2022_), .ZN(new_n2032_));
  OAI22_X1   g01776(.A1(new_n364_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n320_), .ZN(new_n2033_));
  NAND2_X1   g01777(.A1(new_n594_), .A2(\b[22] ), .ZN(new_n2034_));
  AOI21_X1   g01778(.A1(new_n2033_), .A2(new_n2034_), .B(new_n312_), .ZN(new_n2035_));
  NAND2_X1   g01779(.A1(new_n1708_), .A2(new_n2035_), .ZN(new_n2036_));
  XOR2_X1    g01780(.A1(new_n2036_), .A2(\a[5] ), .Z(new_n2037_));
  XNOR2_X1   g01781(.A1(new_n2032_), .A2(new_n2037_), .ZN(new_n2038_));
  INV_X1     g01782(.I(\b[27] ), .ZN(new_n2039_));
  XOR2_X1    g01783(.A1(new_n1921_), .A2(\b[25] ), .Z(new_n2040_));
  NAND2_X1   g01784(.A1(new_n2040_), .A2(new_n1923_), .ZN(new_n2041_));
  XOR2_X1    g01785(.A1(new_n2041_), .A2(new_n2039_), .Z(new_n2042_));
  OAI22_X1   g01786(.A1(new_n405_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n404_), .ZN(new_n2043_));
  NAND2_X1   g01787(.A1(new_n279_), .A2(\b[25] ), .ZN(new_n2044_));
  AOI21_X1   g01788(.A1(new_n2043_), .A2(new_n2044_), .B(new_n264_), .ZN(new_n2045_));
  NAND2_X1   g01789(.A1(new_n2042_), .A2(new_n2045_), .ZN(new_n2046_));
  XOR2_X1    g01790(.A1(new_n2046_), .A2(new_n271_), .Z(new_n2047_));
  NOR2_X1    g01791(.A1(new_n1945_), .A2(new_n1941_), .ZN(new_n2048_));
  NOR2_X1    g01792(.A1(new_n1943_), .A2(new_n2048_), .ZN(new_n2049_));
  NOR3_X1    g01793(.A1(new_n1916_), .A2(new_n1934_), .A3(new_n1937_), .ZN(new_n2050_));
  NOR2_X1    g01794(.A1(new_n1917_), .A2(new_n1938_), .ZN(new_n2051_));
  NOR4_X1    g01795(.A1(new_n2049_), .A2(new_n1932_), .A3(new_n2050_), .A4(new_n2051_), .ZN(new_n2052_));
  XOR2_X1    g01796(.A1(new_n2052_), .A2(new_n2047_), .Z(new_n2053_));
  XOR2_X1    g01797(.A1(new_n2053_), .A2(new_n2038_), .Z(\f[27] ));
  NAND2_X1   g01798(.A1(new_n1977_), .A2(new_n1982_), .ZN(new_n2055_));
  XNOR2_X1   g01799(.A1(new_n1977_), .A2(new_n1982_), .ZN(new_n2056_));
  NAND3_X1   g01800(.A1(new_n1984_), .A2(new_n1987_), .A3(new_n2056_), .ZN(new_n2057_));
  XOR2_X1    g01801(.A1(new_n1960_), .A2(new_n1954_), .Z(new_n2058_));
  AND2_X2    g01802(.A1(new_n2058_), .A2(new_n1956_), .Z(new_n2059_));
  NOR2_X1    g01803(.A1(new_n2058_), .A2(new_n1956_), .ZN(new_n2060_));
  NOR3_X1    g01804(.A1(new_n2059_), .A2(new_n2060_), .A3(new_n1952_), .ZN(new_n2061_));
  AOI21_X1   g01805(.A1(new_n2058_), .A2(new_n1860_), .B(new_n1965_), .ZN(new_n2062_));
  NAND2_X1   g01806(.A1(new_n1960_), .A2(new_n1954_), .ZN(new_n2063_));
  NOR2_X1    g01807(.A1(new_n2062_), .A2(new_n2063_), .ZN(new_n2064_));
  NAND2_X1   g01808(.A1(new_n2062_), .A2(new_n2063_), .ZN(new_n2065_));
  INV_X1     g01809(.I(new_n2065_), .ZN(new_n2066_));
  NOR2_X1    g01810(.A1(new_n2066_), .A2(new_n2064_), .ZN(new_n2067_));
  INV_X1     g01811(.I(new_n2067_), .ZN(new_n2068_));
  OAI22_X1   g01812(.A1(new_n1760_), .A2(new_n393_), .B1(new_n290_), .B2(new_n1755_), .ZN(new_n2069_));
  OAI21_X1   g01813(.A1(new_n292_), .A2(new_n1857_), .B(new_n2069_), .ZN(new_n2070_));
  NAND3_X1   g01814(.A1(new_n2070_), .A2(new_n334_), .A3(new_n1762_), .ZN(new_n2071_));
  XOR2_X1    g01815(.A1(new_n2071_), .A2(\a[26] ), .Z(new_n2072_));
  INV_X1     g01816(.I(new_n2072_), .ZN(new_n2073_));
  INV_X1     g01817(.I(\a[29] ), .ZN(new_n2074_));
  INV_X1     g01818(.I(\a[28] ), .ZN(new_n2075_));
  NOR3_X1    g01819(.A1(new_n2075_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n2076_));
  NAND3_X1   g01820(.A1(new_n2075_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n2077_));
  INV_X1     g01821(.I(new_n2077_), .ZN(new_n2078_));
  NOR2_X1    g01822(.A1(new_n2078_), .A2(new_n2076_), .ZN(new_n2079_));
  NOR2_X1    g01823(.A1(new_n2079_), .A2(new_n258_), .ZN(new_n2080_));
  INV_X1     g01824(.I(new_n1953_), .ZN(new_n2081_));
  XNOR2_X1   g01825(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n2082_));
  NOR2_X1    g01826(.A1(new_n2081_), .A2(new_n2082_), .ZN(new_n2083_));
  INV_X1     g01827(.I(new_n2083_), .ZN(new_n2084_));
  NOR2_X1    g01828(.A1(new_n2084_), .A2(new_n267_), .ZN(new_n2085_));
  NOR2_X1    g01829(.A1(new_n1953_), .A2(new_n2082_), .ZN(new_n2086_));
  INV_X1     g01830(.I(new_n2086_), .ZN(new_n2087_));
  NOR4_X1    g01831(.A1(new_n2085_), .A2(new_n261_), .A3(new_n2080_), .A4(new_n2087_), .ZN(new_n2088_));
  XOR2_X1    g01832(.A1(new_n2088_), .A2(new_n2074_), .Z(new_n2089_));
  NOR2_X1    g01833(.A1(new_n1954_), .A2(new_n2074_), .ZN(new_n2090_));
  XNOR2_X1   g01834(.A1(new_n2089_), .A2(new_n2090_), .ZN(new_n2091_));
  XOR2_X1    g01835(.A1(new_n2091_), .A2(new_n2073_), .Z(new_n2092_));
  OR2_X2     g01836(.A1(new_n2091_), .A2(new_n2073_), .Z(new_n2093_));
  NAND2_X1   g01837(.A1(new_n2091_), .A2(new_n2073_), .ZN(new_n2094_));
  AOI21_X1   g01838(.A1(new_n2093_), .A2(new_n2094_), .B(new_n2068_), .ZN(new_n2095_));
  AOI21_X1   g01839(.A1(new_n2068_), .A2(new_n2092_), .B(new_n2095_), .ZN(new_n2096_));
  OAI22_X1   g01840(.A1(new_n1444_), .A2(new_n450_), .B1(new_n403_), .B2(new_n1439_), .ZN(new_n2097_));
  INV_X1     g01841(.I(new_n1548_), .ZN(new_n2098_));
  NAND2_X1   g01842(.A1(new_n2098_), .A2(\b[5] ), .ZN(new_n2099_));
  AOI21_X1   g01843(.A1(new_n2097_), .A2(new_n2099_), .B(new_n1447_), .ZN(new_n2100_));
  NAND2_X1   g01844(.A1(new_n454_), .A2(new_n2100_), .ZN(new_n2101_));
  XOR2_X1    g01845(.A1(new_n2101_), .A2(\a[23] ), .Z(new_n2102_));
  XOR2_X1    g01846(.A1(new_n2096_), .A2(new_n2102_), .Z(new_n2103_));
  AOI21_X1   g01847(.A1(new_n1974_), .A2(new_n2061_), .B(new_n2103_), .ZN(new_n2104_));
  NAND2_X1   g01848(.A1(new_n1974_), .A2(new_n2061_), .ZN(new_n2105_));
  INV_X1     g01849(.I(new_n2102_), .ZN(new_n2106_));
  XOR2_X1    g01850(.A1(new_n2096_), .A2(new_n2106_), .Z(new_n2107_));
  NOR2_X1    g01851(.A1(new_n2105_), .A2(new_n2107_), .ZN(new_n2108_));
  NOR2_X1    g01852(.A1(new_n2108_), .A2(new_n2104_), .ZN(new_n2109_));
  OAI22_X1   g01853(.A1(new_n1168_), .A2(new_n617_), .B1(new_n510_), .B2(new_n1163_), .ZN(new_n2110_));
  NAND2_X1   g01854(.A1(new_n1774_), .A2(\b[8] ), .ZN(new_n2111_));
  AOI21_X1   g01855(.A1(new_n2110_), .A2(new_n2111_), .B(new_n1171_), .ZN(new_n2112_));
  NAND2_X1   g01856(.A1(new_n616_), .A2(new_n2112_), .ZN(new_n2113_));
  XOR2_X1    g01857(.A1(new_n2113_), .A2(\a[20] ), .Z(new_n2114_));
  XOR2_X1    g01858(.A1(new_n2109_), .A2(new_n2114_), .Z(new_n2115_));
  AOI21_X1   g01859(.A1(new_n2057_), .A2(new_n2055_), .B(new_n2115_), .ZN(new_n2116_));
  NAND2_X1   g01860(.A1(new_n2057_), .A2(new_n2055_), .ZN(new_n2117_));
  INV_X1     g01861(.I(new_n2114_), .ZN(new_n2118_));
  XOR2_X1    g01862(.A1(new_n2109_), .A2(new_n2118_), .Z(new_n2119_));
  NOR2_X1    g01863(.A1(new_n2117_), .A2(new_n2119_), .ZN(new_n2120_));
  NOR2_X1    g01864(.A1(new_n2120_), .A2(new_n2116_), .ZN(new_n2121_));
  INV_X1     g01865(.I(new_n2121_), .ZN(new_n2122_));
  OAI22_X1   g01866(.A1(new_n940_), .A2(new_n795_), .B1(new_n717_), .B2(new_n935_), .ZN(new_n2123_));
  NAND2_X1   g01867(.A1(new_n1458_), .A2(\b[11] ), .ZN(new_n2124_));
  AOI21_X1   g01868(.A1(new_n2123_), .A2(new_n2124_), .B(new_n943_), .ZN(new_n2125_));
  NAND2_X1   g01869(.A1(new_n799_), .A2(new_n2125_), .ZN(new_n2126_));
  XOR2_X1    g01870(.A1(new_n2126_), .A2(\a[17] ), .Z(new_n2127_));
  NOR2_X1    g01871(.A1(new_n2122_), .A2(new_n2127_), .ZN(new_n2128_));
  INV_X1     g01872(.I(new_n2127_), .ZN(new_n2129_));
  NOR2_X1    g01873(.A1(new_n2121_), .A2(new_n2129_), .ZN(new_n2130_));
  NOR2_X1    g01874(.A1(new_n2128_), .A2(new_n2130_), .ZN(new_n2131_));
  OAI22_X1   g01875(.A1(new_n757_), .A2(new_n992_), .B1(new_n904_), .B2(new_n752_), .ZN(new_n2132_));
  NAND2_X1   g01876(.A1(new_n1182_), .A2(\b[14] ), .ZN(new_n2133_));
  AOI21_X1   g01877(.A1(new_n2132_), .A2(new_n2133_), .B(new_n760_), .ZN(new_n2134_));
  NAND2_X1   g01878(.A1(new_n991_), .A2(new_n2134_), .ZN(new_n2135_));
  XOR2_X1    g01879(.A1(new_n2135_), .A2(\a[14] ), .Z(new_n2136_));
  XNOR2_X1   g01880(.A1(new_n2131_), .A2(new_n2136_), .ZN(new_n2137_));
  INV_X1     g01881(.I(new_n2137_), .ZN(new_n2138_));
  OAI22_X1   g01882(.A1(new_n582_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n577_), .ZN(new_n2139_));
  NAND2_X1   g01883(.A1(new_n960_), .A2(\b[17] ), .ZN(new_n2140_));
  AOI21_X1   g01884(.A1(new_n2139_), .A2(new_n2140_), .B(new_n585_), .ZN(new_n2141_));
  NAND2_X1   g01885(.A1(new_n1225_), .A2(new_n2141_), .ZN(new_n2142_));
  XOR2_X1    g01886(.A1(new_n2142_), .A2(\a[11] ), .Z(new_n2143_));
  NOR2_X1    g01887(.A1(new_n2138_), .A2(new_n2143_), .ZN(new_n2144_));
  NAND2_X1   g01888(.A1(new_n2138_), .A2(new_n2143_), .ZN(new_n2145_));
  INV_X1     g01889(.I(new_n2145_), .ZN(new_n2146_));
  NOR2_X1    g01890(.A1(new_n2146_), .A2(new_n2144_), .ZN(new_n2147_));
  OAI22_X1   g01891(.A1(new_n437_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n431_), .ZN(new_n2148_));
  NAND2_X1   g01892(.A1(new_n775_), .A2(\b[20] ), .ZN(new_n2149_));
  AOI21_X1   g01893(.A1(new_n2148_), .A2(new_n2149_), .B(new_n440_), .ZN(new_n2150_));
  NAND2_X1   g01894(.A1(new_n1517_), .A2(new_n2150_), .ZN(new_n2151_));
  XOR2_X1    g01895(.A1(new_n2151_), .A2(\a[8] ), .Z(new_n2152_));
  XOR2_X1    g01896(.A1(new_n2147_), .A2(new_n2152_), .Z(new_n2153_));
  OAI22_X1   g01897(.A1(new_n364_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n320_), .ZN(new_n2154_));
  NAND2_X1   g01898(.A1(new_n594_), .A2(\b[23] ), .ZN(new_n2155_));
  AOI21_X1   g01899(.A1(new_n2154_), .A2(new_n2155_), .B(new_n312_), .ZN(new_n2156_));
  NAND2_X1   g01900(.A1(new_n1828_), .A2(new_n2156_), .ZN(new_n2157_));
  XOR2_X1    g01901(.A1(new_n2157_), .A2(\a[5] ), .Z(new_n2158_));
  NOR2_X1    g01902(.A1(new_n2153_), .A2(new_n2158_), .ZN(new_n2159_));
  NAND2_X1   g01903(.A1(new_n2153_), .A2(new_n2158_), .ZN(new_n2160_));
  INV_X1     g01904(.I(new_n2160_), .ZN(new_n2161_));
  NOR2_X1    g01905(.A1(new_n2161_), .A2(new_n2159_), .ZN(new_n2162_));
  INV_X1     g01906(.I(new_n2032_), .ZN(new_n2163_));
  NOR2_X1    g01907(.A1(new_n2163_), .A2(new_n2037_), .ZN(new_n2164_));
  XOR2_X1    g01908(.A1(new_n2164_), .A2(new_n2162_), .Z(new_n2165_));
  INV_X1     g01909(.I(new_n1921_), .ZN(new_n2166_));
  OAI21_X1   g01910(.A1(new_n1825_), .A2(new_n2039_), .B(new_n1927_), .ZN(new_n2167_));
  NAND2_X1   g01911(.A1(new_n1825_), .A2(new_n2039_), .ZN(new_n2168_));
  AOI22_X1   g01912(.A1(new_n2166_), .A2(new_n2167_), .B1(\b[26] ), .B2(new_n2168_), .ZN(new_n2169_));
  XNOR2_X1   g01913(.A1(\b[27] ), .A2(\b[28] ), .ZN(new_n2170_));
  NOR2_X1    g01914(.A1(new_n2169_), .A2(new_n2170_), .ZN(new_n2171_));
  XNOR2_X1   g01915(.A1(\b[27] ), .A2(\b[28] ), .ZN(new_n2172_));
  AOI21_X1   g01916(.A1(new_n2169_), .A2(new_n2172_), .B(new_n2171_), .ZN(new_n2173_));
  INV_X1     g01917(.I(new_n2173_), .ZN(new_n2174_));
  INV_X1     g01918(.I(\b[28] ), .ZN(new_n2175_));
  OAI22_X1   g01919(.A1(new_n405_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n404_), .ZN(new_n2176_));
  NAND2_X1   g01920(.A1(new_n279_), .A2(\b[26] ), .ZN(new_n2177_));
  AOI21_X1   g01921(.A1(new_n2176_), .A2(new_n2177_), .B(new_n264_), .ZN(new_n2178_));
  NAND2_X1   g01922(.A1(new_n2174_), .A2(new_n2178_), .ZN(new_n2179_));
  XOR2_X1    g01923(.A1(new_n2179_), .A2(\a[2] ), .Z(new_n2180_));
  INV_X1     g01924(.I(new_n2180_), .ZN(new_n2181_));
  NAND2_X1   g01925(.A1(new_n2165_), .A2(new_n2181_), .ZN(new_n2182_));
  OR2_X2     g01926(.A1(new_n2165_), .A2(new_n2181_), .Z(new_n2183_));
  NAND2_X1   g01927(.A1(new_n2183_), .A2(new_n2182_), .ZN(\f[28] ));
  OAI22_X1   g01928(.A1(new_n437_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n431_), .ZN(new_n2185_));
  NAND2_X1   g01929(.A1(new_n775_), .A2(\b[21] ), .ZN(new_n2186_));
  AOI21_X1   g01930(.A1(new_n2185_), .A2(new_n2186_), .B(new_n440_), .ZN(new_n2187_));
  NAND2_X1   g01931(.A1(new_n1604_), .A2(new_n2187_), .ZN(new_n2188_));
  XOR2_X1    g01932(.A1(new_n2188_), .A2(new_n429_), .Z(new_n2189_));
  OAI22_X1   g01933(.A1(new_n582_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n577_), .ZN(new_n2190_));
  NAND2_X1   g01934(.A1(new_n960_), .A2(\b[18] ), .ZN(new_n2191_));
  AOI21_X1   g01935(.A1(new_n2190_), .A2(new_n2191_), .B(new_n585_), .ZN(new_n2192_));
  NAND2_X1   g01936(.A1(new_n1304_), .A2(new_n2192_), .ZN(new_n2193_));
  XOR2_X1    g01937(.A1(new_n2193_), .A2(\a[11] ), .Z(new_n2194_));
  INV_X1     g01938(.I(new_n2194_), .ZN(new_n2195_));
  NOR2_X1    g01939(.A1(new_n2138_), .A2(new_n2143_), .ZN(new_n2196_));
  OAI22_X1   g01940(.A1(new_n1760_), .A2(new_n347_), .B1(new_n393_), .B2(new_n1755_), .ZN(new_n2197_));
  OAI21_X1   g01941(.A1(new_n290_), .A2(new_n1857_), .B(new_n2197_), .ZN(new_n2198_));
  AOI21_X1   g01942(.A1(new_n352_), .A2(new_n1762_), .B(new_n2198_), .ZN(new_n2199_));
  XOR2_X1    g01943(.A1(new_n2199_), .A2(new_n1750_), .Z(new_n2200_));
  INV_X1     g01944(.I(new_n2200_), .ZN(new_n2201_));
  OAI22_X1   g01945(.A1(new_n1444_), .A2(new_n495_), .B1(new_n450_), .B2(new_n1439_), .ZN(new_n2202_));
  NAND2_X1   g01946(.A1(new_n2098_), .A2(\b[6] ), .ZN(new_n2203_));
  AOI21_X1   g01947(.A1(new_n2202_), .A2(new_n2203_), .B(new_n1447_), .ZN(new_n2204_));
  NAND2_X1   g01948(.A1(new_n494_), .A2(new_n2204_), .ZN(new_n2205_));
  XOR2_X1    g01949(.A1(new_n2205_), .A2(\a[23] ), .Z(new_n2206_));
  NAND2_X1   g01950(.A1(new_n2068_), .A2(new_n2093_), .ZN(new_n2207_));
  NAND2_X1   g01951(.A1(new_n2207_), .A2(new_n2094_), .ZN(new_n2208_));
  NAND2_X1   g01952(.A1(new_n2089_), .A2(new_n2090_), .ZN(new_n2209_));
  NOR2_X1    g01953(.A1(new_n2087_), .A2(new_n278_), .ZN(new_n2210_));
  XNOR2_X1   g01954(.A1(\a[26] ), .A2(\a[28] ), .ZN(new_n2211_));
  NAND2_X1   g01955(.A1(new_n1953_), .A2(new_n2211_), .ZN(new_n2212_));
  XNOR2_X1   g01956(.A1(\a[26] ), .A2(\a[29] ), .ZN(new_n2213_));
  NAND2_X1   g01957(.A1(new_n2212_), .A2(new_n2213_), .ZN(new_n2214_));
  OAI22_X1   g01958(.A1(new_n2084_), .A2(new_n292_), .B1(new_n267_), .B2(new_n2079_), .ZN(new_n2215_));
  NOR4_X1    g01959(.A1(new_n2215_), .A2(new_n258_), .A3(new_n2210_), .A4(new_n2214_), .ZN(new_n2216_));
  XOR2_X1    g01960(.A1(new_n2216_), .A2(new_n2074_), .Z(new_n2217_));
  XOR2_X1    g01961(.A1(new_n2209_), .A2(new_n2217_), .Z(new_n2218_));
  INV_X1     g01962(.I(new_n2218_), .ZN(new_n2219_));
  XOR2_X1    g01963(.A1(new_n2208_), .A2(new_n2219_), .Z(new_n2220_));
  XOR2_X1    g01964(.A1(new_n2220_), .A2(new_n2206_), .Z(new_n2221_));
  XOR2_X1    g01965(.A1(new_n2221_), .A2(new_n2201_), .Z(new_n2222_));
  INV_X1     g01966(.I(new_n2222_), .ZN(new_n2223_));
  XOR2_X1    g01967(.A1(new_n2105_), .A2(new_n2106_), .Z(new_n2224_));
  NAND2_X1   g01968(.A1(new_n2224_), .A2(new_n2096_), .ZN(new_n2225_));
  XOR2_X1    g01969(.A1(new_n2225_), .A2(new_n2223_), .Z(new_n2226_));
  NAND2_X1   g01970(.A1(new_n2105_), .A2(new_n2106_), .ZN(new_n2227_));
  XNOR2_X1   g01971(.A1(new_n2226_), .A2(new_n2227_), .ZN(new_n2228_));
  OAI22_X1   g01972(.A1(new_n1168_), .A2(new_n659_), .B1(new_n617_), .B2(new_n1163_), .ZN(new_n2229_));
  NAND2_X1   g01973(.A1(new_n1774_), .A2(\b[9] ), .ZN(new_n2230_));
  AOI21_X1   g01974(.A1(new_n2229_), .A2(new_n2230_), .B(new_n1171_), .ZN(new_n2231_));
  NAND2_X1   g01975(.A1(new_n663_), .A2(new_n2231_), .ZN(new_n2232_));
  XOR2_X1    g01976(.A1(new_n2232_), .A2(\a[20] ), .Z(new_n2233_));
  XOR2_X1    g01977(.A1(new_n2228_), .A2(new_n2233_), .Z(new_n2234_));
  XOR2_X1    g01978(.A1(new_n2117_), .A2(new_n2114_), .Z(new_n2235_));
  NOR3_X1    g01979(.A1(new_n2235_), .A2(new_n2104_), .A3(new_n2108_), .ZN(new_n2236_));
  XOR2_X1    g01980(.A1(new_n2236_), .A2(new_n2234_), .Z(new_n2237_));
  NAND2_X1   g01981(.A1(new_n2117_), .A2(new_n2118_), .ZN(new_n2238_));
  XNOR2_X1   g01982(.A1(new_n2237_), .A2(new_n2238_), .ZN(new_n2239_));
  INV_X1     g01983(.I(new_n2239_), .ZN(new_n2240_));
  OAI22_X1   g01984(.A1(new_n940_), .A2(new_n848_), .B1(new_n795_), .B2(new_n935_), .ZN(new_n2241_));
  NAND2_X1   g01985(.A1(new_n1458_), .A2(\b[12] ), .ZN(new_n2242_));
  AOI21_X1   g01986(.A1(new_n2241_), .A2(new_n2242_), .B(new_n943_), .ZN(new_n2243_));
  NAND2_X1   g01987(.A1(new_n847_), .A2(new_n2243_), .ZN(new_n2244_));
  XOR2_X1    g01988(.A1(new_n2244_), .A2(\a[17] ), .Z(new_n2245_));
  NOR2_X1    g01989(.A1(new_n2240_), .A2(new_n2245_), .ZN(new_n2246_));
  NAND2_X1   g01990(.A1(new_n2240_), .A2(new_n2245_), .ZN(new_n2247_));
  INV_X1     g01991(.I(new_n2247_), .ZN(new_n2248_));
  NOR2_X1    g01992(.A1(new_n2248_), .A2(new_n2246_), .ZN(new_n2249_));
  NOR2_X1    g01993(.A1(new_n2122_), .A2(new_n2127_), .ZN(new_n2250_));
  XOR2_X1    g01994(.A1(new_n2249_), .A2(new_n2250_), .Z(new_n2251_));
  OAI22_X1   g01995(.A1(new_n757_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n752_), .ZN(new_n2252_));
  NAND2_X1   g01996(.A1(new_n1182_), .A2(\b[15] ), .ZN(new_n2253_));
  AOI21_X1   g01997(.A1(new_n2252_), .A2(new_n2253_), .B(new_n760_), .ZN(new_n2254_));
  NAND2_X1   g01998(.A1(new_n1047_), .A2(new_n2254_), .ZN(new_n2255_));
  XOR2_X1    g01999(.A1(new_n2255_), .A2(\a[14] ), .Z(new_n2256_));
  XOR2_X1    g02000(.A1(new_n2251_), .A2(new_n2256_), .Z(new_n2257_));
  NOR3_X1    g02001(.A1(new_n2128_), .A2(new_n2130_), .A3(new_n2136_), .ZN(new_n2258_));
  XNOR2_X1   g02002(.A1(new_n2257_), .A2(new_n2258_), .ZN(new_n2259_));
  XOR2_X1    g02003(.A1(new_n2259_), .A2(new_n2196_), .Z(new_n2260_));
  XOR2_X1    g02004(.A1(new_n2260_), .A2(new_n2195_), .Z(new_n2261_));
  XOR2_X1    g02005(.A1(new_n2261_), .A2(new_n2189_), .Z(new_n2262_));
  INV_X1     g02006(.I(new_n2147_), .ZN(new_n2263_));
  NOR2_X1    g02007(.A1(new_n2263_), .A2(new_n2152_), .ZN(new_n2264_));
  XOR2_X1    g02008(.A1(new_n2262_), .A2(new_n2264_), .Z(new_n2265_));
  OAI22_X1   g02009(.A1(new_n364_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n320_), .ZN(new_n2266_));
  NAND2_X1   g02010(.A1(new_n594_), .A2(\b[24] ), .ZN(new_n2267_));
  AOI21_X1   g02011(.A1(new_n2266_), .A2(new_n2267_), .B(new_n312_), .ZN(new_n2268_));
  NAND2_X1   g02012(.A1(new_n1926_), .A2(new_n2268_), .ZN(new_n2269_));
  XOR2_X1    g02013(.A1(new_n2269_), .A2(\a[5] ), .Z(new_n2270_));
  XOR2_X1    g02014(.A1(new_n2265_), .A2(new_n2270_), .Z(new_n2271_));
  INV_X1     g02015(.I(\b[29] ), .ZN(new_n2272_));
  INV_X1     g02016(.I(new_n2170_), .ZN(new_n2273_));
  XOR2_X1    g02017(.A1(new_n2169_), .A2(new_n2039_), .Z(new_n2274_));
  NAND2_X1   g02018(.A1(new_n2274_), .A2(new_n2273_), .ZN(new_n2275_));
  XOR2_X1    g02019(.A1(new_n2275_), .A2(new_n2272_), .Z(new_n2276_));
  NAND2_X1   g02020(.A1(new_n283_), .A2(\b[29] ), .ZN(new_n2277_));
  NAND2_X1   g02021(.A1(new_n279_), .A2(\b[27] ), .ZN(new_n2278_));
  AOI21_X1   g02022(.A1(\b[28] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n2279_));
  NAND4_X1   g02023(.A1(new_n2276_), .A2(new_n2277_), .A3(new_n2278_), .A4(new_n2279_), .ZN(new_n2280_));
  XOR2_X1    g02024(.A1(new_n2280_), .A2(\a[2] ), .Z(new_n2281_));
  NAND2_X1   g02025(.A1(new_n2163_), .A2(new_n2037_), .ZN(new_n2282_));
  NOR2_X1    g02026(.A1(new_n2161_), .A2(new_n2159_), .ZN(new_n2283_));
  NAND2_X1   g02027(.A1(new_n2282_), .A2(new_n2283_), .ZN(new_n2284_));
  XOR2_X1    g02028(.A1(new_n2284_), .A2(new_n2281_), .Z(new_n2285_));
  XOR2_X1    g02029(.A1(new_n2285_), .A2(new_n2271_), .Z(new_n2286_));
  NAND2_X1   g02030(.A1(new_n2165_), .A2(new_n2181_), .ZN(new_n2287_));
  XOR2_X1    g02031(.A1(new_n2286_), .A2(new_n2287_), .Z(\f[29] ));
  INV_X1     g02032(.I(new_n1755_), .ZN(new_n2289_));
  AOI22_X1   g02033(.A1(\b[6] ), .A2(new_n1759_), .B1(new_n2289_), .B2(\b[5] ), .ZN(new_n2290_));
  NOR2_X1    g02034(.A1(new_n1857_), .A2(new_n393_), .ZN(new_n2291_));
  OAI21_X1   g02035(.A1(new_n2290_), .A2(new_n2291_), .B(new_n1762_), .ZN(new_n2292_));
  NOR2_X1    g02036(.A1(new_n524_), .A2(new_n2292_), .ZN(new_n2293_));
  XOR2_X1    g02037(.A1(new_n2293_), .A2(\a[26] ), .Z(new_n2294_));
  XNOR2_X1   g02038(.A1(\a[29] ), .A2(\a[30] ), .ZN(new_n2295_));
  NOR2_X1    g02039(.A1(new_n2295_), .A2(new_n258_), .ZN(new_n2296_));
  INV_X1     g02040(.I(new_n2217_), .ZN(new_n2297_));
  NOR2_X1    g02041(.A1(new_n2297_), .A2(new_n2209_), .ZN(new_n2298_));
  NOR2_X1    g02042(.A1(new_n2214_), .A2(new_n267_), .ZN(new_n2299_));
  OAI22_X1   g02043(.A1(new_n2084_), .A2(new_n290_), .B1(new_n292_), .B2(new_n2079_), .ZN(new_n2300_));
  NOR4_X1    g02044(.A1(new_n2300_), .A2(new_n677_), .A3(new_n2087_), .A4(new_n2299_), .ZN(new_n2301_));
  XOR2_X1    g02045(.A1(new_n2301_), .A2(new_n2074_), .Z(new_n2302_));
  XOR2_X1    g02046(.A1(new_n2298_), .A2(new_n2302_), .Z(new_n2303_));
  XOR2_X1    g02047(.A1(new_n2303_), .A2(new_n2296_), .Z(new_n2304_));
  XOR2_X1    g02048(.A1(new_n2304_), .A2(new_n2294_), .Z(new_n2305_));
  XOR2_X1    g02049(.A1(new_n2067_), .A2(new_n2072_), .Z(new_n2306_));
  INV_X1     g02050(.I(new_n2209_), .ZN(new_n2307_));
  NOR2_X1    g02051(.A1(new_n2307_), .A2(new_n2217_), .ZN(new_n2308_));
  NOR2_X1    g02052(.A1(new_n2308_), .A2(new_n2298_), .ZN(new_n2309_));
  XOR2_X1    g02053(.A1(new_n2309_), .A2(\a[26] ), .Z(new_n2310_));
  OAI21_X1   g02054(.A1(new_n2310_), .A2(new_n2199_), .B(new_n2073_), .ZN(new_n2311_));
  AOI21_X1   g02055(.A1(new_n2199_), .A2(new_n2310_), .B(new_n2311_), .ZN(new_n2312_));
  NAND2_X1   g02056(.A1(new_n2312_), .A2(new_n2068_), .ZN(new_n2313_));
  NAND3_X1   g02057(.A1(new_n2313_), .A2(new_n2091_), .A3(new_n2306_), .ZN(new_n2314_));
  OAI21_X1   g02058(.A1(new_n2201_), .A2(new_n2218_), .B(new_n2314_), .ZN(new_n2315_));
  NAND2_X1   g02059(.A1(new_n2315_), .A2(new_n2305_), .ZN(new_n2316_));
  AOI21_X1   g02060(.A1(new_n2200_), .A2(new_n2219_), .B(new_n2305_), .ZN(new_n2317_));
  NAND2_X1   g02061(.A1(new_n2317_), .A2(new_n2314_), .ZN(new_n2318_));
  NAND2_X1   g02062(.A1(new_n2316_), .A2(new_n2318_), .ZN(new_n2319_));
  OAI22_X1   g02063(.A1(new_n1444_), .A2(new_n510_), .B1(new_n495_), .B2(new_n1439_), .ZN(new_n2320_));
  NAND2_X1   g02064(.A1(new_n2098_), .A2(\b[7] ), .ZN(new_n2321_));
  AOI21_X1   g02065(.A1(new_n2320_), .A2(new_n2321_), .B(new_n1447_), .ZN(new_n2322_));
  NAND2_X1   g02066(.A1(new_n518_), .A2(new_n2322_), .ZN(new_n2323_));
  XOR2_X1    g02067(.A1(new_n2323_), .A2(\a[23] ), .Z(new_n2324_));
  NOR2_X1    g02068(.A1(new_n2223_), .A2(new_n2227_), .ZN(new_n2325_));
  XOR2_X1    g02069(.A1(new_n2218_), .A2(new_n2200_), .Z(new_n2326_));
  XOR2_X1    g02070(.A1(new_n2208_), .A2(new_n2326_), .Z(new_n2327_));
  NAND2_X1   g02071(.A1(new_n2327_), .A2(new_n2206_), .ZN(new_n2328_));
  OAI21_X1   g02072(.A1(new_n2325_), .A2(new_n2225_), .B(new_n2328_), .ZN(new_n2329_));
  XOR2_X1    g02073(.A1(new_n2329_), .A2(new_n2324_), .Z(new_n2330_));
  XOR2_X1    g02074(.A1(new_n2330_), .A2(new_n2319_), .Z(new_n2331_));
  OAI22_X1   g02075(.A1(new_n1168_), .A2(new_n717_), .B1(new_n659_), .B2(new_n1163_), .ZN(new_n2332_));
  NAND2_X1   g02076(.A1(new_n1774_), .A2(\b[10] ), .ZN(new_n2333_));
  AOI21_X1   g02077(.A1(new_n2332_), .A2(new_n2333_), .B(new_n1171_), .ZN(new_n2334_));
  NAND2_X1   g02078(.A1(new_n716_), .A2(new_n2334_), .ZN(new_n2335_));
  XOR2_X1    g02079(.A1(new_n2335_), .A2(\a[20] ), .Z(new_n2336_));
  INV_X1     g02080(.I(new_n2234_), .ZN(new_n2337_));
  OAI21_X1   g02081(.A1(new_n2337_), .A2(new_n2238_), .B(new_n2236_), .ZN(new_n2338_));
  INV_X1     g02082(.I(new_n2228_), .ZN(new_n2339_));
  NAND2_X1   g02083(.A1(new_n2339_), .A2(new_n2233_), .ZN(new_n2340_));
  NAND2_X1   g02084(.A1(new_n2338_), .A2(new_n2340_), .ZN(new_n2341_));
  XOR2_X1    g02085(.A1(new_n2341_), .A2(new_n2336_), .Z(new_n2342_));
  XNOR2_X1   g02086(.A1(new_n2342_), .A2(new_n2331_), .ZN(new_n2343_));
  OAI22_X1   g02087(.A1(new_n940_), .A2(new_n904_), .B1(new_n848_), .B2(new_n935_), .ZN(new_n2344_));
  NAND2_X1   g02088(.A1(new_n1458_), .A2(\b[13] ), .ZN(new_n2345_));
  AOI21_X1   g02089(.A1(new_n2344_), .A2(new_n2345_), .B(new_n943_), .ZN(new_n2346_));
  NAND2_X1   g02090(.A1(new_n907_), .A2(new_n2346_), .ZN(new_n2347_));
  XOR2_X1    g02091(.A1(new_n2347_), .A2(new_n930_), .Z(new_n2348_));
  NOR3_X1    g02092(.A1(new_n2248_), .A2(new_n2130_), .A3(new_n2246_), .ZN(new_n2349_));
  XOR2_X1    g02093(.A1(new_n2349_), .A2(new_n2348_), .Z(new_n2350_));
  XNOR2_X1   g02094(.A1(new_n2350_), .A2(new_n2343_), .ZN(new_n2351_));
  OAI22_X1   g02095(.A1(new_n757_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n752_), .ZN(new_n2352_));
  NAND2_X1   g02096(.A1(new_n1182_), .A2(\b[16] ), .ZN(new_n2353_));
  AOI21_X1   g02097(.A1(new_n2352_), .A2(new_n2353_), .B(new_n760_), .ZN(new_n2354_));
  NAND2_X1   g02098(.A1(new_n1123_), .A2(new_n2354_), .ZN(new_n2355_));
  XOR2_X1    g02099(.A1(new_n2355_), .A2(new_n747_), .Z(new_n2356_));
  INV_X1     g02100(.I(new_n2256_), .ZN(new_n2357_));
  NOR2_X1    g02101(.A1(new_n2251_), .A2(new_n2357_), .ZN(new_n2358_));
  NOR3_X1    g02102(.A1(new_n2257_), .A2(new_n2358_), .A3(new_n2258_), .ZN(new_n2359_));
  XOR2_X1    g02103(.A1(new_n2359_), .A2(new_n2356_), .Z(new_n2360_));
  XNOR2_X1   g02104(.A1(new_n2360_), .A2(new_n2351_), .ZN(new_n2361_));
  OAI22_X1   g02105(.A1(new_n582_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n577_), .ZN(new_n2362_));
  NAND2_X1   g02106(.A1(new_n960_), .A2(\b[19] ), .ZN(new_n2363_));
  AOI21_X1   g02107(.A1(new_n2362_), .A2(new_n2363_), .B(new_n585_), .ZN(new_n2364_));
  NAND2_X1   g02108(.A1(new_n1396_), .A2(new_n2364_), .ZN(new_n2365_));
  XOR2_X1    g02109(.A1(new_n2365_), .A2(\a[11] ), .Z(new_n2366_));
  NAND2_X1   g02110(.A1(new_n2259_), .A2(new_n2194_), .ZN(new_n2367_));
  OR2_X2     g02111(.A1(new_n2259_), .A2(new_n2194_), .Z(new_n2368_));
  NAND3_X1   g02112(.A1(new_n2368_), .A2(new_n2367_), .A3(new_n2196_), .ZN(new_n2369_));
  OAI21_X1   g02113(.A1(new_n2195_), .A2(new_n2259_), .B(new_n2369_), .ZN(new_n2370_));
  XOR2_X1    g02114(.A1(new_n2370_), .A2(new_n2366_), .Z(new_n2371_));
  XNOR2_X1   g02115(.A1(new_n2371_), .A2(new_n2361_), .ZN(new_n2372_));
  INV_X1     g02116(.I(new_n2372_), .ZN(new_n2373_));
  OAI22_X1   g02117(.A1(new_n437_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n431_), .ZN(new_n2374_));
  NAND2_X1   g02118(.A1(new_n775_), .A2(\b[22] ), .ZN(new_n2375_));
  AOI21_X1   g02119(.A1(new_n2374_), .A2(new_n2375_), .B(new_n440_), .ZN(new_n2376_));
  NAND2_X1   g02120(.A1(new_n1708_), .A2(new_n2376_), .ZN(new_n2377_));
  XOR2_X1    g02121(.A1(new_n2377_), .A2(\a[8] ), .Z(new_n2378_));
  NAND2_X1   g02122(.A1(new_n2263_), .A2(new_n2152_), .ZN(new_n2379_));
  NAND2_X1   g02123(.A1(new_n2262_), .A2(new_n2379_), .ZN(new_n2380_));
  XOR2_X1    g02124(.A1(new_n2259_), .A2(new_n2195_), .Z(new_n2381_));
  XOR2_X1    g02125(.A1(new_n2381_), .A2(new_n2196_), .Z(new_n2382_));
  NOR2_X1    g02126(.A1(new_n2382_), .A2(new_n2189_), .ZN(new_n2383_));
  NOR2_X1    g02127(.A1(new_n2380_), .A2(new_n2383_), .ZN(new_n2384_));
  XNOR2_X1   g02128(.A1(new_n2384_), .A2(new_n2378_), .ZN(new_n2385_));
  XOR2_X1    g02129(.A1(new_n2385_), .A2(new_n2373_), .Z(new_n2386_));
  INV_X1     g02130(.I(new_n2386_), .ZN(new_n2387_));
  OAI22_X1   g02131(.A1(new_n364_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n320_), .ZN(new_n2388_));
  NAND2_X1   g02132(.A1(new_n594_), .A2(\b[25] ), .ZN(new_n2389_));
  AOI21_X1   g02133(.A1(new_n2388_), .A2(new_n2389_), .B(new_n312_), .ZN(new_n2390_));
  NAND2_X1   g02134(.A1(new_n2042_), .A2(new_n2390_), .ZN(new_n2391_));
  XOR2_X1    g02135(.A1(new_n2391_), .A2(\a[5] ), .Z(new_n2392_));
  NOR2_X1    g02136(.A1(new_n2387_), .A2(new_n2392_), .ZN(new_n2393_));
  INV_X1     g02137(.I(new_n2392_), .ZN(new_n2394_));
  NOR2_X1    g02138(.A1(new_n2386_), .A2(new_n2394_), .ZN(new_n2395_));
  NOR2_X1    g02139(.A1(new_n2393_), .A2(new_n2395_), .ZN(new_n2396_));
  OAI21_X1   g02140(.A1(new_n2039_), .A2(new_n2272_), .B(new_n2175_), .ZN(new_n2397_));
  NAND2_X1   g02141(.A1(new_n2169_), .A2(new_n2397_), .ZN(new_n2398_));
  OAI21_X1   g02142(.A1(\b[27] ), .A2(\b[29] ), .B(\b[28] ), .ZN(new_n2399_));
  NAND2_X1   g02143(.A1(new_n2398_), .A2(new_n2399_), .ZN(new_n2400_));
  XOR2_X1    g02144(.A1(\b[29] ), .A2(\b[30] ), .Z(new_n2401_));
  NAND2_X1   g02145(.A1(new_n2400_), .A2(new_n2401_), .ZN(new_n2402_));
  XOR2_X1    g02146(.A1(\b[29] ), .A2(\b[30] ), .Z(new_n2403_));
  OAI21_X1   g02147(.A1(new_n2400_), .A2(new_n2403_), .B(new_n2402_), .ZN(new_n2404_));
  INV_X1     g02148(.I(\b[30] ), .ZN(new_n2405_));
  OAI22_X1   g02149(.A1(new_n405_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n404_), .ZN(new_n2406_));
  NAND2_X1   g02150(.A1(new_n279_), .A2(\b[28] ), .ZN(new_n2407_));
  AOI21_X1   g02151(.A1(new_n2406_), .A2(new_n2407_), .B(new_n264_), .ZN(new_n2408_));
  NAND2_X1   g02152(.A1(new_n2404_), .A2(new_n2408_), .ZN(new_n2409_));
  XOR2_X1    g02153(.A1(new_n2409_), .A2(\a[2] ), .Z(new_n2410_));
  INV_X1     g02154(.I(new_n2410_), .ZN(new_n2411_));
  XOR2_X1    g02155(.A1(new_n2396_), .A2(new_n2411_), .Z(new_n2412_));
  INV_X1     g02156(.I(new_n2284_), .ZN(new_n2413_));
  OAI21_X1   g02157(.A1(new_n2271_), .A2(new_n2413_), .B(new_n2281_), .ZN(new_n2414_));
  AOI21_X1   g02158(.A1(new_n2271_), .A2(new_n2413_), .B(new_n2414_), .ZN(new_n2415_));
  NAND3_X1   g02159(.A1(new_n2286_), .A2(new_n2415_), .A3(new_n2183_), .ZN(new_n2416_));
  XOR2_X1    g02160(.A1(new_n2412_), .A2(new_n2416_), .Z(\f[30] ));
  NAND2_X1   g02161(.A1(new_n2373_), .A2(new_n2378_), .ZN(new_n2418_));
  XOR2_X1    g02162(.A1(new_n2372_), .A2(new_n2378_), .Z(new_n2419_));
  NAND2_X1   g02163(.A1(new_n2419_), .A2(new_n2384_), .ZN(new_n2420_));
  NAND2_X1   g02164(.A1(new_n2420_), .A2(new_n2418_), .ZN(new_n2421_));
  INV_X1     g02165(.I(new_n2324_), .ZN(new_n2422_));
  XOR2_X1    g02166(.A1(new_n2319_), .A2(new_n2422_), .Z(new_n2423_));
  NOR2_X1    g02167(.A1(new_n2325_), .A2(new_n2225_), .ZN(new_n2424_));
  NAND2_X1   g02168(.A1(new_n2423_), .A2(new_n2328_), .ZN(new_n2425_));
  NOR2_X1    g02169(.A1(new_n2424_), .A2(new_n2425_), .ZN(new_n2426_));
  AOI21_X1   g02170(.A1(new_n2324_), .A2(new_n2423_), .B(new_n2426_), .ZN(new_n2427_));
  XOR2_X1    g02171(.A1(new_n2302_), .A2(new_n2296_), .Z(new_n2428_));
  AND2_X2    g02172(.A1(new_n2428_), .A2(new_n2298_), .Z(new_n2429_));
  NOR2_X1    g02173(.A1(new_n2428_), .A2(new_n2298_), .ZN(new_n2430_));
  NOR3_X1    g02174(.A1(new_n2429_), .A2(new_n2430_), .A3(new_n2294_), .ZN(new_n2431_));
  AOI21_X1   g02175(.A1(new_n2428_), .A2(new_n2217_), .B(new_n2307_), .ZN(new_n2432_));
  NAND2_X1   g02176(.A1(new_n2302_), .A2(new_n2296_), .ZN(new_n2433_));
  NOR2_X1    g02177(.A1(new_n2432_), .A2(new_n2433_), .ZN(new_n2434_));
  NAND2_X1   g02178(.A1(new_n2432_), .A2(new_n2433_), .ZN(new_n2435_));
  INV_X1     g02179(.I(new_n2435_), .ZN(new_n2436_));
  NOR2_X1    g02180(.A1(new_n2436_), .A2(new_n2434_), .ZN(new_n2437_));
  OAI22_X1   g02181(.A1(new_n2084_), .A2(new_n393_), .B1(new_n290_), .B2(new_n2079_), .ZN(new_n2438_));
  OAI21_X1   g02182(.A1(new_n292_), .A2(new_n2214_), .B(new_n2438_), .ZN(new_n2439_));
  NAND3_X1   g02183(.A1(new_n2439_), .A2(new_n334_), .A3(new_n2086_), .ZN(new_n2440_));
  XOR2_X1    g02184(.A1(new_n2440_), .A2(\a[29] ), .Z(new_n2441_));
  INV_X1     g02185(.I(\a[32] ), .ZN(new_n2442_));
  INV_X1     g02186(.I(\a[31] ), .ZN(new_n2443_));
  NOR3_X1    g02187(.A1(new_n2443_), .A2(\a[29] ), .A3(\a[30] ), .ZN(new_n2444_));
  NAND3_X1   g02188(.A1(new_n2443_), .A2(\a[29] ), .A3(\a[30] ), .ZN(new_n2445_));
  INV_X1     g02189(.I(new_n2445_), .ZN(new_n2446_));
  NOR2_X1    g02190(.A1(new_n2446_), .A2(new_n2444_), .ZN(new_n2447_));
  NOR2_X1    g02191(.A1(new_n2447_), .A2(new_n258_), .ZN(new_n2448_));
  INV_X1     g02192(.I(new_n2295_), .ZN(new_n2449_));
  XNOR2_X1   g02193(.A1(\a[31] ), .A2(\a[32] ), .ZN(new_n2450_));
  NOR2_X1    g02194(.A1(new_n2449_), .A2(new_n2450_), .ZN(new_n2451_));
  INV_X1     g02195(.I(new_n2451_), .ZN(new_n2452_));
  NOR2_X1    g02196(.A1(new_n2452_), .A2(new_n267_), .ZN(new_n2453_));
  NOR2_X1    g02197(.A1(new_n2295_), .A2(new_n2450_), .ZN(new_n2454_));
  INV_X1     g02198(.I(new_n2454_), .ZN(new_n2455_));
  NOR4_X1    g02199(.A1(new_n2453_), .A2(new_n261_), .A3(new_n2448_), .A4(new_n2455_), .ZN(new_n2456_));
  XOR2_X1    g02200(.A1(new_n2456_), .A2(new_n2442_), .Z(new_n2457_));
  NOR2_X1    g02201(.A1(new_n2296_), .A2(new_n2442_), .ZN(new_n2458_));
  XNOR2_X1   g02202(.A1(new_n2457_), .A2(new_n2458_), .ZN(new_n2459_));
  XOR2_X1    g02203(.A1(new_n2459_), .A2(new_n2441_), .Z(new_n2460_));
  NOR2_X1    g02204(.A1(new_n2437_), .A2(new_n2460_), .ZN(new_n2461_));
  INV_X1     g02205(.I(new_n2437_), .ZN(new_n2462_));
  INV_X1     g02206(.I(new_n2441_), .ZN(new_n2463_));
  NOR2_X1    g02207(.A1(new_n2459_), .A2(new_n2463_), .ZN(new_n2464_));
  AND2_X2    g02208(.A1(new_n2459_), .A2(new_n2463_), .Z(new_n2465_));
  NOR2_X1    g02209(.A1(new_n2465_), .A2(new_n2464_), .ZN(new_n2466_));
  NOR2_X1    g02210(.A1(new_n2462_), .A2(new_n2466_), .ZN(new_n2467_));
  NOR2_X1    g02211(.A1(new_n2467_), .A2(new_n2461_), .ZN(new_n2468_));
  OAI22_X1   g02212(.A1(new_n1760_), .A2(new_n450_), .B1(new_n403_), .B2(new_n1755_), .ZN(new_n2469_));
  INV_X1     g02213(.I(new_n1857_), .ZN(new_n2470_));
  NAND2_X1   g02214(.A1(new_n2470_), .A2(\b[5] ), .ZN(new_n2471_));
  AOI21_X1   g02215(.A1(new_n2469_), .A2(new_n2471_), .B(new_n1763_), .ZN(new_n2472_));
  NAND2_X1   g02216(.A1(new_n454_), .A2(new_n2472_), .ZN(new_n2473_));
  XOR2_X1    g02217(.A1(new_n2473_), .A2(\a[26] ), .Z(new_n2474_));
  XOR2_X1    g02218(.A1(new_n2468_), .A2(new_n2474_), .Z(new_n2475_));
  AOI21_X1   g02219(.A1(new_n2316_), .A2(new_n2431_), .B(new_n2475_), .ZN(new_n2476_));
  NAND2_X1   g02220(.A1(new_n2316_), .A2(new_n2431_), .ZN(new_n2477_));
  INV_X1     g02221(.I(new_n2474_), .ZN(new_n2478_));
  NAND2_X1   g02222(.A1(new_n2468_), .A2(new_n2478_), .ZN(new_n2479_));
  NOR2_X1    g02223(.A1(new_n2468_), .A2(new_n2478_), .ZN(new_n2480_));
  INV_X1     g02224(.I(new_n2480_), .ZN(new_n2481_));
  AOI21_X1   g02225(.A1(new_n2479_), .A2(new_n2481_), .B(new_n2477_), .ZN(new_n2482_));
  NOR2_X1    g02226(.A1(new_n2482_), .A2(new_n2476_), .ZN(new_n2483_));
  OAI22_X1   g02227(.A1(new_n1444_), .A2(new_n617_), .B1(new_n510_), .B2(new_n1439_), .ZN(new_n2484_));
  NAND2_X1   g02228(.A1(new_n2098_), .A2(\b[8] ), .ZN(new_n2485_));
  AOI21_X1   g02229(.A1(new_n2484_), .A2(new_n2485_), .B(new_n1447_), .ZN(new_n2486_));
  NAND2_X1   g02230(.A1(new_n616_), .A2(new_n2486_), .ZN(new_n2487_));
  XOR2_X1    g02231(.A1(new_n2487_), .A2(\a[23] ), .Z(new_n2488_));
  XOR2_X1    g02232(.A1(new_n2483_), .A2(new_n2488_), .Z(new_n2489_));
  INV_X1     g02233(.I(new_n2483_), .ZN(new_n2490_));
  NOR2_X1    g02234(.A1(new_n2490_), .A2(new_n2488_), .ZN(new_n2491_));
  INV_X1     g02235(.I(new_n2488_), .ZN(new_n2492_));
  NOR2_X1    g02236(.A1(new_n2483_), .A2(new_n2492_), .ZN(new_n2493_));
  OAI21_X1   g02237(.A1(new_n2491_), .A2(new_n2493_), .B(new_n2427_), .ZN(new_n2494_));
  OAI21_X1   g02238(.A1(new_n2427_), .A2(new_n2489_), .B(new_n2494_), .ZN(new_n2495_));
  OAI22_X1   g02239(.A1(new_n1168_), .A2(new_n795_), .B1(new_n717_), .B2(new_n1163_), .ZN(new_n2496_));
  NAND2_X1   g02240(.A1(new_n1774_), .A2(\b[11] ), .ZN(new_n2497_));
  AOI21_X1   g02241(.A1(new_n2496_), .A2(new_n2497_), .B(new_n1171_), .ZN(new_n2498_));
  NAND2_X1   g02242(.A1(new_n799_), .A2(new_n2498_), .ZN(new_n2499_));
  XOR2_X1    g02243(.A1(new_n2499_), .A2(\a[20] ), .Z(new_n2500_));
  XNOR2_X1   g02244(.A1(new_n2495_), .A2(new_n2500_), .ZN(new_n2501_));
  OAI22_X1   g02245(.A1(new_n940_), .A2(new_n992_), .B1(new_n904_), .B2(new_n935_), .ZN(new_n2502_));
  NAND2_X1   g02246(.A1(new_n1458_), .A2(\b[14] ), .ZN(new_n2503_));
  AOI21_X1   g02247(.A1(new_n2502_), .A2(new_n2503_), .B(new_n943_), .ZN(new_n2504_));
  NAND2_X1   g02248(.A1(new_n991_), .A2(new_n2504_), .ZN(new_n2505_));
  XOR2_X1    g02249(.A1(new_n2505_), .A2(\a[17] ), .Z(new_n2506_));
  NOR2_X1    g02250(.A1(new_n2501_), .A2(new_n2506_), .ZN(new_n2507_));
  AND2_X2    g02251(.A1(new_n2501_), .A2(new_n2506_), .Z(new_n2508_));
  NOR2_X1    g02252(.A1(new_n2508_), .A2(new_n2507_), .ZN(new_n2509_));
  OAI22_X1   g02253(.A1(new_n757_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n752_), .ZN(new_n2510_));
  NAND2_X1   g02254(.A1(new_n1182_), .A2(\b[17] ), .ZN(new_n2511_));
  AOI21_X1   g02255(.A1(new_n2510_), .A2(new_n2511_), .B(new_n760_), .ZN(new_n2512_));
  NAND2_X1   g02256(.A1(new_n1225_), .A2(new_n2512_), .ZN(new_n2513_));
  XOR2_X1    g02257(.A1(new_n2513_), .A2(\a[14] ), .Z(new_n2514_));
  XNOR2_X1   g02258(.A1(new_n2509_), .A2(new_n2514_), .ZN(new_n2515_));
  OAI22_X1   g02259(.A1(new_n582_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n577_), .ZN(new_n2516_));
  NAND2_X1   g02260(.A1(new_n960_), .A2(\b[20] ), .ZN(new_n2517_));
  AOI21_X1   g02261(.A1(new_n2516_), .A2(new_n2517_), .B(new_n585_), .ZN(new_n2518_));
  NAND2_X1   g02262(.A1(new_n1517_), .A2(new_n2518_), .ZN(new_n2519_));
  XOR2_X1    g02263(.A1(new_n2519_), .A2(\a[11] ), .Z(new_n2520_));
  INV_X1     g02264(.I(new_n2520_), .ZN(new_n2521_));
  XOR2_X1    g02265(.A1(new_n2515_), .A2(new_n2521_), .Z(new_n2522_));
  OAI22_X1   g02266(.A1(new_n437_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n431_), .ZN(new_n2523_));
  NAND2_X1   g02267(.A1(new_n775_), .A2(\b[23] ), .ZN(new_n2524_));
  AOI21_X1   g02268(.A1(new_n2523_), .A2(new_n2524_), .B(new_n440_), .ZN(new_n2525_));
  NAND2_X1   g02269(.A1(new_n1828_), .A2(new_n2525_), .ZN(new_n2526_));
  XOR2_X1    g02270(.A1(new_n2526_), .A2(\a[8] ), .Z(new_n2527_));
  INV_X1     g02271(.I(new_n2527_), .ZN(new_n2528_));
  NAND2_X1   g02272(.A1(new_n2522_), .A2(new_n2528_), .ZN(new_n2529_));
  OR2_X2     g02273(.A1(new_n2522_), .A2(new_n2528_), .Z(new_n2530_));
  NAND2_X1   g02274(.A1(new_n2530_), .A2(new_n2529_), .ZN(new_n2531_));
  OAI22_X1   g02275(.A1(new_n364_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n320_), .ZN(new_n2532_));
  NAND2_X1   g02276(.A1(new_n594_), .A2(\b[26] ), .ZN(new_n2533_));
  AOI21_X1   g02277(.A1(new_n2532_), .A2(new_n2533_), .B(new_n312_), .ZN(new_n2534_));
  NAND2_X1   g02278(.A1(new_n2174_), .A2(new_n2534_), .ZN(new_n2535_));
  XOR2_X1    g02279(.A1(new_n2535_), .A2(\a[5] ), .Z(new_n2536_));
  XOR2_X1    g02280(.A1(new_n2531_), .A2(new_n2536_), .Z(new_n2537_));
  NAND2_X1   g02281(.A1(new_n2421_), .A2(new_n2537_), .ZN(new_n2538_));
  XOR2_X1    g02282(.A1(new_n2531_), .A2(new_n2536_), .Z(new_n2539_));
  OAI21_X1   g02283(.A1(new_n2421_), .A2(new_n2539_), .B(new_n2538_), .ZN(new_n2540_));
  NOR2_X1    g02284(.A1(new_n2387_), .A2(new_n2392_), .ZN(new_n2541_));
  XNOR2_X1   g02285(.A1(new_n2541_), .A2(new_n2540_), .ZN(new_n2542_));
  INV_X1     g02286(.I(\b[31] ), .ZN(new_n2543_));
  XOR2_X1    g02287(.A1(new_n2400_), .A2(\b[29] ), .Z(new_n2544_));
  NAND2_X1   g02288(.A1(new_n2544_), .A2(new_n2401_), .ZN(new_n2545_));
  XOR2_X1    g02289(.A1(new_n2545_), .A2(new_n2543_), .Z(new_n2546_));
  NAND2_X1   g02290(.A1(new_n283_), .A2(\b[31] ), .ZN(new_n2547_));
  NAND2_X1   g02291(.A1(new_n279_), .A2(\b[29] ), .ZN(new_n2548_));
  AOI21_X1   g02292(.A1(\b[30] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n2549_));
  NAND4_X1   g02293(.A1(new_n2546_), .A2(new_n2547_), .A3(new_n2548_), .A4(new_n2549_), .ZN(new_n2550_));
  XOR2_X1    g02294(.A1(new_n2550_), .A2(new_n271_), .Z(new_n2551_));
  NOR2_X1    g02295(.A1(new_n2542_), .A2(new_n2551_), .ZN(new_n2552_));
  XOR2_X1    g02296(.A1(new_n2550_), .A2(new_n271_), .Z(new_n2553_));
  AOI21_X1   g02297(.A1(new_n2542_), .A2(new_n2553_), .B(new_n2552_), .ZN(new_n2554_));
  NOR2_X1    g02298(.A1(new_n2396_), .A2(new_n2411_), .ZN(new_n2555_));
  AOI21_X1   g02299(.A1(new_n2412_), .A2(new_n2416_), .B(new_n2555_), .ZN(new_n2556_));
  XOR2_X1    g02300(.A1(new_n2554_), .A2(new_n2556_), .Z(\f[31] ));
  INV_X1     g02301(.I(new_n2542_), .ZN(new_n2558_));
  XOR2_X1    g02302(.A1(new_n2556_), .A2(new_n2553_), .Z(new_n2559_));
  AOI21_X1   g02303(.A1(new_n2558_), .A2(new_n2553_), .B(new_n2559_), .ZN(new_n2560_));
  OAI22_X1   g02304(.A1(new_n582_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n577_), .ZN(new_n2561_));
  NAND2_X1   g02305(.A1(new_n960_), .A2(\b[21] ), .ZN(new_n2562_));
  AOI21_X1   g02306(.A1(new_n2561_), .A2(new_n2562_), .B(new_n585_), .ZN(new_n2563_));
  NAND2_X1   g02307(.A1(new_n1604_), .A2(new_n2563_), .ZN(new_n2564_));
  XOR2_X1    g02308(.A1(new_n2564_), .A2(\a[11] ), .Z(new_n2565_));
  INV_X1     g02309(.I(new_n2565_), .ZN(new_n2566_));
  OAI22_X1   g02310(.A1(new_n757_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n752_), .ZN(new_n2567_));
  NAND2_X1   g02311(.A1(new_n1182_), .A2(\b[18] ), .ZN(new_n2568_));
  AOI21_X1   g02312(.A1(new_n2567_), .A2(new_n2568_), .B(new_n760_), .ZN(new_n2569_));
  NAND2_X1   g02313(.A1(new_n1304_), .A2(new_n2569_), .ZN(new_n2570_));
  XOR2_X1    g02314(.A1(new_n2570_), .A2(\a[14] ), .Z(new_n2571_));
  INV_X1     g02315(.I(new_n2571_), .ZN(new_n2572_));
  NOR3_X1    g02316(.A1(new_n2508_), .A2(new_n2507_), .A3(new_n2514_), .ZN(new_n2573_));
  OAI22_X1   g02317(.A1(new_n1168_), .A2(new_n848_), .B1(new_n795_), .B2(new_n1163_), .ZN(new_n2574_));
  NAND2_X1   g02318(.A1(new_n1774_), .A2(\b[12] ), .ZN(new_n2575_));
  AOI21_X1   g02319(.A1(new_n2574_), .A2(new_n2575_), .B(new_n1171_), .ZN(new_n2576_));
  NAND2_X1   g02320(.A1(new_n847_), .A2(new_n2576_), .ZN(new_n2577_));
  XOR2_X1    g02321(.A1(new_n2577_), .A2(\a[20] ), .Z(new_n2578_));
  OAI22_X1   g02322(.A1(new_n1444_), .A2(new_n659_), .B1(new_n617_), .B2(new_n1439_), .ZN(new_n2579_));
  NAND2_X1   g02323(.A1(new_n2098_), .A2(\b[9] ), .ZN(new_n2580_));
  AOI21_X1   g02324(.A1(new_n2579_), .A2(new_n2580_), .B(new_n1447_), .ZN(new_n2581_));
  NAND2_X1   g02325(.A1(new_n663_), .A2(new_n2581_), .ZN(new_n2582_));
  XOR2_X1    g02326(.A1(new_n2582_), .A2(\a[23] ), .Z(new_n2583_));
  INV_X1     g02327(.I(new_n2491_), .ZN(new_n2584_));
  OAI21_X1   g02328(.A1(new_n2427_), .A2(new_n2493_), .B(new_n2584_), .ZN(new_n2585_));
  OAI22_X1   g02329(.A1(new_n2084_), .A2(new_n347_), .B1(new_n393_), .B2(new_n2079_), .ZN(new_n2586_));
  OAI21_X1   g02330(.A1(new_n290_), .A2(new_n2214_), .B(new_n2586_), .ZN(new_n2587_));
  AOI21_X1   g02331(.A1(new_n352_), .A2(new_n2086_), .B(new_n2587_), .ZN(new_n2588_));
  XOR2_X1    g02332(.A1(new_n2588_), .A2(new_n2074_), .Z(new_n2589_));
  OAI22_X1   g02333(.A1(new_n1760_), .A2(new_n495_), .B1(new_n450_), .B2(new_n1755_), .ZN(new_n2590_));
  NAND2_X1   g02334(.A1(new_n2470_), .A2(\b[6] ), .ZN(new_n2591_));
  AOI21_X1   g02335(.A1(new_n2590_), .A2(new_n2591_), .B(new_n1763_), .ZN(new_n2592_));
  NAND2_X1   g02336(.A1(new_n494_), .A2(new_n2592_), .ZN(new_n2593_));
  XOR2_X1    g02337(.A1(new_n2593_), .A2(\a[26] ), .Z(new_n2594_));
  INV_X1     g02338(.I(new_n2465_), .ZN(new_n2595_));
  OAI21_X1   g02339(.A1(new_n2437_), .A2(new_n2464_), .B(new_n2595_), .ZN(new_n2596_));
  NAND2_X1   g02340(.A1(new_n2457_), .A2(new_n2458_), .ZN(new_n2597_));
  NOR2_X1    g02341(.A1(new_n2455_), .A2(new_n278_), .ZN(new_n2598_));
  XNOR2_X1   g02342(.A1(\a[29] ), .A2(\a[31] ), .ZN(new_n2599_));
  NAND2_X1   g02343(.A1(new_n2295_), .A2(new_n2599_), .ZN(new_n2600_));
  XNOR2_X1   g02344(.A1(\a[29] ), .A2(\a[32] ), .ZN(new_n2601_));
  NAND2_X1   g02345(.A1(new_n2600_), .A2(new_n2601_), .ZN(new_n2602_));
  OAI22_X1   g02346(.A1(new_n2452_), .A2(new_n292_), .B1(new_n267_), .B2(new_n2447_), .ZN(new_n2603_));
  NOR4_X1    g02347(.A1(new_n2603_), .A2(new_n258_), .A3(new_n2598_), .A4(new_n2602_), .ZN(new_n2604_));
  XOR2_X1    g02348(.A1(new_n2604_), .A2(new_n2442_), .Z(new_n2605_));
  XOR2_X1    g02349(.A1(new_n2597_), .A2(new_n2605_), .Z(new_n2606_));
  XOR2_X1    g02350(.A1(new_n2596_), .A2(new_n2606_), .Z(new_n2607_));
  XNOR2_X1   g02351(.A1(new_n2607_), .A2(new_n2594_), .ZN(new_n2608_));
  XOR2_X1    g02352(.A1(new_n2608_), .A2(new_n2589_), .Z(new_n2609_));
  OAI21_X1   g02353(.A1(new_n2477_), .A2(new_n2468_), .B(new_n2478_), .ZN(new_n2610_));
  XOR2_X1    g02354(.A1(new_n2609_), .A2(new_n2610_), .Z(new_n2611_));
  XOR2_X1    g02355(.A1(new_n2585_), .A2(new_n2611_), .Z(new_n2612_));
  XOR2_X1    g02356(.A1(new_n2612_), .A2(new_n2583_), .Z(new_n2613_));
  XOR2_X1    g02357(.A1(new_n2613_), .A2(new_n2578_), .Z(new_n2614_));
  NOR2_X1    g02358(.A1(new_n2495_), .A2(new_n2500_), .ZN(new_n2615_));
  XOR2_X1    g02359(.A1(new_n2614_), .A2(new_n2615_), .Z(new_n2616_));
  OAI22_X1   g02360(.A1(new_n940_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n935_), .ZN(new_n2617_));
  NAND2_X1   g02361(.A1(new_n1458_), .A2(\b[15] ), .ZN(new_n2618_));
  AOI21_X1   g02362(.A1(new_n2617_), .A2(new_n2618_), .B(new_n943_), .ZN(new_n2619_));
  NAND2_X1   g02363(.A1(new_n1047_), .A2(new_n2619_), .ZN(new_n2620_));
  XOR2_X1    g02364(.A1(new_n2620_), .A2(\a[17] ), .Z(new_n2621_));
  XOR2_X1    g02365(.A1(new_n2616_), .A2(new_n2621_), .Z(new_n2622_));
  NOR2_X1    g02366(.A1(new_n2501_), .A2(new_n2506_), .ZN(new_n2623_));
  INV_X1     g02367(.I(new_n2623_), .ZN(new_n2624_));
  XOR2_X1    g02368(.A1(new_n2622_), .A2(new_n2624_), .Z(new_n2625_));
  XOR2_X1    g02369(.A1(new_n2625_), .A2(new_n2573_), .Z(new_n2626_));
  XOR2_X1    g02370(.A1(new_n2626_), .A2(new_n2572_), .Z(new_n2627_));
  XOR2_X1    g02371(.A1(new_n2627_), .A2(new_n2566_), .Z(new_n2628_));
  NAND2_X1   g02372(.A1(new_n2515_), .A2(new_n2521_), .ZN(new_n2629_));
  XNOR2_X1   g02373(.A1(new_n2628_), .A2(new_n2629_), .ZN(new_n2630_));
  OAI22_X1   g02374(.A1(new_n437_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n431_), .ZN(new_n2631_));
  NAND2_X1   g02375(.A1(new_n775_), .A2(\b[24] ), .ZN(new_n2632_));
  AOI21_X1   g02376(.A1(new_n2631_), .A2(new_n2632_), .B(new_n440_), .ZN(new_n2633_));
  NAND2_X1   g02377(.A1(new_n1926_), .A2(new_n2633_), .ZN(new_n2634_));
  XOR2_X1    g02378(.A1(new_n2634_), .A2(\a[8] ), .Z(new_n2635_));
  INV_X1     g02379(.I(new_n2635_), .ZN(new_n2636_));
  XOR2_X1    g02380(.A1(new_n2630_), .A2(new_n2636_), .Z(new_n2637_));
  INV_X1     g02381(.I(new_n2637_), .ZN(new_n2638_));
  OAI21_X1   g02382(.A1(new_n2421_), .A2(new_n2531_), .B(new_n2530_), .ZN(new_n2639_));
  XOR2_X1    g02383(.A1(new_n2639_), .A2(new_n2638_), .Z(new_n2640_));
  OAI22_X1   g02384(.A1(new_n364_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n320_), .ZN(new_n2641_));
  NAND2_X1   g02385(.A1(new_n594_), .A2(\b[27] ), .ZN(new_n2642_));
  AOI21_X1   g02386(.A1(new_n2641_), .A2(new_n2642_), .B(new_n312_), .ZN(new_n2643_));
  NAND2_X1   g02387(.A1(new_n2276_), .A2(new_n2643_), .ZN(new_n2644_));
  XOR2_X1    g02388(.A1(new_n2644_), .A2(\a[5] ), .Z(new_n2645_));
  XOR2_X1    g02389(.A1(new_n2421_), .A2(new_n2531_), .Z(new_n2646_));
  NAND2_X1   g02390(.A1(new_n2646_), .A2(new_n2536_), .ZN(new_n2647_));
  NOR2_X1    g02391(.A1(new_n2540_), .A2(new_n2395_), .ZN(new_n2648_));
  NAND2_X1   g02392(.A1(new_n2647_), .A2(new_n2648_), .ZN(new_n2649_));
  XOR2_X1    g02393(.A1(new_n2649_), .A2(new_n2645_), .Z(new_n2650_));
  XNOR2_X1   g02394(.A1(new_n2650_), .A2(new_n2640_), .ZN(new_n2651_));
  OAI21_X1   g02395(.A1(new_n2272_), .A2(new_n2543_), .B(new_n2405_), .ZN(new_n2652_));
  NAND3_X1   g02396(.A1(new_n2398_), .A2(new_n2399_), .A3(new_n2652_), .ZN(new_n2653_));
  OAI21_X1   g02397(.A1(\b[29] ), .A2(\b[31] ), .B(\b[30] ), .ZN(new_n2654_));
  NAND2_X1   g02398(.A1(new_n2653_), .A2(new_n2654_), .ZN(new_n2655_));
  XOR2_X1    g02399(.A1(\b[31] ), .A2(\b[32] ), .Z(new_n2656_));
  NAND2_X1   g02400(.A1(new_n2655_), .A2(new_n2656_), .ZN(new_n2657_));
  XOR2_X1    g02401(.A1(\b[31] ), .A2(\b[32] ), .Z(new_n2658_));
  OAI21_X1   g02402(.A1(new_n2655_), .A2(new_n2658_), .B(new_n2657_), .ZN(new_n2659_));
  INV_X1     g02403(.I(\b[32] ), .ZN(new_n2660_));
  OAI22_X1   g02404(.A1(new_n405_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n404_), .ZN(new_n2661_));
  NAND2_X1   g02405(.A1(new_n279_), .A2(\b[30] ), .ZN(new_n2662_));
  AOI21_X1   g02406(.A1(new_n2661_), .A2(new_n2662_), .B(new_n264_), .ZN(new_n2663_));
  NAND2_X1   g02407(.A1(new_n2659_), .A2(new_n2663_), .ZN(new_n2664_));
  XOR2_X1    g02408(.A1(new_n2664_), .A2(new_n271_), .Z(new_n2665_));
  XNOR2_X1   g02409(.A1(new_n2651_), .A2(new_n2665_), .ZN(new_n2666_));
  NAND2_X1   g02410(.A1(new_n2666_), .A2(new_n2560_), .ZN(new_n2667_));
  XNOR2_X1   g02411(.A1(new_n2651_), .A2(new_n2665_), .ZN(new_n2668_));
  OAI21_X1   g02412(.A1(new_n2560_), .A2(new_n2668_), .B(new_n2667_), .ZN(\f[32] ));
  INV_X1     g02413(.I(new_n2079_), .ZN(new_n2670_));
  AOI22_X1   g02414(.A1(\b[6] ), .A2(new_n2083_), .B1(new_n2670_), .B2(\b[5] ), .ZN(new_n2671_));
  NOR2_X1    g02415(.A1(new_n2214_), .A2(new_n393_), .ZN(new_n2672_));
  OAI21_X1   g02416(.A1(new_n2671_), .A2(new_n2672_), .B(new_n2086_), .ZN(new_n2673_));
  NOR2_X1    g02417(.A1(new_n524_), .A2(new_n2673_), .ZN(new_n2674_));
  XOR2_X1    g02418(.A1(new_n2674_), .A2(\a[29] ), .Z(new_n2675_));
  XNOR2_X1   g02419(.A1(\a[32] ), .A2(\a[33] ), .ZN(new_n2676_));
  NOR2_X1    g02420(.A1(new_n2676_), .A2(new_n258_), .ZN(new_n2677_));
  INV_X1     g02421(.I(new_n2605_), .ZN(new_n2678_));
  NOR2_X1    g02422(.A1(new_n2678_), .A2(new_n2597_), .ZN(new_n2679_));
  NOR2_X1    g02423(.A1(new_n2602_), .A2(new_n267_), .ZN(new_n2680_));
  OAI22_X1   g02424(.A1(new_n2452_), .A2(new_n290_), .B1(new_n292_), .B2(new_n2447_), .ZN(new_n2681_));
  NOR4_X1    g02425(.A1(new_n2681_), .A2(new_n677_), .A3(new_n2455_), .A4(new_n2680_), .ZN(new_n2682_));
  XOR2_X1    g02426(.A1(new_n2682_), .A2(new_n2442_), .Z(new_n2683_));
  XOR2_X1    g02427(.A1(new_n2679_), .A2(new_n2683_), .Z(new_n2684_));
  XOR2_X1    g02428(.A1(new_n2684_), .A2(new_n2677_), .Z(new_n2685_));
  XOR2_X1    g02429(.A1(new_n2685_), .A2(new_n2675_), .Z(new_n2686_));
  INV_X1     g02430(.I(new_n2589_), .ZN(new_n2687_));
  XOR2_X1    g02431(.A1(new_n2437_), .A2(new_n2441_), .Z(new_n2688_));
  INV_X1     g02432(.I(new_n2597_), .ZN(new_n2689_));
  NOR2_X1    g02433(.A1(new_n2689_), .A2(new_n2605_), .ZN(new_n2690_));
  NOR2_X1    g02434(.A1(new_n2690_), .A2(new_n2679_), .ZN(new_n2691_));
  XOR2_X1    g02435(.A1(new_n2691_), .A2(\a[29] ), .Z(new_n2692_));
  OAI21_X1   g02436(.A1(new_n2692_), .A2(new_n2588_), .B(new_n2463_), .ZN(new_n2693_));
  AOI21_X1   g02437(.A1(new_n2588_), .A2(new_n2692_), .B(new_n2693_), .ZN(new_n2694_));
  NAND2_X1   g02438(.A1(new_n2694_), .A2(new_n2462_), .ZN(new_n2695_));
  NAND3_X1   g02439(.A1(new_n2695_), .A2(new_n2459_), .A3(new_n2688_), .ZN(new_n2696_));
  OAI21_X1   g02440(.A1(new_n2687_), .A2(new_n2606_), .B(new_n2696_), .ZN(new_n2697_));
  NAND2_X1   g02441(.A1(new_n2697_), .A2(new_n2686_), .ZN(new_n2698_));
  NOR2_X1    g02442(.A1(new_n2687_), .A2(new_n2606_), .ZN(new_n2699_));
  NOR2_X1    g02443(.A1(new_n2686_), .A2(new_n2699_), .ZN(new_n2700_));
  NAND2_X1   g02444(.A1(new_n2696_), .A2(new_n2700_), .ZN(new_n2701_));
  NAND2_X1   g02445(.A1(new_n2698_), .A2(new_n2701_), .ZN(new_n2702_));
  OAI22_X1   g02446(.A1(new_n1760_), .A2(new_n510_), .B1(new_n495_), .B2(new_n1755_), .ZN(new_n2703_));
  NAND2_X1   g02447(.A1(new_n2470_), .A2(\b[7] ), .ZN(new_n2704_));
  AOI21_X1   g02448(.A1(new_n2703_), .A2(new_n2704_), .B(new_n1763_), .ZN(new_n2705_));
  NAND2_X1   g02449(.A1(new_n518_), .A2(new_n2705_), .ZN(new_n2706_));
  XOR2_X1    g02450(.A1(new_n2706_), .A2(\a[26] ), .Z(new_n2707_));
  NOR2_X1    g02451(.A1(new_n2477_), .A2(new_n2481_), .ZN(new_n2708_));
  NOR3_X1    g02452(.A1(new_n2609_), .A2(new_n2708_), .A3(new_n2480_), .ZN(new_n2709_));
  XOR2_X1    g02453(.A1(new_n2606_), .A2(new_n2589_), .Z(new_n2710_));
  XOR2_X1    g02454(.A1(new_n2596_), .A2(new_n2710_), .Z(new_n2711_));
  NAND2_X1   g02455(.A1(new_n2711_), .A2(new_n2594_), .ZN(new_n2712_));
  NAND2_X1   g02456(.A1(new_n2709_), .A2(new_n2712_), .ZN(new_n2713_));
  XOR2_X1    g02457(.A1(new_n2713_), .A2(new_n2707_), .Z(new_n2714_));
  XOR2_X1    g02458(.A1(new_n2714_), .A2(new_n2702_), .Z(new_n2715_));
  OAI22_X1   g02459(.A1(new_n1444_), .A2(new_n717_), .B1(new_n659_), .B2(new_n1439_), .ZN(new_n2716_));
  NAND2_X1   g02460(.A1(new_n2098_), .A2(\b[10] ), .ZN(new_n2717_));
  AOI21_X1   g02461(.A1(new_n2716_), .A2(new_n2717_), .B(new_n1447_), .ZN(new_n2718_));
  NAND2_X1   g02462(.A1(new_n716_), .A2(new_n2718_), .ZN(new_n2719_));
  XOR2_X1    g02463(.A1(new_n2719_), .A2(\a[23] ), .Z(new_n2720_));
  INV_X1     g02464(.I(new_n2583_), .ZN(new_n2721_));
  XOR2_X1    g02465(.A1(new_n2427_), .A2(new_n2492_), .Z(new_n2722_));
  XOR2_X1    g02466(.A1(new_n2611_), .A2(new_n2721_), .Z(new_n2723_));
  OR3_X2     g02467(.A1(new_n2427_), .A2(new_n2488_), .A3(new_n2723_), .Z(new_n2724_));
  NAND2_X1   g02468(.A1(new_n2724_), .A2(new_n2483_), .ZN(new_n2725_));
  OAI22_X1   g02469(.A1(new_n2725_), .A2(new_n2722_), .B1(new_n2721_), .B2(new_n2611_), .ZN(new_n2726_));
  XOR2_X1    g02470(.A1(new_n2726_), .A2(new_n2720_), .Z(new_n2727_));
  XNOR2_X1   g02471(.A1(new_n2727_), .A2(new_n2715_), .ZN(new_n2728_));
  OAI22_X1   g02472(.A1(new_n1168_), .A2(new_n904_), .B1(new_n848_), .B2(new_n1163_), .ZN(new_n2729_));
  NAND2_X1   g02473(.A1(new_n1774_), .A2(\b[13] ), .ZN(new_n2730_));
  AOI21_X1   g02474(.A1(new_n2729_), .A2(new_n2730_), .B(new_n1171_), .ZN(new_n2731_));
  NAND2_X1   g02475(.A1(new_n907_), .A2(new_n2731_), .ZN(new_n2732_));
  XOR2_X1    g02476(.A1(new_n2732_), .A2(new_n1158_), .Z(new_n2733_));
  XOR2_X1    g02477(.A1(new_n2611_), .A2(new_n2583_), .Z(new_n2734_));
  XOR2_X1    g02478(.A1(new_n2585_), .A2(new_n2734_), .Z(new_n2735_));
  AOI21_X1   g02479(.A1(new_n2578_), .A2(new_n2735_), .B(new_n2615_), .ZN(new_n2736_));
  XOR2_X1    g02480(.A1(new_n2736_), .A2(new_n2733_), .Z(new_n2737_));
  XNOR2_X1   g02481(.A1(new_n2728_), .A2(new_n2737_), .ZN(new_n2738_));
  OAI22_X1   g02482(.A1(new_n940_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n935_), .ZN(new_n2739_));
  NAND2_X1   g02483(.A1(new_n1458_), .A2(\b[16] ), .ZN(new_n2740_));
  AOI21_X1   g02484(.A1(new_n2739_), .A2(new_n2740_), .B(new_n943_), .ZN(new_n2741_));
  NAND2_X1   g02485(.A1(new_n1123_), .A2(new_n2741_), .ZN(new_n2742_));
  XOR2_X1    g02486(.A1(new_n2742_), .A2(\a[17] ), .Z(new_n2743_));
  INV_X1     g02487(.I(new_n2621_), .ZN(new_n2744_));
  NOR2_X1    g02488(.A1(new_n2616_), .A2(new_n2744_), .ZN(new_n2745_));
  NOR3_X1    g02489(.A1(new_n2622_), .A2(new_n2745_), .A3(new_n2623_), .ZN(new_n2746_));
  XOR2_X1    g02490(.A1(new_n2746_), .A2(new_n2743_), .Z(new_n2747_));
  XOR2_X1    g02491(.A1(new_n2747_), .A2(new_n2738_), .Z(new_n2748_));
  OAI22_X1   g02492(.A1(new_n757_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n752_), .ZN(new_n2749_));
  NAND2_X1   g02493(.A1(new_n1182_), .A2(\b[19] ), .ZN(new_n2750_));
  AOI21_X1   g02494(.A1(new_n2749_), .A2(new_n2750_), .B(new_n760_), .ZN(new_n2751_));
  NAND2_X1   g02495(.A1(new_n1396_), .A2(new_n2751_), .ZN(new_n2752_));
  XOR2_X1    g02496(.A1(new_n2752_), .A2(\a[14] ), .Z(new_n2753_));
  NAND2_X1   g02497(.A1(new_n2625_), .A2(new_n2571_), .ZN(new_n2754_));
  OR2_X2     g02498(.A1(new_n2625_), .A2(new_n2571_), .Z(new_n2755_));
  NAND3_X1   g02499(.A1(new_n2755_), .A2(new_n2754_), .A3(new_n2573_), .ZN(new_n2756_));
  OAI21_X1   g02500(.A1(new_n2572_), .A2(new_n2625_), .B(new_n2756_), .ZN(new_n2757_));
  XOR2_X1    g02501(.A1(new_n2757_), .A2(new_n2753_), .Z(new_n2758_));
  XNOR2_X1   g02502(.A1(new_n2758_), .A2(new_n2748_), .ZN(new_n2759_));
  INV_X1     g02503(.I(new_n2759_), .ZN(new_n2760_));
  OAI22_X1   g02504(.A1(new_n582_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n577_), .ZN(new_n2761_));
  NAND2_X1   g02505(.A1(new_n960_), .A2(\b[22] ), .ZN(new_n2762_));
  AOI21_X1   g02506(.A1(new_n2761_), .A2(new_n2762_), .B(new_n585_), .ZN(new_n2763_));
  NAND2_X1   g02507(.A1(new_n1708_), .A2(new_n2763_), .ZN(new_n2764_));
  XOR2_X1    g02508(.A1(new_n2764_), .A2(\a[11] ), .Z(new_n2765_));
  INV_X1     g02509(.I(new_n2628_), .ZN(new_n2766_));
  NOR2_X1    g02510(.A1(new_n2766_), .A2(new_n2629_), .ZN(new_n2767_));
  INV_X1     g02511(.I(new_n2767_), .ZN(new_n2768_));
  XOR2_X1    g02512(.A1(new_n2625_), .A2(new_n2572_), .Z(new_n2769_));
  XOR2_X1    g02513(.A1(new_n2769_), .A2(new_n2573_), .Z(new_n2770_));
  OAI21_X1   g02514(.A1(new_n2566_), .A2(new_n2770_), .B(new_n2768_), .ZN(new_n2771_));
  XOR2_X1    g02515(.A1(new_n2771_), .A2(new_n2765_), .Z(new_n2772_));
  XOR2_X1    g02516(.A1(new_n2772_), .A2(new_n2760_), .Z(new_n2773_));
  OAI22_X1   g02517(.A1(new_n437_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n431_), .ZN(new_n2774_));
  NAND2_X1   g02518(.A1(new_n775_), .A2(\b[25] ), .ZN(new_n2775_));
  AOI21_X1   g02519(.A1(new_n2774_), .A2(new_n2775_), .B(new_n440_), .ZN(new_n2776_));
  NAND2_X1   g02520(.A1(new_n2042_), .A2(new_n2776_), .ZN(new_n2777_));
  XOR2_X1    g02521(.A1(new_n2777_), .A2(\a[8] ), .Z(new_n2778_));
  NOR2_X1    g02522(.A1(new_n2630_), .A2(new_n2636_), .ZN(new_n2779_));
  NOR2_X1    g02523(.A1(new_n2638_), .A2(new_n2779_), .ZN(new_n2780_));
  NAND2_X1   g02524(.A1(new_n2639_), .A2(new_n2780_), .ZN(new_n2781_));
  XOR2_X1    g02525(.A1(new_n2781_), .A2(new_n2778_), .Z(new_n2782_));
  XNOR2_X1   g02526(.A1(new_n2782_), .A2(new_n2773_), .ZN(new_n2783_));
  INV_X1     g02527(.I(new_n2783_), .ZN(new_n2784_));
  OAI22_X1   g02528(.A1(new_n364_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n320_), .ZN(new_n2785_));
  NAND2_X1   g02529(.A1(new_n594_), .A2(\b[28] ), .ZN(new_n2786_));
  AOI21_X1   g02530(.A1(new_n2785_), .A2(new_n2786_), .B(new_n312_), .ZN(new_n2787_));
  NAND2_X1   g02531(.A1(new_n2404_), .A2(new_n2787_), .ZN(new_n2788_));
  XOR2_X1    g02532(.A1(new_n2788_), .A2(\a[5] ), .Z(new_n2789_));
  NOR2_X1    g02533(.A1(new_n2784_), .A2(new_n2789_), .ZN(new_n2790_));
  INV_X1     g02534(.I(new_n2790_), .ZN(new_n2791_));
  NAND2_X1   g02535(.A1(new_n2784_), .A2(new_n2789_), .ZN(new_n2792_));
  NAND2_X1   g02536(.A1(new_n2791_), .A2(new_n2792_), .ZN(new_n2793_));
  INV_X1     g02537(.I(\b[33] ), .ZN(new_n2794_));
  XOR2_X1    g02538(.A1(new_n2655_), .A2(\b[31] ), .Z(new_n2795_));
  NAND2_X1   g02539(.A1(new_n2795_), .A2(new_n2656_), .ZN(new_n2796_));
  XOR2_X1    g02540(.A1(new_n2796_), .A2(new_n2794_), .Z(new_n2797_));
  NAND2_X1   g02541(.A1(new_n283_), .A2(\b[33] ), .ZN(new_n2798_));
  NAND2_X1   g02542(.A1(new_n279_), .A2(\b[31] ), .ZN(new_n2799_));
  AOI21_X1   g02543(.A1(\b[32] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n2800_));
  NAND4_X1   g02544(.A1(new_n2797_), .A2(new_n2798_), .A3(new_n2799_), .A4(new_n2800_), .ZN(new_n2801_));
  XOR2_X1    g02545(.A1(new_n2801_), .A2(\a[2] ), .Z(new_n2802_));
  XNOR2_X1   g02546(.A1(new_n2793_), .A2(new_n2802_), .ZN(new_n2803_));
  INV_X1     g02547(.I(new_n2651_), .ZN(new_n2804_));
  NAND2_X1   g02548(.A1(new_n2560_), .A2(new_n2804_), .ZN(new_n2805_));
  XOR2_X1    g02549(.A1(new_n2803_), .A2(new_n2805_), .Z(new_n2806_));
  XOR2_X1    g02550(.A1(new_n2560_), .A2(new_n2804_), .Z(new_n2807_));
  NAND2_X1   g02551(.A1(new_n2807_), .A2(new_n2665_), .ZN(new_n2808_));
  XNOR2_X1   g02552(.A1(new_n2806_), .A2(new_n2808_), .ZN(\f[33] ));
  NAND2_X1   g02553(.A1(new_n2760_), .A2(new_n2765_), .ZN(new_n2810_));
  INV_X1     g02554(.I(new_n2771_), .ZN(new_n2811_));
  XOR2_X1    g02555(.A1(new_n2759_), .A2(new_n2765_), .Z(new_n2812_));
  NAND2_X1   g02556(.A1(new_n2811_), .A2(new_n2812_), .ZN(new_n2813_));
  NAND2_X1   g02557(.A1(new_n2813_), .A2(new_n2810_), .ZN(new_n2814_));
  INV_X1     g02558(.I(new_n2814_), .ZN(new_n2815_));
  XNOR2_X1   g02559(.A1(new_n2738_), .A2(new_n2743_), .ZN(new_n2816_));
  INV_X1     g02560(.I(new_n2816_), .ZN(new_n2817_));
  OAI21_X1   g02561(.A1(new_n2746_), .A2(new_n2743_), .B(new_n2817_), .ZN(new_n2818_));
  NAND2_X1   g02562(.A1(new_n2702_), .A2(new_n2707_), .ZN(new_n2819_));
  XNOR2_X1   g02563(.A1(new_n2702_), .A2(new_n2707_), .ZN(new_n2820_));
  NAND3_X1   g02564(.A1(new_n2820_), .A2(new_n2709_), .A3(new_n2712_), .ZN(new_n2821_));
  XOR2_X1    g02565(.A1(new_n2683_), .A2(new_n2677_), .Z(new_n2822_));
  AND2_X2    g02566(.A1(new_n2822_), .A2(new_n2679_), .Z(new_n2823_));
  NOR2_X1    g02567(.A1(new_n2822_), .A2(new_n2679_), .ZN(new_n2824_));
  NOR3_X1    g02568(.A1(new_n2823_), .A2(new_n2824_), .A3(new_n2675_), .ZN(new_n2825_));
  AOI21_X1   g02569(.A1(new_n2822_), .A2(new_n2605_), .B(new_n2689_), .ZN(new_n2826_));
  NAND2_X1   g02570(.A1(new_n2683_), .A2(new_n2677_), .ZN(new_n2827_));
  NOR2_X1    g02571(.A1(new_n2826_), .A2(new_n2827_), .ZN(new_n2828_));
  NAND2_X1   g02572(.A1(new_n2826_), .A2(new_n2827_), .ZN(new_n2829_));
  INV_X1     g02573(.I(new_n2829_), .ZN(new_n2830_));
  NOR2_X1    g02574(.A1(new_n2830_), .A2(new_n2828_), .ZN(new_n2831_));
  OAI22_X1   g02575(.A1(new_n2452_), .A2(new_n393_), .B1(new_n290_), .B2(new_n2447_), .ZN(new_n2832_));
  OAI21_X1   g02576(.A1(new_n292_), .A2(new_n2602_), .B(new_n2832_), .ZN(new_n2833_));
  NAND3_X1   g02577(.A1(new_n2833_), .A2(new_n334_), .A3(new_n2454_), .ZN(new_n2834_));
  XOR2_X1    g02578(.A1(new_n2834_), .A2(\a[32] ), .Z(new_n2835_));
  INV_X1     g02579(.I(\a[35] ), .ZN(new_n2836_));
  INV_X1     g02580(.I(\a[34] ), .ZN(new_n2837_));
  NOR3_X1    g02581(.A1(new_n2837_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n2838_));
  NAND3_X1   g02582(.A1(new_n2837_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n2839_));
  INV_X1     g02583(.I(new_n2839_), .ZN(new_n2840_));
  NOR2_X1    g02584(.A1(new_n2840_), .A2(new_n2838_), .ZN(new_n2841_));
  NOR2_X1    g02585(.A1(new_n2841_), .A2(new_n258_), .ZN(new_n2842_));
  INV_X1     g02586(.I(new_n2676_), .ZN(new_n2843_));
  XNOR2_X1   g02587(.A1(\a[34] ), .A2(\a[35] ), .ZN(new_n2844_));
  NOR2_X1    g02588(.A1(new_n2843_), .A2(new_n2844_), .ZN(new_n2845_));
  INV_X1     g02589(.I(new_n2845_), .ZN(new_n2846_));
  NOR2_X1    g02590(.A1(new_n2846_), .A2(new_n267_), .ZN(new_n2847_));
  NOR2_X1    g02591(.A1(new_n2676_), .A2(new_n2844_), .ZN(new_n2848_));
  INV_X1     g02592(.I(new_n2848_), .ZN(new_n2849_));
  NOR4_X1    g02593(.A1(new_n2847_), .A2(new_n261_), .A3(new_n2842_), .A4(new_n2849_), .ZN(new_n2850_));
  XOR2_X1    g02594(.A1(new_n2850_), .A2(new_n2836_), .Z(new_n2851_));
  NOR2_X1    g02595(.A1(new_n2677_), .A2(new_n2836_), .ZN(new_n2852_));
  XNOR2_X1   g02596(.A1(new_n2851_), .A2(new_n2852_), .ZN(new_n2853_));
  XOR2_X1    g02597(.A1(new_n2853_), .A2(new_n2835_), .Z(new_n2854_));
  NOR2_X1    g02598(.A1(new_n2831_), .A2(new_n2854_), .ZN(new_n2855_));
  INV_X1     g02599(.I(new_n2831_), .ZN(new_n2856_));
  INV_X1     g02600(.I(new_n2835_), .ZN(new_n2857_));
  NOR2_X1    g02601(.A1(new_n2853_), .A2(new_n2857_), .ZN(new_n2858_));
  AND2_X2    g02602(.A1(new_n2853_), .A2(new_n2857_), .Z(new_n2859_));
  NOR2_X1    g02603(.A1(new_n2859_), .A2(new_n2858_), .ZN(new_n2860_));
  NOR2_X1    g02604(.A1(new_n2856_), .A2(new_n2860_), .ZN(new_n2861_));
  NOR2_X1    g02605(.A1(new_n2861_), .A2(new_n2855_), .ZN(new_n2862_));
  OAI22_X1   g02606(.A1(new_n2084_), .A2(new_n450_), .B1(new_n403_), .B2(new_n2079_), .ZN(new_n2863_));
  INV_X1     g02607(.I(new_n2214_), .ZN(new_n2864_));
  NAND2_X1   g02608(.A1(new_n2864_), .A2(\b[5] ), .ZN(new_n2865_));
  AOI21_X1   g02609(.A1(new_n2863_), .A2(new_n2865_), .B(new_n2087_), .ZN(new_n2866_));
  NAND2_X1   g02610(.A1(new_n454_), .A2(new_n2866_), .ZN(new_n2867_));
  XOR2_X1    g02611(.A1(new_n2867_), .A2(\a[29] ), .Z(new_n2868_));
  XOR2_X1    g02612(.A1(new_n2862_), .A2(new_n2868_), .Z(new_n2869_));
  AOI21_X1   g02613(.A1(new_n2698_), .A2(new_n2825_), .B(new_n2869_), .ZN(new_n2870_));
  NAND2_X1   g02614(.A1(new_n2698_), .A2(new_n2825_), .ZN(new_n2871_));
  INV_X1     g02615(.I(new_n2868_), .ZN(new_n2872_));
  NAND2_X1   g02616(.A1(new_n2862_), .A2(new_n2872_), .ZN(new_n2873_));
  NOR2_X1    g02617(.A1(new_n2862_), .A2(new_n2872_), .ZN(new_n2874_));
  INV_X1     g02618(.I(new_n2874_), .ZN(new_n2875_));
  AOI21_X1   g02619(.A1(new_n2873_), .A2(new_n2875_), .B(new_n2871_), .ZN(new_n2876_));
  NOR2_X1    g02620(.A1(new_n2876_), .A2(new_n2870_), .ZN(new_n2877_));
  OAI22_X1   g02621(.A1(new_n1760_), .A2(new_n617_), .B1(new_n510_), .B2(new_n1755_), .ZN(new_n2878_));
  NAND2_X1   g02622(.A1(new_n2470_), .A2(\b[8] ), .ZN(new_n2879_));
  AOI21_X1   g02623(.A1(new_n2878_), .A2(new_n2879_), .B(new_n1763_), .ZN(new_n2880_));
  NAND2_X1   g02624(.A1(new_n616_), .A2(new_n2880_), .ZN(new_n2881_));
  XOR2_X1    g02625(.A1(new_n2881_), .A2(\a[26] ), .Z(new_n2882_));
  XOR2_X1    g02626(.A1(new_n2877_), .A2(new_n2882_), .Z(new_n2883_));
  AOI21_X1   g02627(.A1(new_n2819_), .A2(new_n2821_), .B(new_n2883_), .ZN(new_n2884_));
  NAND2_X1   g02628(.A1(new_n2821_), .A2(new_n2819_), .ZN(new_n2885_));
  INV_X1     g02629(.I(new_n2882_), .ZN(new_n2886_));
  NAND2_X1   g02630(.A1(new_n2877_), .A2(new_n2886_), .ZN(new_n2887_));
  OAI21_X1   g02631(.A1(new_n2876_), .A2(new_n2870_), .B(new_n2882_), .ZN(new_n2888_));
  AOI21_X1   g02632(.A1(new_n2887_), .A2(new_n2888_), .B(new_n2885_), .ZN(new_n2889_));
  NOR2_X1    g02633(.A1(new_n2884_), .A2(new_n2889_), .ZN(new_n2890_));
  OAI22_X1   g02634(.A1(new_n1444_), .A2(new_n795_), .B1(new_n717_), .B2(new_n1439_), .ZN(new_n2891_));
  NAND2_X1   g02635(.A1(new_n2098_), .A2(\b[11] ), .ZN(new_n2892_));
  AOI21_X1   g02636(.A1(new_n2891_), .A2(new_n2892_), .B(new_n1447_), .ZN(new_n2893_));
  NAND2_X1   g02637(.A1(new_n799_), .A2(new_n2893_), .ZN(new_n2894_));
  XOR2_X1    g02638(.A1(new_n2894_), .A2(\a[23] ), .Z(new_n2895_));
  XOR2_X1    g02639(.A1(new_n2890_), .A2(new_n2895_), .Z(new_n2896_));
  OAI22_X1   g02640(.A1(new_n1168_), .A2(new_n992_), .B1(new_n904_), .B2(new_n1163_), .ZN(new_n2897_));
  NAND2_X1   g02641(.A1(new_n1774_), .A2(\b[14] ), .ZN(new_n2898_));
  AOI21_X1   g02642(.A1(new_n2897_), .A2(new_n2898_), .B(new_n1171_), .ZN(new_n2899_));
  NAND2_X1   g02643(.A1(new_n991_), .A2(new_n2899_), .ZN(new_n2900_));
  XOR2_X1    g02644(.A1(new_n2900_), .A2(\a[20] ), .Z(new_n2901_));
  NOR2_X1    g02645(.A1(new_n2896_), .A2(new_n2901_), .ZN(new_n2902_));
  INV_X1     g02646(.I(new_n2902_), .ZN(new_n2903_));
  NAND2_X1   g02647(.A1(new_n2896_), .A2(new_n2901_), .ZN(new_n2904_));
  NAND2_X1   g02648(.A1(new_n2903_), .A2(new_n2904_), .ZN(new_n2905_));
  OAI22_X1   g02649(.A1(new_n940_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n935_), .ZN(new_n2906_));
  NAND2_X1   g02650(.A1(new_n1458_), .A2(\b[17] ), .ZN(new_n2907_));
  AOI21_X1   g02651(.A1(new_n2906_), .A2(new_n2907_), .B(new_n943_), .ZN(new_n2908_));
  NAND2_X1   g02652(.A1(new_n1225_), .A2(new_n2908_), .ZN(new_n2909_));
  XOR2_X1    g02653(.A1(new_n2909_), .A2(\a[17] ), .Z(new_n2910_));
  XNOR2_X1   g02654(.A1(new_n2905_), .A2(new_n2910_), .ZN(new_n2911_));
  OAI22_X1   g02655(.A1(new_n757_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n752_), .ZN(new_n2912_));
  NAND2_X1   g02656(.A1(new_n1182_), .A2(\b[20] ), .ZN(new_n2913_));
  AOI21_X1   g02657(.A1(new_n2912_), .A2(new_n2913_), .B(new_n760_), .ZN(new_n2914_));
  NAND2_X1   g02658(.A1(new_n1517_), .A2(new_n2914_), .ZN(new_n2915_));
  XOR2_X1    g02659(.A1(new_n2915_), .A2(\a[14] ), .Z(new_n2916_));
  INV_X1     g02660(.I(new_n2916_), .ZN(new_n2917_));
  XOR2_X1    g02661(.A1(new_n2911_), .A2(new_n2917_), .Z(new_n2918_));
  NOR2_X1    g02662(.A1(new_n2818_), .A2(new_n2918_), .ZN(new_n2919_));
  INV_X1     g02663(.I(new_n2818_), .ZN(new_n2920_));
  XOR2_X1    g02664(.A1(new_n2911_), .A2(new_n2916_), .Z(new_n2921_));
  NOR2_X1    g02665(.A1(new_n2920_), .A2(new_n2921_), .ZN(new_n2922_));
  NOR2_X1    g02666(.A1(new_n2922_), .A2(new_n2919_), .ZN(new_n2923_));
  INV_X1     g02667(.I(new_n2923_), .ZN(new_n2924_));
  OAI22_X1   g02668(.A1(new_n582_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n577_), .ZN(new_n2925_));
  NAND2_X1   g02669(.A1(new_n960_), .A2(\b[23] ), .ZN(new_n2926_));
  AOI21_X1   g02670(.A1(new_n2925_), .A2(new_n2926_), .B(new_n585_), .ZN(new_n2927_));
  NAND2_X1   g02671(.A1(new_n1828_), .A2(new_n2927_), .ZN(new_n2928_));
  XOR2_X1    g02672(.A1(new_n2928_), .A2(\a[11] ), .Z(new_n2929_));
  NOR2_X1    g02673(.A1(new_n2924_), .A2(new_n2929_), .ZN(new_n2930_));
  INV_X1     g02674(.I(new_n2929_), .ZN(new_n2931_));
  NOR2_X1    g02675(.A1(new_n2923_), .A2(new_n2931_), .ZN(new_n2932_));
  NOR2_X1    g02676(.A1(new_n2930_), .A2(new_n2932_), .ZN(new_n2933_));
  NOR2_X1    g02677(.A1(new_n2815_), .A2(new_n2933_), .ZN(new_n2934_));
  XOR2_X1    g02678(.A1(new_n2923_), .A2(new_n2929_), .Z(new_n2935_));
  NOR2_X1    g02679(.A1(new_n2814_), .A2(new_n2935_), .ZN(new_n2936_));
  NOR2_X1    g02680(.A1(new_n2934_), .A2(new_n2936_), .ZN(new_n2937_));
  OAI22_X1   g02681(.A1(new_n437_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n431_), .ZN(new_n2938_));
  NAND2_X1   g02682(.A1(new_n775_), .A2(\b[26] ), .ZN(new_n2939_));
  AOI21_X1   g02683(.A1(new_n2938_), .A2(new_n2939_), .B(new_n440_), .ZN(new_n2940_));
  NAND2_X1   g02684(.A1(new_n2174_), .A2(new_n2940_), .ZN(new_n2941_));
  XOR2_X1    g02685(.A1(new_n2941_), .A2(\a[8] ), .Z(new_n2942_));
  XNOR2_X1   g02686(.A1(new_n2937_), .A2(new_n2942_), .ZN(new_n2943_));
  OAI22_X1   g02687(.A1(new_n364_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n320_), .ZN(new_n2944_));
  NAND2_X1   g02688(.A1(new_n594_), .A2(\b[29] ), .ZN(new_n2945_));
  AOI21_X1   g02689(.A1(new_n2944_), .A2(new_n2945_), .B(new_n312_), .ZN(new_n2946_));
  NAND2_X1   g02690(.A1(new_n2546_), .A2(new_n2946_), .ZN(new_n2947_));
  XOR2_X1    g02691(.A1(new_n2947_), .A2(\a[5] ), .Z(new_n2948_));
  XOR2_X1    g02692(.A1(new_n2943_), .A2(new_n2948_), .Z(new_n2949_));
  NOR2_X1    g02693(.A1(new_n2791_), .A2(new_n2949_), .ZN(new_n2950_));
  XNOR2_X1   g02694(.A1(new_n2943_), .A2(new_n2948_), .ZN(new_n2951_));
  NOR2_X1    g02695(.A1(new_n2790_), .A2(new_n2951_), .ZN(new_n2952_));
  NOR2_X1    g02696(.A1(new_n2950_), .A2(new_n2952_), .ZN(new_n2953_));
  OAI21_X1   g02697(.A1(new_n2543_), .A2(new_n2794_), .B(new_n2660_), .ZN(new_n2954_));
  NAND3_X1   g02698(.A1(new_n2653_), .A2(new_n2654_), .A3(new_n2954_), .ZN(new_n2955_));
  OAI21_X1   g02699(.A1(\b[31] ), .A2(\b[33] ), .B(\b[32] ), .ZN(new_n2956_));
  NAND2_X1   g02700(.A1(new_n2955_), .A2(new_n2956_), .ZN(new_n2957_));
  INV_X1     g02701(.I(new_n2957_), .ZN(new_n2958_));
  XNOR2_X1   g02702(.A1(\b[33] ), .A2(\b[34] ), .ZN(new_n2959_));
  NOR2_X1    g02703(.A1(new_n2958_), .A2(new_n2959_), .ZN(new_n2960_));
  XNOR2_X1   g02704(.A1(\b[33] ), .A2(\b[34] ), .ZN(new_n2961_));
  AOI21_X1   g02705(.A1(new_n2958_), .A2(new_n2961_), .B(new_n2960_), .ZN(new_n2962_));
  INV_X1     g02706(.I(new_n2962_), .ZN(new_n2963_));
  INV_X1     g02707(.I(\b[34] ), .ZN(new_n2964_));
  OAI22_X1   g02708(.A1(new_n405_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n404_), .ZN(new_n2965_));
  NAND2_X1   g02709(.A1(new_n279_), .A2(\b[32] ), .ZN(new_n2966_));
  AOI21_X1   g02710(.A1(new_n2965_), .A2(new_n2966_), .B(new_n264_), .ZN(new_n2967_));
  NAND2_X1   g02711(.A1(new_n2963_), .A2(new_n2967_), .ZN(new_n2968_));
  XOR2_X1    g02712(.A1(new_n2968_), .A2(\a[2] ), .Z(new_n2969_));
  NAND2_X1   g02713(.A1(new_n2793_), .A2(new_n2802_), .ZN(new_n2970_));
  NAND2_X1   g02714(.A1(new_n2803_), .A2(new_n2665_), .ZN(new_n2971_));
  NAND3_X1   g02715(.A1(new_n2971_), .A2(new_n2560_), .A3(new_n2804_), .ZN(new_n2972_));
  NAND2_X1   g02716(.A1(new_n2972_), .A2(new_n2970_), .ZN(new_n2973_));
  XOR2_X1    g02717(.A1(new_n2973_), .A2(new_n2969_), .Z(new_n2974_));
  XOR2_X1    g02718(.A1(new_n2974_), .A2(new_n2953_), .Z(\f[34] ));
  XOR2_X1    g02719(.A1(new_n2953_), .A2(new_n2969_), .Z(new_n2976_));
  NAND2_X1   g02720(.A1(new_n2976_), .A2(new_n2969_), .ZN(new_n2977_));
  NAND3_X1   g02721(.A1(new_n2972_), .A2(new_n2970_), .A3(new_n2976_), .ZN(new_n2978_));
  NAND2_X1   g02722(.A1(new_n2978_), .A2(new_n2977_), .ZN(new_n2979_));
  NOR2_X1    g02723(.A1(new_n2937_), .A2(new_n2942_), .ZN(new_n2980_));
  INV_X1     g02724(.I(new_n2932_), .ZN(new_n2981_));
  AOI21_X1   g02725(.A1(new_n2814_), .A2(new_n2981_), .B(new_n2930_), .ZN(new_n2982_));
  OAI22_X1   g02726(.A1(new_n757_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n752_), .ZN(new_n2983_));
  NAND2_X1   g02727(.A1(new_n1182_), .A2(\b[21] ), .ZN(new_n2984_));
  AOI21_X1   g02728(.A1(new_n2983_), .A2(new_n2984_), .B(new_n760_), .ZN(new_n2985_));
  NAND2_X1   g02729(.A1(new_n1604_), .A2(new_n2985_), .ZN(new_n2986_));
  XOR2_X1    g02730(.A1(new_n2986_), .A2(\a[14] ), .Z(new_n2987_));
  INV_X1     g02731(.I(new_n2987_), .ZN(new_n2988_));
  OAI22_X1   g02732(.A1(new_n940_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n935_), .ZN(new_n2989_));
  NAND2_X1   g02733(.A1(new_n1458_), .A2(\b[18] ), .ZN(new_n2990_));
  AOI21_X1   g02734(.A1(new_n2989_), .A2(new_n2990_), .B(new_n943_), .ZN(new_n2991_));
  NAND2_X1   g02735(.A1(new_n1304_), .A2(new_n2991_), .ZN(new_n2992_));
  XOR2_X1    g02736(.A1(new_n2992_), .A2(\a[17] ), .Z(new_n2993_));
  INV_X1     g02737(.I(new_n2993_), .ZN(new_n2994_));
  NAND2_X1   g02738(.A1(new_n2905_), .A2(new_n2910_), .ZN(new_n2995_));
  OAI21_X1   g02739(.A1(new_n2920_), .A2(new_n2911_), .B(new_n2995_), .ZN(new_n2996_));
  NOR3_X1    g02740(.A1(new_n2884_), .A2(new_n2889_), .A3(new_n2895_), .ZN(new_n2997_));
  INV_X1     g02741(.I(new_n2997_), .ZN(new_n2998_));
  OAI22_X1   g02742(.A1(new_n2452_), .A2(new_n347_), .B1(new_n393_), .B2(new_n2447_), .ZN(new_n2999_));
  OAI21_X1   g02743(.A1(new_n290_), .A2(new_n2602_), .B(new_n2999_), .ZN(new_n3000_));
  AOI21_X1   g02744(.A1(new_n352_), .A2(new_n2454_), .B(new_n3000_), .ZN(new_n3001_));
  XOR2_X1    g02745(.A1(new_n3001_), .A2(new_n2442_), .Z(new_n3002_));
  OAI22_X1   g02746(.A1(new_n2084_), .A2(new_n495_), .B1(new_n450_), .B2(new_n2079_), .ZN(new_n3003_));
  NAND2_X1   g02747(.A1(new_n2864_), .A2(\b[6] ), .ZN(new_n3004_));
  AOI21_X1   g02748(.A1(new_n3003_), .A2(new_n3004_), .B(new_n2087_), .ZN(new_n3005_));
  NAND2_X1   g02749(.A1(new_n494_), .A2(new_n3005_), .ZN(new_n3006_));
  XOR2_X1    g02750(.A1(new_n3006_), .A2(\a[29] ), .Z(new_n3007_));
  INV_X1     g02751(.I(new_n2859_), .ZN(new_n3008_));
  OAI21_X1   g02752(.A1(new_n2831_), .A2(new_n2858_), .B(new_n3008_), .ZN(new_n3009_));
  NAND2_X1   g02753(.A1(new_n2851_), .A2(new_n2852_), .ZN(new_n3010_));
  NOR2_X1    g02754(.A1(new_n2849_), .A2(new_n278_), .ZN(new_n3011_));
  XNOR2_X1   g02755(.A1(\a[32] ), .A2(\a[34] ), .ZN(new_n3012_));
  NAND2_X1   g02756(.A1(new_n2676_), .A2(new_n3012_), .ZN(new_n3013_));
  XNOR2_X1   g02757(.A1(\a[32] ), .A2(\a[35] ), .ZN(new_n3014_));
  NAND2_X1   g02758(.A1(new_n3013_), .A2(new_n3014_), .ZN(new_n3015_));
  OAI22_X1   g02759(.A1(new_n2846_), .A2(new_n292_), .B1(new_n267_), .B2(new_n2841_), .ZN(new_n3016_));
  NOR4_X1    g02760(.A1(new_n3016_), .A2(new_n258_), .A3(new_n3011_), .A4(new_n3015_), .ZN(new_n3017_));
  XOR2_X1    g02761(.A1(new_n3017_), .A2(new_n2836_), .Z(new_n3018_));
  XOR2_X1    g02762(.A1(new_n3010_), .A2(new_n3018_), .Z(new_n3019_));
  XOR2_X1    g02763(.A1(new_n3009_), .A2(new_n3019_), .Z(new_n3020_));
  XNOR2_X1   g02764(.A1(new_n3020_), .A2(new_n3007_), .ZN(new_n3021_));
  XOR2_X1    g02765(.A1(new_n3021_), .A2(new_n3002_), .Z(new_n3022_));
  OAI21_X1   g02766(.A1(new_n2871_), .A2(new_n2862_), .B(new_n2872_), .ZN(new_n3023_));
  XNOR2_X1   g02767(.A1(new_n3022_), .A2(new_n3023_), .ZN(new_n3024_));
  OAI22_X1   g02768(.A1(new_n1760_), .A2(new_n659_), .B1(new_n617_), .B2(new_n1755_), .ZN(new_n3025_));
  NAND2_X1   g02769(.A1(new_n2470_), .A2(\b[9] ), .ZN(new_n3026_));
  AOI21_X1   g02770(.A1(new_n3025_), .A2(new_n3026_), .B(new_n1763_), .ZN(new_n3027_));
  NAND2_X1   g02771(.A1(new_n663_), .A2(new_n3027_), .ZN(new_n3028_));
  XOR2_X1    g02772(.A1(new_n3028_), .A2(\a[26] ), .Z(new_n3029_));
  XOR2_X1    g02773(.A1(new_n3024_), .A2(new_n3029_), .Z(new_n3030_));
  XOR2_X1    g02774(.A1(new_n2885_), .A2(new_n2886_), .Z(new_n3031_));
  NAND2_X1   g02775(.A1(new_n3031_), .A2(new_n2877_), .ZN(new_n3032_));
  XNOR2_X1   g02776(.A1(new_n3032_), .A2(new_n3030_), .ZN(new_n3033_));
  NAND2_X1   g02777(.A1(new_n2885_), .A2(new_n2886_), .ZN(new_n3034_));
  XNOR2_X1   g02778(.A1(new_n3033_), .A2(new_n3034_), .ZN(new_n3035_));
  OAI22_X1   g02779(.A1(new_n1444_), .A2(new_n848_), .B1(new_n795_), .B2(new_n1439_), .ZN(new_n3036_));
  NAND2_X1   g02780(.A1(new_n2098_), .A2(\b[12] ), .ZN(new_n3037_));
  AOI21_X1   g02781(.A1(new_n3036_), .A2(new_n3037_), .B(new_n1447_), .ZN(new_n3038_));
  NAND2_X1   g02782(.A1(new_n847_), .A2(new_n3038_), .ZN(new_n3039_));
  XOR2_X1    g02783(.A1(new_n3039_), .A2(\a[23] ), .Z(new_n3040_));
  XOR2_X1    g02784(.A1(new_n3035_), .A2(new_n3040_), .Z(new_n3041_));
  OAI22_X1   g02785(.A1(new_n1168_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n1163_), .ZN(new_n3042_));
  NAND2_X1   g02786(.A1(new_n1774_), .A2(\b[15] ), .ZN(new_n3043_));
  AOI21_X1   g02787(.A1(new_n3042_), .A2(new_n3043_), .B(new_n1171_), .ZN(new_n3044_));
  NAND2_X1   g02788(.A1(new_n1047_), .A2(new_n3044_), .ZN(new_n3045_));
  XOR2_X1    g02789(.A1(new_n3045_), .A2(\a[20] ), .Z(new_n3046_));
  XOR2_X1    g02790(.A1(new_n3041_), .A2(new_n3046_), .Z(new_n3047_));
  NOR2_X1    g02791(.A1(new_n3047_), .A2(new_n2998_), .ZN(new_n3048_));
  INV_X1     g02792(.I(new_n3046_), .ZN(new_n3049_));
  XOR2_X1    g02793(.A1(new_n3041_), .A2(new_n3049_), .Z(new_n3050_));
  NOR2_X1    g02794(.A1(new_n3050_), .A2(new_n2997_), .ZN(new_n3051_));
  NOR2_X1    g02795(.A1(new_n3048_), .A2(new_n3051_), .ZN(new_n3052_));
  INV_X1     g02796(.I(new_n3052_), .ZN(new_n3053_));
  NOR2_X1    g02797(.A1(new_n3053_), .A2(new_n2903_), .ZN(new_n3054_));
  NOR2_X1    g02798(.A1(new_n3052_), .A2(new_n2902_), .ZN(new_n3055_));
  NOR2_X1    g02799(.A1(new_n3054_), .A2(new_n3055_), .ZN(new_n3056_));
  INV_X1     g02800(.I(new_n3056_), .ZN(new_n3057_));
  XOR2_X1    g02801(.A1(new_n2996_), .A2(new_n3057_), .Z(new_n3058_));
  XOR2_X1    g02802(.A1(new_n3058_), .A2(new_n2994_), .Z(new_n3059_));
  XOR2_X1    g02803(.A1(new_n3059_), .A2(new_n2988_), .Z(new_n3060_));
  XOR2_X1    g02804(.A1(new_n2818_), .A2(new_n2911_), .Z(new_n3061_));
  OAI21_X1   g02805(.A1(new_n3061_), .A2(new_n2917_), .B(new_n2924_), .ZN(new_n3062_));
  INV_X1     g02806(.I(new_n3062_), .ZN(new_n3063_));
  AND2_X2    g02807(.A1(new_n3060_), .A2(new_n3063_), .Z(new_n3064_));
  NOR2_X1    g02808(.A1(new_n3060_), .A2(new_n3063_), .ZN(new_n3065_));
  NOR2_X1    g02809(.A1(new_n3064_), .A2(new_n3065_), .ZN(new_n3066_));
  OAI22_X1   g02810(.A1(new_n582_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n577_), .ZN(new_n3067_));
  NAND2_X1   g02811(.A1(new_n960_), .A2(\b[24] ), .ZN(new_n3068_));
  AOI21_X1   g02812(.A1(new_n3067_), .A2(new_n3068_), .B(new_n585_), .ZN(new_n3069_));
  NAND2_X1   g02813(.A1(new_n1926_), .A2(new_n3069_), .ZN(new_n3070_));
  XOR2_X1    g02814(.A1(new_n3070_), .A2(\a[11] ), .Z(new_n3071_));
  NOR2_X1    g02815(.A1(new_n3066_), .A2(new_n3071_), .ZN(new_n3072_));
  NAND2_X1   g02816(.A1(new_n3066_), .A2(new_n3071_), .ZN(new_n3073_));
  INV_X1     g02817(.I(new_n3073_), .ZN(new_n3074_));
  NOR2_X1    g02818(.A1(new_n3074_), .A2(new_n3072_), .ZN(new_n3075_));
  OAI22_X1   g02819(.A1(new_n437_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n431_), .ZN(new_n3076_));
  NAND2_X1   g02820(.A1(new_n775_), .A2(\b[27] ), .ZN(new_n3077_));
  AOI21_X1   g02821(.A1(new_n3076_), .A2(new_n3077_), .B(new_n440_), .ZN(new_n3078_));
  NAND2_X1   g02822(.A1(new_n2276_), .A2(new_n3078_), .ZN(new_n3079_));
  XOR2_X1    g02823(.A1(new_n3079_), .A2(\a[8] ), .Z(new_n3080_));
  INV_X1     g02824(.I(new_n3080_), .ZN(new_n3081_));
  XOR2_X1    g02825(.A1(new_n3075_), .A2(new_n3081_), .Z(new_n3082_));
  NOR2_X1    g02826(.A1(new_n3082_), .A2(new_n2982_), .ZN(new_n3083_));
  INV_X1     g02827(.I(new_n2982_), .ZN(new_n3084_));
  XOR2_X1    g02828(.A1(new_n3075_), .A2(new_n3080_), .Z(new_n3085_));
  NOR2_X1    g02829(.A1(new_n3085_), .A2(new_n3084_), .ZN(new_n3086_));
  NOR2_X1    g02830(.A1(new_n3083_), .A2(new_n3086_), .ZN(new_n3087_));
  XOR2_X1    g02831(.A1(new_n3087_), .A2(new_n2980_), .Z(new_n3088_));
  OAI22_X1   g02832(.A1(new_n364_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n320_), .ZN(new_n3089_));
  NAND2_X1   g02833(.A1(new_n594_), .A2(\b[30] ), .ZN(new_n3090_));
  AOI21_X1   g02834(.A1(new_n3089_), .A2(new_n3090_), .B(new_n312_), .ZN(new_n3091_));
  NAND2_X1   g02835(.A1(new_n2659_), .A2(new_n3091_), .ZN(new_n3092_));
  XOR2_X1    g02836(.A1(new_n3092_), .A2(new_n308_), .Z(new_n3093_));
  AOI21_X1   g02837(.A1(new_n2943_), .A2(new_n2948_), .B(new_n2790_), .ZN(new_n3094_));
  XOR2_X1    g02838(.A1(new_n3094_), .A2(new_n3093_), .Z(new_n3095_));
  XNOR2_X1   g02839(.A1(new_n3095_), .A2(new_n3088_), .ZN(new_n3096_));
  INV_X1     g02840(.I(\b[35] ), .ZN(new_n3097_));
  INV_X1     g02841(.I(new_n2959_), .ZN(new_n3098_));
  XOR2_X1    g02842(.A1(new_n2957_), .A2(\b[33] ), .Z(new_n3099_));
  NAND2_X1   g02843(.A1(new_n3099_), .A2(new_n3098_), .ZN(new_n3100_));
  XOR2_X1    g02844(.A1(new_n3100_), .A2(new_n3097_), .Z(new_n3101_));
  OAI22_X1   g02845(.A1(new_n405_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n404_), .ZN(new_n3102_));
  NAND2_X1   g02846(.A1(new_n279_), .A2(\b[33] ), .ZN(new_n3103_));
  AOI21_X1   g02847(.A1(new_n3102_), .A2(new_n3103_), .B(new_n264_), .ZN(new_n3104_));
  NAND2_X1   g02848(.A1(new_n3101_), .A2(new_n3104_), .ZN(new_n3105_));
  XOR2_X1    g02849(.A1(new_n3105_), .A2(\a[2] ), .Z(new_n3106_));
  XOR2_X1    g02850(.A1(new_n3096_), .A2(new_n3106_), .Z(new_n3107_));
  NOR2_X1    g02851(.A1(new_n3096_), .A2(new_n3106_), .ZN(new_n3108_));
  INV_X1     g02852(.I(new_n3108_), .ZN(new_n3109_));
  NAND2_X1   g02853(.A1(new_n3096_), .A2(new_n3106_), .ZN(new_n3110_));
  NAND2_X1   g02854(.A1(new_n3109_), .A2(new_n3110_), .ZN(new_n3111_));
  MUX2_X1    g02855(.I0(new_n3111_), .I1(new_n3107_), .S(new_n2979_), .Z(\f[35] ));
  XOR2_X1    g02856(.A1(new_n3075_), .A2(new_n2982_), .Z(new_n3113_));
  NOR2_X1    g02857(.A1(new_n3113_), .A2(new_n3081_), .ZN(new_n3114_));
  NOR4_X1    g02858(.A1(new_n3114_), .A2(new_n3083_), .A3(new_n3086_), .A4(new_n2980_), .ZN(new_n3115_));
  INV_X1     g02859(.I(new_n2447_), .ZN(new_n3116_));
  AOI22_X1   g02860(.A1(\b[6] ), .A2(new_n2451_), .B1(new_n3116_), .B2(\b[5] ), .ZN(new_n3117_));
  NOR2_X1    g02861(.A1(new_n2602_), .A2(new_n393_), .ZN(new_n3118_));
  OAI21_X1   g02862(.A1(new_n3117_), .A2(new_n3118_), .B(new_n2454_), .ZN(new_n3119_));
  NOR2_X1    g02863(.A1(new_n524_), .A2(new_n3119_), .ZN(new_n3120_));
  XOR2_X1    g02864(.A1(new_n3120_), .A2(\a[32] ), .Z(new_n3121_));
  XNOR2_X1   g02865(.A1(\a[35] ), .A2(\a[36] ), .ZN(new_n3122_));
  NOR2_X1    g02866(.A1(new_n3122_), .A2(new_n258_), .ZN(new_n3123_));
  INV_X1     g02867(.I(new_n3018_), .ZN(new_n3124_));
  NOR2_X1    g02868(.A1(new_n3124_), .A2(new_n3010_), .ZN(new_n3125_));
  NOR2_X1    g02869(.A1(new_n3015_), .A2(new_n267_), .ZN(new_n3126_));
  OAI22_X1   g02870(.A1(new_n2846_), .A2(new_n290_), .B1(new_n292_), .B2(new_n2841_), .ZN(new_n3127_));
  NOR4_X1    g02871(.A1(new_n3127_), .A2(new_n677_), .A3(new_n2849_), .A4(new_n3126_), .ZN(new_n3128_));
  XOR2_X1    g02872(.A1(new_n3128_), .A2(new_n2836_), .Z(new_n3129_));
  XOR2_X1    g02873(.A1(new_n3125_), .A2(new_n3129_), .Z(new_n3130_));
  XOR2_X1    g02874(.A1(new_n3130_), .A2(new_n3123_), .Z(new_n3131_));
  XOR2_X1    g02875(.A1(new_n3131_), .A2(new_n3121_), .Z(new_n3132_));
  INV_X1     g02876(.I(new_n3002_), .ZN(new_n3133_));
  XOR2_X1    g02877(.A1(new_n2831_), .A2(new_n2835_), .Z(new_n3134_));
  INV_X1     g02878(.I(new_n3010_), .ZN(new_n3135_));
  NOR2_X1    g02879(.A1(new_n3135_), .A2(new_n3018_), .ZN(new_n3136_));
  NOR2_X1    g02880(.A1(new_n3136_), .A2(new_n3125_), .ZN(new_n3137_));
  XOR2_X1    g02881(.A1(new_n3137_), .A2(\a[32] ), .Z(new_n3138_));
  OAI21_X1   g02882(.A1(new_n3138_), .A2(new_n3001_), .B(new_n2857_), .ZN(new_n3139_));
  AOI21_X1   g02883(.A1(new_n3001_), .A2(new_n3138_), .B(new_n3139_), .ZN(new_n3140_));
  NAND2_X1   g02884(.A1(new_n3140_), .A2(new_n2856_), .ZN(new_n3141_));
  NAND3_X1   g02885(.A1(new_n3141_), .A2(new_n2853_), .A3(new_n3134_), .ZN(new_n3142_));
  OAI21_X1   g02886(.A1(new_n3133_), .A2(new_n3019_), .B(new_n3142_), .ZN(new_n3143_));
  NAND2_X1   g02887(.A1(new_n3143_), .A2(new_n3132_), .ZN(new_n3144_));
  NOR2_X1    g02888(.A1(new_n3133_), .A2(new_n3019_), .ZN(new_n3145_));
  NOR2_X1    g02889(.A1(new_n3132_), .A2(new_n3145_), .ZN(new_n3146_));
  NAND2_X1   g02890(.A1(new_n3142_), .A2(new_n3146_), .ZN(new_n3147_));
  NAND2_X1   g02891(.A1(new_n3144_), .A2(new_n3147_), .ZN(new_n3148_));
  OAI22_X1   g02892(.A1(new_n2084_), .A2(new_n510_), .B1(new_n495_), .B2(new_n2079_), .ZN(new_n3149_));
  NAND2_X1   g02893(.A1(new_n2864_), .A2(\b[7] ), .ZN(new_n3150_));
  AOI21_X1   g02894(.A1(new_n3149_), .A2(new_n3150_), .B(new_n2087_), .ZN(new_n3151_));
  NAND2_X1   g02895(.A1(new_n518_), .A2(new_n3151_), .ZN(new_n3152_));
  XOR2_X1    g02896(.A1(new_n3152_), .A2(\a[29] ), .Z(new_n3153_));
  NOR2_X1    g02897(.A1(new_n2871_), .A2(new_n2875_), .ZN(new_n3154_));
  NOR3_X1    g02898(.A1(new_n3022_), .A2(new_n3154_), .A3(new_n2874_), .ZN(new_n3155_));
  XOR2_X1    g02899(.A1(new_n3019_), .A2(new_n3002_), .Z(new_n3156_));
  XOR2_X1    g02900(.A1(new_n3009_), .A2(new_n3156_), .Z(new_n3157_));
  NAND2_X1   g02901(.A1(new_n3157_), .A2(new_n3007_), .ZN(new_n3158_));
  NAND2_X1   g02902(.A1(new_n3155_), .A2(new_n3158_), .ZN(new_n3159_));
  XOR2_X1    g02903(.A1(new_n3159_), .A2(new_n3153_), .Z(new_n3160_));
  XOR2_X1    g02904(.A1(new_n3160_), .A2(new_n3148_), .Z(new_n3161_));
  OAI22_X1   g02905(.A1(new_n1760_), .A2(new_n717_), .B1(new_n659_), .B2(new_n1755_), .ZN(new_n3162_));
  NAND2_X1   g02906(.A1(new_n2470_), .A2(\b[10] ), .ZN(new_n3163_));
  AOI21_X1   g02907(.A1(new_n3162_), .A2(new_n3163_), .B(new_n1763_), .ZN(new_n3164_));
  NAND2_X1   g02908(.A1(new_n716_), .A2(new_n3164_), .ZN(new_n3165_));
  XOR2_X1    g02909(.A1(new_n3165_), .A2(\a[26] ), .Z(new_n3166_));
  NAND2_X1   g02910(.A1(new_n3024_), .A2(new_n3029_), .ZN(new_n3167_));
  OR2_X2     g02911(.A1(new_n2885_), .A2(new_n2888_), .Z(new_n3168_));
  NAND4_X1   g02912(.A1(new_n3168_), .A2(new_n3030_), .A3(new_n2888_), .A4(new_n3167_), .ZN(new_n3169_));
  XOR2_X1    g02913(.A1(new_n3169_), .A2(new_n3166_), .Z(new_n3170_));
  XNOR2_X1   g02914(.A1(new_n3170_), .A2(new_n3161_), .ZN(new_n3171_));
  OAI22_X1   g02915(.A1(new_n1444_), .A2(new_n904_), .B1(new_n848_), .B2(new_n1439_), .ZN(new_n3172_));
  NAND2_X1   g02916(.A1(new_n2098_), .A2(\b[13] ), .ZN(new_n3173_));
  AOI21_X1   g02917(.A1(new_n3172_), .A2(new_n3173_), .B(new_n1447_), .ZN(new_n3174_));
  NAND2_X1   g02918(.A1(new_n907_), .A2(new_n3174_), .ZN(new_n3175_));
  XOR2_X1    g02919(.A1(new_n3175_), .A2(new_n1434_), .Z(new_n3176_));
  AOI21_X1   g02920(.A1(new_n3035_), .A2(new_n3040_), .B(new_n2997_), .ZN(new_n3177_));
  XOR2_X1    g02921(.A1(new_n3177_), .A2(new_n3176_), .Z(new_n3178_));
  XNOR2_X1   g02922(.A1(new_n3178_), .A2(new_n3171_), .ZN(new_n3179_));
  OAI22_X1   g02923(.A1(new_n1168_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n1163_), .ZN(new_n3180_));
  NAND2_X1   g02924(.A1(new_n1774_), .A2(\b[16] ), .ZN(new_n3181_));
  AOI21_X1   g02925(.A1(new_n3180_), .A2(new_n3181_), .B(new_n1171_), .ZN(new_n3182_));
  NAND2_X1   g02926(.A1(new_n1123_), .A2(new_n3182_), .ZN(new_n3183_));
  XOR2_X1    g02927(.A1(new_n3183_), .A2(\a[20] ), .Z(new_n3184_));
  INV_X1     g02928(.I(new_n3184_), .ZN(new_n3185_));
  NOR2_X1    g02929(.A1(new_n3053_), .A2(new_n2902_), .ZN(new_n3186_));
  XOR2_X1    g02930(.A1(new_n3041_), .A2(new_n2997_), .Z(new_n3187_));
  OAI21_X1   g02931(.A1(new_n3049_), .A2(new_n3187_), .B(new_n3186_), .ZN(new_n3188_));
  XOR2_X1    g02932(.A1(new_n3188_), .A2(new_n3185_), .Z(new_n3189_));
  XOR2_X1    g02933(.A1(new_n3189_), .A2(new_n3179_), .Z(new_n3190_));
  OAI22_X1   g02934(.A1(new_n940_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n935_), .ZN(new_n3191_));
  NAND2_X1   g02935(.A1(new_n1458_), .A2(\b[19] ), .ZN(new_n3192_));
  AOI21_X1   g02936(.A1(new_n3191_), .A2(new_n3192_), .B(new_n943_), .ZN(new_n3193_));
  NAND2_X1   g02937(.A1(new_n1396_), .A2(new_n3193_), .ZN(new_n3194_));
  XOR2_X1    g02938(.A1(new_n3194_), .A2(\a[17] ), .Z(new_n3195_));
  XOR2_X1    g02939(.A1(new_n3056_), .A2(new_n2994_), .Z(new_n3196_));
  NAND2_X1   g02940(.A1(new_n3057_), .A2(new_n2993_), .ZN(new_n3197_));
  OAI21_X1   g02941(.A1(new_n2996_), .A2(new_n3196_), .B(new_n3197_), .ZN(new_n3198_));
  XOR2_X1    g02942(.A1(new_n3198_), .A2(new_n3195_), .Z(new_n3199_));
  XNOR2_X1   g02943(.A1(new_n3199_), .A2(new_n3190_), .ZN(new_n3200_));
  OAI22_X1   g02944(.A1(new_n757_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n752_), .ZN(new_n3201_));
  NAND2_X1   g02945(.A1(new_n1182_), .A2(\b[22] ), .ZN(new_n3202_));
  AOI21_X1   g02946(.A1(new_n3201_), .A2(new_n3202_), .B(new_n760_), .ZN(new_n3203_));
  NAND2_X1   g02947(.A1(new_n1708_), .A2(new_n3203_), .ZN(new_n3204_));
  XOR2_X1    g02948(.A1(new_n3204_), .A2(\a[14] ), .Z(new_n3205_));
  NAND2_X1   g02949(.A1(new_n3056_), .A2(new_n2994_), .ZN(new_n3206_));
  NAND2_X1   g02950(.A1(new_n3197_), .A2(new_n3206_), .ZN(new_n3207_));
  XNOR2_X1   g02951(.A1(new_n2996_), .A2(new_n3207_), .ZN(new_n3208_));
  AOI21_X1   g02952(.A1(new_n2987_), .A2(new_n3208_), .B(new_n3064_), .ZN(new_n3209_));
  XOR2_X1    g02953(.A1(new_n3209_), .A2(new_n3205_), .Z(new_n3210_));
  XOR2_X1    g02954(.A1(new_n3210_), .A2(new_n3200_), .Z(new_n3211_));
  OAI22_X1   g02955(.A1(new_n582_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n577_), .ZN(new_n3212_));
  NAND2_X1   g02956(.A1(new_n960_), .A2(\b[25] ), .ZN(new_n3213_));
  AOI21_X1   g02957(.A1(new_n3212_), .A2(new_n3213_), .B(new_n585_), .ZN(new_n3214_));
  NAND2_X1   g02958(.A1(new_n2042_), .A2(new_n3214_), .ZN(new_n3215_));
  XOR2_X1    g02959(.A1(new_n3215_), .A2(\a[11] ), .Z(new_n3216_));
  INV_X1     g02960(.I(new_n3071_), .ZN(new_n3217_));
  NOR4_X1    g02961(.A1(new_n2815_), .A2(new_n2929_), .A3(new_n3074_), .A4(new_n3072_), .ZN(new_n3218_));
  XOR2_X1    g02962(.A1(new_n2814_), .A2(new_n2931_), .Z(new_n3219_));
  NAND2_X1   g02963(.A1(new_n3219_), .A2(new_n2923_), .ZN(new_n3220_));
  OAI22_X1   g02964(.A1(new_n3220_), .A2(new_n3218_), .B1(new_n3066_), .B2(new_n3217_), .ZN(new_n3221_));
  XOR2_X1    g02965(.A1(new_n3221_), .A2(new_n3216_), .Z(new_n3222_));
  XNOR2_X1   g02966(.A1(new_n3222_), .A2(new_n3211_), .ZN(new_n3223_));
  OAI22_X1   g02967(.A1(new_n437_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n431_), .ZN(new_n3224_));
  NAND2_X1   g02968(.A1(new_n775_), .A2(\b[28] ), .ZN(new_n3225_));
  AOI21_X1   g02969(.A1(new_n3224_), .A2(new_n3225_), .B(new_n440_), .ZN(new_n3226_));
  NAND2_X1   g02970(.A1(new_n2404_), .A2(new_n3226_), .ZN(new_n3227_));
  XOR2_X1    g02971(.A1(new_n3227_), .A2(\a[8] ), .Z(new_n3228_));
  XOR2_X1    g02972(.A1(new_n3223_), .A2(new_n3228_), .Z(new_n3229_));
  OAI22_X1   g02973(.A1(new_n364_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n320_), .ZN(new_n3230_));
  NAND2_X1   g02974(.A1(new_n594_), .A2(\b[31] ), .ZN(new_n3231_));
  AOI21_X1   g02975(.A1(new_n3230_), .A2(new_n3231_), .B(new_n312_), .ZN(new_n3232_));
  NAND2_X1   g02976(.A1(new_n2797_), .A2(new_n3232_), .ZN(new_n3233_));
  XOR2_X1    g02977(.A1(new_n3233_), .A2(\a[5] ), .Z(new_n3234_));
  XOR2_X1    g02978(.A1(new_n3229_), .A2(new_n3234_), .Z(new_n3235_));
  NAND2_X1   g02979(.A1(new_n3235_), .A2(new_n3115_), .ZN(new_n3236_));
  XOR2_X1    g02980(.A1(new_n3229_), .A2(new_n3234_), .Z(new_n3237_));
  OAI21_X1   g02981(.A1(new_n3115_), .A2(new_n3237_), .B(new_n3236_), .ZN(new_n3238_));
  OAI21_X1   g02982(.A1(new_n2794_), .A2(new_n3097_), .B(new_n2964_), .ZN(new_n3239_));
  NAND2_X1   g02983(.A1(new_n2958_), .A2(new_n3239_), .ZN(new_n3240_));
  OAI21_X1   g02984(.A1(\b[33] ), .A2(\b[35] ), .B(\b[34] ), .ZN(new_n3241_));
  NAND2_X1   g02985(.A1(new_n3240_), .A2(new_n3241_), .ZN(new_n3242_));
  XOR2_X1    g02986(.A1(\b[35] ), .A2(\b[36] ), .Z(new_n3243_));
  NAND2_X1   g02987(.A1(new_n3242_), .A2(new_n3243_), .ZN(new_n3244_));
  XOR2_X1    g02988(.A1(\b[35] ), .A2(\b[36] ), .Z(new_n3245_));
  OAI21_X1   g02989(.A1(new_n3242_), .A2(new_n3245_), .B(new_n3244_), .ZN(new_n3246_));
  INV_X1     g02990(.I(\b[36] ), .ZN(new_n3247_));
  OAI22_X1   g02991(.A1(new_n405_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n404_), .ZN(new_n3248_));
  NAND2_X1   g02992(.A1(new_n279_), .A2(\b[34] ), .ZN(new_n3249_));
  AOI21_X1   g02993(.A1(new_n3248_), .A2(new_n3249_), .B(new_n264_), .ZN(new_n3250_));
  NAND2_X1   g02994(.A1(new_n3246_), .A2(new_n3250_), .ZN(new_n3251_));
  XOR2_X1    g02995(.A1(new_n3251_), .A2(\a[2] ), .Z(new_n3252_));
  INV_X1     g02996(.I(new_n3252_), .ZN(new_n3253_));
  XOR2_X1    g02997(.A1(new_n3238_), .A2(new_n3253_), .Z(new_n3254_));
  AOI21_X1   g02998(.A1(new_n2978_), .A2(new_n2977_), .B(new_n3096_), .ZN(new_n3255_));
  XNOR2_X1   g02999(.A1(new_n3255_), .A2(new_n3254_), .ZN(new_n3256_));
  XOR2_X1    g03000(.A1(new_n2979_), .A2(new_n3096_), .Z(new_n3257_));
  NOR2_X1    g03001(.A1(new_n3257_), .A2(new_n3106_), .ZN(new_n3258_));
  XOR2_X1    g03002(.A1(new_n3258_), .A2(new_n3256_), .Z(\f[36] ));
  NAND2_X1   g03003(.A1(new_n3229_), .A2(new_n3228_), .ZN(new_n3260_));
  NAND2_X1   g03004(.A1(new_n3229_), .A2(new_n3115_), .ZN(new_n3261_));
  NAND2_X1   g03005(.A1(new_n3261_), .A2(new_n3260_), .ZN(new_n3262_));
  XOR2_X1    g03006(.A1(new_n3200_), .A2(new_n3205_), .Z(new_n3263_));
  NAND2_X1   g03007(.A1(new_n3263_), .A2(new_n3205_), .ZN(new_n3264_));
  NAND2_X1   g03008(.A1(new_n3209_), .A2(new_n3263_), .ZN(new_n3265_));
  NAND2_X1   g03009(.A1(new_n3265_), .A2(new_n3264_), .ZN(new_n3266_));
  XOR2_X1    g03010(.A1(new_n3179_), .A2(new_n3185_), .Z(new_n3267_));
  AOI21_X1   g03011(.A1(new_n3188_), .A2(new_n3185_), .B(new_n3267_), .ZN(new_n3268_));
  NAND2_X1   g03012(.A1(new_n3148_), .A2(new_n3153_), .ZN(new_n3269_));
  XNOR2_X1   g03013(.A1(new_n3148_), .A2(new_n3153_), .ZN(new_n3270_));
  NAND3_X1   g03014(.A1(new_n3270_), .A2(new_n3155_), .A3(new_n3158_), .ZN(new_n3271_));
  NAND2_X1   g03015(.A1(new_n3271_), .A2(new_n3269_), .ZN(new_n3272_));
  INV_X1     g03016(.I(new_n3272_), .ZN(new_n3273_));
  XOR2_X1    g03017(.A1(new_n3129_), .A2(new_n3123_), .Z(new_n3274_));
  AND2_X2    g03018(.A1(new_n3274_), .A2(new_n3125_), .Z(new_n3275_));
  NOR2_X1    g03019(.A1(new_n3274_), .A2(new_n3125_), .ZN(new_n3276_));
  NOR3_X1    g03020(.A1(new_n3275_), .A2(new_n3276_), .A3(new_n3121_), .ZN(new_n3277_));
  NAND2_X1   g03021(.A1(new_n3144_), .A2(new_n3277_), .ZN(new_n3278_));
  AOI21_X1   g03022(.A1(new_n3274_), .A2(new_n3018_), .B(new_n3135_), .ZN(new_n3279_));
  NAND2_X1   g03023(.A1(new_n3129_), .A2(new_n3123_), .ZN(new_n3280_));
  XOR2_X1    g03024(.A1(new_n3279_), .A2(new_n3280_), .Z(new_n3281_));
  INV_X1     g03025(.I(new_n3281_), .ZN(new_n3282_));
  OAI22_X1   g03026(.A1(new_n2846_), .A2(new_n393_), .B1(new_n290_), .B2(new_n2841_), .ZN(new_n3283_));
  OAI21_X1   g03027(.A1(new_n292_), .A2(new_n3015_), .B(new_n3283_), .ZN(new_n3284_));
  NAND3_X1   g03028(.A1(new_n3284_), .A2(new_n334_), .A3(new_n2848_), .ZN(new_n3285_));
  XOR2_X1    g03029(.A1(new_n3285_), .A2(\a[35] ), .Z(new_n3286_));
  INV_X1     g03030(.I(new_n3286_), .ZN(new_n3287_));
  INV_X1     g03031(.I(\a[38] ), .ZN(new_n3288_));
  INV_X1     g03032(.I(\a[37] ), .ZN(new_n3289_));
  NOR3_X1    g03033(.A1(new_n3289_), .A2(\a[35] ), .A3(\a[36] ), .ZN(new_n3290_));
  NAND3_X1   g03034(.A1(new_n3289_), .A2(\a[35] ), .A3(\a[36] ), .ZN(new_n3291_));
  INV_X1     g03035(.I(new_n3291_), .ZN(new_n3292_));
  NOR2_X1    g03036(.A1(new_n3292_), .A2(new_n3290_), .ZN(new_n3293_));
  NOR2_X1    g03037(.A1(new_n3293_), .A2(new_n258_), .ZN(new_n3294_));
  INV_X1     g03038(.I(new_n3122_), .ZN(new_n3295_));
  XNOR2_X1   g03039(.A1(\a[37] ), .A2(\a[38] ), .ZN(new_n3296_));
  NOR2_X1    g03040(.A1(new_n3295_), .A2(new_n3296_), .ZN(new_n3297_));
  INV_X1     g03041(.I(new_n3297_), .ZN(new_n3298_));
  NOR2_X1    g03042(.A1(new_n3298_), .A2(new_n267_), .ZN(new_n3299_));
  NOR2_X1    g03043(.A1(new_n3122_), .A2(new_n3296_), .ZN(new_n3300_));
  INV_X1     g03044(.I(new_n3300_), .ZN(new_n3301_));
  NOR4_X1    g03045(.A1(new_n3299_), .A2(new_n261_), .A3(new_n3294_), .A4(new_n3301_), .ZN(new_n3302_));
  XOR2_X1    g03046(.A1(new_n3302_), .A2(new_n3288_), .Z(new_n3303_));
  NOR2_X1    g03047(.A1(new_n3123_), .A2(new_n3288_), .ZN(new_n3304_));
  XNOR2_X1   g03048(.A1(new_n3303_), .A2(new_n3304_), .ZN(new_n3305_));
  XOR2_X1    g03049(.A1(new_n3305_), .A2(new_n3287_), .Z(new_n3306_));
  OR2_X2     g03050(.A1(new_n3305_), .A2(new_n3287_), .Z(new_n3307_));
  NAND2_X1   g03051(.A1(new_n3305_), .A2(new_n3287_), .ZN(new_n3308_));
  AOI21_X1   g03052(.A1(new_n3307_), .A2(new_n3308_), .B(new_n3282_), .ZN(new_n3309_));
  AOI21_X1   g03053(.A1(new_n3282_), .A2(new_n3306_), .B(new_n3309_), .ZN(new_n3310_));
  OAI22_X1   g03054(.A1(new_n2452_), .A2(new_n450_), .B1(new_n403_), .B2(new_n2447_), .ZN(new_n3311_));
  INV_X1     g03055(.I(new_n2602_), .ZN(new_n3312_));
  NAND2_X1   g03056(.A1(new_n3312_), .A2(\b[5] ), .ZN(new_n3313_));
  AOI21_X1   g03057(.A1(new_n3311_), .A2(new_n3313_), .B(new_n2455_), .ZN(new_n3314_));
  NAND2_X1   g03058(.A1(new_n454_), .A2(new_n3314_), .ZN(new_n3315_));
  XOR2_X1    g03059(.A1(new_n3315_), .A2(\a[32] ), .Z(new_n3316_));
  XOR2_X1    g03060(.A1(new_n3310_), .A2(new_n3316_), .Z(new_n3317_));
  INV_X1     g03061(.I(new_n3317_), .ZN(new_n3318_));
  INV_X1     g03062(.I(new_n3316_), .ZN(new_n3319_));
  XOR2_X1    g03063(.A1(new_n3310_), .A2(new_n3319_), .Z(new_n3320_));
  NOR2_X1    g03064(.A1(new_n3278_), .A2(new_n3320_), .ZN(new_n3321_));
  AOI21_X1   g03065(.A1(new_n3278_), .A2(new_n3318_), .B(new_n3321_), .ZN(new_n3322_));
  OAI22_X1   g03066(.A1(new_n2084_), .A2(new_n617_), .B1(new_n510_), .B2(new_n2079_), .ZN(new_n3323_));
  NAND2_X1   g03067(.A1(new_n2864_), .A2(\b[8] ), .ZN(new_n3324_));
  AOI21_X1   g03068(.A1(new_n3323_), .A2(new_n3324_), .B(new_n2087_), .ZN(new_n3325_));
  NAND2_X1   g03069(.A1(new_n616_), .A2(new_n3325_), .ZN(new_n3326_));
  XOR2_X1    g03070(.A1(new_n3326_), .A2(\a[29] ), .Z(new_n3327_));
  XOR2_X1    g03071(.A1(new_n3322_), .A2(new_n3327_), .Z(new_n3328_));
  NOR2_X1    g03072(.A1(new_n3273_), .A2(new_n3328_), .ZN(new_n3329_));
  INV_X1     g03073(.I(new_n3327_), .ZN(new_n3330_));
  NAND2_X1   g03074(.A1(new_n3322_), .A2(new_n3330_), .ZN(new_n3331_));
  NOR2_X1    g03075(.A1(new_n3322_), .A2(new_n3330_), .ZN(new_n3332_));
  INV_X1     g03076(.I(new_n3332_), .ZN(new_n3333_));
  AOI21_X1   g03077(.A1(new_n3331_), .A2(new_n3333_), .B(new_n3272_), .ZN(new_n3334_));
  NOR2_X1    g03078(.A1(new_n3329_), .A2(new_n3334_), .ZN(new_n3335_));
  OAI22_X1   g03079(.A1(new_n1760_), .A2(new_n795_), .B1(new_n717_), .B2(new_n1755_), .ZN(new_n3336_));
  NAND2_X1   g03080(.A1(new_n2470_), .A2(\b[11] ), .ZN(new_n3337_));
  AOI21_X1   g03081(.A1(new_n3336_), .A2(new_n3337_), .B(new_n1763_), .ZN(new_n3338_));
  NAND2_X1   g03082(.A1(new_n799_), .A2(new_n3338_), .ZN(new_n3339_));
  XOR2_X1    g03083(.A1(new_n3339_), .A2(\a[26] ), .Z(new_n3340_));
  XOR2_X1    g03084(.A1(new_n3335_), .A2(new_n3340_), .Z(new_n3341_));
  OAI22_X1   g03085(.A1(new_n1444_), .A2(new_n992_), .B1(new_n904_), .B2(new_n1439_), .ZN(new_n3342_));
  NAND2_X1   g03086(.A1(new_n2098_), .A2(\b[14] ), .ZN(new_n3343_));
  AOI21_X1   g03087(.A1(new_n3342_), .A2(new_n3343_), .B(new_n1447_), .ZN(new_n3344_));
  NAND2_X1   g03088(.A1(new_n991_), .A2(new_n3344_), .ZN(new_n3345_));
  XOR2_X1    g03089(.A1(new_n3345_), .A2(\a[23] ), .Z(new_n3346_));
  XOR2_X1    g03090(.A1(new_n3341_), .A2(new_n3346_), .Z(new_n3347_));
  INV_X1     g03091(.I(new_n3347_), .ZN(new_n3348_));
  OAI22_X1   g03092(.A1(new_n1168_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n1163_), .ZN(new_n3349_));
  NAND2_X1   g03093(.A1(new_n1774_), .A2(\b[17] ), .ZN(new_n3350_));
  AOI21_X1   g03094(.A1(new_n3349_), .A2(new_n3350_), .B(new_n1171_), .ZN(new_n3351_));
  NAND2_X1   g03095(.A1(new_n1225_), .A2(new_n3351_), .ZN(new_n3352_));
  XOR2_X1    g03096(.A1(new_n3352_), .A2(\a[20] ), .Z(new_n3353_));
  NOR2_X1    g03097(.A1(new_n3348_), .A2(new_n3353_), .ZN(new_n3354_));
  NAND2_X1   g03098(.A1(new_n3348_), .A2(new_n3353_), .ZN(new_n3355_));
  INV_X1     g03099(.I(new_n3355_), .ZN(new_n3356_));
  NOR2_X1    g03100(.A1(new_n3356_), .A2(new_n3354_), .ZN(new_n3357_));
  OAI22_X1   g03101(.A1(new_n940_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n935_), .ZN(new_n3358_));
  NAND2_X1   g03102(.A1(new_n1458_), .A2(\b[20] ), .ZN(new_n3359_));
  AOI21_X1   g03103(.A1(new_n3358_), .A2(new_n3359_), .B(new_n943_), .ZN(new_n3360_));
  NAND2_X1   g03104(.A1(new_n1517_), .A2(new_n3360_), .ZN(new_n3361_));
  XOR2_X1    g03105(.A1(new_n3361_), .A2(\a[17] ), .Z(new_n3362_));
  INV_X1     g03106(.I(new_n3362_), .ZN(new_n3363_));
  XOR2_X1    g03107(.A1(new_n3357_), .A2(new_n3363_), .Z(new_n3364_));
  XOR2_X1    g03108(.A1(new_n3357_), .A2(new_n3363_), .Z(new_n3365_));
  NOR2_X1    g03109(.A1(new_n3268_), .A2(new_n3365_), .ZN(new_n3366_));
  AOI21_X1   g03110(.A1(new_n3268_), .A2(new_n3364_), .B(new_n3366_), .ZN(new_n3367_));
  OAI22_X1   g03111(.A1(new_n757_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n752_), .ZN(new_n3368_));
  NAND2_X1   g03112(.A1(new_n1182_), .A2(\b[23] ), .ZN(new_n3369_));
  AOI21_X1   g03113(.A1(new_n3368_), .A2(new_n3369_), .B(new_n760_), .ZN(new_n3370_));
  NAND2_X1   g03114(.A1(new_n1828_), .A2(new_n3370_), .ZN(new_n3371_));
  XOR2_X1    g03115(.A1(new_n3371_), .A2(\a[14] ), .Z(new_n3372_));
  INV_X1     g03116(.I(new_n3372_), .ZN(new_n3373_));
  XOR2_X1    g03117(.A1(new_n3367_), .A2(new_n3373_), .Z(new_n3374_));
  INV_X1     g03118(.I(new_n3374_), .ZN(new_n3375_));
  XOR2_X1    g03119(.A1(new_n3367_), .A2(new_n3372_), .Z(new_n3376_));
  NOR2_X1    g03120(.A1(new_n3266_), .A2(new_n3376_), .ZN(new_n3377_));
  AOI21_X1   g03121(.A1(new_n3266_), .A2(new_n3375_), .B(new_n3377_), .ZN(new_n3378_));
  OAI22_X1   g03122(.A1(new_n582_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n577_), .ZN(new_n3379_));
  NAND2_X1   g03123(.A1(new_n960_), .A2(\b[26] ), .ZN(new_n3380_));
  AOI21_X1   g03124(.A1(new_n3379_), .A2(new_n3380_), .B(new_n585_), .ZN(new_n3381_));
  NAND2_X1   g03125(.A1(new_n2174_), .A2(new_n3381_), .ZN(new_n3382_));
  XOR2_X1    g03126(.A1(new_n3382_), .A2(\a[11] ), .Z(new_n3383_));
  NOR2_X1    g03127(.A1(new_n3378_), .A2(new_n3383_), .ZN(new_n3384_));
  INV_X1     g03128(.I(new_n3384_), .ZN(new_n3385_));
  NAND2_X1   g03129(.A1(new_n3378_), .A2(new_n3383_), .ZN(new_n3386_));
  NAND2_X1   g03130(.A1(new_n3385_), .A2(new_n3386_), .ZN(new_n3387_));
  OAI22_X1   g03131(.A1(new_n437_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n431_), .ZN(new_n3388_));
  NAND2_X1   g03132(.A1(new_n775_), .A2(\b[29] ), .ZN(new_n3389_));
  AOI21_X1   g03133(.A1(new_n3388_), .A2(new_n3389_), .B(new_n440_), .ZN(new_n3390_));
  NAND2_X1   g03134(.A1(new_n2546_), .A2(new_n3390_), .ZN(new_n3391_));
  XOR2_X1    g03135(.A1(new_n3391_), .A2(\a[8] ), .Z(new_n3392_));
  INV_X1     g03136(.I(new_n3392_), .ZN(new_n3393_));
  XOR2_X1    g03137(.A1(new_n3387_), .A2(new_n3393_), .Z(new_n3394_));
  OAI22_X1   g03138(.A1(new_n364_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n320_), .ZN(new_n3395_));
  NAND2_X1   g03139(.A1(new_n594_), .A2(\b[32] ), .ZN(new_n3396_));
  AOI21_X1   g03140(.A1(new_n3395_), .A2(new_n3396_), .B(new_n312_), .ZN(new_n3397_));
  NAND2_X1   g03141(.A1(new_n2963_), .A2(new_n3397_), .ZN(new_n3398_));
  XOR2_X1    g03142(.A1(new_n3398_), .A2(\a[5] ), .Z(new_n3399_));
  XOR2_X1    g03143(.A1(new_n3394_), .A2(new_n3399_), .Z(new_n3400_));
  NAND2_X1   g03144(.A1(new_n3262_), .A2(new_n3400_), .ZN(new_n3401_));
  XOR2_X1    g03145(.A1(new_n3394_), .A2(new_n3399_), .Z(new_n3402_));
  OAI21_X1   g03146(.A1(new_n3262_), .A2(new_n3402_), .B(new_n3401_), .ZN(new_n3403_));
  XOR2_X1    g03147(.A1(new_n3229_), .A2(new_n3115_), .Z(new_n3404_));
  INV_X1     g03148(.I(new_n3404_), .ZN(new_n3405_));
  NOR2_X1    g03149(.A1(new_n3405_), .A2(new_n3234_), .ZN(new_n3406_));
  XNOR2_X1   g03150(.A1(new_n3403_), .A2(new_n3406_), .ZN(new_n3407_));
  INV_X1     g03151(.I(\b[37] ), .ZN(new_n3408_));
  XOR2_X1    g03152(.A1(new_n3242_), .A2(\b[35] ), .Z(new_n3409_));
  NAND2_X1   g03153(.A1(new_n3409_), .A2(new_n3243_), .ZN(new_n3410_));
  XOR2_X1    g03154(.A1(new_n3410_), .A2(new_n3408_), .Z(new_n3411_));
  OAI22_X1   g03155(.A1(new_n405_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n404_), .ZN(new_n3412_));
  NAND2_X1   g03156(.A1(new_n279_), .A2(\b[35] ), .ZN(new_n3413_));
  AOI21_X1   g03157(.A1(new_n3412_), .A2(new_n3413_), .B(new_n264_), .ZN(new_n3414_));
  NAND2_X1   g03158(.A1(new_n3411_), .A2(new_n3414_), .ZN(new_n3415_));
  XOR2_X1    g03159(.A1(new_n3415_), .A2(\a[2] ), .Z(new_n3416_));
  OR2_X2     g03160(.A1(new_n3238_), .A2(new_n3253_), .Z(new_n3417_));
  NAND2_X1   g03161(.A1(new_n2979_), .A2(new_n3110_), .ZN(new_n3418_));
  NAND4_X1   g03162(.A1(new_n3418_), .A2(new_n3109_), .A3(new_n3417_), .A4(new_n3254_), .ZN(new_n3419_));
  XOR2_X1    g03163(.A1(new_n3419_), .A2(new_n3416_), .Z(new_n3420_));
  XOR2_X1    g03164(.A1(new_n3420_), .A2(new_n3407_), .Z(\f[37] ));
  OAI22_X1   g03165(.A1(new_n757_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n752_), .ZN(new_n3422_));
  NAND2_X1   g03166(.A1(new_n1182_), .A2(\b[24] ), .ZN(new_n3423_));
  AOI21_X1   g03167(.A1(new_n3422_), .A2(new_n3423_), .B(new_n760_), .ZN(new_n3424_));
  NAND2_X1   g03168(.A1(new_n1926_), .A2(new_n3424_), .ZN(new_n3425_));
  XOR2_X1    g03169(.A1(new_n3425_), .A2(\a[14] ), .Z(new_n3426_));
  OAI22_X1   g03170(.A1(new_n940_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n935_), .ZN(new_n3427_));
  NAND2_X1   g03171(.A1(new_n1458_), .A2(\b[21] ), .ZN(new_n3428_));
  AOI21_X1   g03172(.A1(new_n3427_), .A2(new_n3428_), .B(new_n943_), .ZN(new_n3429_));
  NAND2_X1   g03173(.A1(new_n1604_), .A2(new_n3429_), .ZN(new_n3430_));
  XOR2_X1    g03174(.A1(new_n3430_), .A2(\a[17] ), .Z(new_n3431_));
  INV_X1     g03175(.I(new_n3431_), .ZN(new_n3432_));
  INV_X1     g03176(.I(new_n3357_), .ZN(new_n3433_));
  XOR2_X1    g03177(.A1(new_n3268_), .A2(new_n3433_), .Z(new_n3434_));
  AOI21_X1   g03178(.A1(new_n3362_), .A2(new_n3434_), .B(new_n3367_), .ZN(new_n3435_));
  NAND2_X1   g03179(.A1(new_n3282_), .A2(new_n3307_), .ZN(new_n3436_));
  NAND2_X1   g03180(.A1(new_n3436_), .A2(new_n3308_), .ZN(new_n3437_));
  OAI22_X1   g03181(.A1(new_n2846_), .A2(new_n347_), .B1(new_n393_), .B2(new_n2841_), .ZN(new_n3438_));
  OAI21_X1   g03182(.A1(new_n290_), .A2(new_n3015_), .B(new_n3438_), .ZN(new_n3439_));
  AOI21_X1   g03183(.A1(new_n352_), .A2(new_n2848_), .B(new_n3439_), .ZN(new_n3440_));
  NAND2_X1   g03184(.A1(new_n3303_), .A2(new_n3304_), .ZN(new_n3441_));
  INV_X1     g03185(.I(new_n3441_), .ZN(new_n3442_));
  NOR2_X1    g03186(.A1(new_n3301_), .A2(new_n278_), .ZN(new_n3443_));
  XNOR2_X1   g03187(.A1(\a[35] ), .A2(\a[37] ), .ZN(new_n3444_));
  NAND2_X1   g03188(.A1(new_n3122_), .A2(new_n3444_), .ZN(new_n3445_));
  XNOR2_X1   g03189(.A1(\a[35] ), .A2(\a[38] ), .ZN(new_n3446_));
  NAND2_X1   g03190(.A1(new_n3445_), .A2(new_n3446_), .ZN(new_n3447_));
  OAI22_X1   g03191(.A1(new_n3298_), .A2(new_n292_), .B1(new_n267_), .B2(new_n3293_), .ZN(new_n3448_));
  NOR4_X1    g03192(.A1(new_n3448_), .A2(new_n258_), .A3(new_n3443_), .A4(new_n3447_), .ZN(new_n3449_));
  XOR2_X1    g03193(.A1(new_n3449_), .A2(new_n3288_), .Z(new_n3450_));
  NOR2_X1    g03194(.A1(new_n3442_), .A2(new_n3450_), .ZN(new_n3451_));
  INV_X1     g03195(.I(new_n3450_), .ZN(new_n3452_));
  NOR2_X1    g03196(.A1(new_n3452_), .A2(new_n3441_), .ZN(new_n3453_));
  NOR2_X1    g03197(.A1(new_n3451_), .A2(new_n3453_), .ZN(new_n3454_));
  XOR2_X1    g03198(.A1(new_n3454_), .A2(\a[35] ), .Z(new_n3455_));
  NOR2_X1    g03199(.A1(new_n3455_), .A2(new_n3440_), .ZN(new_n3456_));
  NAND2_X1   g03200(.A1(new_n3455_), .A2(new_n3440_), .ZN(new_n3457_));
  INV_X1     g03201(.I(new_n3457_), .ZN(new_n3458_));
  NOR2_X1    g03202(.A1(new_n3458_), .A2(new_n3456_), .ZN(new_n3459_));
  OAI22_X1   g03203(.A1(new_n2452_), .A2(new_n495_), .B1(new_n450_), .B2(new_n2447_), .ZN(new_n3460_));
  NAND2_X1   g03204(.A1(new_n3312_), .A2(\b[6] ), .ZN(new_n3461_));
  AOI21_X1   g03205(.A1(new_n3460_), .A2(new_n3461_), .B(new_n2455_), .ZN(new_n3462_));
  NAND2_X1   g03206(.A1(new_n494_), .A2(new_n3462_), .ZN(new_n3463_));
  XOR2_X1    g03207(.A1(new_n3463_), .A2(\a[32] ), .Z(new_n3464_));
  XOR2_X1    g03208(.A1(new_n3459_), .A2(new_n3464_), .Z(new_n3465_));
  NAND2_X1   g03209(.A1(new_n3465_), .A2(new_n3437_), .ZN(new_n3466_));
  XOR2_X1    g03210(.A1(new_n3459_), .A2(new_n3464_), .Z(new_n3467_));
  OAI21_X1   g03211(.A1(new_n3437_), .A2(new_n3467_), .B(new_n3466_), .ZN(new_n3468_));
  XOR2_X1    g03212(.A1(new_n3278_), .A2(new_n3319_), .Z(new_n3469_));
  NAND2_X1   g03213(.A1(new_n3469_), .A2(new_n3310_), .ZN(new_n3470_));
  XOR2_X1    g03214(.A1(new_n3470_), .A2(new_n3468_), .Z(new_n3471_));
  NAND2_X1   g03215(.A1(new_n3278_), .A2(new_n3319_), .ZN(new_n3472_));
  XNOR2_X1   g03216(.A1(new_n3471_), .A2(new_n3472_), .ZN(new_n3473_));
  OAI22_X1   g03217(.A1(new_n2084_), .A2(new_n659_), .B1(new_n617_), .B2(new_n2079_), .ZN(new_n3474_));
  NAND2_X1   g03218(.A1(new_n2864_), .A2(\b[9] ), .ZN(new_n3475_));
  AOI21_X1   g03219(.A1(new_n3474_), .A2(new_n3475_), .B(new_n2087_), .ZN(new_n3476_));
  NAND2_X1   g03220(.A1(new_n663_), .A2(new_n3476_), .ZN(new_n3477_));
  XOR2_X1    g03221(.A1(new_n3477_), .A2(\a[29] ), .Z(new_n3478_));
  XNOR2_X1   g03222(.A1(new_n3473_), .A2(new_n3478_), .ZN(new_n3479_));
  XOR2_X1    g03223(.A1(new_n3272_), .A2(new_n3330_), .Z(new_n3480_));
  NAND2_X1   g03224(.A1(new_n3480_), .A2(new_n3322_), .ZN(new_n3481_));
  XNOR2_X1   g03225(.A1(new_n3479_), .A2(new_n3481_), .ZN(new_n3482_));
  NOR2_X1    g03226(.A1(new_n3273_), .A2(new_n3327_), .ZN(new_n3483_));
  XOR2_X1    g03227(.A1(new_n3482_), .A2(new_n3483_), .Z(new_n3484_));
  OAI22_X1   g03228(.A1(new_n1760_), .A2(new_n848_), .B1(new_n795_), .B2(new_n1755_), .ZN(new_n3485_));
  NAND2_X1   g03229(.A1(new_n2470_), .A2(\b[12] ), .ZN(new_n3486_));
  AOI21_X1   g03230(.A1(new_n3485_), .A2(new_n3486_), .B(new_n1763_), .ZN(new_n3487_));
  NAND2_X1   g03231(.A1(new_n847_), .A2(new_n3487_), .ZN(new_n3488_));
  XOR2_X1    g03232(.A1(new_n3488_), .A2(\a[26] ), .Z(new_n3489_));
  XNOR2_X1   g03233(.A1(new_n3484_), .A2(new_n3489_), .ZN(new_n3490_));
  NOR3_X1    g03234(.A1(new_n3329_), .A2(new_n3334_), .A3(new_n3340_), .ZN(new_n3491_));
  XOR2_X1    g03235(.A1(new_n3490_), .A2(new_n3491_), .Z(new_n3492_));
  INV_X1     g03236(.I(new_n3492_), .ZN(new_n3493_));
  OAI22_X1   g03237(.A1(new_n1444_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n1439_), .ZN(new_n3494_));
  NAND2_X1   g03238(.A1(new_n2098_), .A2(\b[15] ), .ZN(new_n3495_));
  AOI21_X1   g03239(.A1(new_n3494_), .A2(new_n3495_), .B(new_n1447_), .ZN(new_n3496_));
  NAND2_X1   g03240(.A1(new_n1047_), .A2(new_n3496_), .ZN(new_n3497_));
  XOR2_X1    g03241(.A1(new_n3497_), .A2(\a[23] ), .Z(new_n3498_));
  NOR2_X1    g03242(.A1(new_n3493_), .A2(new_n3498_), .ZN(new_n3499_));
  NAND2_X1   g03243(.A1(new_n3493_), .A2(new_n3498_), .ZN(new_n3500_));
  INV_X1     g03244(.I(new_n3500_), .ZN(new_n3501_));
  NOR2_X1    g03245(.A1(new_n3501_), .A2(new_n3499_), .ZN(new_n3502_));
  NOR2_X1    g03246(.A1(new_n3341_), .A2(new_n3346_), .ZN(new_n3503_));
  XOR2_X1    g03247(.A1(new_n3502_), .A2(new_n3503_), .Z(new_n3504_));
  OAI22_X1   g03248(.A1(new_n1168_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n1163_), .ZN(new_n3505_));
  NAND2_X1   g03249(.A1(new_n1774_), .A2(\b[18] ), .ZN(new_n3506_));
  AOI21_X1   g03250(.A1(new_n3505_), .A2(new_n3506_), .B(new_n1171_), .ZN(new_n3507_));
  NAND2_X1   g03251(.A1(new_n1304_), .A2(new_n3507_), .ZN(new_n3508_));
  XOR2_X1    g03252(.A1(new_n3508_), .A2(\a[20] ), .Z(new_n3509_));
  INV_X1     g03253(.I(new_n3509_), .ZN(new_n3510_));
  XOR2_X1    g03254(.A1(new_n3504_), .A2(new_n3510_), .Z(new_n3511_));
  INV_X1     g03255(.I(new_n3511_), .ZN(new_n3512_));
  OAI21_X1   g03256(.A1(new_n3268_), .A2(new_n3433_), .B(new_n3355_), .ZN(new_n3513_));
  NOR2_X1    g03257(.A1(new_n3512_), .A2(new_n3513_), .ZN(new_n3514_));
  NAND2_X1   g03258(.A1(new_n3512_), .A2(new_n3513_), .ZN(new_n3515_));
  INV_X1     g03259(.I(new_n3515_), .ZN(new_n3516_));
  NOR2_X1    g03260(.A1(new_n3516_), .A2(new_n3514_), .ZN(new_n3517_));
  XOR2_X1    g03261(.A1(new_n3517_), .A2(new_n3435_), .Z(new_n3518_));
  XOR2_X1    g03262(.A1(new_n3518_), .A2(new_n3432_), .Z(new_n3519_));
  XOR2_X1    g03263(.A1(new_n3519_), .A2(new_n3426_), .Z(new_n3520_));
  XOR2_X1    g03264(.A1(new_n3266_), .A2(new_n3373_), .Z(new_n3521_));
  NAND2_X1   g03265(.A1(new_n3521_), .A2(new_n3367_), .ZN(new_n3522_));
  XOR2_X1    g03266(.A1(new_n3522_), .A2(new_n3520_), .Z(new_n3523_));
  NAND2_X1   g03267(.A1(new_n3266_), .A2(new_n3373_), .ZN(new_n3524_));
  XNOR2_X1   g03268(.A1(new_n3523_), .A2(new_n3524_), .ZN(new_n3525_));
  OAI22_X1   g03269(.A1(new_n582_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n577_), .ZN(new_n3526_));
  NAND2_X1   g03270(.A1(new_n960_), .A2(\b[27] ), .ZN(new_n3527_));
  AOI21_X1   g03271(.A1(new_n3526_), .A2(new_n3527_), .B(new_n585_), .ZN(new_n3528_));
  NAND2_X1   g03272(.A1(new_n2276_), .A2(new_n3528_), .ZN(new_n3529_));
  XOR2_X1    g03273(.A1(new_n3529_), .A2(\a[11] ), .Z(new_n3530_));
  XOR2_X1    g03274(.A1(new_n3525_), .A2(new_n3530_), .Z(new_n3531_));
  XOR2_X1    g03275(.A1(new_n3531_), .A2(new_n3384_), .Z(new_n3532_));
  OAI22_X1   g03276(.A1(new_n437_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n431_), .ZN(new_n3533_));
  NAND2_X1   g03277(.A1(new_n775_), .A2(\b[30] ), .ZN(new_n3534_));
  AOI21_X1   g03278(.A1(new_n3533_), .A2(new_n3534_), .B(new_n440_), .ZN(new_n3535_));
  NAND2_X1   g03279(.A1(new_n2659_), .A2(new_n3535_), .ZN(new_n3536_));
  XOR2_X1    g03280(.A1(new_n3536_), .A2(\a[8] ), .Z(new_n3537_));
  XOR2_X1    g03281(.A1(new_n3532_), .A2(new_n3537_), .Z(new_n3538_));
  INV_X1     g03282(.I(new_n3538_), .ZN(new_n3539_));
  XOR2_X1    g03283(.A1(new_n3262_), .A2(new_n3393_), .Z(new_n3540_));
  NAND3_X1   g03284(.A1(new_n3540_), .A2(new_n3385_), .A3(new_n3386_), .ZN(new_n3541_));
  XOR2_X1    g03285(.A1(new_n3541_), .A2(new_n3539_), .Z(new_n3542_));
  NAND2_X1   g03286(.A1(new_n3262_), .A2(new_n3393_), .ZN(new_n3543_));
  XNOR2_X1   g03287(.A1(new_n3542_), .A2(new_n3543_), .ZN(new_n3544_));
  OAI22_X1   g03288(.A1(new_n364_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n320_), .ZN(new_n3545_));
  NAND2_X1   g03289(.A1(new_n594_), .A2(\b[33] ), .ZN(new_n3546_));
  AOI21_X1   g03290(.A1(new_n3545_), .A2(new_n3546_), .B(new_n312_), .ZN(new_n3547_));
  NAND2_X1   g03291(.A1(new_n3101_), .A2(new_n3547_), .ZN(new_n3548_));
  XOR2_X1    g03292(.A1(new_n3548_), .A2(\a[5] ), .Z(new_n3549_));
  XOR2_X1    g03293(.A1(new_n3262_), .A2(new_n3394_), .Z(new_n3550_));
  NAND2_X1   g03294(.A1(new_n3550_), .A2(new_n3399_), .ZN(new_n3551_));
  AOI21_X1   g03295(.A1(new_n3234_), .A2(new_n3405_), .B(new_n3403_), .ZN(new_n3552_));
  NAND2_X1   g03296(.A1(new_n3552_), .A2(new_n3551_), .ZN(new_n3553_));
  XOR2_X1    g03297(.A1(new_n3553_), .A2(new_n3549_), .Z(new_n3554_));
  XNOR2_X1   g03298(.A1(new_n3544_), .A2(new_n3554_), .ZN(new_n3555_));
  OAI21_X1   g03299(.A1(new_n3097_), .A2(new_n3408_), .B(new_n3247_), .ZN(new_n3556_));
  NAND3_X1   g03300(.A1(new_n3240_), .A2(new_n3241_), .A3(new_n3556_), .ZN(new_n3557_));
  OAI21_X1   g03301(.A1(\b[35] ), .A2(\b[37] ), .B(\b[36] ), .ZN(new_n3558_));
  NAND2_X1   g03302(.A1(new_n3557_), .A2(new_n3558_), .ZN(new_n3559_));
  INV_X1     g03303(.I(new_n3559_), .ZN(new_n3560_));
  XNOR2_X1   g03304(.A1(\b[37] ), .A2(\b[38] ), .ZN(new_n3561_));
  NOR2_X1    g03305(.A1(new_n3560_), .A2(new_n3561_), .ZN(new_n3562_));
  XNOR2_X1   g03306(.A1(\b[37] ), .A2(\b[38] ), .ZN(new_n3563_));
  AOI21_X1   g03307(.A1(new_n3560_), .A2(new_n3563_), .B(new_n3562_), .ZN(new_n3564_));
  INV_X1     g03308(.I(new_n3564_), .ZN(new_n3565_));
  INV_X1     g03309(.I(\b[38] ), .ZN(new_n3566_));
  OAI22_X1   g03310(.A1(new_n405_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n404_), .ZN(new_n3567_));
  NAND2_X1   g03311(.A1(new_n279_), .A2(\b[36] ), .ZN(new_n3568_));
  AOI21_X1   g03312(.A1(new_n3567_), .A2(new_n3568_), .B(new_n264_), .ZN(new_n3569_));
  NAND2_X1   g03313(.A1(new_n3565_), .A2(new_n3569_), .ZN(new_n3570_));
  XOR2_X1    g03314(.A1(new_n3570_), .A2(\a[2] ), .Z(new_n3571_));
  INV_X1     g03315(.I(new_n3571_), .ZN(new_n3572_));
  NAND2_X1   g03316(.A1(new_n3555_), .A2(new_n3572_), .ZN(new_n3573_));
  OR2_X2     g03317(.A1(new_n3555_), .A2(new_n3572_), .Z(new_n3574_));
  NAND2_X1   g03318(.A1(new_n3574_), .A2(new_n3573_), .ZN(\f[38] ));
  INV_X1     g03319(.I(new_n3530_), .ZN(new_n3576_));
  NOR2_X1    g03320(.A1(new_n3447_), .A2(new_n267_), .ZN(new_n3577_));
  OAI22_X1   g03321(.A1(new_n3298_), .A2(new_n290_), .B1(new_n292_), .B2(new_n3293_), .ZN(new_n3578_));
  NOR4_X1    g03322(.A1(new_n3578_), .A2(new_n677_), .A3(new_n3301_), .A4(new_n3577_), .ZN(new_n3579_));
  XOR2_X1    g03323(.A1(new_n3579_), .A2(new_n3288_), .Z(new_n3580_));
  XNOR2_X1   g03324(.A1(\a[38] ), .A2(\a[39] ), .ZN(new_n3581_));
  NOR2_X1    g03325(.A1(new_n3581_), .A2(new_n258_), .ZN(new_n3582_));
  XOR2_X1    g03326(.A1(new_n3580_), .A2(new_n3582_), .Z(new_n3583_));
  XOR2_X1    g03327(.A1(new_n3583_), .A2(new_n3453_), .Z(new_n3584_));
  INV_X1     g03328(.I(new_n2841_), .ZN(new_n3585_));
  AOI22_X1   g03329(.A1(\b[6] ), .A2(new_n2845_), .B1(new_n3585_), .B2(\b[5] ), .ZN(new_n3586_));
  NOR2_X1    g03330(.A1(new_n3015_), .A2(new_n393_), .ZN(new_n3587_));
  OAI21_X1   g03331(.A1(new_n3586_), .A2(new_n3587_), .B(new_n2848_), .ZN(new_n3588_));
  NOR2_X1    g03332(.A1(new_n524_), .A2(new_n3588_), .ZN(new_n3589_));
  XOR2_X1    g03333(.A1(new_n3589_), .A2(\a[35] ), .Z(new_n3590_));
  NOR2_X1    g03334(.A1(new_n3282_), .A2(new_n3307_), .ZN(new_n3591_));
  NAND2_X1   g03335(.A1(new_n3440_), .A2(new_n2836_), .ZN(new_n3592_));
  OR2_X2     g03336(.A1(new_n3440_), .A2(new_n2836_), .Z(new_n3593_));
  NAND4_X1   g03337(.A1(new_n3307_), .A2(new_n3454_), .A3(new_n3592_), .A4(new_n3593_), .ZN(new_n3594_));
  NOR4_X1    g03338(.A1(new_n3591_), .A2(new_n3456_), .A3(new_n3458_), .A4(new_n3594_), .ZN(new_n3595_));
  XOR2_X1    g03339(.A1(new_n3595_), .A2(new_n3590_), .Z(new_n3596_));
  XNOR2_X1   g03340(.A1(new_n3596_), .A2(new_n3584_), .ZN(new_n3597_));
  OAI22_X1   g03341(.A1(new_n2452_), .A2(new_n510_), .B1(new_n495_), .B2(new_n2447_), .ZN(new_n3598_));
  NAND2_X1   g03342(.A1(new_n3312_), .A2(\b[7] ), .ZN(new_n3599_));
  AOI21_X1   g03343(.A1(new_n3598_), .A2(new_n3599_), .B(new_n2455_), .ZN(new_n3600_));
  NAND2_X1   g03344(.A1(new_n518_), .A2(new_n3600_), .ZN(new_n3601_));
  XOR2_X1    g03345(.A1(new_n3601_), .A2(\a[32] ), .Z(new_n3602_));
  NOR2_X1    g03346(.A1(new_n3472_), .A2(new_n3468_), .ZN(new_n3603_));
  XNOR2_X1   g03347(.A1(new_n3437_), .A2(new_n3459_), .ZN(new_n3604_));
  NAND2_X1   g03348(.A1(new_n3604_), .A2(new_n3464_), .ZN(new_n3605_));
  OAI21_X1   g03349(.A1(new_n3470_), .A2(new_n3603_), .B(new_n3605_), .ZN(new_n3606_));
  XOR2_X1    g03350(.A1(new_n3606_), .A2(new_n3602_), .Z(new_n3607_));
  XNOR2_X1   g03351(.A1(new_n3607_), .A2(new_n3597_), .ZN(new_n3608_));
  OAI22_X1   g03352(.A1(new_n2084_), .A2(new_n717_), .B1(new_n659_), .B2(new_n2079_), .ZN(new_n3609_));
  NAND2_X1   g03353(.A1(new_n2864_), .A2(\b[10] ), .ZN(new_n3610_));
  AOI21_X1   g03354(.A1(new_n3609_), .A2(new_n3610_), .B(new_n2087_), .ZN(new_n3611_));
  NAND2_X1   g03355(.A1(new_n716_), .A2(new_n3611_), .ZN(new_n3612_));
  XOR2_X1    g03356(.A1(new_n3612_), .A2(\a[29] ), .Z(new_n3613_));
  INV_X1     g03357(.I(new_n3473_), .ZN(new_n3614_));
  NAND2_X1   g03358(.A1(new_n3614_), .A2(new_n3478_), .ZN(new_n3615_));
  NAND2_X1   g03359(.A1(new_n3273_), .A2(new_n3332_), .ZN(new_n3616_));
  NAND4_X1   g03360(.A1(new_n3479_), .A2(new_n3333_), .A3(new_n3615_), .A4(new_n3616_), .ZN(new_n3617_));
  XOR2_X1    g03361(.A1(new_n3617_), .A2(new_n3613_), .Z(new_n3618_));
  XNOR2_X1   g03362(.A1(new_n3618_), .A2(new_n3608_), .ZN(new_n3619_));
  OAI22_X1   g03363(.A1(new_n1760_), .A2(new_n904_), .B1(new_n848_), .B2(new_n1755_), .ZN(new_n3620_));
  NAND2_X1   g03364(.A1(new_n2470_), .A2(\b[13] ), .ZN(new_n3621_));
  AOI21_X1   g03365(.A1(new_n3620_), .A2(new_n3621_), .B(new_n1763_), .ZN(new_n3622_));
  NAND2_X1   g03366(.A1(new_n907_), .A2(new_n3622_), .ZN(new_n3623_));
  XOR2_X1    g03367(.A1(new_n3623_), .A2(new_n1750_), .Z(new_n3624_));
  AOI21_X1   g03368(.A1(new_n3484_), .A2(new_n3489_), .B(new_n3491_), .ZN(new_n3625_));
  XOR2_X1    g03369(.A1(new_n3625_), .A2(new_n3624_), .Z(new_n3626_));
  XNOR2_X1   g03370(.A1(new_n3626_), .A2(new_n3619_), .ZN(new_n3627_));
  OAI22_X1   g03371(.A1(new_n1444_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n1439_), .ZN(new_n3628_));
  NAND2_X1   g03372(.A1(new_n2098_), .A2(\b[16] ), .ZN(new_n3629_));
  AOI21_X1   g03373(.A1(new_n3628_), .A2(new_n3629_), .B(new_n1447_), .ZN(new_n3630_));
  NAND2_X1   g03374(.A1(new_n1123_), .A2(new_n3630_), .ZN(new_n3631_));
  XOR2_X1    g03375(.A1(new_n3631_), .A2(\a[23] ), .Z(new_n3632_));
  NOR3_X1    g03376(.A1(new_n3501_), .A2(new_n3499_), .A3(new_n3503_), .ZN(new_n3633_));
  XOR2_X1    g03377(.A1(new_n3633_), .A2(new_n3632_), .Z(new_n3634_));
  XOR2_X1    g03378(.A1(new_n3634_), .A2(new_n3627_), .Z(new_n3635_));
  OAI22_X1   g03379(.A1(new_n1168_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n1163_), .ZN(new_n3636_));
  NAND2_X1   g03380(.A1(new_n1774_), .A2(\b[19] ), .ZN(new_n3637_));
  AOI21_X1   g03381(.A1(new_n3636_), .A2(new_n3637_), .B(new_n1171_), .ZN(new_n3638_));
  NAND2_X1   g03382(.A1(new_n1396_), .A2(new_n3638_), .ZN(new_n3639_));
  XOR2_X1    g03383(.A1(new_n3639_), .A2(\a[20] ), .Z(new_n3640_));
  NOR2_X1    g03384(.A1(new_n3504_), .A2(new_n3510_), .ZN(new_n3641_));
  NOR2_X1    g03385(.A1(new_n3512_), .A2(new_n3641_), .ZN(new_n3642_));
  NAND2_X1   g03386(.A1(new_n3642_), .A2(new_n3513_), .ZN(new_n3643_));
  XOR2_X1    g03387(.A1(new_n3643_), .A2(new_n3640_), .Z(new_n3644_));
  XNOR2_X1   g03388(.A1(new_n3644_), .A2(new_n3635_), .ZN(new_n3645_));
  OAI22_X1   g03389(.A1(new_n940_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n935_), .ZN(new_n3646_));
  NAND2_X1   g03390(.A1(new_n1458_), .A2(\b[22] ), .ZN(new_n3647_));
  AOI21_X1   g03391(.A1(new_n3646_), .A2(new_n3647_), .B(new_n943_), .ZN(new_n3648_));
  NAND2_X1   g03392(.A1(new_n1708_), .A2(new_n3648_), .ZN(new_n3649_));
  XOR2_X1    g03393(.A1(new_n3649_), .A2(\a[17] ), .Z(new_n3650_));
  NAND2_X1   g03394(.A1(new_n3517_), .A2(new_n3431_), .ZN(new_n3651_));
  OAI21_X1   g03395(.A1(new_n3516_), .A2(new_n3514_), .B(new_n3432_), .ZN(new_n3652_));
  NAND3_X1   g03396(.A1(new_n3651_), .A2(new_n3435_), .A3(new_n3652_), .ZN(new_n3653_));
  OAI21_X1   g03397(.A1(new_n3432_), .A2(new_n3517_), .B(new_n3653_), .ZN(new_n3654_));
  XOR2_X1    g03398(.A1(new_n3654_), .A2(new_n3650_), .Z(new_n3655_));
  XNOR2_X1   g03399(.A1(new_n3655_), .A2(new_n3645_), .ZN(new_n3656_));
  OAI22_X1   g03400(.A1(new_n757_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n752_), .ZN(new_n3657_));
  NAND2_X1   g03401(.A1(new_n1182_), .A2(\b[25] ), .ZN(new_n3658_));
  AOI21_X1   g03402(.A1(new_n3657_), .A2(new_n3658_), .B(new_n760_), .ZN(new_n3659_));
  NAND2_X1   g03403(.A1(new_n2042_), .A2(new_n3659_), .ZN(new_n3660_));
  XOR2_X1    g03404(.A1(new_n3660_), .A2(\a[14] ), .Z(new_n3661_));
  NOR2_X1    g03405(.A1(new_n3520_), .A2(new_n3524_), .ZN(new_n3662_));
  XOR2_X1    g03406(.A1(new_n3517_), .A2(new_n3431_), .Z(new_n3663_));
  XOR2_X1    g03407(.A1(new_n3663_), .A2(new_n3435_), .Z(new_n3664_));
  NAND2_X1   g03408(.A1(new_n3664_), .A2(new_n3426_), .ZN(new_n3665_));
  OAI21_X1   g03409(.A1(new_n3522_), .A2(new_n3662_), .B(new_n3665_), .ZN(new_n3666_));
  XOR2_X1    g03410(.A1(new_n3666_), .A2(new_n3661_), .Z(new_n3667_));
  XNOR2_X1   g03411(.A1(new_n3667_), .A2(new_n3656_), .ZN(new_n3668_));
  OAI22_X1   g03412(.A1(new_n582_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n577_), .ZN(new_n3669_));
  NAND2_X1   g03413(.A1(new_n960_), .A2(\b[28] ), .ZN(new_n3670_));
  AOI21_X1   g03414(.A1(new_n3669_), .A2(new_n3670_), .B(new_n585_), .ZN(new_n3671_));
  NAND2_X1   g03415(.A1(new_n2404_), .A2(new_n3671_), .ZN(new_n3672_));
  XOR2_X1    g03416(.A1(new_n3672_), .A2(\a[11] ), .Z(new_n3673_));
  XNOR2_X1   g03417(.A1(new_n3668_), .A2(new_n3673_), .ZN(new_n3674_));
  INV_X1     g03418(.I(new_n3674_), .ZN(new_n3675_));
  OR3_X2     g03419(.A1(new_n3675_), .A2(new_n3525_), .A3(new_n3576_), .Z(new_n3676_));
  OAI21_X1   g03420(.A1(new_n3525_), .A2(new_n3576_), .B(new_n3675_), .ZN(new_n3677_));
  NAND2_X1   g03421(.A1(new_n3676_), .A2(new_n3677_), .ZN(new_n3678_));
  OAI22_X1   g03422(.A1(new_n437_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n431_), .ZN(new_n3679_));
  NAND2_X1   g03423(.A1(new_n775_), .A2(\b[31] ), .ZN(new_n3680_));
  AOI21_X1   g03424(.A1(new_n3679_), .A2(new_n3680_), .B(new_n440_), .ZN(new_n3681_));
  NAND2_X1   g03425(.A1(new_n2797_), .A2(new_n3681_), .ZN(new_n3682_));
  XOR2_X1    g03426(.A1(new_n3682_), .A2(new_n429_), .Z(new_n3683_));
  NOR2_X1    g03427(.A1(new_n3539_), .A2(new_n3543_), .ZN(new_n3684_));
  INV_X1     g03428(.I(new_n3532_), .ZN(new_n3685_));
  NAND2_X1   g03429(.A1(new_n3685_), .A2(new_n3537_), .ZN(new_n3686_));
  OAI21_X1   g03430(.A1(new_n3684_), .A2(new_n3541_), .B(new_n3686_), .ZN(new_n3687_));
  XOR2_X1    g03431(.A1(new_n3687_), .A2(new_n3683_), .Z(new_n3688_));
  XOR2_X1    g03432(.A1(new_n3688_), .A2(new_n3678_), .Z(new_n3689_));
  OAI22_X1   g03433(.A1(new_n364_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n320_), .ZN(new_n3690_));
  NAND2_X1   g03434(.A1(new_n594_), .A2(\b[34] ), .ZN(new_n3691_));
  AOI21_X1   g03435(.A1(new_n3690_), .A2(new_n3691_), .B(new_n312_), .ZN(new_n3692_));
  NAND2_X1   g03436(.A1(new_n3246_), .A2(new_n3692_), .ZN(new_n3693_));
  XOR2_X1    g03437(.A1(new_n3693_), .A2(new_n308_), .Z(new_n3694_));
  XNOR2_X1   g03438(.A1(new_n3689_), .A2(new_n3694_), .ZN(new_n3695_));
  INV_X1     g03439(.I(\b[39] ), .ZN(new_n3696_));
  INV_X1     g03440(.I(new_n3561_), .ZN(new_n3697_));
  XOR2_X1    g03441(.A1(new_n3559_), .A2(\b[37] ), .Z(new_n3698_));
  NAND2_X1   g03442(.A1(new_n3698_), .A2(new_n3697_), .ZN(new_n3699_));
  XOR2_X1    g03443(.A1(new_n3699_), .A2(new_n3696_), .Z(new_n3700_));
  NAND2_X1   g03444(.A1(new_n283_), .A2(\b[39] ), .ZN(new_n3701_));
  NAND2_X1   g03445(.A1(new_n279_), .A2(\b[37] ), .ZN(new_n3702_));
  AOI21_X1   g03446(.A1(\b[38] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n3703_));
  NAND4_X1   g03447(.A1(new_n3700_), .A2(new_n3701_), .A3(new_n3702_), .A4(new_n3703_), .ZN(new_n3704_));
  XOR2_X1    g03448(.A1(new_n3704_), .A2(\a[2] ), .Z(new_n3705_));
  NOR2_X1    g03449(.A1(new_n3695_), .A2(new_n3705_), .ZN(new_n3706_));
  INV_X1     g03450(.I(new_n3695_), .ZN(new_n3707_));
  INV_X1     g03451(.I(new_n3705_), .ZN(new_n3708_));
  NOR2_X1    g03452(.A1(new_n3707_), .A2(new_n3708_), .ZN(new_n3709_));
  NOR2_X1    g03453(.A1(new_n3709_), .A2(new_n3706_), .ZN(new_n3710_));
  NAND2_X1   g03454(.A1(new_n3555_), .A2(new_n3572_), .ZN(new_n3711_));
  XOR2_X1    g03455(.A1(new_n3710_), .A2(new_n3711_), .Z(\f[39] ));
  NAND2_X1   g03456(.A1(new_n3689_), .A2(new_n3694_), .ZN(new_n3713_));
  NAND2_X1   g03457(.A1(new_n3675_), .A2(new_n3673_), .ZN(new_n3714_));
  NAND2_X1   g03458(.A1(new_n3677_), .A2(new_n3714_), .ZN(new_n3715_));
  XNOR2_X1   g03459(.A1(new_n3627_), .A2(new_n3632_), .ZN(new_n3716_));
  INV_X1     g03460(.I(new_n3716_), .ZN(new_n3717_));
  OAI21_X1   g03461(.A1(new_n3632_), .A2(new_n3633_), .B(new_n3717_), .ZN(new_n3718_));
  AOI21_X1   g03462(.A1(new_n3583_), .A2(new_n3450_), .B(new_n3442_), .ZN(new_n3719_));
  NAND2_X1   g03463(.A1(new_n3580_), .A2(new_n3582_), .ZN(new_n3720_));
  XOR2_X1    g03464(.A1(new_n3719_), .A2(new_n3720_), .Z(new_n3721_));
  OAI22_X1   g03465(.A1(new_n3298_), .A2(new_n393_), .B1(new_n290_), .B2(new_n3293_), .ZN(new_n3722_));
  OAI21_X1   g03466(.A1(new_n292_), .A2(new_n3447_), .B(new_n3722_), .ZN(new_n3723_));
  NAND3_X1   g03467(.A1(new_n3723_), .A2(new_n334_), .A3(new_n3300_), .ZN(new_n3724_));
  XOR2_X1    g03468(.A1(new_n3724_), .A2(\a[38] ), .Z(new_n3725_));
  INV_X1     g03469(.I(\a[41] ), .ZN(new_n3726_));
  INV_X1     g03470(.I(\a[40] ), .ZN(new_n3727_));
  NOR3_X1    g03471(.A1(new_n3727_), .A2(\a[38] ), .A3(\a[39] ), .ZN(new_n3728_));
  NAND3_X1   g03472(.A1(new_n3727_), .A2(\a[38] ), .A3(\a[39] ), .ZN(new_n3729_));
  INV_X1     g03473(.I(new_n3729_), .ZN(new_n3730_));
  NOR2_X1    g03474(.A1(new_n3730_), .A2(new_n3728_), .ZN(new_n3731_));
  NOR2_X1    g03475(.A1(new_n3731_), .A2(new_n258_), .ZN(new_n3732_));
  INV_X1     g03476(.I(new_n3581_), .ZN(new_n3733_));
  XNOR2_X1   g03477(.A1(\a[40] ), .A2(\a[41] ), .ZN(new_n3734_));
  NOR2_X1    g03478(.A1(new_n3733_), .A2(new_n3734_), .ZN(new_n3735_));
  INV_X1     g03479(.I(new_n3735_), .ZN(new_n3736_));
  NOR2_X1    g03480(.A1(new_n3736_), .A2(new_n267_), .ZN(new_n3737_));
  NOR2_X1    g03481(.A1(new_n3581_), .A2(new_n3734_), .ZN(new_n3738_));
  INV_X1     g03482(.I(new_n3738_), .ZN(new_n3739_));
  NOR4_X1    g03483(.A1(new_n3737_), .A2(new_n261_), .A3(new_n3732_), .A4(new_n3739_), .ZN(new_n3740_));
  XOR2_X1    g03484(.A1(new_n3740_), .A2(new_n3726_), .Z(new_n3741_));
  NOR2_X1    g03485(.A1(new_n3582_), .A2(new_n3726_), .ZN(new_n3742_));
  XNOR2_X1   g03486(.A1(new_n3741_), .A2(new_n3742_), .ZN(new_n3743_));
  XOR2_X1    g03487(.A1(new_n3743_), .A2(new_n3725_), .Z(new_n3744_));
  NOR2_X1    g03488(.A1(new_n3721_), .A2(new_n3744_), .ZN(new_n3745_));
  INV_X1     g03489(.I(new_n3721_), .ZN(new_n3746_));
  INV_X1     g03490(.I(new_n3725_), .ZN(new_n3747_));
  NOR2_X1    g03491(.A1(new_n3743_), .A2(new_n3747_), .ZN(new_n3748_));
  INV_X1     g03492(.I(new_n3748_), .ZN(new_n3749_));
  NAND2_X1   g03493(.A1(new_n3743_), .A2(new_n3747_), .ZN(new_n3750_));
  AOI21_X1   g03494(.A1(new_n3749_), .A2(new_n3750_), .B(new_n3746_), .ZN(new_n3751_));
  NOR2_X1    g03495(.A1(new_n3751_), .A2(new_n3745_), .ZN(new_n3752_));
  INV_X1     g03496(.I(new_n3752_), .ZN(new_n3753_));
  OAI22_X1   g03497(.A1(new_n2846_), .A2(new_n450_), .B1(new_n403_), .B2(new_n2841_), .ZN(new_n3754_));
  INV_X1     g03498(.I(new_n3015_), .ZN(new_n3755_));
  NAND2_X1   g03499(.A1(new_n3755_), .A2(\b[5] ), .ZN(new_n3756_));
  AOI21_X1   g03500(.A1(new_n3754_), .A2(new_n3756_), .B(new_n2849_), .ZN(new_n3757_));
  NAND2_X1   g03501(.A1(new_n454_), .A2(new_n3757_), .ZN(new_n3758_));
  XOR2_X1    g03502(.A1(new_n3758_), .A2(\a[35] ), .Z(new_n3759_));
  NOR2_X1    g03503(.A1(new_n3753_), .A2(new_n3759_), .ZN(new_n3760_));
  INV_X1     g03504(.I(new_n3760_), .ZN(new_n3761_));
  NAND2_X1   g03505(.A1(new_n3753_), .A2(new_n3759_), .ZN(new_n3762_));
  NAND2_X1   g03506(.A1(new_n3761_), .A2(new_n3762_), .ZN(new_n3763_));
  OAI22_X1   g03507(.A1(new_n2452_), .A2(new_n617_), .B1(new_n510_), .B2(new_n2447_), .ZN(new_n3764_));
  NAND2_X1   g03508(.A1(new_n3312_), .A2(\b[8] ), .ZN(new_n3765_));
  AOI21_X1   g03509(.A1(new_n3764_), .A2(new_n3765_), .B(new_n2455_), .ZN(new_n3766_));
  NAND2_X1   g03510(.A1(new_n616_), .A2(new_n3766_), .ZN(new_n3767_));
  XOR2_X1    g03511(.A1(new_n3767_), .A2(\a[32] ), .Z(new_n3768_));
  XNOR2_X1   g03512(.A1(new_n3763_), .A2(new_n3768_), .ZN(new_n3769_));
  OAI22_X1   g03513(.A1(new_n2084_), .A2(new_n795_), .B1(new_n717_), .B2(new_n2079_), .ZN(new_n3770_));
  NAND2_X1   g03514(.A1(new_n2864_), .A2(\b[11] ), .ZN(new_n3771_));
  AOI21_X1   g03515(.A1(new_n3770_), .A2(new_n3771_), .B(new_n2087_), .ZN(new_n3772_));
  NAND2_X1   g03516(.A1(new_n799_), .A2(new_n3772_), .ZN(new_n3773_));
  XOR2_X1    g03517(.A1(new_n3773_), .A2(\a[29] ), .Z(new_n3774_));
  NOR2_X1    g03518(.A1(new_n3769_), .A2(new_n3774_), .ZN(new_n3775_));
  INV_X1     g03519(.I(new_n3775_), .ZN(new_n3776_));
  NAND2_X1   g03520(.A1(new_n3769_), .A2(new_n3774_), .ZN(new_n3777_));
  NAND2_X1   g03521(.A1(new_n3776_), .A2(new_n3777_), .ZN(new_n3778_));
  OAI22_X1   g03522(.A1(new_n1760_), .A2(new_n992_), .B1(new_n904_), .B2(new_n1755_), .ZN(new_n3779_));
  NAND2_X1   g03523(.A1(new_n2470_), .A2(\b[14] ), .ZN(new_n3780_));
  AOI21_X1   g03524(.A1(new_n3779_), .A2(new_n3780_), .B(new_n1763_), .ZN(new_n3781_));
  NAND2_X1   g03525(.A1(new_n991_), .A2(new_n3781_), .ZN(new_n3782_));
  XOR2_X1    g03526(.A1(new_n3782_), .A2(\a[26] ), .Z(new_n3783_));
  XOR2_X1    g03527(.A1(new_n3778_), .A2(new_n3783_), .Z(new_n3784_));
  OAI22_X1   g03528(.A1(new_n1444_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n1439_), .ZN(new_n3785_));
  NAND2_X1   g03529(.A1(new_n2098_), .A2(\b[17] ), .ZN(new_n3786_));
  AOI21_X1   g03530(.A1(new_n3785_), .A2(new_n3786_), .B(new_n1447_), .ZN(new_n3787_));
  NAND2_X1   g03531(.A1(new_n1225_), .A2(new_n3787_), .ZN(new_n3788_));
  XOR2_X1    g03532(.A1(new_n3788_), .A2(\a[23] ), .Z(new_n3789_));
  XNOR2_X1   g03533(.A1(new_n3784_), .A2(new_n3789_), .ZN(new_n3790_));
  OAI22_X1   g03534(.A1(new_n1168_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n1163_), .ZN(new_n3791_));
  NAND2_X1   g03535(.A1(new_n1774_), .A2(\b[20] ), .ZN(new_n3792_));
  AOI21_X1   g03536(.A1(new_n3791_), .A2(new_n3792_), .B(new_n1171_), .ZN(new_n3793_));
  NAND2_X1   g03537(.A1(new_n1517_), .A2(new_n3793_), .ZN(new_n3794_));
  XOR2_X1    g03538(.A1(new_n3794_), .A2(\a[20] ), .Z(new_n3795_));
  XOR2_X1    g03539(.A1(new_n3790_), .A2(new_n3795_), .Z(new_n3796_));
  NOR2_X1    g03540(.A1(new_n3718_), .A2(new_n3796_), .ZN(new_n3797_));
  INV_X1     g03541(.I(new_n3718_), .ZN(new_n3798_));
  INV_X1     g03542(.I(new_n3795_), .ZN(new_n3799_));
  XOR2_X1    g03543(.A1(new_n3790_), .A2(new_n3799_), .Z(new_n3800_));
  NOR2_X1    g03544(.A1(new_n3798_), .A2(new_n3800_), .ZN(new_n3801_));
  NOR2_X1    g03545(.A1(new_n3801_), .A2(new_n3797_), .ZN(new_n3802_));
  OAI22_X1   g03546(.A1(new_n940_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n935_), .ZN(new_n3803_));
  NAND2_X1   g03547(.A1(new_n1458_), .A2(\b[23] ), .ZN(new_n3804_));
  AOI21_X1   g03548(.A1(new_n3803_), .A2(new_n3804_), .B(new_n943_), .ZN(new_n3805_));
  NAND2_X1   g03549(.A1(new_n1828_), .A2(new_n3805_), .ZN(new_n3806_));
  XOR2_X1    g03550(.A1(new_n3806_), .A2(\a[17] ), .Z(new_n3807_));
  XNOR2_X1   g03551(.A1(new_n3802_), .A2(new_n3807_), .ZN(new_n3808_));
  OAI22_X1   g03552(.A1(new_n757_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n752_), .ZN(new_n3809_));
  NAND2_X1   g03553(.A1(new_n1182_), .A2(\b[26] ), .ZN(new_n3810_));
  AOI21_X1   g03554(.A1(new_n3809_), .A2(new_n3810_), .B(new_n760_), .ZN(new_n3811_));
  NAND2_X1   g03555(.A1(new_n2174_), .A2(new_n3811_), .ZN(new_n3812_));
  XOR2_X1    g03556(.A1(new_n3812_), .A2(\a[14] ), .Z(new_n3813_));
  XNOR2_X1   g03557(.A1(new_n3808_), .A2(new_n3813_), .ZN(new_n3814_));
  OAI22_X1   g03558(.A1(new_n582_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n577_), .ZN(new_n3815_));
  NAND2_X1   g03559(.A1(new_n960_), .A2(\b[29] ), .ZN(new_n3816_));
  AOI21_X1   g03560(.A1(new_n3815_), .A2(new_n3816_), .B(new_n585_), .ZN(new_n3817_));
  NAND2_X1   g03561(.A1(new_n2546_), .A2(new_n3817_), .ZN(new_n3818_));
  XOR2_X1    g03562(.A1(new_n3818_), .A2(new_n572_), .Z(new_n3819_));
  XNOR2_X1   g03563(.A1(new_n3814_), .A2(new_n3819_), .ZN(new_n3820_));
  INV_X1     g03564(.I(new_n3820_), .ZN(new_n3821_));
  XOR2_X1    g03565(.A1(new_n3814_), .A2(new_n3819_), .Z(new_n3822_));
  NOR2_X1    g03566(.A1(new_n3715_), .A2(new_n3822_), .ZN(new_n3823_));
  AOI21_X1   g03567(.A1(new_n3715_), .A2(new_n3821_), .B(new_n3823_), .ZN(new_n3824_));
  OAI22_X1   g03568(.A1(new_n437_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n431_), .ZN(new_n3825_));
  NAND2_X1   g03569(.A1(new_n775_), .A2(\b[32] ), .ZN(new_n3826_));
  AOI21_X1   g03570(.A1(new_n3825_), .A2(new_n3826_), .B(new_n440_), .ZN(new_n3827_));
  NAND2_X1   g03571(.A1(new_n2963_), .A2(new_n3827_), .ZN(new_n3828_));
  XOR2_X1    g03572(.A1(new_n3828_), .A2(\a[8] ), .Z(new_n3829_));
  XOR2_X1    g03573(.A1(new_n3824_), .A2(new_n3829_), .Z(new_n3830_));
  OAI22_X1   g03574(.A1(new_n364_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n320_), .ZN(new_n3831_));
  NAND2_X1   g03575(.A1(new_n594_), .A2(\b[35] ), .ZN(new_n3832_));
  AOI21_X1   g03576(.A1(new_n3831_), .A2(new_n3832_), .B(new_n312_), .ZN(new_n3833_));
  NAND2_X1   g03577(.A1(new_n3411_), .A2(new_n3833_), .ZN(new_n3834_));
  XOR2_X1    g03578(.A1(new_n3834_), .A2(\a[5] ), .Z(new_n3835_));
  XOR2_X1    g03579(.A1(new_n3830_), .A2(new_n3835_), .Z(new_n3836_));
  OAI21_X1   g03580(.A1(new_n3408_), .A2(new_n3696_), .B(new_n3566_), .ZN(new_n3837_));
  NAND2_X1   g03581(.A1(new_n3560_), .A2(new_n3837_), .ZN(new_n3838_));
  OAI21_X1   g03582(.A1(\b[37] ), .A2(\b[39] ), .B(\b[38] ), .ZN(new_n3839_));
  NAND2_X1   g03583(.A1(new_n3838_), .A2(new_n3839_), .ZN(new_n3840_));
  XOR2_X1    g03584(.A1(\b[39] ), .A2(\b[40] ), .Z(new_n3841_));
  NAND2_X1   g03585(.A1(new_n3840_), .A2(new_n3841_), .ZN(new_n3842_));
  XOR2_X1    g03586(.A1(\b[39] ), .A2(\b[40] ), .Z(new_n3843_));
  OAI21_X1   g03587(.A1(new_n3840_), .A2(new_n3843_), .B(new_n3842_), .ZN(new_n3844_));
  INV_X1     g03588(.I(\b[40] ), .ZN(new_n3845_));
  OAI22_X1   g03589(.A1(new_n405_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n404_), .ZN(new_n3846_));
  NAND2_X1   g03590(.A1(new_n279_), .A2(\b[38] ), .ZN(new_n3847_));
  AOI21_X1   g03591(.A1(new_n3846_), .A2(new_n3847_), .B(new_n264_), .ZN(new_n3848_));
  NAND2_X1   g03592(.A1(new_n3844_), .A2(new_n3848_), .ZN(new_n3849_));
  XOR2_X1    g03593(.A1(new_n3849_), .A2(\a[2] ), .Z(new_n3850_));
  INV_X1     g03594(.I(new_n3850_), .ZN(new_n3851_));
  XOR2_X1    g03595(.A1(new_n3836_), .A2(new_n3851_), .Z(new_n3852_));
  NOR2_X1    g03596(.A1(new_n3852_), .A2(new_n3713_), .ZN(new_n3853_));
  XOR2_X1    g03597(.A1(new_n3836_), .A2(new_n3850_), .Z(new_n3854_));
  AOI21_X1   g03598(.A1(new_n3689_), .A2(new_n3694_), .B(new_n3854_), .ZN(new_n3855_));
  NOR2_X1    g03599(.A1(new_n3855_), .A2(new_n3853_), .ZN(new_n3856_));
  INV_X1     g03600(.I(new_n3856_), .ZN(new_n3857_));
  NAND2_X1   g03601(.A1(new_n3710_), .A2(new_n3574_), .ZN(new_n3858_));
  NOR2_X1    g03602(.A1(new_n3858_), .A2(new_n3709_), .ZN(new_n3859_));
  OAI21_X1   g03603(.A1(new_n3707_), .A2(new_n3708_), .B(new_n3857_), .ZN(new_n3860_));
  OAI22_X1   g03604(.A1(new_n3859_), .A2(new_n3857_), .B1(new_n3858_), .B2(new_n3860_), .ZN(\f[40] ));
  XNOR2_X1   g03605(.A1(new_n3713_), .A2(new_n3836_), .ZN(new_n3862_));
  OAI22_X1   g03606(.A1(new_n3859_), .A2(new_n3856_), .B1(new_n3851_), .B2(new_n3862_), .ZN(new_n3863_));
  INV_X1     g03607(.I(new_n3829_), .ZN(new_n3864_));
  NAND2_X1   g03608(.A1(new_n3824_), .A2(new_n3864_), .ZN(new_n3865_));
  OAI22_X1   g03609(.A1(new_n940_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n935_), .ZN(new_n3866_));
  NAND2_X1   g03610(.A1(new_n1458_), .A2(\b[24] ), .ZN(new_n3867_));
  AOI21_X1   g03611(.A1(new_n3866_), .A2(new_n3867_), .B(new_n943_), .ZN(new_n3868_));
  NAND2_X1   g03612(.A1(new_n1926_), .A2(new_n3868_), .ZN(new_n3869_));
  XOR2_X1    g03613(.A1(new_n3869_), .A2(\a[17] ), .Z(new_n3870_));
  OAI22_X1   g03614(.A1(new_n1168_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n1163_), .ZN(new_n3871_));
  NAND2_X1   g03615(.A1(new_n1774_), .A2(\b[21] ), .ZN(new_n3872_));
  AOI21_X1   g03616(.A1(new_n3871_), .A2(new_n3872_), .B(new_n1171_), .ZN(new_n3873_));
  NAND2_X1   g03617(.A1(new_n1604_), .A2(new_n3873_), .ZN(new_n3874_));
  XOR2_X1    g03618(.A1(new_n3874_), .A2(\a[20] ), .Z(new_n3875_));
  INV_X1     g03619(.I(new_n3875_), .ZN(new_n3876_));
  INV_X1     g03620(.I(new_n3802_), .ZN(new_n3877_));
  XNOR2_X1   g03621(.A1(new_n3718_), .A2(new_n3790_), .ZN(new_n3878_));
  OAI21_X1   g03622(.A1(new_n3799_), .A2(new_n3878_), .B(new_n3877_), .ZN(new_n3879_));
  NOR2_X1    g03623(.A1(new_n3763_), .A2(new_n3768_), .ZN(new_n3880_));
  OAI22_X1   g03624(.A1(new_n3298_), .A2(new_n347_), .B1(new_n393_), .B2(new_n3293_), .ZN(new_n3881_));
  OAI21_X1   g03625(.A1(new_n290_), .A2(new_n3447_), .B(new_n3881_), .ZN(new_n3882_));
  AOI21_X1   g03626(.A1(new_n352_), .A2(new_n3300_), .B(new_n3882_), .ZN(new_n3883_));
  NAND2_X1   g03627(.A1(new_n3741_), .A2(new_n3742_), .ZN(new_n3884_));
  NOR2_X1    g03628(.A1(new_n3739_), .A2(new_n278_), .ZN(new_n3885_));
  XNOR2_X1   g03629(.A1(\a[38] ), .A2(\a[40] ), .ZN(new_n3886_));
  NAND2_X1   g03630(.A1(new_n3581_), .A2(new_n3886_), .ZN(new_n3887_));
  XNOR2_X1   g03631(.A1(\a[38] ), .A2(\a[41] ), .ZN(new_n3888_));
  NAND2_X1   g03632(.A1(new_n3887_), .A2(new_n3888_), .ZN(new_n3889_));
  OAI22_X1   g03633(.A1(new_n3736_), .A2(new_n292_), .B1(new_n267_), .B2(new_n3731_), .ZN(new_n3890_));
  NOR4_X1    g03634(.A1(new_n3890_), .A2(new_n258_), .A3(new_n3885_), .A4(new_n3889_), .ZN(new_n3891_));
  XOR2_X1    g03635(.A1(new_n3891_), .A2(new_n3726_), .Z(new_n3892_));
  XNOR2_X1   g03636(.A1(new_n3884_), .A2(new_n3892_), .ZN(new_n3893_));
  XOR2_X1    g03637(.A1(new_n3893_), .A2(\a[38] ), .Z(new_n3894_));
  XOR2_X1    g03638(.A1(new_n3894_), .A2(new_n3883_), .Z(new_n3895_));
  OAI21_X1   g03639(.A1(new_n3746_), .A2(new_n3743_), .B(new_n3747_), .ZN(new_n3896_));
  XNOR2_X1   g03640(.A1(new_n3895_), .A2(new_n3896_), .ZN(new_n3897_));
  OAI22_X1   g03641(.A1(new_n2846_), .A2(new_n495_), .B1(new_n450_), .B2(new_n2841_), .ZN(new_n3898_));
  NAND2_X1   g03642(.A1(new_n3755_), .A2(\b[6] ), .ZN(new_n3899_));
  AOI21_X1   g03643(.A1(new_n3898_), .A2(new_n3899_), .B(new_n2849_), .ZN(new_n3900_));
  NAND2_X1   g03644(.A1(new_n494_), .A2(new_n3900_), .ZN(new_n3901_));
  XOR2_X1    g03645(.A1(new_n3901_), .A2(\a[35] ), .Z(new_n3902_));
  XNOR2_X1   g03646(.A1(new_n3897_), .A2(new_n3902_), .ZN(new_n3903_));
  XOR2_X1    g03647(.A1(new_n3903_), .A2(new_n3760_), .Z(new_n3904_));
  OAI22_X1   g03648(.A1(new_n2452_), .A2(new_n659_), .B1(new_n617_), .B2(new_n2447_), .ZN(new_n3905_));
  NAND2_X1   g03649(.A1(new_n3312_), .A2(\b[9] ), .ZN(new_n3906_));
  AOI21_X1   g03650(.A1(new_n3905_), .A2(new_n3906_), .B(new_n2455_), .ZN(new_n3907_));
  NAND2_X1   g03651(.A1(new_n663_), .A2(new_n3907_), .ZN(new_n3908_));
  XOR2_X1    g03652(.A1(new_n3908_), .A2(\a[32] ), .Z(new_n3909_));
  XNOR2_X1   g03653(.A1(new_n3904_), .A2(new_n3909_), .ZN(new_n3910_));
  OAI22_X1   g03654(.A1(new_n2084_), .A2(new_n848_), .B1(new_n795_), .B2(new_n2079_), .ZN(new_n3911_));
  NAND2_X1   g03655(.A1(new_n2864_), .A2(\b[12] ), .ZN(new_n3912_));
  AOI21_X1   g03656(.A1(new_n3911_), .A2(new_n3912_), .B(new_n2087_), .ZN(new_n3913_));
  NAND2_X1   g03657(.A1(new_n847_), .A2(new_n3913_), .ZN(new_n3914_));
  XOR2_X1    g03658(.A1(new_n3914_), .A2(\a[29] ), .Z(new_n3915_));
  XNOR2_X1   g03659(.A1(new_n3910_), .A2(new_n3915_), .ZN(new_n3916_));
  XOR2_X1    g03660(.A1(new_n3910_), .A2(new_n3915_), .Z(new_n3917_));
  MUX2_X1    g03661(.I0(new_n3917_), .I1(new_n3916_), .S(new_n3880_), .Z(new_n3918_));
  XOR2_X1    g03662(.A1(new_n3918_), .A2(new_n3776_), .Z(new_n3919_));
  OAI22_X1   g03663(.A1(new_n1760_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n1755_), .ZN(new_n3920_));
  NAND2_X1   g03664(.A1(new_n2470_), .A2(\b[15] ), .ZN(new_n3921_));
  AOI21_X1   g03665(.A1(new_n3920_), .A2(new_n3921_), .B(new_n1763_), .ZN(new_n3922_));
  NAND2_X1   g03666(.A1(new_n1047_), .A2(new_n3922_), .ZN(new_n3923_));
  XOR2_X1    g03667(.A1(new_n3923_), .A2(\a[26] ), .Z(new_n3924_));
  XOR2_X1    g03668(.A1(new_n3919_), .A2(new_n3924_), .Z(new_n3925_));
  NOR2_X1    g03669(.A1(new_n3778_), .A2(new_n3783_), .ZN(new_n3926_));
  XOR2_X1    g03670(.A1(new_n3925_), .A2(new_n3926_), .Z(new_n3927_));
  OAI22_X1   g03671(.A1(new_n1444_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n1439_), .ZN(new_n3928_));
  NAND2_X1   g03672(.A1(new_n2098_), .A2(\b[18] ), .ZN(new_n3929_));
  AOI21_X1   g03673(.A1(new_n3928_), .A2(new_n3929_), .B(new_n1447_), .ZN(new_n3930_));
  NAND2_X1   g03674(.A1(new_n1304_), .A2(new_n3930_), .ZN(new_n3931_));
  XOR2_X1    g03675(.A1(new_n3931_), .A2(\a[23] ), .Z(new_n3932_));
  INV_X1     g03676(.I(new_n3932_), .ZN(new_n3933_));
  XOR2_X1    g03677(.A1(new_n3927_), .A2(new_n3933_), .Z(new_n3934_));
  INV_X1     g03678(.I(new_n3934_), .ZN(new_n3935_));
  INV_X1     g03679(.I(new_n3789_), .ZN(new_n3936_));
  NAND2_X1   g03680(.A1(new_n3718_), .A2(new_n3790_), .ZN(new_n3937_));
  OAI21_X1   g03681(.A1(new_n3784_), .A2(new_n3936_), .B(new_n3937_), .ZN(new_n3938_));
  NOR2_X1    g03682(.A1(new_n3938_), .A2(new_n3935_), .ZN(new_n3939_));
  NAND2_X1   g03683(.A1(new_n3938_), .A2(new_n3935_), .ZN(new_n3940_));
  INV_X1     g03684(.I(new_n3940_), .ZN(new_n3941_));
  NOR2_X1    g03685(.A1(new_n3941_), .A2(new_n3939_), .ZN(new_n3942_));
  XOR2_X1    g03686(.A1(new_n3942_), .A2(new_n3879_), .Z(new_n3943_));
  XOR2_X1    g03687(.A1(new_n3943_), .A2(new_n3876_), .Z(new_n3944_));
  XOR2_X1    g03688(.A1(new_n3944_), .A2(new_n3870_), .Z(new_n3945_));
  NOR2_X1    g03689(.A1(new_n3877_), .A2(new_n3807_), .ZN(new_n3946_));
  XOR2_X1    g03690(.A1(new_n3945_), .A2(new_n3946_), .Z(new_n3947_));
  OAI22_X1   g03691(.A1(new_n757_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n752_), .ZN(new_n3948_));
  NAND2_X1   g03692(.A1(new_n1182_), .A2(\b[27] ), .ZN(new_n3949_));
  AOI21_X1   g03693(.A1(new_n3948_), .A2(new_n3949_), .B(new_n760_), .ZN(new_n3950_));
  NAND2_X1   g03694(.A1(new_n2276_), .A2(new_n3950_), .ZN(new_n3951_));
  XOR2_X1    g03695(.A1(new_n3951_), .A2(\a[14] ), .Z(new_n3952_));
  XOR2_X1    g03696(.A1(new_n3947_), .A2(new_n3952_), .Z(new_n3953_));
  INV_X1     g03697(.I(new_n3953_), .ZN(new_n3954_));
  INV_X1     g03698(.I(new_n3808_), .ZN(new_n3955_));
  NOR2_X1    g03699(.A1(new_n3955_), .A2(new_n3813_), .ZN(new_n3956_));
  INV_X1     g03700(.I(new_n3956_), .ZN(new_n3957_));
  NOR2_X1    g03701(.A1(new_n3954_), .A2(new_n3957_), .ZN(new_n3958_));
  INV_X1     g03702(.I(new_n3958_), .ZN(new_n3959_));
  NAND2_X1   g03703(.A1(new_n3954_), .A2(new_n3957_), .ZN(new_n3960_));
  NAND2_X1   g03704(.A1(new_n3959_), .A2(new_n3960_), .ZN(new_n3961_));
  OAI22_X1   g03705(.A1(new_n582_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n577_), .ZN(new_n3962_));
  NAND2_X1   g03706(.A1(new_n960_), .A2(\b[30] ), .ZN(new_n3963_));
  AOI21_X1   g03707(.A1(new_n3962_), .A2(new_n3963_), .B(new_n585_), .ZN(new_n3964_));
  NAND2_X1   g03708(.A1(new_n2659_), .A2(new_n3964_), .ZN(new_n3965_));
  XOR2_X1    g03709(.A1(new_n3965_), .A2(\a[11] ), .Z(new_n3966_));
  XNOR2_X1   g03710(.A1(new_n3961_), .A2(new_n3966_), .ZN(new_n3967_));
  NAND2_X1   g03711(.A1(new_n3715_), .A2(new_n3814_), .ZN(new_n3968_));
  XOR2_X1    g03712(.A1(new_n3968_), .A2(new_n3967_), .Z(new_n3969_));
  XOR2_X1    g03713(.A1(new_n3715_), .A2(new_n3814_), .Z(new_n3970_));
  NAND2_X1   g03714(.A1(new_n3970_), .A2(new_n3819_), .ZN(new_n3971_));
  XOR2_X1    g03715(.A1(new_n3969_), .A2(new_n3971_), .Z(new_n3972_));
  OAI22_X1   g03716(.A1(new_n437_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n431_), .ZN(new_n3973_));
  NAND2_X1   g03717(.A1(new_n775_), .A2(\b[33] ), .ZN(new_n3974_));
  AOI21_X1   g03718(.A1(new_n3973_), .A2(new_n3974_), .B(new_n440_), .ZN(new_n3975_));
  NAND2_X1   g03719(.A1(new_n3101_), .A2(new_n3975_), .ZN(new_n3976_));
  XOR2_X1    g03720(.A1(new_n3976_), .A2(\a[8] ), .Z(new_n3977_));
  XOR2_X1    g03721(.A1(new_n3972_), .A2(new_n3977_), .Z(new_n3978_));
  OAI22_X1   g03722(.A1(new_n364_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n320_), .ZN(new_n3979_));
  NAND2_X1   g03723(.A1(new_n594_), .A2(\b[36] ), .ZN(new_n3980_));
  AOI21_X1   g03724(.A1(new_n3979_), .A2(new_n3980_), .B(new_n312_), .ZN(new_n3981_));
  NAND2_X1   g03725(.A1(new_n3565_), .A2(new_n3981_), .ZN(new_n3982_));
  XOR2_X1    g03726(.A1(new_n3982_), .A2(\a[5] ), .Z(new_n3983_));
  XOR2_X1    g03727(.A1(new_n3978_), .A2(new_n3983_), .Z(new_n3984_));
  XOR2_X1    g03728(.A1(new_n3978_), .A2(new_n3983_), .Z(new_n3985_));
  NAND2_X1   g03729(.A1(new_n3985_), .A2(new_n3865_), .ZN(new_n3986_));
  OAI21_X1   g03730(.A1(new_n3865_), .A2(new_n3984_), .B(new_n3986_), .ZN(new_n3987_));
  NAND2_X1   g03731(.A1(new_n3830_), .A2(new_n3835_), .ZN(new_n3988_));
  NAND3_X1   g03732(.A1(new_n3713_), .A2(new_n3988_), .A3(new_n3836_), .ZN(new_n3989_));
  XNOR2_X1   g03733(.A1(new_n3987_), .A2(new_n3989_), .ZN(new_n3990_));
  XOR2_X1    g03734(.A1(new_n3840_), .A2(\b[39] ), .Z(new_n3991_));
  NAND2_X1   g03735(.A1(new_n3991_), .A2(new_n3841_), .ZN(new_n3992_));
  NOR2_X1    g03736(.A1(new_n3992_), .A2(\b[41] ), .ZN(new_n3993_));
  INV_X1     g03737(.I(new_n3993_), .ZN(new_n3994_));
  NAND2_X1   g03738(.A1(new_n3992_), .A2(\b[41] ), .ZN(new_n3995_));
  NAND2_X1   g03739(.A1(new_n3994_), .A2(new_n3995_), .ZN(new_n3996_));
  INV_X1     g03740(.I(\b[41] ), .ZN(new_n3997_));
  OAI22_X1   g03741(.A1(new_n405_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n404_), .ZN(new_n3998_));
  NAND2_X1   g03742(.A1(new_n279_), .A2(\b[39] ), .ZN(new_n3999_));
  AOI21_X1   g03743(.A1(new_n3998_), .A2(new_n3999_), .B(new_n264_), .ZN(new_n4000_));
  NAND2_X1   g03744(.A1(new_n3996_), .A2(new_n4000_), .ZN(new_n4001_));
  XOR2_X1    g03745(.A1(new_n4001_), .A2(\a[2] ), .Z(new_n4002_));
  INV_X1     g03746(.I(new_n4002_), .ZN(new_n4003_));
  XOR2_X1    g03747(.A1(new_n3990_), .A2(new_n4003_), .Z(new_n4004_));
  NAND2_X1   g03748(.A1(new_n3990_), .A2(new_n4003_), .ZN(new_n4005_));
  NOR2_X1    g03749(.A1(new_n3990_), .A2(new_n4003_), .ZN(new_n4006_));
  INV_X1     g03750(.I(new_n4006_), .ZN(new_n4007_));
  NAND2_X1   g03751(.A1(new_n4007_), .A2(new_n4005_), .ZN(new_n4008_));
  MUX2_X1    g03752(.I0(new_n4008_), .I1(new_n4004_), .S(new_n3863_), .Z(\f[41] ));
  OAI21_X1   g03753(.A1(new_n3696_), .A2(new_n3997_), .B(new_n3845_), .ZN(new_n4010_));
  NAND3_X1   g03754(.A1(new_n3838_), .A2(new_n3839_), .A3(new_n4010_), .ZN(new_n4011_));
  OAI21_X1   g03755(.A1(\b[39] ), .A2(\b[41] ), .B(\b[40] ), .ZN(new_n4012_));
  NAND2_X1   g03756(.A1(new_n4011_), .A2(new_n4012_), .ZN(new_n4013_));
  XOR2_X1    g03757(.A1(\b[41] ), .A2(\b[42] ), .Z(new_n4014_));
  NAND2_X1   g03758(.A1(new_n4013_), .A2(new_n4014_), .ZN(new_n4015_));
  XOR2_X1    g03759(.A1(\b[41] ), .A2(\b[42] ), .Z(new_n4016_));
  OAI21_X1   g03760(.A1(new_n4013_), .A2(new_n4016_), .B(new_n4015_), .ZN(new_n4017_));
  INV_X1     g03761(.I(\b[42] ), .ZN(new_n4018_));
  OAI22_X1   g03762(.A1(new_n405_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n404_), .ZN(new_n4019_));
  NAND2_X1   g03763(.A1(new_n279_), .A2(\b[40] ), .ZN(new_n4020_));
  AOI21_X1   g03764(.A1(new_n4019_), .A2(new_n4020_), .B(new_n264_), .ZN(new_n4021_));
  NAND2_X1   g03765(.A1(new_n4017_), .A2(new_n4021_), .ZN(new_n4022_));
  XOR2_X1    g03766(.A1(new_n4022_), .A2(\a[2] ), .Z(new_n4023_));
  OAI22_X1   g03767(.A1(new_n364_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n320_), .ZN(new_n4024_));
  NAND2_X1   g03768(.A1(new_n594_), .A2(\b[37] ), .ZN(new_n4025_));
  AOI21_X1   g03769(.A1(new_n4024_), .A2(new_n4025_), .B(new_n312_), .ZN(new_n4026_));
  NAND2_X1   g03770(.A1(new_n3700_), .A2(new_n4026_), .ZN(new_n4027_));
  XOR2_X1    g03771(.A1(new_n4027_), .A2(\a[5] ), .Z(new_n4028_));
  INV_X1     g03772(.I(new_n4028_), .ZN(new_n4029_));
  XNOR2_X1   g03773(.A1(new_n3978_), .A2(new_n3865_), .ZN(new_n4030_));
  NAND2_X1   g03774(.A1(new_n4030_), .A2(new_n3983_), .ZN(new_n4031_));
  NAND2_X1   g03775(.A1(new_n3987_), .A2(new_n3989_), .ZN(new_n4032_));
  NAND2_X1   g03776(.A1(new_n4032_), .A2(new_n4031_), .ZN(new_n4033_));
  INV_X1     g03777(.I(new_n3884_), .ZN(new_n4034_));
  NAND2_X1   g03778(.A1(new_n4034_), .A2(new_n3892_), .ZN(new_n4035_));
  NOR2_X1    g03779(.A1(new_n3889_), .A2(new_n267_), .ZN(new_n4036_));
  OAI22_X1   g03780(.A1(new_n3736_), .A2(new_n290_), .B1(new_n292_), .B2(new_n3731_), .ZN(new_n4037_));
  NOR4_X1    g03781(.A1(new_n4037_), .A2(new_n677_), .A3(new_n3739_), .A4(new_n4036_), .ZN(new_n4038_));
  XOR2_X1    g03782(.A1(new_n4038_), .A2(new_n3726_), .Z(new_n4039_));
  XNOR2_X1   g03783(.A1(\a[41] ), .A2(\a[42] ), .ZN(new_n4040_));
  NOR2_X1    g03784(.A1(new_n4040_), .A2(new_n258_), .ZN(new_n4041_));
  XOR2_X1    g03785(.A1(new_n4039_), .A2(new_n4041_), .Z(new_n4042_));
  XNOR2_X1   g03786(.A1(new_n4042_), .A2(new_n4035_), .ZN(new_n4043_));
  INV_X1     g03787(.I(new_n3293_), .ZN(new_n4044_));
  AOI22_X1   g03788(.A1(\b[6] ), .A2(new_n3297_), .B1(new_n4044_), .B2(\b[5] ), .ZN(new_n4045_));
  NOR2_X1    g03789(.A1(new_n3447_), .A2(new_n393_), .ZN(new_n4046_));
  OAI21_X1   g03790(.A1(new_n4045_), .A2(new_n4046_), .B(new_n3300_), .ZN(new_n4047_));
  NOR2_X1    g03791(.A1(new_n524_), .A2(new_n4047_), .ZN(new_n4048_));
  XOR2_X1    g03792(.A1(new_n4048_), .A2(new_n3288_), .Z(new_n4049_));
  NAND2_X1   g03793(.A1(new_n3721_), .A2(new_n3748_), .ZN(new_n4050_));
  NAND2_X1   g03794(.A1(new_n3883_), .A2(new_n3288_), .ZN(new_n4051_));
  NOR2_X1    g03795(.A1(new_n3883_), .A2(new_n3288_), .ZN(new_n4052_));
  NAND2_X1   g03796(.A1(new_n3749_), .A2(new_n3893_), .ZN(new_n4053_));
  NOR2_X1    g03797(.A1(new_n4053_), .A2(new_n4052_), .ZN(new_n4054_));
  NAND4_X1   g03798(.A1(new_n3895_), .A2(new_n4050_), .A3(new_n4051_), .A4(new_n4054_), .ZN(new_n4055_));
  XOR2_X1    g03799(.A1(new_n4055_), .A2(new_n4049_), .Z(new_n4056_));
  XNOR2_X1   g03800(.A1(new_n4056_), .A2(new_n4043_), .ZN(new_n4057_));
  OAI22_X1   g03801(.A1(new_n2846_), .A2(new_n510_), .B1(new_n495_), .B2(new_n2841_), .ZN(new_n4058_));
  NAND2_X1   g03802(.A1(new_n3755_), .A2(\b[7] ), .ZN(new_n4059_));
  AOI21_X1   g03803(.A1(new_n4058_), .A2(new_n4059_), .B(new_n2849_), .ZN(new_n4060_));
  NAND2_X1   g03804(.A1(new_n518_), .A2(new_n4060_), .ZN(new_n4061_));
  XOR2_X1    g03805(.A1(new_n4061_), .A2(\a[35] ), .Z(new_n4062_));
  INV_X1     g03806(.I(new_n3897_), .ZN(new_n4063_));
  NAND2_X1   g03807(.A1(new_n4063_), .A2(new_n3902_), .ZN(new_n4064_));
  NAND3_X1   g03808(.A1(new_n3903_), .A2(new_n3762_), .A3(new_n4064_), .ZN(new_n4065_));
  XOR2_X1    g03809(.A1(new_n4065_), .A2(new_n4062_), .Z(new_n4066_));
  XNOR2_X1   g03810(.A1(new_n4066_), .A2(new_n4057_), .ZN(new_n4067_));
  OAI22_X1   g03811(.A1(new_n2452_), .A2(new_n717_), .B1(new_n659_), .B2(new_n2447_), .ZN(new_n4068_));
  NAND2_X1   g03812(.A1(new_n3312_), .A2(\b[10] ), .ZN(new_n4069_));
  AOI21_X1   g03813(.A1(new_n4068_), .A2(new_n4069_), .B(new_n2455_), .ZN(new_n4070_));
  NAND2_X1   g03814(.A1(new_n716_), .A2(new_n4070_), .ZN(new_n4071_));
  XOR2_X1    g03815(.A1(new_n4071_), .A2(new_n2442_), .Z(new_n4072_));
  AOI21_X1   g03816(.A1(new_n3904_), .A2(new_n3909_), .B(new_n3880_), .ZN(new_n4073_));
  XOR2_X1    g03817(.A1(new_n4073_), .A2(new_n4072_), .Z(new_n4074_));
  XNOR2_X1   g03818(.A1(new_n4067_), .A2(new_n4074_), .ZN(new_n4075_));
  OAI22_X1   g03819(.A1(new_n2084_), .A2(new_n904_), .B1(new_n848_), .B2(new_n2079_), .ZN(new_n4076_));
  NAND2_X1   g03820(.A1(new_n2864_), .A2(\b[13] ), .ZN(new_n4077_));
  AOI21_X1   g03821(.A1(new_n4076_), .A2(new_n4077_), .B(new_n2087_), .ZN(new_n4078_));
  NAND2_X1   g03822(.A1(new_n907_), .A2(new_n4078_), .ZN(new_n4079_));
  XOR2_X1    g03823(.A1(new_n4079_), .A2(\a[29] ), .Z(new_n4080_));
  XOR2_X1    g03824(.A1(new_n3910_), .A2(new_n3880_), .Z(new_n4081_));
  NAND2_X1   g03825(.A1(new_n4081_), .A2(new_n3915_), .ZN(new_n4082_));
  XOR2_X1    g03826(.A1(new_n4082_), .A2(new_n4080_), .Z(new_n4083_));
  XOR2_X1    g03827(.A1(new_n4083_), .A2(new_n4075_), .Z(new_n4084_));
  OAI22_X1   g03828(.A1(new_n1760_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n1755_), .ZN(new_n4085_));
  NAND2_X1   g03829(.A1(new_n2470_), .A2(\b[16] ), .ZN(new_n4086_));
  AOI21_X1   g03830(.A1(new_n4085_), .A2(new_n4086_), .B(new_n1763_), .ZN(new_n4087_));
  NAND2_X1   g03831(.A1(new_n1123_), .A2(new_n4087_), .ZN(new_n4088_));
  XOR2_X1    g03832(.A1(new_n4088_), .A2(\a[26] ), .Z(new_n4089_));
  INV_X1     g03833(.I(new_n4089_), .ZN(new_n4090_));
  INV_X1     g03834(.I(new_n3924_), .ZN(new_n4091_));
  NAND2_X1   g03835(.A1(new_n3925_), .A2(new_n3926_), .ZN(new_n4092_));
  OAI21_X1   g03836(.A1(new_n3919_), .A2(new_n4091_), .B(new_n4092_), .ZN(new_n4093_));
  XOR2_X1    g03837(.A1(new_n4093_), .A2(new_n4090_), .Z(new_n4094_));
  XOR2_X1    g03838(.A1(new_n4094_), .A2(new_n4084_), .Z(new_n4095_));
  OAI22_X1   g03839(.A1(new_n1444_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n1439_), .ZN(new_n4096_));
  NAND2_X1   g03840(.A1(new_n2098_), .A2(\b[19] ), .ZN(new_n4097_));
  AOI21_X1   g03841(.A1(new_n4096_), .A2(new_n4097_), .B(new_n1447_), .ZN(new_n4098_));
  NAND2_X1   g03842(.A1(new_n1396_), .A2(new_n4098_), .ZN(new_n4099_));
  XOR2_X1    g03843(.A1(new_n4099_), .A2(\a[23] ), .Z(new_n4100_));
  NOR2_X1    g03844(.A1(new_n3927_), .A2(new_n3933_), .ZN(new_n4101_));
  NOR2_X1    g03845(.A1(new_n3935_), .A2(new_n4101_), .ZN(new_n4102_));
  NAND2_X1   g03846(.A1(new_n3938_), .A2(new_n4102_), .ZN(new_n4103_));
  XOR2_X1    g03847(.A1(new_n4103_), .A2(new_n4100_), .Z(new_n4104_));
  XNOR2_X1   g03848(.A1(new_n4104_), .A2(new_n4095_), .ZN(new_n4105_));
  OAI22_X1   g03849(.A1(new_n1168_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n1163_), .ZN(new_n4106_));
  NAND2_X1   g03850(.A1(new_n1774_), .A2(\b[22] ), .ZN(new_n4107_));
  AOI21_X1   g03851(.A1(new_n4106_), .A2(new_n4107_), .B(new_n1171_), .ZN(new_n4108_));
  NAND2_X1   g03852(.A1(new_n1708_), .A2(new_n4108_), .ZN(new_n4109_));
  XOR2_X1    g03853(.A1(new_n4109_), .A2(new_n1158_), .Z(new_n4110_));
  NAND2_X1   g03854(.A1(new_n3942_), .A2(new_n3875_), .ZN(new_n4111_));
  NOR2_X1    g03855(.A1(new_n3942_), .A2(new_n3875_), .ZN(new_n4112_));
  NOR2_X1    g03856(.A1(new_n4112_), .A2(new_n3879_), .ZN(new_n4113_));
  NOR2_X1    g03857(.A1(new_n3942_), .A2(new_n3876_), .ZN(new_n4114_));
  AOI21_X1   g03858(.A1(new_n4113_), .A2(new_n4111_), .B(new_n4114_), .ZN(new_n4115_));
  XOR2_X1    g03859(.A1(new_n4115_), .A2(new_n4110_), .Z(new_n4116_));
  XNOR2_X1   g03860(.A1(new_n4116_), .A2(new_n4105_), .ZN(new_n4117_));
  OAI22_X1   g03861(.A1(new_n940_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n935_), .ZN(new_n4118_));
  NAND2_X1   g03862(.A1(new_n1458_), .A2(\b[25] ), .ZN(new_n4119_));
  AOI21_X1   g03863(.A1(new_n4118_), .A2(new_n4119_), .B(new_n943_), .ZN(new_n4120_));
  NAND2_X1   g03864(.A1(new_n2042_), .A2(new_n4120_), .ZN(new_n4121_));
  XOR2_X1    g03865(.A1(new_n4121_), .A2(new_n930_), .Z(new_n4122_));
  XOR2_X1    g03866(.A1(new_n3942_), .A2(new_n3876_), .Z(new_n4123_));
  XOR2_X1    g03867(.A1(new_n4123_), .A2(new_n3879_), .Z(new_n4124_));
  AOI22_X1   g03868(.A1(new_n3945_), .A2(new_n3946_), .B1(new_n3870_), .B2(new_n4124_), .ZN(new_n4125_));
  XOR2_X1    g03869(.A1(new_n4125_), .A2(new_n4122_), .Z(new_n4126_));
  XNOR2_X1   g03870(.A1(new_n4126_), .A2(new_n4117_), .ZN(new_n4127_));
  INV_X1     g03871(.I(new_n4127_), .ZN(new_n4128_));
  OAI22_X1   g03872(.A1(new_n757_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n752_), .ZN(new_n4129_));
  NAND2_X1   g03873(.A1(new_n1182_), .A2(\b[28] ), .ZN(new_n4130_));
  AOI21_X1   g03874(.A1(new_n4129_), .A2(new_n4130_), .B(new_n760_), .ZN(new_n4131_));
  NAND2_X1   g03875(.A1(new_n2404_), .A2(new_n4131_), .ZN(new_n4132_));
  XOR2_X1    g03876(.A1(new_n4132_), .A2(\a[14] ), .Z(new_n4133_));
  INV_X1     g03877(.I(new_n3952_), .ZN(new_n4134_));
  OAI21_X1   g03878(.A1(new_n3947_), .A2(new_n4134_), .B(new_n3959_), .ZN(new_n4135_));
  XOR2_X1    g03879(.A1(new_n4135_), .A2(new_n4133_), .Z(new_n4136_));
  XOR2_X1    g03880(.A1(new_n4136_), .A2(new_n4128_), .Z(new_n4137_));
  OAI22_X1   g03881(.A1(new_n582_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n577_), .ZN(new_n4138_));
  NAND2_X1   g03882(.A1(new_n960_), .A2(\b[31] ), .ZN(new_n4139_));
  AOI21_X1   g03883(.A1(new_n4138_), .A2(new_n4139_), .B(new_n585_), .ZN(new_n4140_));
  NAND2_X1   g03884(.A1(new_n2797_), .A2(new_n4140_), .ZN(new_n4141_));
  XOR2_X1    g03885(.A1(new_n4141_), .A2(\a[11] ), .Z(new_n4142_));
  NAND2_X1   g03886(.A1(new_n3967_), .A2(new_n3819_), .ZN(new_n4143_));
  NAND3_X1   g03887(.A1(new_n3715_), .A2(new_n3814_), .A3(new_n4143_), .ZN(new_n4144_));
  NAND2_X1   g03888(.A1(new_n3961_), .A2(new_n3966_), .ZN(new_n4145_));
  NAND2_X1   g03889(.A1(new_n4144_), .A2(new_n4145_), .ZN(new_n4146_));
  XOR2_X1    g03890(.A1(new_n4146_), .A2(new_n4142_), .Z(new_n4147_));
  XNOR2_X1   g03891(.A1(new_n4147_), .A2(new_n4137_), .ZN(new_n4148_));
  OAI22_X1   g03892(.A1(new_n437_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n431_), .ZN(new_n4149_));
  NAND2_X1   g03893(.A1(new_n775_), .A2(\b[34] ), .ZN(new_n4150_));
  AOI21_X1   g03894(.A1(new_n4149_), .A2(new_n4150_), .B(new_n440_), .ZN(new_n4151_));
  NAND2_X1   g03895(.A1(new_n3246_), .A2(new_n4151_), .ZN(new_n4152_));
  XOR2_X1    g03896(.A1(new_n4152_), .A2(\a[8] ), .Z(new_n4153_));
  INV_X1     g03897(.I(new_n3977_), .ZN(new_n4154_));
  NOR2_X1    g03898(.A1(new_n3972_), .A2(new_n4154_), .ZN(new_n4155_));
  NOR2_X1    g03899(.A1(new_n3824_), .A2(new_n3864_), .ZN(new_n4156_));
  NOR3_X1    g03900(.A1(new_n3978_), .A2(new_n4155_), .A3(new_n4156_), .ZN(new_n4157_));
  XNOR2_X1   g03901(.A1(new_n4157_), .A2(new_n4153_), .ZN(new_n4158_));
  XNOR2_X1   g03902(.A1(new_n4158_), .A2(new_n4148_), .ZN(new_n4159_));
  XOR2_X1    g03903(.A1(new_n4033_), .A2(new_n4159_), .Z(new_n4160_));
  XOR2_X1    g03904(.A1(new_n4160_), .A2(new_n4029_), .Z(new_n4161_));
  XOR2_X1    g03905(.A1(new_n4161_), .A2(new_n4023_), .Z(new_n4162_));
  OAI21_X1   g03906(.A1(new_n3863_), .A2(new_n3990_), .B(new_n4003_), .ZN(new_n4163_));
  XNOR2_X1   g03907(.A1(new_n4162_), .A2(new_n4163_), .ZN(\f[42] ));
  OAI22_X1   g03908(.A1(new_n364_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n320_), .ZN(new_n4165_));
  NAND2_X1   g03909(.A1(new_n594_), .A2(\b[38] ), .ZN(new_n4166_));
  AOI21_X1   g03910(.A1(new_n4165_), .A2(new_n4166_), .B(new_n312_), .ZN(new_n4167_));
  NAND2_X1   g03911(.A1(new_n3844_), .A2(new_n4167_), .ZN(new_n4168_));
  XOR2_X1    g03912(.A1(new_n4168_), .A2(\a[5] ), .Z(new_n4169_));
  OAI22_X1   g03913(.A1(new_n437_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n431_), .ZN(new_n4170_));
  NAND2_X1   g03914(.A1(new_n775_), .A2(\b[35] ), .ZN(new_n4171_));
  AOI21_X1   g03915(.A1(new_n4170_), .A2(new_n4171_), .B(new_n440_), .ZN(new_n4172_));
  NAND2_X1   g03916(.A1(new_n3411_), .A2(new_n4172_), .ZN(new_n4173_));
  XOR2_X1    g03917(.A1(new_n4173_), .A2(\a[8] ), .Z(new_n4174_));
  XOR2_X1    g03918(.A1(new_n4148_), .A2(new_n4153_), .Z(new_n4175_));
  NAND2_X1   g03919(.A1(new_n4175_), .A2(new_n4153_), .ZN(new_n4176_));
  NAND2_X1   g03920(.A1(new_n4157_), .A2(new_n4175_), .ZN(new_n4177_));
  NAND2_X1   g03921(.A1(new_n4177_), .A2(new_n4176_), .ZN(new_n4178_));
  NAND2_X1   g03922(.A1(new_n4128_), .A2(new_n4133_), .ZN(new_n4179_));
  INV_X1     g03923(.I(new_n4135_), .ZN(new_n4180_));
  XOR2_X1    g03924(.A1(new_n4127_), .A2(new_n4133_), .Z(new_n4181_));
  NAND2_X1   g03925(.A1(new_n4180_), .A2(new_n4181_), .ZN(new_n4182_));
  XOR2_X1    g03926(.A1(new_n4084_), .A2(new_n4090_), .Z(new_n4183_));
  AOI21_X1   g03927(.A1(new_n4093_), .A2(new_n4090_), .B(new_n4183_), .ZN(new_n4184_));
  INV_X1     g03928(.I(new_n4184_), .ZN(new_n4185_));
  XOR2_X1    g03929(.A1(new_n4075_), .A2(new_n4080_), .Z(new_n4186_));
  NAND2_X1   g03930(.A1(new_n4186_), .A2(new_n4080_), .ZN(new_n4187_));
  NAND2_X1   g03931(.A1(new_n4186_), .A2(new_n4082_), .ZN(new_n4188_));
  NAND2_X1   g03932(.A1(new_n4188_), .A2(new_n4187_), .ZN(new_n4189_));
  NAND2_X1   g03933(.A1(new_n4042_), .A2(new_n3892_), .ZN(new_n4190_));
  NAND2_X1   g03934(.A1(new_n4190_), .A2(new_n3884_), .ZN(new_n4191_));
  NAND2_X1   g03935(.A1(new_n4039_), .A2(new_n4041_), .ZN(new_n4192_));
  XNOR2_X1   g03936(.A1(new_n4191_), .A2(new_n4192_), .ZN(new_n4193_));
  OAI22_X1   g03937(.A1(new_n3736_), .A2(new_n393_), .B1(new_n290_), .B2(new_n3731_), .ZN(new_n4194_));
  OAI21_X1   g03938(.A1(new_n292_), .A2(new_n3889_), .B(new_n4194_), .ZN(new_n4195_));
  NAND3_X1   g03939(.A1(new_n4195_), .A2(new_n334_), .A3(new_n3738_), .ZN(new_n4196_));
  XOR2_X1    g03940(.A1(new_n4196_), .A2(\a[41] ), .Z(new_n4197_));
  INV_X1     g03941(.I(\a[44] ), .ZN(new_n4198_));
  INV_X1     g03942(.I(\a[43] ), .ZN(new_n4199_));
  NOR3_X1    g03943(.A1(new_n4199_), .A2(\a[41] ), .A3(\a[42] ), .ZN(new_n4200_));
  NAND3_X1   g03944(.A1(new_n4199_), .A2(\a[41] ), .A3(\a[42] ), .ZN(new_n4201_));
  INV_X1     g03945(.I(new_n4201_), .ZN(new_n4202_));
  NOR2_X1    g03946(.A1(new_n4202_), .A2(new_n4200_), .ZN(new_n4203_));
  NOR2_X1    g03947(.A1(new_n4203_), .A2(new_n258_), .ZN(new_n4204_));
  INV_X1     g03948(.I(new_n4040_), .ZN(new_n4205_));
  XNOR2_X1   g03949(.A1(\a[43] ), .A2(\a[44] ), .ZN(new_n4206_));
  NOR2_X1    g03950(.A1(new_n4205_), .A2(new_n4206_), .ZN(new_n4207_));
  INV_X1     g03951(.I(new_n4207_), .ZN(new_n4208_));
  NOR2_X1    g03952(.A1(new_n4208_), .A2(new_n267_), .ZN(new_n4209_));
  NOR2_X1    g03953(.A1(new_n4040_), .A2(new_n4206_), .ZN(new_n4210_));
  INV_X1     g03954(.I(new_n4210_), .ZN(new_n4211_));
  NOR4_X1    g03955(.A1(new_n4209_), .A2(new_n261_), .A3(new_n4204_), .A4(new_n4211_), .ZN(new_n4212_));
  XOR2_X1    g03956(.A1(new_n4212_), .A2(new_n4198_), .Z(new_n4213_));
  NOR2_X1    g03957(.A1(new_n4041_), .A2(new_n4198_), .ZN(new_n4214_));
  XNOR2_X1   g03958(.A1(new_n4213_), .A2(new_n4214_), .ZN(new_n4215_));
  XOR2_X1    g03959(.A1(new_n4215_), .A2(new_n4197_), .Z(new_n4216_));
  NOR2_X1    g03960(.A1(new_n4193_), .A2(new_n4216_), .ZN(new_n4217_));
  INV_X1     g03961(.I(new_n4193_), .ZN(new_n4218_));
  INV_X1     g03962(.I(new_n4197_), .ZN(new_n4219_));
  NOR2_X1    g03963(.A1(new_n4215_), .A2(new_n4219_), .ZN(new_n4220_));
  INV_X1     g03964(.I(new_n4220_), .ZN(new_n4221_));
  NAND2_X1   g03965(.A1(new_n4215_), .A2(new_n4219_), .ZN(new_n4222_));
  AOI21_X1   g03966(.A1(new_n4221_), .A2(new_n4222_), .B(new_n4218_), .ZN(new_n4223_));
  NOR2_X1    g03967(.A1(new_n4223_), .A2(new_n4217_), .ZN(new_n4224_));
  INV_X1     g03968(.I(new_n4224_), .ZN(new_n4225_));
  OAI22_X1   g03969(.A1(new_n3298_), .A2(new_n450_), .B1(new_n403_), .B2(new_n3293_), .ZN(new_n4226_));
  INV_X1     g03970(.I(new_n3447_), .ZN(new_n4227_));
  NAND2_X1   g03971(.A1(new_n4227_), .A2(\b[5] ), .ZN(new_n4228_));
  AOI21_X1   g03972(.A1(new_n4226_), .A2(new_n4228_), .B(new_n3301_), .ZN(new_n4229_));
  NAND2_X1   g03973(.A1(new_n454_), .A2(new_n4229_), .ZN(new_n4230_));
  XOR2_X1    g03974(.A1(new_n4230_), .A2(\a[38] ), .Z(new_n4231_));
  NOR2_X1    g03975(.A1(new_n4225_), .A2(new_n4231_), .ZN(new_n4232_));
  INV_X1     g03976(.I(new_n4232_), .ZN(new_n4233_));
  NAND2_X1   g03977(.A1(new_n4225_), .A2(new_n4231_), .ZN(new_n4234_));
  NAND2_X1   g03978(.A1(new_n4233_), .A2(new_n4234_), .ZN(new_n4235_));
  OAI22_X1   g03979(.A1(new_n2846_), .A2(new_n617_), .B1(new_n510_), .B2(new_n2841_), .ZN(new_n4236_));
  NAND2_X1   g03980(.A1(new_n3755_), .A2(\b[8] ), .ZN(new_n4237_));
  AOI21_X1   g03981(.A1(new_n4236_), .A2(new_n4237_), .B(new_n2849_), .ZN(new_n4238_));
  NAND2_X1   g03982(.A1(new_n616_), .A2(new_n4238_), .ZN(new_n4239_));
  XOR2_X1    g03983(.A1(new_n4239_), .A2(\a[35] ), .Z(new_n4240_));
  XNOR2_X1   g03984(.A1(new_n4235_), .A2(new_n4240_), .ZN(new_n4241_));
  OAI22_X1   g03985(.A1(new_n2452_), .A2(new_n795_), .B1(new_n717_), .B2(new_n2447_), .ZN(new_n4242_));
  NAND2_X1   g03986(.A1(new_n3312_), .A2(\b[11] ), .ZN(new_n4243_));
  AOI21_X1   g03987(.A1(new_n4242_), .A2(new_n4243_), .B(new_n2455_), .ZN(new_n4244_));
  NAND2_X1   g03988(.A1(new_n799_), .A2(new_n4244_), .ZN(new_n4245_));
  XOR2_X1    g03989(.A1(new_n4245_), .A2(\a[32] ), .Z(new_n4246_));
  XNOR2_X1   g03990(.A1(new_n4241_), .A2(new_n4246_), .ZN(new_n4247_));
  OAI22_X1   g03991(.A1(new_n2084_), .A2(new_n992_), .B1(new_n904_), .B2(new_n2079_), .ZN(new_n4248_));
  NAND2_X1   g03992(.A1(new_n2864_), .A2(\b[14] ), .ZN(new_n4249_));
  AOI21_X1   g03993(.A1(new_n4248_), .A2(new_n4249_), .B(new_n2087_), .ZN(new_n4250_));
  NAND2_X1   g03994(.A1(new_n991_), .A2(new_n4250_), .ZN(new_n4251_));
  XOR2_X1    g03995(.A1(new_n4251_), .A2(\a[29] ), .Z(new_n4252_));
  XNOR2_X1   g03996(.A1(new_n4247_), .A2(new_n4252_), .ZN(new_n4253_));
  OAI22_X1   g03997(.A1(new_n1760_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n1755_), .ZN(new_n4254_));
  NAND2_X1   g03998(.A1(new_n2470_), .A2(\b[17] ), .ZN(new_n4255_));
  AOI21_X1   g03999(.A1(new_n4254_), .A2(new_n4255_), .B(new_n1763_), .ZN(new_n4256_));
  NAND2_X1   g04000(.A1(new_n1225_), .A2(new_n4256_), .ZN(new_n4257_));
  XOR2_X1    g04001(.A1(new_n4257_), .A2(\a[26] ), .Z(new_n4258_));
  XNOR2_X1   g04002(.A1(new_n4253_), .A2(new_n4258_), .ZN(new_n4259_));
  INV_X1     g04003(.I(new_n4259_), .ZN(new_n4260_));
  XOR2_X1    g04004(.A1(new_n4253_), .A2(new_n4258_), .Z(new_n4261_));
  NOR2_X1    g04005(.A1(new_n4189_), .A2(new_n4261_), .ZN(new_n4262_));
  AOI21_X1   g04006(.A1(new_n4189_), .A2(new_n4260_), .B(new_n4262_), .ZN(new_n4263_));
  OAI22_X1   g04007(.A1(new_n1444_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n1439_), .ZN(new_n4264_));
  NAND2_X1   g04008(.A1(new_n2098_), .A2(\b[20] ), .ZN(new_n4265_));
  AOI21_X1   g04009(.A1(new_n4264_), .A2(new_n4265_), .B(new_n1447_), .ZN(new_n4266_));
  NAND2_X1   g04010(.A1(new_n1517_), .A2(new_n4266_), .ZN(new_n4267_));
  XOR2_X1    g04011(.A1(new_n4267_), .A2(\a[23] ), .Z(new_n4268_));
  XOR2_X1    g04012(.A1(new_n4263_), .A2(new_n4268_), .Z(new_n4269_));
  XOR2_X1    g04013(.A1(new_n4263_), .A2(new_n4268_), .Z(new_n4270_));
  NAND2_X1   g04014(.A1(new_n4185_), .A2(new_n4270_), .ZN(new_n4271_));
  OAI21_X1   g04015(.A1(new_n4185_), .A2(new_n4269_), .B(new_n4271_), .ZN(new_n4272_));
  OAI22_X1   g04016(.A1(new_n1168_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n1163_), .ZN(new_n4273_));
  NAND2_X1   g04017(.A1(new_n1774_), .A2(\b[23] ), .ZN(new_n4274_));
  AOI21_X1   g04018(.A1(new_n4273_), .A2(new_n4274_), .B(new_n1171_), .ZN(new_n4275_));
  NAND2_X1   g04019(.A1(new_n1828_), .A2(new_n4275_), .ZN(new_n4276_));
  XOR2_X1    g04020(.A1(new_n4276_), .A2(\a[20] ), .Z(new_n4277_));
  XOR2_X1    g04021(.A1(new_n4272_), .A2(new_n4277_), .Z(new_n4278_));
  INV_X1     g04022(.I(new_n4278_), .ZN(new_n4279_));
  OAI22_X1   g04023(.A1(new_n940_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n935_), .ZN(new_n4280_));
  NAND2_X1   g04024(.A1(new_n1458_), .A2(\b[26] ), .ZN(new_n4281_));
  AOI21_X1   g04025(.A1(new_n4280_), .A2(new_n4281_), .B(new_n943_), .ZN(new_n4282_));
  NAND2_X1   g04026(.A1(new_n2174_), .A2(new_n4282_), .ZN(new_n4283_));
  XOR2_X1    g04027(.A1(new_n4283_), .A2(\a[17] ), .Z(new_n4284_));
  NOR2_X1    g04028(.A1(new_n4279_), .A2(new_n4284_), .ZN(new_n4285_));
  NAND2_X1   g04029(.A1(new_n4279_), .A2(new_n4284_), .ZN(new_n4286_));
  INV_X1     g04030(.I(new_n4286_), .ZN(new_n4287_));
  NOR2_X1    g04031(.A1(new_n4287_), .A2(new_n4285_), .ZN(new_n4288_));
  OAI22_X1   g04032(.A1(new_n757_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n752_), .ZN(new_n4289_));
  NAND2_X1   g04033(.A1(new_n1182_), .A2(\b[29] ), .ZN(new_n4290_));
  AOI21_X1   g04034(.A1(new_n4289_), .A2(new_n4290_), .B(new_n760_), .ZN(new_n4291_));
  NAND2_X1   g04035(.A1(new_n2546_), .A2(new_n4291_), .ZN(new_n4292_));
  XOR2_X1    g04036(.A1(new_n4292_), .A2(\a[14] ), .Z(new_n4293_));
  XOR2_X1    g04037(.A1(new_n4288_), .A2(new_n4293_), .Z(new_n4294_));
  OAI22_X1   g04038(.A1(new_n582_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n577_), .ZN(new_n4295_));
  NAND2_X1   g04039(.A1(new_n960_), .A2(\b[32] ), .ZN(new_n4296_));
  AOI21_X1   g04040(.A1(new_n4295_), .A2(new_n4296_), .B(new_n585_), .ZN(new_n4297_));
  NAND2_X1   g04041(.A1(new_n2963_), .A2(new_n4297_), .ZN(new_n4298_));
  XOR2_X1    g04042(.A1(new_n4298_), .A2(\a[11] ), .Z(new_n4299_));
  INV_X1     g04043(.I(new_n4299_), .ZN(new_n4300_));
  XOR2_X1    g04044(.A1(new_n4294_), .A2(new_n4300_), .Z(new_n4301_));
  AOI21_X1   g04045(.A1(new_n4182_), .A2(new_n4179_), .B(new_n4301_), .ZN(new_n4302_));
  NAND2_X1   g04046(.A1(new_n4182_), .A2(new_n4179_), .ZN(new_n4303_));
  XOR2_X1    g04047(.A1(new_n4294_), .A2(new_n4299_), .Z(new_n4304_));
  NOR2_X1    g04048(.A1(new_n4303_), .A2(new_n4304_), .ZN(new_n4305_));
  NOR2_X1    g04049(.A1(new_n4305_), .A2(new_n4302_), .ZN(new_n4306_));
  XOR2_X1    g04050(.A1(new_n4178_), .A2(new_n4306_), .Z(new_n4307_));
  XOR2_X1    g04051(.A1(new_n4307_), .A2(new_n4174_), .Z(new_n4308_));
  XOR2_X1    g04052(.A1(new_n4308_), .A2(new_n4169_), .Z(new_n4309_));
  XOR2_X1    g04053(.A1(new_n4033_), .A2(new_n4029_), .Z(new_n4310_));
  NAND2_X1   g04054(.A1(new_n4310_), .A2(new_n4159_), .ZN(new_n4311_));
  XOR2_X1    g04055(.A1(new_n4309_), .A2(new_n4311_), .Z(new_n4312_));
  INV_X1     g04056(.I(new_n4033_), .ZN(new_n4313_));
  NOR2_X1    g04057(.A1(new_n4313_), .A2(new_n4028_), .ZN(new_n4314_));
  XOR2_X1    g04058(.A1(new_n4312_), .A2(new_n4314_), .Z(new_n4315_));
  INV_X1     g04059(.I(\b[43] ), .ZN(new_n4316_));
  XOR2_X1    g04060(.A1(new_n4013_), .A2(\b[41] ), .Z(new_n4317_));
  AND3_X2    g04061(.A1(new_n4317_), .A2(new_n4316_), .A3(new_n4014_), .Z(new_n4318_));
  AOI21_X1   g04062(.A1(new_n4317_), .A2(new_n4014_), .B(new_n4316_), .ZN(new_n4319_));
  OR2_X2     g04063(.A1(new_n4318_), .A2(new_n4319_), .Z(new_n4320_));
  OAI22_X1   g04064(.A1(new_n405_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n404_), .ZN(new_n4321_));
  NAND2_X1   g04065(.A1(new_n279_), .A2(\b[41] ), .ZN(new_n4322_));
  AOI21_X1   g04066(.A1(new_n4321_), .A2(new_n4322_), .B(new_n264_), .ZN(new_n4323_));
  NAND2_X1   g04067(.A1(new_n4320_), .A2(new_n4323_), .ZN(new_n4324_));
  XOR2_X1    g04068(.A1(new_n4324_), .A2(new_n271_), .Z(new_n4325_));
  XOR2_X1    g04069(.A1(new_n4315_), .A2(new_n4325_), .Z(new_n4326_));
  XOR2_X1    g04070(.A1(new_n4159_), .A2(new_n4029_), .Z(new_n4327_));
  XOR2_X1    g04071(.A1(new_n4159_), .A2(new_n4029_), .Z(new_n4328_));
  OAI21_X1   g04072(.A1(new_n4328_), .A2(new_n4313_), .B(new_n4023_), .ZN(new_n4329_));
  AOI21_X1   g04073(.A1(new_n4313_), .A2(new_n4327_), .B(new_n4329_), .ZN(new_n4330_));
  NOR2_X1    g04074(.A1(new_n4007_), .A2(new_n3863_), .ZN(new_n4331_));
  NOR4_X1    g04075(.A1(new_n4162_), .A2(new_n4006_), .A3(new_n4330_), .A4(new_n4331_), .ZN(new_n4332_));
  XOR2_X1    g04076(.A1(new_n4326_), .A2(new_n4332_), .Z(\f[43] ));
  INV_X1     g04077(.I(new_n4174_), .ZN(new_n4334_));
  NAND2_X1   g04078(.A1(new_n4306_), .A2(new_n4334_), .ZN(new_n4335_));
  NOR2_X1    g04079(.A1(new_n4306_), .A2(new_n4334_), .ZN(new_n4336_));
  INV_X1     g04080(.I(new_n4336_), .ZN(new_n4337_));
  NAND2_X1   g04081(.A1(new_n4178_), .A2(new_n4337_), .ZN(new_n4338_));
  OAI22_X1   g04082(.A1(new_n1168_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n1163_), .ZN(new_n4339_));
  NAND2_X1   g04083(.A1(new_n1774_), .A2(\b[24] ), .ZN(new_n4340_));
  AOI21_X1   g04084(.A1(new_n4339_), .A2(new_n4340_), .B(new_n1171_), .ZN(new_n4341_));
  NAND2_X1   g04085(.A1(new_n1926_), .A2(new_n4341_), .ZN(new_n4342_));
  XOR2_X1    g04086(.A1(new_n4342_), .A2(\a[20] ), .Z(new_n4343_));
  OAI22_X1   g04087(.A1(new_n1444_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n1439_), .ZN(new_n4344_));
  NAND2_X1   g04088(.A1(new_n2098_), .A2(\b[21] ), .ZN(new_n4345_));
  AOI21_X1   g04089(.A1(new_n4344_), .A2(new_n4345_), .B(new_n1447_), .ZN(new_n4346_));
  NAND2_X1   g04090(.A1(new_n1604_), .A2(new_n4346_), .ZN(new_n4347_));
  XOR2_X1    g04091(.A1(new_n4347_), .A2(\a[23] ), .Z(new_n4348_));
  INV_X1     g04092(.I(new_n4348_), .ZN(new_n4349_));
  XNOR2_X1   g04093(.A1(new_n4184_), .A2(new_n4263_), .ZN(new_n4350_));
  NAND2_X1   g04094(.A1(new_n4350_), .A2(new_n4268_), .ZN(new_n4351_));
  NAND2_X1   g04095(.A1(new_n4351_), .A2(new_n4272_), .ZN(new_n4352_));
  NOR2_X1    g04096(.A1(new_n4235_), .A2(new_n4240_), .ZN(new_n4353_));
  OAI22_X1   g04097(.A1(new_n3736_), .A2(new_n347_), .B1(new_n393_), .B2(new_n3731_), .ZN(new_n4354_));
  OAI21_X1   g04098(.A1(new_n290_), .A2(new_n3889_), .B(new_n4354_), .ZN(new_n4355_));
  AOI21_X1   g04099(.A1(new_n352_), .A2(new_n3738_), .B(new_n4355_), .ZN(new_n4356_));
  NAND2_X1   g04100(.A1(new_n4213_), .A2(new_n4214_), .ZN(new_n4357_));
  NOR2_X1    g04101(.A1(new_n4211_), .A2(new_n278_), .ZN(new_n4358_));
  XNOR2_X1   g04102(.A1(\a[41] ), .A2(\a[43] ), .ZN(new_n4359_));
  NAND2_X1   g04103(.A1(new_n4040_), .A2(new_n4359_), .ZN(new_n4360_));
  XNOR2_X1   g04104(.A1(\a[41] ), .A2(\a[44] ), .ZN(new_n4361_));
  NAND2_X1   g04105(.A1(new_n4360_), .A2(new_n4361_), .ZN(new_n4362_));
  OAI22_X1   g04106(.A1(new_n4208_), .A2(new_n292_), .B1(new_n267_), .B2(new_n4203_), .ZN(new_n4363_));
  NOR4_X1    g04107(.A1(new_n4363_), .A2(new_n258_), .A3(new_n4358_), .A4(new_n4362_), .ZN(new_n4364_));
  XOR2_X1    g04108(.A1(new_n4364_), .A2(new_n4198_), .Z(new_n4365_));
  XNOR2_X1   g04109(.A1(new_n4357_), .A2(new_n4365_), .ZN(new_n4366_));
  XOR2_X1    g04110(.A1(new_n4366_), .A2(\a[41] ), .Z(new_n4367_));
  XOR2_X1    g04111(.A1(new_n4367_), .A2(new_n4356_), .Z(new_n4368_));
  OAI21_X1   g04112(.A1(new_n4218_), .A2(new_n4215_), .B(new_n4219_), .ZN(new_n4369_));
  XNOR2_X1   g04113(.A1(new_n4369_), .A2(new_n4368_), .ZN(new_n4370_));
  OAI22_X1   g04114(.A1(new_n3298_), .A2(new_n495_), .B1(new_n450_), .B2(new_n3293_), .ZN(new_n4371_));
  NAND2_X1   g04115(.A1(new_n4227_), .A2(\b[6] ), .ZN(new_n4372_));
  AOI21_X1   g04116(.A1(new_n4371_), .A2(new_n4372_), .B(new_n3301_), .ZN(new_n4373_));
  NAND2_X1   g04117(.A1(new_n494_), .A2(new_n4373_), .ZN(new_n4374_));
  XOR2_X1    g04118(.A1(new_n4374_), .A2(\a[38] ), .Z(new_n4375_));
  XNOR2_X1   g04119(.A1(new_n4370_), .A2(new_n4375_), .ZN(new_n4376_));
  XOR2_X1    g04120(.A1(new_n4376_), .A2(new_n4232_), .Z(new_n4377_));
  OAI22_X1   g04121(.A1(new_n2846_), .A2(new_n659_), .B1(new_n617_), .B2(new_n2841_), .ZN(new_n4378_));
  NAND2_X1   g04122(.A1(new_n3755_), .A2(\b[9] ), .ZN(new_n4379_));
  AOI21_X1   g04123(.A1(new_n4378_), .A2(new_n4379_), .B(new_n2849_), .ZN(new_n4380_));
  NAND2_X1   g04124(.A1(new_n663_), .A2(new_n4380_), .ZN(new_n4381_));
  XOR2_X1    g04125(.A1(new_n4381_), .A2(\a[35] ), .Z(new_n4382_));
  XNOR2_X1   g04126(.A1(new_n4377_), .A2(new_n4382_), .ZN(new_n4383_));
  OAI22_X1   g04127(.A1(new_n2452_), .A2(new_n848_), .B1(new_n795_), .B2(new_n2447_), .ZN(new_n4384_));
  NAND2_X1   g04128(.A1(new_n3312_), .A2(\b[12] ), .ZN(new_n4385_));
  AOI21_X1   g04129(.A1(new_n4384_), .A2(new_n4385_), .B(new_n2455_), .ZN(new_n4386_));
  NAND2_X1   g04130(.A1(new_n847_), .A2(new_n4386_), .ZN(new_n4387_));
  XOR2_X1    g04131(.A1(new_n4387_), .A2(\a[32] ), .Z(new_n4388_));
  XNOR2_X1   g04132(.A1(new_n4383_), .A2(new_n4388_), .ZN(new_n4389_));
  XOR2_X1    g04133(.A1(new_n4383_), .A2(new_n4388_), .Z(new_n4390_));
  MUX2_X1    g04134(.I0(new_n4390_), .I1(new_n4389_), .S(new_n4353_), .Z(new_n4391_));
  NOR2_X1    g04135(.A1(new_n4241_), .A2(new_n4246_), .ZN(new_n4392_));
  XOR2_X1    g04136(.A1(new_n4391_), .A2(new_n4392_), .Z(new_n4393_));
  OAI22_X1   g04137(.A1(new_n2084_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n2079_), .ZN(new_n4394_));
  NAND2_X1   g04138(.A1(new_n2864_), .A2(\b[15] ), .ZN(new_n4395_));
  AOI21_X1   g04139(.A1(new_n4394_), .A2(new_n4395_), .B(new_n2087_), .ZN(new_n4396_));
  NAND2_X1   g04140(.A1(new_n1047_), .A2(new_n4396_), .ZN(new_n4397_));
  XOR2_X1    g04141(.A1(new_n4397_), .A2(\a[29] ), .Z(new_n4398_));
  XOR2_X1    g04142(.A1(new_n4393_), .A2(new_n4398_), .Z(new_n4399_));
  NAND2_X1   g04143(.A1(new_n4247_), .A2(new_n4252_), .ZN(new_n4400_));
  OAI21_X1   g04144(.A1(new_n4189_), .A2(new_n4253_), .B(new_n4400_), .ZN(new_n4401_));
  XOR2_X1    g04145(.A1(new_n4399_), .A2(new_n4401_), .Z(new_n4402_));
  INV_X1     g04146(.I(new_n4402_), .ZN(new_n4403_));
  OAI22_X1   g04147(.A1(new_n1760_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n1755_), .ZN(new_n4404_));
  NAND2_X1   g04148(.A1(new_n2470_), .A2(\b[18] ), .ZN(new_n4405_));
  AOI21_X1   g04149(.A1(new_n4404_), .A2(new_n4405_), .B(new_n1763_), .ZN(new_n4406_));
  NAND2_X1   g04150(.A1(new_n1304_), .A2(new_n4406_), .ZN(new_n4407_));
  XOR2_X1    g04151(.A1(new_n4407_), .A2(\a[26] ), .Z(new_n4408_));
  NOR2_X1    g04152(.A1(new_n4403_), .A2(new_n4408_), .ZN(new_n4409_));
  NAND2_X1   g04153(.A1(new_n4403_), .A2(new_n4408_), .ZN(new_n4410_));
  INV_X1     g04154(.I(new_n4410_), .ZN(new_n4411_));
  NOR2_X1    g04155(.A1(new_n4411_), .A2(new_n4409_), .ZN(new_n4412_));
  INV_X1     g04156(.I(new_n4412_), .ZN(new_n4413_));
  XOR2_X1    g04157(.A1(new_n4189_), .A2(new_n4253_), .Z(new_n4414_));
  NAND2_X1   g04158(.A1(new_n4414_), .A2(new_n4258_), .ZN(new_n4415_));
  NAND2_X1   g04159(.A1(new_n4185_), .A2(new_n4263_), .ZN(new_n4416_));
  NAND2_X1   g04160(.A1(new_n4416_), .A2(new_n4415_), .ZN(new_n4417_));
  NOR2_X1    g04161(.A1(new_n4413_), .A2(new_n4417_), .ZN(new_n4418_));
  NAND2_X1   g04162(.A1(new_n4413_), .A2(new_n4417_), .ZN(new_n4419_));
  INV_X1     g04163(.I(new_n4419_), .ZN(new_n4420_));
  NOR2_X1    g04164(.A1(new_n4420_), .A2(new_n4418_), .ZN(new_n4421_));
  XOR2_X1    g04165(.A1(new_n4421_), .A2(new_n4352_), .Z(new_n4422_));
  XOR2_X1    g04166(.A1(new_n4422_), .A2(new_n4349_), .Z(new_n4423_));
  XOR2_X1    g04167(.A1(new_n4423_), .A2(new_n4343_), .Z(new_n4424_));
  NOR2_X1    g04168(.A1(new_n4272_), .A2(new_n4277_), .ZN(new_n4425_));
  XOR2_X1    g04169(.A1(new_n4424_), .A2(new_n4425_), .Z(new_n4426_));
  OAI22_X1   g04170(.A1(new_n940_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n935_), .ZN(new_n4427_));
  NAND2_X1   g04171(.A1(new_n1458_), .A2(\b[27] ), .ZN(new_n4428_));
  AOI21_X1   g04172(.A1(new_n4427_), .A2(new_n4428_), .B(new_n943_), .ZN(new_n4429_));
  NAND2_X1   g04173(.A1(new_n2276_), .A2(new_n4429_), .ZN(new_n4430_));
  XOR2_X1    g04174(.A1(new_n4430_), .A2(\a[17] ), .Z(new_n4431_));
  XOR2_X1    g04175(.A1(new_n4426_), .A2(new_n4431_), .Z(new_n4432_));
  INV_X1     g04176(.I(new_n4432_), .ZN(new_n4433_));
  NOR2_X1    g04177(.A1(new_n4279_), .A2(new_n4284_), .ZN(new_n4434_));
  INV_X1     g04178(.I(new_n4434_), .ZN(new_n4435_));
  NOR2_X1    g04179(.A1(new_n4433_), .A2(new_n4435_), .ZN(new_n4436_));
  INV_X1     g04180(.I(new_n4436_), .ZN(new_n4437_));
  NAND2_X1   g04181(.A1(new_n4433_), .A2(new_n4435_), .ZN(new_n4438_));
  NAND2_X1   g04182(.A1(new_n4437_), .A2(new_n4438_), .ZN(new_n4439_));
  OAI22_X1   g04183(.A1(new_n757_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n752_), .ZN(new_n4440_));
  NAND2_X1   g04184(.A1(new_n1182_), .A2(\b[30] ), .ZN(new_n4441_));
  AOI21_X1   g04185(.A1(new_n4440_), .A2(new_n4441_), .B(new_n760_), .ZN(new_n4442_));
  NAND2_X1   g04186(.A1(new_n2659_), .A2(new_n4442_), .ZN(new_n4443_));
  XOR2_X1    g04187(.A1(new_n4443_), .A2(\a[14] ), .Z(new_n4444_));
  XNOR2_X1   g04188(.A1(new_n4439_), .A2(new_n4444_), .ZN(new_n4445_));
  NAND2_X1   g04189(.A1(new_n4303_), .A2(new_n4288_), .ZN(new_n4446_));
  XOR2_X1    g04190(.A1(new_n4446_), .A2(new_n4445_), .Z(new_n4447_));
  INV_X1     g04191(.I(new_n4293_), .ZN(new_n4448_));
  XOR2_X1    g04192(.A1(new_n4303_), .A2(new_n4288_), .Z(new_n4449_));
  NAND2_X1   g04193(.A1(new_n4449_), .A2(new_n4448_), .ZN(new_n4450_));
  XOR2_X1    g04194(.A1(new_n4447_), .A2(new_n4450_), .Z(new_n4451_));
  OAI22_X1   g04195(.A1(new_n582_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n577_), .ZN(new_n4452_));
  NAND2_X1   g04196(.A1(new_n960_), .A2(\b[33] ), .ZN(new_n4453_));
  AOI21_X1   g04197(.A1(new_n4452_), .A2(new_n4453_), .B(new_n585_), .ZN(new_n4454_));
  NAND2_X1   g04198(.A1(new_n3101_), .A2(new_n4454_), .ZN(new_n4455_));
  XOR2_X1    g04199(.A1(new_n4455_), .A2(\a[11] ), .Z(new_n4456_));
  XOR2_X1    g04200(.A1(new_n4451_), .A2(new_n4456_), .Z(new_n4457_));
  XNOR2_X1   g04201(.A1(new_n4303_), .A2(new_n4294_), .ZN(new_n4458_));
  OAI22_X1   g04202(.A1(new_n4458_), .A2(new_n4300_), .B1(new_n4302_), .B2(new_n4305_), .ZN(new_n4459_));
  XOR2_X1    g04203(.A1(new_n4457_), .A2(new_n4459_), .Z(new_n4460_));
  OAI22_X1   g04204(.A1(new_n437_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n431_), .ZN(new_n4461_));
  NAND2_X1   g04205(.A1(new_n775_), .A2(\b[36] ), .ZN(new_n4462_));
  AOI21_X1   g04206(.A1(new_n4461_), .A2(new_n4462_), .B(new_n440_), .ZN(new_n4463_));
  NAND2_X1   g04207(.A1(new_n3565_), .A2(new_n4463_), .ZN(new_n4464_));
  XOR2_X1    g04208(.A1(new_n4464_), .A2(\a[8] ), .Z(new_n4465_));
  INV_X1     g04209(.I(new_n4465_), .ZN(new_n4466_));
  AND2_X2    g04210(.A1(new_n4460_), .A2(new_n4466_), .Z(new_n4467_));
  NOR2_X1    g04211(.A1(new_n4460_), .A2(new_n4466_), .ZN(new_n4468_));
  NOR2_X1    g04212(.A1(new_n4467_), .A2(new_n4468_), .ZN(new_n4469_));
  OAI22_X1   g04213(.A1(new_n364_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n320_), .ZN(new_n4470_));
  NAND2_X1   g04214(.A1(new_n594_), .A2(\b[39] ), .ZN(new_n4471_));
  AOI21_X1   g04215(.A1(new_n4470_), .A2(new_n4471_), .B(new_n312_), .ZN(new_n4472_));
  NAND2_X1   g04216(.A1(new_n3996_), .A2(new_n4472_), .ZN(new_n4473_));
  XOR2_X1    g04217(.A1(new_n4473_), .A2(\a[5] ), .Z(new_n4474_));
  XOR2_X1    g04218(.A1(new_n4469_), .A2(new_n4474_), .Z(new_n4475_));
  AOI21_X1   g04219(.A1(new_n4335_), .A2(new_n4338_), .B(new_n4475_), .ZN(new_n4476_));
  NAND2_X1   g04220(.A1(new_n4338_), .A2(new_n4335_), .ZN(new_n4477_));
  XNOR2_X1   g04221(.A1(new_n4469_), .A2(new_n4474_), .ZN(new_n4478_));
  NOR2_X1    g04222(.A1(new_n4477_), .A2(new_n4478_), .ZN(new_n4479_));
  NOR2_X1    g04223(.A1(new_n4479_), .A2(new_n4476_), .ZN(new_n4480_));
  NAND2_X1   g04224(.A1(new_n4309_), .A2(new_n4314_), .ZN(new_n4481_));
  NAND3_X1   g04225(.A1(new_n4481_), .A2(new_n4159_), .A3(new_n4310_), .ZN(new_n4482_));
  NAND2_X1   g04226(.A1(new_n4337_), .A2(new_n4335_), .ZN(new_n4483_));
  XOR2_X1    g04227(.A1(new_n4178_), .A2(new_n4483_), .Z(new_n4484_));
  NAND2_X1   g04228(.A1(new_n4484_), .A2(new_n4169_), .ZN(new_n4485_));
  NAND2_X1   g04229(.A1(new_n4482_), .A2(new_n4485_), .ZN(new_n4486_));
  NAND2_X1   g04230(.A1(new_n4486_), .A2(new_n4480_), .ZN(new_n4487_));
  INV_X1     g04231(.I(new_n4480_), .ZN(new_n4488_));
  NAND3_X1   g04232(.A1(new_n4482_), .A2(new_n4488_), .A3(new_n4485_), .ZN(new_n4489_));
  NAND2_X1   g04233(.A1(new_n4487_), .A2(new_n4489_), .ZN(new_n4490_));
  OAI21_X1   g04234(.A1(new_n3997_), .A2(new_n4316_), .B(new_n4018_), .ZN(new_n4491_));
  NAND3_X1   g04235(.A1(new_n4011_), .A2(new_n4012_), .A3(new_n4491_), .ZN(new_n4492_));
  OAI21_X1   g04236(.A1(\b[41] ), .A2(\b[43] ), .B(\b[42] ), .ZN(new_n4493_));
  NAND2_X1   g04237(.A1(new_n4492_), .A2(new_n4493_), .ZN(new_n4494_));
  INV_X1     g04238(.I(new_n4494_), .ZN(new_n4495_));
  XNOR2_X1   g04239(.A1(\b[43] ), .A2(\b[44] ), .ZN(new_n4496_));
  NOR2_X1    g04240(.A1(new_n4495_), .A2(new_n4496_), .ZN(new_n4497_));
  XNOR2_X1   g04241(.A1(\b[43] ), .A2(\b[44] ), .ZN(new_n4498_));
  AOI21_X1   g04242(.A1(new_n4495_), .A2(new_n4498_), .B(new_n4497_), .ZN(new_n4499_));
  INV_X1     g04243(.I(new_n4499_), .ZN(new_n4500_));
  INV_X1     g04244(.I(\b[44] ), .ZN(new_n4501_));
  OAI22_X1   g04245(.A1(new_n405_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n404_), .ZN(new_n4502_));
  NAND2_X1   g04246(.A1(new_n279_), .A2(\b[42] ), .ZN(new_n4503_));
  AOI21_X1   g04247(.A1(new_n4502_), .A2(new_n4503_), .B(new_n264_), .ZN(new_n4504_));
  NAND2_X1   g04248(.A1(new_n4500_), .A2(new_n4504_), .ZN(new_n4505_));
  XOR2_X1    g04249(.A1(new_n4505_), .A2(\a[2] ), .Z(new_n4506_));
  XOR2_X1    g04250(.A1(new_n4490_), .A2(new_n4506_), .Z(\f[44] ));
  AOI21_X1   g04251(.A1(new_n4487_), .A2(new_n4489_), .B(new_n4506_), .ZN(new_n4508_));
  INV_X1     g04252(.I(\b[45] ), .ZN(new_n4509_));
  INV_X1     g04253(.I(new_n4496_), .ZN(new_n4510_));
  XOR2_X1    g04254(.A1(new_n4494_), .A2(\b[43] ), .Z(new_n4511_));
  NAND2_X1   g04255(.A1(new_n4511_), .A2(new_n4510_), .ZN(new_n4512_));
  XOR2_X1    g04256(.A1(new_n4512_), .A2(new_n4509_), .Z(new_n4513_));
  NOR2_X1    g04257(.A1(new_n405_), .A2(new_n4509_), .ZN(new_n4514_));
  NOR2_X1    g04258(.A1(new_n280_), .A2(new_n4316_), .ZN(new_n4515_));
  NOR2_X1    g04259(.A1(new_n404_), .A2(new_n4501_), .ZN(new_n4516_));
  NOR4_X1    g04260(.A1(new_n4514_), .A2(new_n264_), .A3(new_n4515_), .A4(new_n4516_), .ZN(new_n4517_));
  NAND2_X1   g04261(.A1(new_n4513_), .A2(new_n4517_), .ZN(new_n4518_));
  INV_X1     g04262(.I(new_n4357_), .ZN(new_n4519_));
  NAND2_X1   g04263(.A1(new_n4519_), .A2(new_n4365_), .ZN(new_n4520_));
  NOR2_X1    g04264(.A1(new_n4362_), .A2(new_n267_), .ZN(new_n4521_));
  OAI22_X1   g04265(.A1(new_n4208_), .A2(new_n290_), .B1(new_n292_), .B2(new_n4203_), .ZN(new_n4522_));
  NOR4_X1    g04266(.A1(new_n4522_), .A2(new_n677_), .A3(new_n4211_), .A4(new_n4521_), .ZN(new_n4523_));
  XOR2_X1    g04267(.A1(new_n4523_), .A2(new_n4198_), .Z(new_n4524_));
  XNOR2_X1   g04268(.A1(\a[44] ), .A2(\a[45] ), .ZN(new_n4525_));
  NOR2_X1    g04269(.A1(new_n4525_), .A2(new_n258_), .ZN(new_n4526_));
  XOR2_X1    g04270(.A1(new_n4524_), .A2(new_n4526_), .Z(new_n4527_));
  XNOR2_X1   g04271(.A1(new_n4527_), .A2(new_n4520_), .ZN(new_n4528_));
  INV_X1     g04272(.I(new_n3731_), .ZN(new_n4529_));
  AOI22_X1   g04273(.A1(\b[6] ), .A2(new_n3735_), .B1(new_n4529_), .B2(\b[5] ), .ZN(new_n4530_));
  NOR2_X1    g04274(.A1(new_n3889_), .A2(new_n393_), .ZN(new_n4531_));
  OAI21_X1   g04275(.A1(new_n4530_), .A2(new_n4531_), .B(new_n3738_), .ZN(new_n4532_));
  NOR2_X1    g04276(.A1(new_n524_), .A2(new_n4532_), .ZN(new_n4533_));
  XOR2_X1    g04277(.A1(new_n4533_), .A2(new_n3726_), .Z(new_n4534_));
  NAND2_X1   g04278(.A1(new_n4193_), .A2(new_n4220_), .ZN(new_n4535_));
  NAND2_X1   g04279(.A1(new_n4356_), .A2(new_n3726_), .ZN(new_n4536_));
  NOR2_X1    g04280(.A1(new_n4356_), .A2(new_n3726_), .ZN(new_n4537_));
  NAND2_X1   g04281(.A1(new_n4221_), .A2(new_n4366_), .ZN(new_n4538_));
  NOR2_X1    g04282(.A1(new_n4538_), .A2(new_n4537_), .ZN(new_n4539_));
  NAND4_X1   g04283(.A1(new_n4368_), .A2(new_n4535_), .A3(new_n4536_), .A4(new_n4539_), .ZN(new_n4540_));
  XOR2_X1    g04284(.A1(new_n4540_), .A2(new_n4534_), .Z(new_n4541_));
  XNOR2_X1   g04285(.A1(new_n4541_), .A2(new_n4528_), .ZN(new_n4542_));
  OAI22_X1   g04286(.A1(new_n3298_), .A2(new_n510_), .B1(new_n495_), .B2(new_n3293_), .ZN(new_n4543_));
  NAND2_X1   g04287(.A1(new_n4227_), .A2(\b[7] ), .ZN(new_n4544_));
  AOI21_X1   g04288(.A1(new_n4543_), .A2(new_n4544_), .B(new_n3301_), .ZN(new_n4545_));
  NAND2_X1   g04289(.A1(new_n518_), .A2(new_n4545_), .ZN(new_n4546_));
  XOR2_X1    g04290(.A1(new_n4546_), .A2(\a[38] ), .Z(new_n4547_));
  INV_X1     g04291(.I(new_n4370_), .ZN(new_n4548_));
  NAND2_X1   g04292(.A1(new_n4548_), .A2(new_n4375_), .ZN(new_n4549_));
  NAND3_X1   g04293(.A1(new_n4376_), .A2(new_n4234_), .A3(new_n4549_), .ZN(new_n4550_));
  XOR2_X1    g04294(.A1(new_n4550_), .A2(new_n4547_), .Z(new_n4551_));
  XNOR2_X1   g04295(.A1(new_n4551_), .A2(new_n4542_), .ZN(new_n4552_));
  OAI22_X1   g04296(.A1(new_n2846_), .A2(new_n717_), .B1(new_n659_), .B2(new_n2841_), .ZN(new_n4553_));
  NAND2_X1   g04297(.A1(new_n3755_), .A2(\b[10] ), .ZN(new_n4554_));
  AOI21_X1   g04298(.A1(new_n4553_), .A2(new_n4554_), .B(new_n2849_), .ZN(new_n4555_));
  NAND2_X1   g04299(.A1(new_n716_), .A2(new_n4555_), .ZN(new_n4556_));
  XOR2_X1    g04300(.A1(new_n4556_), .A2(new_n2836_), .Z(new_n4557_));
  AOI21_X1   g04301(.A1(new_n4377_), .A2(new_n4382_), .B(new_n4353_), .ZN(new_n4558_));
  XOR2_X1    g04302(.A1(new_n4558_), .A2(new_n4557_), .Z(new_n4559_));
  XNOR2_X1   g04303(.A1(new_n4552_), .A2(new_n4559_), .ZN(new_n4560_));
  OAI22_X1   g04304(.A1(new_n2452_), .A2(new_n904_), .B1(new_n848_), .B2(new_n2447_), .ZN(new_n4561_));
  NAND2_X1   g04305(.A1(new_n3312_), .A2(\b[13] ), .ZN(new_n4562_));
  AOI21_X1   g04306(.A1(new_n4561_), .A2(new_n4562_), .B(new_n2455_), .ZN(new_n4563_));
  NAND2_X1   g04307(.A1(new_n907_), .A2(new_n4563_), .ZN(new_n4564_));
  XOR2_X1    g04308(.A1(new_n4564_), .A2(\a[32] ), .Z(new_n4565_));
  XOR2_X1    g04309(.A1(new_n4383_), .A2(new_n4353_), .Z(new_n4566_));
  NAND2_X1   g04310(.A1(new_n4566_), .A2(new_n4388_), .ZN(new_n4567_));
  XOR2_X1    g04311(.A1(new_n4567_), .A2(new_n4565_), .Z(new_n4568_));
  XOR2_X1    g04312(.A1(new_n4568_), .A2(new_n4560_), .Z(new_n4569_));
  INV_X1     g04313(.I(new_n4569_), .ZN(new_n4570_));
  OAI22_X1   g04314(.A1(new_n2084_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n2079_), .ZN(new_n4571_));
  NAND2_X1   g04315(.A1(new_n2864_), .A2(\b[16] ), .ZN(new_n4572_));
  AOI21_X1   g04316(.A1(new_n4571_), .A2(new_n4572_), .B(new_n2087_), .ZN(new_n4573_));
  NAND2_X1   g04317(.A1(new_n1123_), .A2(new_n4573_), .ZN(new_n4574_));
  XOR2_X1    g04318(.A1(new_n4574_), .A2(\a[29] ), .Z(new_n4575_));
  OR2_X2     g04319(.A1(new_n4399_), .A2(new_n4401_), .Z(new_n4576_));
  NAND2_X1   g04320(.A1(new_n4393_), .A2(new_n4398_), .ZN(new_n4577_));
  NAND2_X1   g04321(.A1(new_n4576_), .A2(new_n4577_), .ZN(new_n4578_));
  XOR2_X1    g04322(.A1(new_n4578_), .A2(new_n4575_), .Z(new_n4579_));
  XOR2_X1    g04323(.A1(new_n4579_), .A2(new_n4570_), .Z(new_n4580_));
  OAI22_X1   g04324(.A1(new_n1760_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n1755_), .ZN(new_n4581_));
  NAND2_X1   g04325(.A1(new_n2470_), .A2(\b[19] ), .ZN(new_n4582_));
  AOI21_X1   g04326(.A1(new_n4581_), .A2(new_n4582_), .B(new_n1763_), .ZN(new_n4583_));
  NAND2_X1   g04327(.A1(new_n1396_), .A2(new_n4583_), .ZN(new_n4584_));
  XOR2_X1    g04328(.A1(new_n4584_), .A2(\a[26] ), .Z(new_n4585_));
  NAND3_X1   g04329(.A1(new_n4412_), .A2(new_n4410_), .A3(new_n4417_), .ZN(new_n4586_));
  XOR2_X1    g04330(.A1(new_n4586_), .A2(new_n4585_), .Z(new_n4587_));
  XNOR2_X1   g04331(.A1(new_n4587_), .A2(new_n4580_), .ZN(new_n4588_));
  OAI22_X1   g04332(.A1(new_n1444_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n1439_), .ZN(new_n4589_));
  NAND2_X1   g04333(.A1(new_n2098_), .A2(\b[22] ), .ZN(new_n4590_));
  AOI21_X1   g04334(.A1(new_n4589_), .A2(new_n4590_), .B(new_n1447_), .ZN(new_n4591_));
  NAND2_X1   g04335(.A1(new_n1708_), .A2(new_n4591_), .ZN(new_n4592_));
  XOR2_X1    g04336(.A1(new_n4592_), .A2(new_n1434_), .Z(new_n4593_));
  NAND2_X1   g04337(.A1(new_n4421_), .A2(new_n4348_), .ZN(new_n4594_));
  NOR2_X1    g04338(.A1(new_n4421_), .A2(new_n4348_), .ZN(new_n4595_));
  NOR2_X1    g04339(.A1(new_n4595_), .A2(new_n4352_), .ZN(new_n4596_));
  NOR2_X1    g04340(.A1(new_n4421_), .A2(new_n4349_), .ZN(new_n4597_));
  AOI21_X1   g04341(.A1(new_n4596_), .A2(new_n4594_), .B(new_n4597_), .ZN(new_n4598_));
  XOR2_X1    g04342(.A1(new_n4598_), .A2(new_n4593_), .Z(new_n4599_));
  XNOR2_X1   g04343(.A1(new_n4599_), .A2(new_n4588_), .ZN(new_n4600_));
  OAI22_X1   g04344(.A1(new_n1168_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n1163_), .ZN(new_n4601_));
  NAND2_X1   g04345(.A1(new_n1774_), .A2(\b[25] ), .ZN(new_n4602_));
  AOI21_X1   g04346(.A1(new_n4601_), .A2(new_n4602_), .B(new_n1171_), .ZN(new_n4603_));
  NAND2_X1   g04347(.A1(new_n2042_), .A2(new_n4603_), .ZN(new_n4604_));
  XOR2_X1    g04348(.A1(new_n4604_), .A2(new_n1158_), .Z(new_n4605_));
  XOR2_X1    g04349(.A1(new_n4421_), .A2(new_n4349_), .Z(new_n4606_));
  XOR2_X1    g04350(.A1(new_n4606_), .A2(new_n4352_), .Z(new_n4607_));
  AOI22_X1   g04351(.A1(new_n4424_), .A2(new_n4425_), .B1(new_n4343_), .B2(new_n4607_), .ZN(new_n4608_));
  XOR2_X1    g04352(.A1(new_n4608_), .A2(new_n4605_), .Z(new_n4609_));
  XNOR2_X1   g04353(.A1(new_n4609_), .A2(new_n4600_), .ZN(new_n4610_));
  INV_X1     g04354(.I(new_n4610_), .ZN(new_n4611_));
  OAI22_X1   g04355(.A1(new_n940_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n935_), .ZN(new_n4612_));
  NAND2_X1   g04356(.A1(new_n1458_), .A2(\b[28] ), .ZN(new_n4613_));
  AOI21_X1   g04357(.A1(new_n4612_), .A2(new_n4613_), .B(new_n943_), .ZN(new_n4614_));
  NAND2_X1   g04358(.A1(new_n2404_), .A2(new_n4614_), .ZN(new_n4615_));
  XOR2_X1    g04359(.A1(new_n4615_), .A2(\a[17] ), .Z(new_n4616_));
  INV_X1     g04360(.I(new_n4431_), .ZN(new_n4617_));
  OAI21_X1   g04361(.A1(new_n4426_), .A2(new_n4617_), .B(new_n4437_), .ZN(new_n4618_));
  XOR2_X1    g04362(.A1(new_n4618_), .A2(new_n4616_), .Z(new_n4619_));
  XOR2_X1    g04363(.A1(new_n4619_), .A2(new_n4611_), .Z(new_n4620_));
  OAI22_X1   g04364(.A1(new_n757_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n752_), .ZN(new_n4621_));
  NAND2_X1   g04365(.A1(new_n1182_), .A2(\b[31] ), .ZN(new_n4622_));
  AOI21_X1   g04366(.A1(new_n4621_), .A2(new_n4622_), .B(new_n760_), .ZN(new_n4623_));
  NAND2_X1   g04367(.A1(new_n2797_), .A2(new_n4623_), .ZN(new_n4624_));
  XOR2_X1    g04368(.A1(new_n4624_), .A2(\a[14] ), .Z(new_n4625_));
  NAND2_X1   g04369(.A1(new_n4445_), .A2(new_n4448_), .ZN(new_n4626_));
  NAND3_X1   g04370(.A1(new_n4303_), .A2(new_n4288_), .A3(new_n4626_), .ZN(new_n4627_));
  NAND2_X1   g04371(.A1(new_n4439_), .A2(new_n4444_), .ZN(new_n4628_));
  NAND2_X1   g04372(.A1(new_n4627_), .A2(new_n4628_), .ZN(new_n4629_));
  XOR2_X1    g04373(.A1(new_n4629_), .A2(new_n4625_), .Z(new_n4630_));
  XNOR2_X1   g04374(.A1(new_n4630_), .A2(new_n4620_), .ZN(new_n4631_));
  OAI22_X1   g04375(.A1(new_n582_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n577_), .ZN(new_n4632_));
  NAND2_X1   g04376(.A1(new_n960_), .A2(\b[34] ), .ZN(new_n4633_));
  AOI21_X1   g04377(.A1(new_n4632_), .A2(new_n4633_), .B(new_n585_), .ZN(new_n4634_));
  NAND2_X1   g04378(.A1(new_n3246_), .A2(new_n4634_), .ZN(new_n4635_));
  XOR2_X1    g04379(.A1(new_n4635_), .A2(\a[11] ), .Z(new_n4636_));
  INV_X1     g04380(.I(new_n4456_), .ZN(new_n4637_));
  NOR2_X1    g04381(.A1(new_n4451_), .A2(new_n4637_), .ZN(new_n4638_));
  INV_X1     g04382(.I(new_n4459_), .ZN(new_n4639_));
  NOR3_X1    g04383(.A1(new_n4457_), .A2(new_n4638_), .A3(new_n4639_), .ZN(new_n4640_));
  XOR2_X1    g04384(.A1(new_n4640_), .A2(new_n4636_), .Z(new_n4641_));
  XOR2_X1    g04385(.A1(new_n4641_), .A2(new_n4631_), .Z(new_n4642_));
  OAI22_X1   g04386(.A1(new_n437_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n431_), .ZN(new_n4643_));
  NAND2_X1   g04387(.A1(new_n775_), .A2(\b[37] ), .ZN(new_n4644_));
  AOI21_X1   g04388(.A1(new_n4643_), .A2(new_n4644_), .B(new_n440_), .ZN(new_n4645_));
  NAND2_X1   g04389(.A1(new_n3700_), .A2(new_n4645_), .ZN(new_n4646_));
  XOR2_X1    g04390(.A1(new_n4646_), .A2(new_n429_), .Z(new_n4647_));
  NOR2_X1    g04391(.A1(new_n4178_), .A2(new_n4337_), .ZN(new_n4648_));
  NOR4_X1    g04392(.A1(new_n4648_), .A2(new_n4336_), .A3(new_n4467_), .A4(new_n4468_), .ZN(new_n4649_));
  XOR2_X1    g04393(.A1(new_n4649_), .A2(new_n4647_), .Z(new_n4650_));
  XNOR2_X1   g04394(.A1(new_n4650_), .A2(new_n4642_), .ZN(new_n4651_));
  OAI22_X1   g04395(.A1(new_n364_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n320_), .ZN(new_n4652_));
  NAND2_X1   g04396(.A1(new_n594_), .A2(\b[40] ), .ZN(new_n4653_));
  AOI21_X1   g04397(.A1(new_n4652_), .A2(new_n4653_), .B(new_n312_), .ZN(new_n4654_));
  NAND2_X1   g04398(.A1(new_n4017_), .A2(new_n4654_), .ZN(new_n4655_));
  XOR2_X1    g04399(.A1(new_n4655_), .A2(\a[5] ), .Z(new_n4656_));
  INV_X1     g04400(.I(new_n4656_), .ZN(new_n4657_));
  XOR2_X1    g04401(.A1(new_n4651_), .A2(new_n4657_), .Z(new_n4658_));
  XNOR2_X1   g04402(.A1(new_n4477_), .A2(new_n4469_), .ZN(new_n4659_));
  NAND2_X1   g04403(.A1(new_n4659_), .A2(new_n4474_), .ZN(new_n4660_));
  NAND2_X1   g04404(.A1(new_n4487_), .A2(new_n4660_), .ZN(new_n4661_));
  XOR2_X1    g04405(.A1(new_n4661_), .A2(new_n4658_), .Z(new_n4662_));
  XOR2_X1    g04406(.A1(new_n4662_), .A2(\a[2] ), .Z(new_n4663_));
  XOR2_X1    g04407(.A1(new_n4663_), .A2(new_n4518_), .Z(new_n4664_));
  XOR2_X1    g04408(.A1(new_n4664_), .A2(new_n4508_), .Z(\f[45] ));
  OAI22_X1   g04409(.A1(new_n364_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n320_), .ZN(new_n4666_));
  NAND2_X1   g04410(.A1(new_n594_), .A2(\b[41] ), .ZN(new_n4667_));
  AOI21_X1   g04411(.A1(new_n4666_), .A2(new_n4667_), .B(new_n312_), .ZN(new_n4668_));
  NAND2_X1   g04412(.A1(new_n4320_), .A2(new_n4668_), .ZN(new_n4669_));
  XOR2_X1    g04413(.A1(new_n4669_), .A2(\a[5] ), .Z(new_n4670_));
  INV_X1     g04414(.I(new_n4670_), .ZN(new_n4671_));
  OAI22_X1   g04415(.A1(new_n437_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n431_), .ZN(new_n4672_));
  NAND2_X1   g04416(.A1(new_n775_), .A2(\b[38] ), .ZN(new_n4673_));
  AOI21_X1   g04417(.A1(new_n4672_), .A2(new_n4673_), .B(new_n440_), .ZN(new_n4674_));
  NAND2_X1   g04418(.A1(new_n3844_), .A2(new_n4674_), .ZN(new_n4675_));
  XOR2_X1    g04419(.A1(new_n4675_), .A2(\a[8] ), .Z(new_n4676_));
  INV_X1     g04420(.I(new_n4676_), .ZN(new_n4677_));
  XOR2_X1    g04421(.A1(new_n4631_), .A2(new_n4636_), .Z(new_n4678_));
  OAI21_X1   g04422(.A1(new_n4636_), .A2(new_n4640_), .B(new_n4678_), .ZN(new_n4679_));
  NAND2_X1   g04423(.A1(new_n4611_), .A2(new_n4616_), .ZN(new_n4680_));
  INV_X1     g04424(.I(new_n4618_), .ZN(new_n4681_));
  XOR2_X1    g04425(.A1(new_n4610_), .A2(new_n4616_), .Z(new_n4682_));
  NAND2_X1   g04426(.A1(new_n4681_), .A2(new_n4682_), .ZN(new_n4683_));
  NAND2_X1   g04427(.A1(new_n4570_), .A2(new_n4575_), .ZN(new_n4684_));
  XOR2_X1    g04428(.A1(new_n4569_), .A2(new_n4575_), .Z(new_n4685_));
  NAND3_X1   g04429(.A1(new_n4576_), .A2(new_n4577_), .A3(new_n4685_), .ZN(new_n4686_));
  NAND2_X1   g04430(.A1(new_n4686_), .A2(new_n4684_), .ZN(new_n4687_));
  INV_X1     g04431(.I(new_n4687_), .ZN(new_n4688_));
  XOR2_X1    g04432(.A1(new_n4560_), .A2(new_n4565_), .Z(new_n4689_));
  NAND2_X1   g04433(.A1(new_n4689_), .A2(new_n4565_), .ZN(new_n4690_));
  NAND2_X1   g04434(.A1(new_n4689_), .A2(new_n4567_), .ZN(new_n4691_));
  NAND2_X1   g04435(.A1(new_n4691_), .A2(new_n4690_), .ZN(new_n4692_));
  NAND2_X1   g04436(.A1(new_n4527_), .A2(new_n4365_), .ZN(new_n4693_));
  NAND2_X1   g04437(.A1(new_n4693_), .A2(new_n4357_), .ZN(new_n4694_));
  NAND2_X1   g04438(.A1(new_n4524_), .A2(new_n4526_), .ZN(new_n4695_));
  XNOR2_X1   g04439(.A1(new_n4694_), .A2(new_n4695_), .ZN(new_n4696_));
  OAI22_X1   g04440(.A1(new_n4208_), .A2(new_n393_), .B1(new_n290_), .B2(new_n4203_), .ZN(new_n4697_));
  OAI21_X1   g04441(.A1(new_n292_), .A2(new_n4362_), .B(new_n4697_), .ZN(new_n4698_));
  NAND3_X1   g04442(.A1(new_n4698_), .A2(new_n334_), .A3(new_n4210_), .ZN(new_n4699_));
  XOR2_X1    g04443(.A1(new_n4699_), .A2(\a[44] ), .Z(new_n4700_));
  INV_X1     g04444(.I(\a[47] ), .ZN(new_n4701_));
  INV_X1     g04445(.I(\a[46] ), .ZN(new_n4702_));
  NOR3_X1    g04446(.A1(new_n4702_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n4703_));
  NAND3_X1   g04447(.A1(new_n4702_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n4704_));
  INV_X1     g04448(.I(new_n4704_), .ZN(new_n4705_));
  NOR2_X1    g04449(.A1(new_n4705_), .A2(new_n4703_), .ZN(new_n4706_));
  NOR2_X1    g04450(.A1(new_n4706_), .A2(new_n258_), .ZN(new_n4707_));
  INV_X1     g04451(.I(new_n4525_), .ZN(new_n4708_));
  XNOR2_X1   g04452(.A1(\a[46] ), .A2(\a[47] ), .ZN(new_n4709_));
  NOR2_X1    g04453(.A1(new_n4708_), .A2(new_n4709_), .ZN(new_n4710_));
  INV_X1     g04454(.I(new_n4710_), .ZN(new_n4711_));
  NOR2_X1    g04455(.A1(new_n4711_), .A2(new_n267_), .ZN(new_n4712_));
  NOR2_X1    g04456(.A1(new_n4525_), .A2(new_n4709_), .ZN(new_n4713_));
  INV_X1     g04457(.I(new_n4713_), .ZN(new_n4714_));
  NOR4_X1    g04458(.A1(new_n4712_), .A2(new_n261_), .A3(new_n4707_), .A4(new_n4714_), .ZN(new_n4715_));
  XOR2_X1    g04459(.A1(new_n4715_), .A2(new_n4701_), .Z(new_n4716_));
  NOR2_X1    g04460(.A1(new_n4526_), .A2(new_n4701_), .ZN(new_n4717_));
  XNOR2_X1   g04461(.A1(new_n4716_), .A2(new_n4717_), .ZN(new_n4718_));
  XOR2_X1    g04462(.A1(new_n4718_), .A2(new_n4700_), .Z(new_n4719_));
  NOR2_X1    g04463(.A1(new_n4696_), .A2(new_n4719_), .ZN(new_n4720_));
  INV_X1     g04464(.I(new_n4696_), .ZN(new_n4721_));
  INV_X1     g04465(.I(new_n4700_), .ZN(new_n4722_));
  NOR2_X1    g04466(.A1(new_n4718_), .A2(new_n4722_), .ZN(new_n4723_));
  INV_X1     g04467(.I(new_n4723_), .ZN(new_n4724_));
  NAND2_X1   g04468(.A1(new_n4718_), .A2(new_n4722_), .ZN(new_n4725_));
  AOI21_X1   g04469(.A1(new_n4724_), .A2(new_n4725_), .B(new_n4721_), .ZN(new_n4726_));
  NOR2_X1    g04470(.A1(new_n4726_), .A2(new_n4720_), .ZN(new_n4727_));
  INV_X1     g04471(.I(new_n4727_), .ZN(new_n4728_));
  OAI22_X1   g04472(.A1(new_n3736_), .A2(new_n450_), .B1(new_n403_), .B2(new_n3731_), .ZN(new_n4729_));
  INV_X1     g04473(.I(new_n3889_), .ZN(new_n4730_));
  NAND2_X1   g04474(.A1(new_n4730_), .A2(\b[5] ), .ZN(new_n4731_));
  AOI21_X1   g04475(.A1(new_n4729_), .A2(new_n4731_), .B(new_n3739_), .ZN(new_n4732_));
  NAND2_X1   g04476(.A1(new_n454_), .A2(new_n4732_), .ZN(new_n4733_));
  XOR2_X1    g04477(.A1(new_n4733_), .A2(\a[41] ), .Z(new_n4734_));
  NOR2_X1    g04478(.A1(new_n4728_), .A2(new_n4734_), .ZN(new_n4735_));
  INV_X1     g04479(.I(new_n4735_), .ZN(new_n4736_));
  NAND2_X1   g04480(.A1(new_n4728_), .A2(new_n4734_), .ZN(new_n4737_));
  NAND2_X1   g04481(.A1(new_n4736_), .A2(new_n4737_), .ZN(new_n4738_));
  OAI22_X1   g04482(.A1(new_n3298_), .A2(new_n617_), .B1(new_n510_), .B2(new_n3293_), .ZN(new_n4739_));
  NAND2_X1   g04483(.A1(new_n4227_), .A2(\b[8] ), .ZN(new_n4740_));
  AOI21_X1   g04484(.A1(new_n4739_), .A2(new_n4740_), .B(new_n3301_), .ZN(new_n4741_));
  NAND2_X1   g04485(.A1(new_n616_), .A2(new_n4741_), .ZN(new_n4742_));
  XOR2_X1    g04486(.A1(new_n4742_), .A2(\a[38] ), .Z(new_n4743_));
  XNOR2_X1   g04487(.A1(new_n4738_), .A2(new_n4743_), .ZN(new_n4744_));
  OAI22_X1   g04488(.A1(new_n2846_), .A2(new_n795_), .B1(new_n717_), .B2(new_n2841_), .ZN(new_n4745_));
  NAND2_X1   g04489(.A1(new_n3755_), .A2(\b[11] ), .ZN(new_n4746_));
  AOI21_X1   g04490(.A1(new_n4745_), .A2(new_n4746_), .B(new_n2849_), .ZN(new_n4747_));
  NAND2_X1   g04491(.A1(new_n799_), .A2(new_n4747_), .ZN(new_n4748_));
  XOR2_X1    g04492(.A1(new_n4748_), .A2(\a[35] ), .Z(new_n4749_));
  XNOR2_X1   g04493(.A1(new_n4744_), .A2(new_n4749_), .ZN(new_n4750_));
  OAI22_X1   g04494(.A1(new_n2452_), .A2(new_n992_), .B1(new_n904_), .B2(new_n2447_), .ZN(new_n4751_));
  NAND2_X1   g04495(.A1(new_n3312_), .A2(\b[14] ), .ZN(new_n4752_));
  AOI21_X1   g04496(.A1(new_n4751_), .A2(new_n4752_), .B(new_n2455_), .ZN(new_n4753_));
  NAND2_X1   g04497(.A1(new_n991_), .A2(new_n4753_), .ZN(new_n4754_));
  XOR2_X1    g04498(.A1(new_n4754_), .A2(\a[32] ), .Z(new_n4755_));
  XNOR2_X1   g04499(.A1(new_n4750_), .A2(new_n4755_), .ZN(new_n4756_));
  OAI22_X1   g04500(.A1(new_n2084_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n2079_), .ZN(new_n4757_));
  NAND2_X1   g04501(.A1(new_n2864_), .A2(\b[17] ), .ZN(new_n4758_));
  AOI21_X1   g04502(.A1(new_n4757_), .A2(new_n4758_), .B(new_n2087_), .ZN(new_n4759_));
  NAND2_X1   g04503(.A1(new_n1225_), .A2(new_n4759_), .ZN(new_n4760_));
  XOR2_X1    g04504(.A1(new_n4760_), .A2(\a[29] ), .Z(new_n4761_));
  XOR2_X1    g04505(.A1(new_n4756_), .A2(new_n4761_), .Z(new_n4762_));
  XOR2_X1    g04506(.A1(new_n4756_), .A2(new_n4761_), .Z(new_n4763_));
  NOR2_X1    g04507(.A1(new_n4692_), .A2(new_n4763_), .ZN(new_n4764_));
  AOI21_X1   g04508(.A1(new_n4692_), .A2(new_n4762_), .B(new_n4764_), .ZN(new_n4765_));
  OAI22_X1   g04509(.A1(new_n1760_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n1755_), .ZN(new_n4766_));
  NAND2_X1   g04510(.A1(new_n2470_), .A2(\b[20] ), .ZN(new_n4767_));
  AOI21_X1   g04511(.A1(new_n4766_), .A2(new_n4767_), .B(new_n1763_), .ZN(new_n4768_));
  NAND2_X1   g04512(.A1(new_n1517_), .A2(new_n4768_), .ZN(new_n4769_));
  XOR2_X1    g04513(.A1(new_n4769_), .A2(\a[26] ), .Z(new_n4770_));
  XOR2_X1    g04514(.A1(new_n4765_), .A2(new_n4770_), .Z(new_n4771_));
  NOR2_X1    g04515(.A1(new_n4688_), .A2(new_n4771_), .ZN(new_n4772_));
  INV_X1     g04516(.I(new_n4770_), .ZN(new_n4773_));
  XOR2_X1    g04517(.A1(new_n4765_), .A2(new_n4773_), .Z(new_n4774_));
  NOR2_X1    g04518(.A1(new_n4687_), .A2(new_n4774_), .ZN(new_n4775_));
  NOR2_X1    g04519(.A1(new_n4772_), .A2(new_n4775_), .ZN(new_n4776_));
  OAI22_X1   g04520(.A1(new_n1444_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n1439_), .ZN(new_n4777_));
  NAND2_X1   g04521(.A1(new_n2098_), .A2(\b[23] ), .ZN(new_n4778_));
  AOI21_X1   g04522(.A1(new_n4777_), .A2(new_n4778_), .B(new_n1447_), .ZN(new_n4779_));
  NAND2_X1   g04523(.A1(new_n1828_), .A2(new_n4779_), .ZN(new_n4780_));
  XOR2_X1    g04524(.A1(new_n4780_), .A2(\a[23] ), .Z(new_n4781_));
  XNOR2_X1   g04525(.A1(new_n4776_), .A2(new_n4781_), .ZN(new_n4782_));
  INV_X1     g04526(.I(new_n4782_), .ZN(new_n4783_));
  OAI22_X1   g04527(.A1(new_n1168_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n1163_), .ZN(new_n4784_));
  NAND2_X1   g04528(.A1(new_n1774_), .A2(\b[26] ), .ZN(new_n4785_));
  AOI21_X1   g04529(.A1(new_n4784_), .A2(new_n4785_), .B(new_n1171_), .ZN(new_n4786_));
  NAND2_X1   g04530(.A1(new_n2174_), .A2(new_n4786_), .ZN(new_n4787_));
  XOR2_X1    g04531(.A1(new_n4787_), .A2(\a[20] ), .Z(new_n4788_));
  NOR2_X1    g04532(.A1(new_n4783_), .A2(new_n4788_), .ZN(new_n4789_));
  NAND2_X1   g04533(.A1(new_n4783_), .A2(new_n4788_), .ZN(new_n4790_));
  INV_X1     g04534(.I(new_n4790_), .ZN(new_n4791_));
  NOR2_X1    g04535(.A1(new_n4791_), .A2(new_n4789_), .ZN(new_n4792_));
  OAI22_X1   g04536(.A1(new_n940_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n935_), .ZN(new_n4793_));
  NAND2_X1   g04537(.A1(new_n1458_), .A2(\b[29] ), .ZN(new_n4794_));
  AOI21_X1   g04538(.A1(new_n4793_), .A2(new_n4794_), .B(new_n943_), .ZN(new_n4795_));
  NAND2_X1   g04539(.A1(new_n2546_), .A2(new_n4795_), .ZN(new_n4796_));
  XOR2_X1    g04540(.A1(new_n4796_), .A2(\a[17] ), .Z(new_n4797_));
  XOR2_X1    g04541(.A1(new_n4792_), .A2(new_n4797_), .Z(new_n4798_));
  OAI22_X1   g04542(.A1(new_n757_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n752_), .ZN(new_n4799_));
  NAND2_X1   g04543(.A1(new_n1182_), .A2(\b[32] ), .ZN(new_n4800_));
  AOI21_X1   g04544(.A1(new_n4799_), .A2(new_n4800_), .B(new_n760_), .ZN(new_n4801_));
  NAND2_X1   g04545(.A1(new_n2963_), .A2(new_n4801_), .ZN(new_n4802_));
  XOR2_X1    g04546(.A1(new_n4802_), .A2(\a[14] ), .Z(new_n4803_));
  INV_X1     g04547(.I(new_n4803_), .ZN(new_n4804_));
  XOR2_X1    g04548(.A1(new_n4798_), .A2(new_n4804_), .Z(new_n4805_));
  AOI21_X1   g04549(.A1(new_n4683_), .A2(new_n4680_), .B(new_n4805_), .ZN(new_n4806_));
  NAND2_X1   g04550(.A1(new_n4683_), .A2(new_n4680_), .ZN(new_n4807_));
  XOR2_X1    g04551(.A1(new_n4798_), .A2(new_n4803_), .Z(new_n4808_));
  NOR2_X1    g04552(.A1(new_n4807_), .A2(new_n4808_), .ZN(new_n4809_));
  NOR2_X1    g04553(.A1(new_n4809_), .A2(new_n4806_), .ZN(new_n4810_));
  OAI22_X1   g04554(.A1(new_n582_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n577_), .ZN(new_n4811_));
  NAND2_X1   g04555(.A1(new_n960_), .A2(\b[35] ), .ZN(new_n4812_));
  AOI21_X1   g04556(.A1(new_n4811_), .A2(new_n4812_), .B(new_n585_), .ZN(new_n4813_));
  NAND2_X1   g04557(.A1(new_n3411_), .A2(new_n4813_), .ZN(new_n4814_));
  XOR2_X1    g04558(.A1(new_n4814_), .A2(\a[11] ), .Z(new_n4815_));
  XNOR2_X1   g04559(.A1(new_n4810_), .A2(new_n4815_), .ZN(new_n4816_));
  XNOR2_X1   g04560(.A1(new_n4679_), .A2(new_n4816_), .ZN(new_n4817_));
  NOR2_X1    g04561(.A1(new_n4817_), .A2(new_n4677_), .ZN(new_n4818_));
  NAND2_X1   g04562(.A1(new_n4817_), .A2(new_n4677_), .ZN(new_n4819_));
  INV_X1     g04563(.I(new_n4819_), .ZN(new_n4820_));
  NOR2_X1    g04564(.A1(new_n4820_), .A2(new_n4818_), .ZN(new_n4821_));
  XOR2_X1    g04565(.A1(new_n4821_), .A2(new_n4671_), .Z(new_n4822_));
  OAI21_X1   g04566(.A1(new_n4661_), .A2(new_n4651_), .B(new_n4657_), .ZN(new_n4823_));
  XOR2_X1    g04567(.A1(new_n4823_), .A2(new_n4822_), .Z(new_n4824_));
  OAI21_X1   g04568(.A1(new_n4316_), .A2(new_n4509_), .B(new_n4501_), .ZN(new_n4825_));
  NAND2_X1   g04569(.A1(new_n4495_), .A2(new_n4825_), .ZN(new_n4826_));
  OAI21_X1   g04570(.A1(\b[43] ), .A2(\b[45] ), .B(\b[44] ), .ZN(new_n4827_));
  NAND2_X1   g04571(.A1(new_n4826_), .A2(new_n4827_), .ZN(new_n4828_));
  XNOR2_X1   g04572(.A1(\b[45] ), .A2(\b[46] ), .ZN(new_n4829_));
  INV_X1     g04573(.I(new_n4829_), .ZN(new_n4830_));
  NAND2_X1   g04574(.A1(new_n4828_), .A2(new_n4830_), .ZN(new_n4831_));
  XOR2_X1    g04575(.A1(\b[45] ), .A2(\b[46] ), .Z(new_n4832_));
  OAI21_X1   g04576(.A1(new_n4828_), .A2(new_n4832_), .B(new_n4831_), .ZN(new_n4833_));
  INV_X1     g04577(.I(\b[46] ), .ZN(new_n4834_));
  OAI22_X1   g04578(.A1(new_n405_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n404_), .ZN(new_n4835_));
  NAND2_X1   g04579(.A1(new_n279_), .A2(\b[44] ), .ZN(new_n4836_));
  AOI21_X1   g04580(.A1(new_n4835_), .A2(new_n4836_), .B(new_n264_), .ZN(new_n4837_));
  NAND2_X1   g04581(.A1(new_n4833_), .A2(new_n4837_), .ZN(new_n4838_));
  XOR2_X1    g04582(.A1(new_n4838_), .A2(\a[2] ), .Z(new_n4839_));
  XNOR2_X1   g04583(.A1(new_n4824_), .A2(new_n4839_), .ZN(new_n4840_));
  XOR2_X1    g04584(.A1(new_n4518_), .A2(new_n271_), .Z(new_n4841_));
  NAND2_X1   g04585(.A1(new_n4662_), .A2(new_n4841_), .ZN(new_n4842_));
  XOR2_X1    g04586(.A1(new_n4840_), .A2(new_n4842_), .Z(\f[46] ));
  NOR2_X1    g04587(.A1(new_n4821_), .A2(new_n4671_), .ZN(new_n4844_));
  NOR2_X1    g04588(.A1(new_n4651_), .A2(new_n4657_), .ZN(new_n4845_));
  INV_X1     g04589(.I(new_n4845_), .ZN(new_n4846_));
  NAND3_X1   g04590(.A1(new_n4487_), .A2(new_n4845_), .A3(new_n4660_), .ZN(new_n4847_));
  NAND3_X1   g04591(.A1(new_n4847_), .A2(new_n4846_), .A3(new_n4822_), .ZN(new_n4848_));
  NOR2_X1    g04592(.A1(new_n4848_), .A2(new_n4844_), .ZN(new_n4849_));
  OAI22_X1   g04593(.A1(new_n1444_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n1439_), .ZN(new_n4850_));
  NAND2_X1   g04594(.A1(new_n2098_), .A2(\b[24] ), .ZN(new_n4851_));
  AOI21_X1   g04595(.A1(new_n4850_), .A2(new_n4851_), .B(new_n1447_), .ZN(new_n4852_));
  NAND2_X1   g04596(.A1(new_n1926_), .A2(new_n4852_), .ZN(new_n4853_));
  XOR2_X1    g04597(.A1(new_n4853_), .A2(\a[23] ), .Z(new_n4854_));
  OAI22_X1   g04598(.A1(new_n1760_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n1755_), .ZN(new_n4855_));
  NAND2_X1   g04599(.A1(new_n2470_), .A2(\b[21] ), .ZN(new_n4856_));
  AOI21_X1   g04600(.A1(new_n4855_), .A2(new_n4856_), .B(new_n1763_), .ZN(new_n4857_));
  NAND2_X1   g04601(.A1(new_n1604_), .A2(new_n4857_), .ZN(new_n4858_));
  XOR2_X1    g04602(.A1(new_n4858_), .A2(\a[26] ), .Z(new_n4859_));
  INV_X1     g04603(.I(new_n4859_), .ZN(new_n4860_));
  INV_X1     g04604(.I(new_n4776_), .ZN(new_n4861_));
  XOR2_X1    g04605(.A1(new_n4687_), .A2(new_n4765_), .Z(new_n4862_));
  OAI21_X1   g04606(.A1(new_n4773_), .A2(new_n4862_), .B(new_n4861_), .ZN(new_n4863_));
  NOR2_X1    g04607(.A1(new_n4738_), .A2(new_n4743_), .ZN(new_n4864_));
  OAI22_X1   g04608(.A1(new_n4208_), .A2(new_n347_), .B1(new_n393_), .B2(new_n4203_), .ZN(new_n4865_));
  OAI21_X1   g04609(.A1(new_n290_), .A2(new_n4362_), .B(new_n4865_), .ZN(new_n4866_));
  AOI21_X1   g04610(.A1(new_n352_), .A2(new_n4210_), .B(new_n4866_), .ZN(new_n4867_));
  NAND2_X1   g04611(.A1(new_n4716_), .A2(new_n4717_), .ZN(new_n4868_));
  NOR2_X1    g04612(.A1(new_n4714_), .A2(new_n278_), .ZN(new_n4869_));
  XNOR2_X1   g04613(.A1(\a[44] ), .A2(\a[46] ), .ZN(new_n4870_));
  NAND2_X1   g04614(.A1(new_n4525_), .A2(new_n4870_), .ZN(new_n4871_));
  XNOR2_X1   g04615(.A1(\a[44] ), .A2(\a[47] ), .ZN(new_n4872_));
  NAND2_X1   g04616(.A1(new_n4871_), .A2(new_n4872_), .ZN(new_n4873_));
  OAI22_X1   g04617(.A1(new_n4711_), .A2(new_n292_), .B1(new_n267_), .B2(new_n4706_), .ZN(new_n4874_));
  NOR4_X1    g04618(.A1(new_n4874_), .A2(new_n258_), .A3(new_n4869_), .A4(new_n4873_), .ZN(new_n4875_));
  XOR2_X1    g04619(.A1(new_n4875_), .A2(new_n4701_), .Z(new_n4876_));
  XNOR2_X1   g04620(.A1(new_n4868_), .A2(new_n4876_), .ZN(new_n4877_));
  XOR2_X1    g04621(.A1(new_n4877_), .A2(\a[44] ), .Z(new_n4878_));
  XOR2_X1    g04622(.A1(new_n4878_), .A2(new_n4867_), .Z(new_n4879_));
  OAI21_X1   g04623(.A1(new_n4721_), .A2(new_n4718_), .B(new_n4722_), .ZN(new_n4880_));
  XNOR2_X1   g04624(.A1(new_n4880_), .A2(new_n4879_), .ZN(new_n4881_));
  OAI22_X1   g04625(.A1(new_n3736_), .A2(new_n495_), .B1(new_n450_), .B2(new_n3731_), .ZN(new_n4882_));
  NAND2_X1   g04626(.A1(new_n4730_), .A2(\b[6] ), .ZN(new_n4883_));
  AOI21_X1   g04627(.A1(new_n4882_), .A2(new_n4883_), .B(new_n3739_), .ZN(new_n4884_));
  NAND2_X1   g04628(.A1(new_n494_), .A2(new_n4884_), .ZN(new_n4885_));
  XOR2_X1    g04629(.A1(new_n4885_), .A2(\a[41] ), .Z(new_n4886_));
  XNOR2_X1   g04630(.A1(new_n4881_), .A2(new_n4886_), .ZN(new_n4887_));
  XOR2_X1    g04631(.A1(new_n4887_), .A2(new_n4735_), .Z(new_n4888_));
  OAI22_X1   g04632(.A1(new_n3298_), .A2(new_n659_), .B1(new_n617_), .B2(new_n3293_), .ZN(new_n4889_));
  NAND2_X1   g04633(.A1(new_n4227_), .A2(\b[9] ), .ZN(new_n4890_));
  AOI21_X1   g04634(.A1(new_n4889_), .A2(new_n4890_), .B(new_n3301_), .ZN(new_n4891_));
  NAND2_X1   g04635(.A1(new_n663_), .A2(new_n4891_), .ZN(new_n4892_));
  XOR2_X1    g04636(.A1(new_n4892_), .A2(\a[38] ), .Z(new_n4893_));
  XNOR2_X1   g04637(.A1(new_n4888_), .A2(new_n4893_), .ZN(new_n4894_));
  OAI22_X1   g04638(.A1(new_n2846_), .A2(new_n848_), .B1(new_n795_), .B2(new_n2841_), .ZN(new_n4895_));
  NAND2_X1   g04639(.A1(new_n3755_), .A2(\b[12] ), .ZN(new_n4896_));
  AOI21_X1   g04640(.A1(new_n4895_), .A2(new_n4896_), .B(new_n2849_), .ZN(new_n4897_));
  NAND2_X1   g04641(.A1(new_n847_), .A2(new_n4897_), .ZN(new_n4898_));
  XOR2_X1    g04642(.A1(new_n4898_), .A2(\a[35] ), .Z(new_n4899_));
  XOR2_X1    g04643(.A1(new_n4894_), .A2(new_n4899_), .Z(new_n4900_));
  NAND2_X1   g04644(.A1(new_n4900_), .A2(new_n4864_), .ZN(new_n4901_));
  XOR2_X1    g04645(.A1(new_n4894_), .A2(new_n4899_), .Z(new_n4902_));
  OAI21_X1   g04646(.A1(new_n4864_), .A2(new_n4902_), .B(new_n4901_), .ZN(new_n4903_));
  NOR2_X1    g04647(.A1(new_n4744_), .A2(new_n4749_), .ZN(new_n4904_));
  INV_X1     g04648(.I(new_n4904_), .ZN(new_n4905_));
  XOR2_X1    g04649(.A1(new_n4903_), .A2(new_n4905_), .Z(new_n4906_));
  OAI22_X1   g04650(.A1(new_n2452_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n2447_), .ZN(new_n4907_));
  NAND2_X1   g04651(.A1(new_n3312_), .A2(\b[15] ), .ZN(new_n4908_));
  AOI21_X1   g04652(.A1(new_n4907_), .A2(new_n4908_), .B(new_n2455_), .ZN(new_n4909_));
  NAND2_X1   g04653(.A1(new_n1047_), .A2(new_n4909_), .ZN(new_n4910_));
  XOR2_X1    g04654(.A1(new_n4910_), .A2(\a[32] ), .Z(new_n4911_));
  INV_X1     g04655(.I(new_n4911_), .ZN(new_n4912_));
  XOR2_X1    g04656(.A1(new_n4906_), .A2(new_n4912_), .Z(new_n4913_));
  NAND2_X1   g04657(.A1(new_n4750_), .A2(new_n4755_), .ZN(new_n4914_));
  OAI21_X1   g04658(.A1(new_n4692_), .A2(new_n4756_), .B(new_n4914_), .ZN(new_n4915_));
  XNOR2_X1   g04659(.A1(new_n4913_), .A2(new_n4915_), .ZN(new_n4916_));
  OAI22_X1   g04660(.A1(new_n2084_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n2079_), .ZN(new_n4917_));
  NAND2_X1   g04661(.A1(new_n2864_), .A2(\b[18] ), .ZN(new_n4918_));
  AOI21_X1   g04662(.A1(new_n4917_), .A2(new_n4918_), .B(new_n2087_), .ZN(new_n4919_));
  NAND2_X1   g04663(.A1(new_n1304_), .A2(new_n4919_), .ZN(new_n4920_));
  XOR2_X1    g04664(.A1(new_n4920_), .A2(\a[29] ), .Z(new_n4921_));
  XNOR2_X1   g04665(.A1(new_n4916_), .A2(new_n4921_), .ZN(new_n4922_));
  XOR2_X1    g04666(.A1(new_n4692_), .A2(new_n4756_), .Z(new_n4923_));
  NAND2_X1   g04667(.A1(new_n4923_), .A2(new_n4761_), .ZN(new_n4924_));
  NAND2_X1   g04668(.A1(new_n4688_), .A2(new_n4765_), .ZN(new_n4925_));
  NAND2_X1   g04669(.A1(new_n4925_), .A2(new_n4924_), .ZN(new_n4926_));
  NOR2_X1    g04670(.A1(new_n4926_), .A2(new_n4922_), .ZN(new_n4927_));
  NAND2_X1   g04671(.A1(new_n4926_), .A2(new_n4922_), .ZN(new_n4928_));
  INV_X1     g04672(.I(new_n4928_), .ZN(new_n4929_));
  NOR2_X1    g04673(.A1(new_n4929_), .A2(new_n4927_), .ZN(new_n4930_));
  XOR2_X1    g04674(.A1(new_n4930_), .A2(new_n4863_), .Z(new_n4931_));
  XOR2_X1    g04675(.A1(new_n4931_), .A2(new_n4860_), .Z(new_n4932_));
  XOR2_X1    g04676(.A1(new_n4932_), .A2(new_n4854_), .Z(new_n4933_));
  NOR2_X1    g04677(.A1(new_n4861_), .A2(new_n4781_), .ZN(new_n4934_));
  XOR2_X1    g04678(.A1(new_n4933_), .A2(new_n4934_), .Z(new_n4935_));
  OAI22_X1   g04679(.A1(new_n1168_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n1163_), .ZN(new_n4936_));
  NAND2_X1   g04680(.A1(new_n1774_), .A2(\b[27] ), .ZN(new_n4937_));
  AOI21_X1   g04681(.A1(new_n4936_), .A2(new_n4937_), .B(new_n1171_), .ZN(new_n4938_));
  NAND2_X1   g04682(.A1(new_n2276_), .A2(new_n4938_), .ZN(new_n4939_));
  XOR2_X1    g04683(.A1(new_n4939_), .A2(\a[20] ), .Z(new_n4940_));
  XOR2_X1    g04684(.A1(new_n4935_), .A2(new_n4940_), .Z(new_n4941_));
  NOR2_X1    g04685(.A1(new_n4783_), .A2(new_n4788_), .ZN(new_n4942_));
  XNOR2_X1   g04686(.A1(new_n4941_), .A2(new_n4942_), .ZN(new_n4943_));
  OAI22_X1   g04687(.A1(new_n940_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n935_), .ZN(new_n4944_));
  NAND2_X1   g04688(.A1(new_n1458_), .A2(\b[30] ), .ZN(new_n4945_));
  AOI21_X1   g04689(.A1(new_n4944_), .A2(new_n4945_), .B(new_n943_), .ZN(new_n4946_));
  NAND2_X1   g04690(.A1(new_n2659_), .A2(new_n4946_), .ZN(new_n4947_));
  XOR2_X1    g04691(.A1(new_n4947_), .A2(\a[17] ), .Z(new_n4948_));
  XNOR2_X1   g04692(.A1(new_n4943_), .A2(new_n4948_), .ZN(new_n4949_));
  NAND2_X1   g04693(.A1(new_n4807_), .A2(new_n4792_), .ZN(new_n4950_));
  XOR2_X1    g04694(.A1(new_n4950_), .A2(new_n4949_), .Z(new_n4951_));
  INV_X1     g04695(.I(new_n4797_), .ZN(new_n4952_));
  XOR2_X1    g04696(.A1(new_n4807_), .A2(new_n4792_), .Z(new_n4953_));
  NAND2_X1   g04697(.A1(new_n4953_), .A2(new_n4952_), .ZN(new_n4954_));
  XOR2_X1    g04698(.A1(new_n4951_), .A2(new_n4954_), .Z(new_n4955_));
  OAI22_X1   g04699(.A1(new_n757_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n752_), .ZN(new_n4956_));
  NAND2_X1   g04700(.A1(new_n1182_), .A2(\b[33] ), .ZN(new_n4957_));
  AOI21_X1   g04701(.A1(new_n4956_), .A2(new_n4957_), .B(new_n760_), .ZN(new_n4958_));
  NAND2_X1   g04702(.A1(new_n3101_), .A2(new_n4958_), .ZN(new_n4959_));
  XOR2_X1    g04703(.A1(new_n4959_), .A2(\a[14] ), .Z(new_n4960_));
  XOR2_X1    g04704(.A1(new_n4955_), .A2(new_n4960_), .Z(new_n4961_));
  INV_X1     g04705(.I(new_n4810_), .ZN(new_n4962_));
  XNOR2_X1   g04706(.A1(new_n4807_), .A2(new_n4798_), .ZN(new_n4963_));
  OAI21_X1   g04707(.A1(new_n4804_), .A2(new_n4963_), .B(new_n4962_), .ZN(new_n4964_));
  XOR2_X1    g04708(.A1(new_n4961_), .A2(new_n4964_), .Z(new_n4965_));
  OAI22_X1   g04709(.A1(new_n582_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n577_), .ZN(new_n4966_));
  NAND2_X1   g04710(.A1(new_n960_), .A2(\b[36] ), .ZN(new_n4967_));
  AOI21_X1   g04711(.A1(new_n4966_), .A2(new_n4967_), .B(new_n585_), .ZN(new_n4968_));
  NAND2_X1   g04712(.A1(new_n3565_), .A2(new_n4968_), .ZN(new_n4969_));
  XOR2_X1    g04713(.A1(new_n4969_), .A2(\a[11] ), .Z(new_n4970_));
  INV_X1     g04714(.I(new_n4970_), .ZN(new_n4971_));
  XOR2_X1    g04715(.A1(new_n4965_), .A2(new_n4971_), .Z(new_n4972_));
  INV_X1     g04716(.I(new_n4972_), .ZN(new_n4973_));
  NAND2_X1   g04717(.A1(new_n4962_), .A2(new_n4815_), .ZN(new_n4974_));
  NAND2_X1   g04718(.A1(new_n4679_), .A2(new_n4816_), .ZN(new_n4975_));
  NAND2_X1   g04719(.A1(new_n4975_), .A2(new_n4974_), .ZN(new_n4976_));
  XOR2_X1    g04720(.A1(new_n4976_), .A2(new_n4973_), .Z(new_n4977_));
  INV_X1     g04721(.I(new_n4977_), .ZN(new_n4978_));
  OAI22_X1   g04722(.A1(new_n437_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n431_), .ZN(new_n4979_));
  NAND2_X1   g04723(.A1(new_n775_), .A2(\b[39] ), .ZN(new_n4980_));
  AOI21_X1   g04724(.A1(new_n4979_), .A2(new_n4980_), .B(new_n440_), .ZN(new_n4981_));
  NAND2_X1   g04725(.A1(new_n3996_), .A2(new_n4981_), .ZN(new_n4982_));
  XOR2_X1    g04726(.A1(new_n4982_), .A2(\a[8] ), .Z(new_n4983_));
  NOR2_X1    g04727(.A1(new_n4978_), .A2(new_n4983_), .ZN(new_n4984_));
  INV_X1     g04728(.I(new_n4984_), .ZN(new_n4985_));
  NAND2_X1   g04729(.A1(new_n4978_), .A2(new_n4983_), .ZN(new_n4986_));
  AOI21_X1   g04730(.A1(new_n4985_), .A2(new_n4986_), .B(new_n4819_), .ZN(new_n4987_));
  XOR2_X1    g04731(.A1(new_n4977_), .A2(new_n4983_), .Z(new_n4988_));
  NOR2_X1    g04732(.A1(new_n4988_), .A2(new_n4820_), .ZN(new_n4989_));
  NOR2_X1    g04733(.A1(new_n4987_), .A2(new_n4989_), .ZN(new_n4990_));
  OAI22_X1   g04734(.A1(new_n364_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n320_), .ZN(new_n4991_));
  NAND2_X1   g04735(.A1(new_n594_), .A2(\b[42] ), .ZN(new_n4992_));
  AOI21_X1   g04736(.A1(new_n4991_), .A2(new_n4992_), .B(new_n312_), .ZN(new_n4993_));
  NAND2_X1   g04737(.A1(new_n4500_), .A2(new_n4993_), .ZN(new_n4994_));
  XOR2_X1    g04738(.A1(new_n4994_), .A2(\a[5] ), .Z(new_n4995_));
  XNOR2_X1   g04739(.A1(new_n4990_), .A2(new_n4995_), .ZN(new_n4996_));
  INV_X1     g04740(.I(\b[47] ), .ZN(new_n4997_));
  NOR2_X1    g04741(.A1(new_n4828_), .A2(new_n4509_), .ZN(new_n4998_));
  INV_X1     g04742(.I(new_n4828_), .ZN(new_n4999_));
  NOR2_X1    g04743(.A1(new_n4999_), .A2(\b[45] ), .ZN(new_n5000_));
  OR2_X2     g04744(.A1(new_n5000_), .A2(new_n4998_), .Z(new_n5001_));
  AND3_X2    g04745(.A1(new_n5001_), .A2(new_n4997_), .A3(new_n4830_), .Z(new_n5002_));
  AOI21_X1   g04746(.A1(new_n5001_), .A2(new_n4830_), .B(new_n4997_), .ZN(new_n5003_));
  OR2_X2     g04747(.A1(new_n5002_), .A2(new_n5003_), .Z(new_n5004_));
  OAI22_X1   g04748(.A1(new_n405_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n404_), .ZN(new_n5005_));
  NAND2_X1   g04749(.A1(new_n279_), .A2(\b[45] ), .ZN(new_n5006_));
  AOI21_X1   g04750(.A1(new_n5005_), .A2(new_n5006_), .B(new_n264_), .ZN(new_n5007_));
  NAND2_X1   g04751(.A1(new_n5004_), .A2(new_n5007_), .ZN(new_n5008_));
  XOR2_X1    g04752(.A1(new_n5008_), .A2(\a[2] ), .Z(new_n5009_));
  XNOR2_X1   g04753(.A1(new_n4996_), .A2(new_n5009_), .ZN(new_n5010_));
  INV_X1     g04754(.I(new_n5010_), .ZN(new_n5011_));
  XOR2_X1    g04755(.A1(new_n4996_), .A2(new_n5009_), .Z(new_n5012_));
  NOR2_X1    g04756(.A1(new_n4849_), .A2(new_n5012_), .ZN(new_n5013_));
  AOI21_X1   g04757(.A1(new_n4849_), .A2(new_n5011_), .B(new_n5013_), .ZN(new_n5014_));
  INV_X1     g04758(.I(new_n5014_), .ZN(\f[47] ));
  INV_X1     g04759(.I(new_n4995_), .ZN(new_n5016_));
  OR2_X2     g04760(.A1(new_n4996_), .A2(new_n4844_), .Z(new_n5017_));
  OAI22_X1   g04761(.A1(new_n4848_), .A2(new_n5017_), .B1(new_n5016_), .B2(new_n4996_), .ZN(new_n5018_));
  INV_X1     g04762(.I(new_n4868_), .ZN(new_n5019_));
  NAND2_X1   g04763(.A1(new_n5019_), .A2(new_n4876_), .ZN(new_n5020_));
  NOR2_X1    g04764(.A1(new_n4873_), .A2(new_n267_), .ZN(new_n5021_));
  OAI22_X1   g04765(.A1(new_n4711_), .A2(new_n290_), .B1(new_n292_), .B2(new_n4706_), .ZN(new_n5022_));
  NOR4_X1    g04766(.A1(new_n5022_), .A2(new_n677_), .A3(new_n4714_), .A4(new_n5021_), .ZN(new_n5023_));
  XOR2_X1    g04767(.A1(new_n5023_), .A2(new_n4701_), .Z(new_n5024_));
  XNOR2_X1   g04768(.A1(\a[47] ), .A2(\a[48] ), .ZN(new_n5025_));
  NOR2_X1    g04769(.A1(new_n5025_), .A2(new_n258_), .ZN(new_n5026_));
  XOR2_X1    g04770(.A1(new_n5024_), .A2(new_n5026_), .Z(new_n5027_));
  XNOR2_X1   g04771(.A1(new_n5027_), .A2(new_n5020_), .ZN(new_n5028_));
  INV_X1     g04772(.I(new_n4203_), .ZN(new_n5029_));
  AOI22_X1   g04773(.A1(\b[6] ), .A2(new_n4207_), .B1(new_n5029_), .B2(\b[5] ), .ZN(new_n5030_));
  NOR2_X1    g04774(.A1(new_n4362_), .A2(new_n393_), .ZN(new_n5031_));
  OAI21_X1   g04775(.A1(new_n5030_), .A2(new_n5031_), .B(new_n4210_), .ZN(new_n5032_));
  NOR2_X1    g04776(.A1(new_n524_), .A2(new_n5032_), .ZN(new_n5033_));
  XOR2_X1    g04777(.A1(new_n5033_), .A2(new_n4198_), .Z(new_n5034_));
  NAND2_X1   g04778(.A1(new_n4696_), .A2(new_n4723_), .ZN(new_n5035_));
  NAND2_X1   g04779(.A1(new_n4867_), .A2(new_n4198_), .ZN(new_n5036_));
  NOR2_X1    g04780(.A1(new_n4867_), .A2(new_n4198_), .ZN(new_n5037_));
  NAND2_X1   g04781(.A1(new_n4724_), .A2(new_n4877_), .ZN(new_n5038_));
  NOR2_X1    g04782(.A1(new_n5038_), .A2(new_n5037_), .ZN(new_n5039_));
  NAND4_X1   g04783(.A1(new_n4879_), .A2(new_n5035_), .A3(new_n5036_), .A4(new_n5039_), .ZN(new_n5040_));
  XOR2_X1    g04784(.A1(new_n5040_), .A2(new_n5034_), .Z(new_n5041_));
  XNOR2_X1   g04785(.A1(new_n5041_), .A2(new_n5028_), .ZN(new_n5042_));
  OAI22_X1   g04786(.A1(new_n3736_), .A2(new_n510_), .B1(new_n495_), .B2(new_n3731_), .ZN(new_n5043_));
  NAND2_X1   g04787(.A1(new_n4730_), .A2(\b[7] ), .ZN(new_n5044_));
  AOI21_X1   g04788(.A1(new_n5043_), .A2(new_n5044_), .B(new_n3739_), .ZN(new_n5045_));
  NAND2_X1   g04789(.A1(new_n518_), .A2(new_n5045_), .ZN(new_n5046_));
  XOR2_X1    g04790(.A1(new_n5046_), .A2(\a[41] ), .Z(new_n5047_));
  INV_X1     g04791(.I(new_n4881_), .ZN(new_n5048_));
  NAND2_X1   g04792(.A1(new_n5048_), .A2(new_n4886_), .ZN(new_n5049_));
  NAND3_X1   g04793(.A1(new_n4887_), .A2(new_n4737_), .A3(new_n5049_), .ZN(new_n5050_));
  XOR2_X1    g04794(.A1(new_n5050_), .A2(new_n5047_), .Z(new_n5051_));
  XNOR2_X1   g04795(.A1(new_n5051_), .A2(new_n5042_), .ZN(new_n5052_));
  OAI22_X1   g04796(.A1(new_n3298_), .A2(new_n717_), .B1(new_n659_), .B2(new_n3293_), .ZN(new_n5053_));
  NAND2_X1   g04797(.A1(new_n4227_), .A2(\b[10] ), .ZN(new_n5054_));
  AOI21_X1   g04798(.A1(new_n5053_), .A2(new_n5054_), .B(new_n3301_), .ZN(new_n5055_));
  NAND2_X1   g04799(.A1(new_n716_), .A2(new_n5055_), .ZN(new_n5056_));
  XOR2_X1    g04800(.A1(new_n5056_), .A2(new_n3288_), .Z(new_n5057_));
  AOI21_X1   g04801(.A1(new_n4888_), .A2(new_n4893_), .B(new_n4864_), .ZN(new_n5058_));
  XOR2_X1    g04802(.A1(new_n5058_), .A2(new_n5057_), .Z(new_n5059_));
  XNOR2_X1   g04803(.A1(new_n5052_), .A2(new_n5059_), .ZN(new_n5060_));
  OAI22_X1   g04804(.A1(new_n2846_), .A2(new_n904_), .B1(new_n848_), .B2(new_n2841_), .ZN(new_n5061_));
  NAND2_X1   g04805(.A1(new_n3755_), .A2(\b[13] ), .ZN(new_n5062_));
  AOI21_X1   g04806(.A1(new_n5061_), .A2(new_n5062_), .B(new_n2849_), .ZN(new_n5063_));
  NAND2_X1   g04807(.A1(new_n907_), .A2(new_n5063_), .ZN(new_n5064_));
  XOR2_X1    g04808(.A1(new_n5064_), .A2(new_n2836_), .Z(new_n5065_));
  XOR2_X1    g04809(.A1(new_n4894_), .A2(new_n4864_), .Z(new_n5066_));
  NAND2_X1   g04810(.A1(new_n5066_), .A2(new_n4899_), .ZN(new_n5067_));
  NAND2_X1   g04811(.A1(new_n5067_), .A2(new_n4905_), .ZN(new_n5068_));
  NOR2_X1    g04812(.A1(new_n4903_), .A2(new_n5068_), .ZN(new_n5069_));
  XOR2_X1    g04813(.A1(new_n5069_), .A2(new_n5065_), .Z(new_n5070_));
  XNOR2_X1   g04814(.A1(new_n5070_), .A2(new_n5060_), .ZN(new_n5071_));
  OAI22_X1   g04815(.A1(new_n2452_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n2447_), .ZN(new_n5072_));
  NAND2_X1   g04816(.A1(new_n3312_), .A2(\b[16] ), .ZN(new_n5073_));
  AOI21_X1   g04817(.A1(new_n5072_), .A2(new_n5073_), .B(new_n2455_), .ZN(new_n5074_));
  NAND2_X1   g04818(.A1(new_n1123_), .A2(new_n5074_), .ZN(new_n5075_));
  XOR2_X1    g04819(.A1(new_n5075_), .A2(\a[32] ), .Z(new_n5076_));
  XOR2_X1    g04820(.A1(new_n4906_), .A2(new_n4912_), .Z(new_n5077_));
  NAND2_X1   g04821(.A1(new_n5077_), .A2(new_n4915_), .ZN(new_n5078_));
  XOR2_X1    g04822(.A1(new_n5078_), .A2(new_n5076_), .Z(new_n5079_));
  XNOR2_X1   g04823(.A1(new_n5079_), .A2(new_n5071_), .ZN(new_n5080_));
  OAI22_X1   g04824(.A1(new_n2084_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n2079_), .ZN(new_n5081_));
  NAND2_X1   g04825(.A1(new_n2864_), .A2(\b[19] ), .ZN(new_n5082_));
  AOI21_X1   g04826(.A1(new_n5081_), .A2(new_n5082_), .B(new_n2087_), .ZN(new_n5083_));
  NAND2_X1   g04827(.A1(new_n1396_), .A2(new_n5083_), .ZN(new_n5084_));
  XOR2_X1    g04828(.A1(new_n5084_), .A2(\a[29] ), .Z(new_n5085_));
  XOR2_X1    g04829(.A1(new_n4916_), .A2(new_n4921_), .Z(new_n5086_));
  NAND2_X1   g04830(.A1(new_n4926_), .A2(new_n5086_), .ZN(new_n5087_));
  XOR2_X1    g04831(.A1(new_n5087_), .A2(new_n5085_), .Z(new_n5088_));
  XNOR2_X1   g04832(.A1(new_n5088_), .A2(new_n5080_), .ZN(new_n5089_));
  OAI22_X1   g04833(.A1(new_n1760_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n1755_), .ZN(new_n5090_));
  NAND2_X1   g04834(.A1(new_n2470_), .A2(\b[22] ), .ZN(new_n5091_));
  AOI21_X1   g04835(.A1(new_n5090_), .A2(new_n5091_), .B(new_n1763_), .ZN(new_n5092_));
  NAND2_X1   g04836(.A1(new_n1708_), .A2(new_n5092_), .ZN(new_n5093_));
  XOR2_X1    g04837(.A1(new_n5093_), .A2(new_n1750_), .Z(new_n5094_));
  NAND2_X1   g04838(.A1(new_n4930_), .A2(new_n4859_), .ZN(new_n5095_));
  NOR2_X1    g04839(.A1(new_n4930_), .A2(new_n4859_), .ZN(new_n5096_));
  NOR2_X1    g04840(.A1(new_n5096_), .A2(new_n4863_), .ZN(new_n5097_));
  NOR2_X1    g04841(.A1(new_n4930_), .A2(new_n4860_), .ZN(new_n5098_));
  AOI21_X1   g04842(.A1(new_n5097_), .A2(new_n5095_), .B(new_n5098_), .ZN(new_n5099_));
  XOR2_X1    g04843(.A1(new_n5099_), .A2(new_n5094_), .Z(new_n5100_));
  XNOR2_X1   g04844(.A1(new_n5100_), .A2(new_n5089_), .ZN(new_n5101_));
  OAI22_X1   g04845(.A1(new_n1444_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n1439_), .ZN(new_n5102_));
  NAND2_X1   g04846(.A1(new_n2098_), .A2(\b[25] ), .ZN(new_n5103_));
  AOI21_X1   g04847(.A1(new_n5102_), .A2(new_n5103_), .B(new_n1447_), .ZN(new_n5104_));
  NAND2_X1   g04848(.A1(new_n2042_), .A2(new_n5104_), .ZN(new_n5105_));
  XOR2_X1    g04849(.A1(new_n5105_), .A2(new_n1434_), .Z(new_n5106_));
  XOR2_X1    g04850(.A1(new_n4930_), .A2(new_n4860_), .Z(new_n5107_));
  XOR2_X1    g04851(.A1(new_n5107_), .A2(new_n4863_), .Z(new_n5108_));
  AOI22_X1   g04852(.A1(new_n4933_), .A2(new_n4934_), .B1(new_n4854_), .B2(new_n5108_), .ZN(new_n5109_));
  XOR2_X1    g04853(.A1(new_n5109_), .A2(new_n5106_), .Z(new_n5110_));
  XNOR2_X1   g04854(.A1(new_n5110_), .A2(new_n5101_), .ZN(new_n5111_));
  OAI22_X1   g04855(.A1(new_n1168_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n1163_), .ZN(new_n5112_));
  NAND2_X1   g04856(.A1(new_n1774_), .A2(\b[28] ), .ZN(new_n5113_));
  AOI21_X1   g04857(.A1(new_n5112_), .A2(new_n5113_), .B(new_n1171_), .ZN(new_n5114_));
  NAND2_X1   g04858(.A1(new_n2404_), .A2(new_n5114_), .ZN(new_n5115_));
  XOR2_X1    g04859(.A1(new_n5115_), .A2(new_n1158_), .Z(new_n5116_));
  NAND2_X1   g04860(.A1(new_n4941_), .A2(new_n4942_), .ZN(new_n5117_));
  INV_X1     g04861(.I(new_n4935_), .ZN(new_n5118_));
  NAND2_X1   g04862(.A1(new_n5118_), .A2(new_n4940_), .ZN(new_n5119_));
  NAND2_X1   g04863(.A1(new_n5117_), .A2(new_n5119_), .ZN(new_n5120_));
  XOR2_X1    g04864(.A1(new_n5120_), .A2(new_n5116_), .Z(new_n5121_));
  XOR2_X1    g04865(.A1(new_n5121_), .A2(new_n5111_), .Z(new_n5122_));
  OAI22_X1   g04866(.A1(new_n940_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n935_), .ZN(new_n5123_));
  NAND2_X1   g04867(.A1(new_n1458_), .A2(\b[31] ), .ZN(new_n5124_));
  AOI21_X1   g04868(.A1(new_n5123_), .A2(new_n5124_), .B(new_n943_), .ZN(new_n5125_));
  NAND2_X1   g04869(.A1(new_n2797_), .A2(new_n5125_), .ZN(new_n5126_));
  XOR2_X1    g04870(.A1(new_n5126_), .A2(\a[17] ), .Z(new_n5127_));
  NAND2_X1   g04871(.A1(new_n4949_), .A2(new_n4952_), .ZN(new_n5128_));
  NAND3_X1   g04872(.A1(new_n4807_), .A2(new_n4792_), .A3(new_n5128_), .ZN(new_n5129_));
  NAND2_X1   g04873(.A1(new_n4943_), .A2(new_n4948_), .ZN(new_n5130_));
  NAND2_X1   g04874(.A1(new_n5129_), .A2(new_n5130_), .ZN(new_n5131_));
  XOR2_X1    g04875(.A1(new_n5131_), .A2(new_n5127_), .Z(new_n5132_));
  XNOR2_X1   g04876(.A1(new_n5132_), .A2(new_n5122_), .ZN(new_n5133_));
  OAI22_X1   g04877(.A1(new_n757_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n752_), .ZN(new_n5134_));
  NAND2_X1   g04878(.A1(new_n1182_), .A2(\b[34] ), .ZN(new_n5135_));
  AOI21_X1   g04879(.A1(new_n5134_), .A2(new_n5135_), .B(new_n760_), .ZN(new_n5136_));
  NAND2_X1   g04880(.A1(new_n3246_), .A2(new_n5136_), .ZN(new_n5137_));
  XOR2_X1    g04881(.A1(new_n5137_), .A2(\a[14] ), .Z(new_n5138_));
  INV_X1     g04882(.I(new_n4960_), .ZN(new_n5139_));
  NOR2_X1    g04883(.A1(new_n4955_), .A2(new_n5139_), .ZN(new_n5140_));
  INV_X1     g04884(.I(new_n4964_), .ZN(new_n5141_));
  NOR3_X1    g04885(.A1(new_n4961_), .A2(new_n5140_), .A3(new_n5141_), .ZN(new_n5142_));
  XOR2_X1    g04886(.A1(new_n5142_), .A2(new_n5138_), .Z(new_n5143_));
  XOR2_X1    g04887(.A1(new_n5143_), .A2(new_n5133_), .Z(new_n5144_));
  OAI22_X1   g04888(.A1(new_n582_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n577_), .ZN(new_n5145_));
  NAND2_X1   g04889(.A1(new_n960_), .A2(\b[37] ), .ZN(new_n5146_));
  AOI21_X1   g04890(.A1(new_n5145_), .A2(new_n5146_), .B(new_n585_), .ZN(new_n5147_));
  NAND2_X1   g04891(.A1(new_n3700_), .A2(new_n5147_), .ZN(new_n5148_));
  XOR2_X1    g04892(.A1(new_n5148_), .A2(\a[11] ), .Z(new_n5149_));
  NOR2_X1    g04893(.A1(new_n4965_), .A2(new_n4971_), .ZN(new_n5150_));
  NOR2_X1    g04894(.A1(new_n4973_), .A2(new_n5150_), .ZN(new_n5151_));
  NAND2_X1   g04895(.A1(new_n4976_), .A2(new_n5151_), .ZN(new_n5152_));
  XOR2_X1    g04896(.A1(new_n5152_), .A2(new_n5149_), .Z(new_n5153_));
  XNOR2_X1   g04897(.A1(new_n5153_), .A2(new_n5144_), .ZN(new_n5154_));
  OAI22_X1   g04898(.A1(new_n437_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n431_), .ZN(new_n5155_));
  NAND2_X1   g04899(.A1(new_n775_), .A2(\b[40] ), .ZN(new_n5156_));
  AOI21_X1   g04900(.A1(new_n5155_), .A2(new_n5156_), .B(new_n440_), .ZN(new_n5157_));
  NAND2_X1   g04901(.A1(new_n4017_), .A2(new_n5157_), .ZN(new_n5158_));
  XOR2_X1    g04902(.A1(new_n5158_), .A2(\a[8] ), .Z(new_n5159_));
  NAND2_X1   g04903(.A1(new_n4986_), .A2(new_n4819_), .ZN(new_n5160_));
  XOR2_X1    g04904(.A1(new_n5160_), .A2(new_n5159_), .Z(new_n5161_));
  XNOR2_X1   g04905(.A1(new_n5161_), .A2(new_n5154_), .ZN(new_n5162_));
  OAI22_X1   g04906(.A1(new_n364_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n320_), .ZN(new_n5163_));
  NAND2_X1   g04907(.A1(new_n594_), .A2(\b[43] ), .ZN(new_n5164_));
  AOI21_X1   g04908(.A1(new_n5163_), .A2(new_n5164_), .B(new_n312_), .ZN(new_n5165_));
  NAND2_X1   g04909(.A1(new_n4513_), .A2(new_n5165_), .ZN(new_n5166_));
  XOR2_X1    g04910(.A1(new_n5166_), .A2(\a[5] ), .Z(new_n5167_));
  XOR2_X1    g04911(.A1(new_n5162_), .A2(new_n5167_), .Z(new_n5168_));
  OAI21_X1   g04912(.A1(new_n4509_), .A2(new_n4997_), .B(new_n4834_), .ZN(new_n5169_));
  NAND2_X1   g04913(.A1(new_n4999_), .A2(new_n5169_), .ZN(new_n5170_));
  OAI21_X1   g04914(.A1(\b[45] ), .A2(\b[47] ), .B(\b[46] ), .ZN(new_n5171_));
  NAND2_X1   g04915(.A1(new_n5170_), .A2(new_n5171_), .ZN(new_n5172_));
  XNOR2_X1   g04916(.A1(\b[47] ), .A2(\b[48] ), .ZN(new_n5173_));
  INV_X1     g04917(.I(new_n5173_), .ZN(new_n5174_));
  NAND2_X1   g04918(.A1(new_n5172_), .A2(new_n5174_), .ZN(new_n5175_));
  XOR2_X1    g04919(.A1(\b[47] ), .A2(\b[48] ), .Z(new_n5176_));
  OAI21_X1   g04920(.A1(new_n5172_), .A2(new_n5176_), .B(new_n5175_), .ZN(new_n5177_));
  INV_X1     g04921(.I(\b[48] ), .ZN(new_n5178_));
  OAI22_X1   g04922(.A1(new_n405_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n404_), .ZN(new_n5179_));
  NAND2_X1   g04923(.A1(new_n279_), .A2(\b[46] ), .ZN(new_n5180_));
  AOI21_X1   g04924(.A1(new_n5179_), .A2(new_n5180_), .B(new_n264_), .ZN(new_n5181_));
  NAND2_X1   g04925(.A1(new_n5177_), .A2(new_n5181_), .ZN(new_n5182_));
  XOR2_X1    g04926(.A1(new_n5182_), .A2(\a[2] ), .Z(new_n5183_));
  XOR2_X1    g04927(.A1(new_n5168_), .A2(new_n5183_), .Z(new_n5184_));
  XOR2_X1    g04928(.A1(new_n5168_), .A2(new_n5183_), .Z(new_n5185_));
  NOR2_X1    g04929(.A1(new_n5018_), .A2(new_n5185_), .ZN(new_n5186_));
  AOI21_X1   g04930(.A1(new_n5018_), .A2(new_n5184_), .B(new_n5186_), .ZN(new_n5187_));
  XOR2_X1    g04931(.A1(new_n4849_), .A2(new_n4996_), .Z(new_n5188_));
  AOI21_X1   g04932(.A1(new_n5009_), .A2(new_n5188_), .B(new_n5014_), .ZN(new_n5189_));
  XNOR2_X1   g04933(.A1(new_n5189_), .A2(new_n5187_), .ZN(\f[48] ));
  NOR2_X1    g04934(.A1(new_n5172_), .A2(new_n4997_), .ZN(new_n5191_));
  AOI21_X1   g04935(.A1(new_n5170_), .A2(new_n5171_), .B(\b[47] ), .ZN(new_n5192_));
  OAI21_X1   g04936(.A1(new_n5191_), .A2(new_n5192_), .B(new_n5174_), .ZN(new_n5193_));
  NOR2_X1    g04937(.A1(new_n5193_), .A2(\b[49] ), .ZN(new_n5194_));
  AND2_X2    g04938(.A1(new_n5193_), .A2(\b[49] ), .Z(new_n5195_));
  OR2_X2     g04939(.A1(new_n5195_), .A2(new_n5194_), .Z(new_n5196_));
  INV_X1     g04940(.I(\b[49] ), .ZN(new_n5197_));
  OAI22_X1   g04941(.A1(new_n405_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n404_), .ZN(new_n5198_));
  NAND2_X1   g04942(.A1(new_n279_), .A2(\b[47] ), .ZN(new_n5199_));
  AOI21_X1   g04943(.A1(new_n5198_), .A2(new_n5199_), .B(new_n264_), .ZN(new_n5200_));
  NAND2_X1   g04944(.A1(new_n5196_), .A2(new_n5200_), .ZN(new_n5201_));
  XOR2_X1    g04945(.A1(new_n5201_), .A2(\a[2] ), .Z(new_n5202_));
  OAI22_X1   g04946(.A1(new_n364_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n320_), .ZN(new_n5203_));
  NAND2_X1   g04947(.A1(new_n594_), .A2(\b[44] ), .ZN(new_n5204_));
  AOI21_X1   g04948(.A1(new_n5203_), .A2(new_n5204_), .B(new_n312_), .ZN(new_n5205_));
  NAND2_X1   g04949(.A1(new_n4833_), .A2(new_n5205_), .ZN(new_n5206_));
  XOR2_X1    g04950(.A1(new_n5206_), .A2(\a[5] ), .Z(new_n5207_));
  INV_X1     g04951(.I(new_n5207_), .ZN(new_n5208_));
  NAND2_X1   g04952(.A1(new_n5162_), .A2(new_n5167_), .ZN(new_n5209_));
  NAND2_X1   g04953(.A1(new_n5018_), .A2(new_n5209_), .ZN(new_n5210_));
  OAI21_X1   g04954(.A1(new_n5162_), .A2(new_n5167_), .B(new_n5210_), .ZN(new_n5211_));
  NAND2_X1   g04955(.A1(new_n5027_), .A2(new_n4876_), .ZN(new_n5212_));
  NAND2_X1   g04956(.A1(new_n5212_), .A2(new_n4868_), .ZN(new_n5213_));
  NAND2_X1   g04957(.A1(new_n5024_), .A2(new_n5026_), .ZN(new_n5214_));
  XNOR2_X1   g04958(.A1(new_n5213_), .A2(new_n5214_), .ZN(new_n5215_));
  OAI22_X1   g04959(.A1(new_n4711_), .A2(new_n393_), .B1(new_n290_), .B2(new_n4706_), .ZN(new_n5216_));
  OAI21_X1   g04960(.A1(new_n292_), .A2(new_n4873_), .B(new_n5216_), .ZN(new_n5217_));
  NAND3_X1   g04961(.A1(new_n5217_), .A2(new_n334_), .A3(new_n4713_), .ZN(new_n5218_));
  XOR2_X1    g04962(.A1(new_n5218_), .A2(\a[47] ), .Z(new_n5219_));
  INV_X1     g04963(.I(\a[50] ), .ZN(new_n5220_));
  INV_X1     g04964(.I(\a[49] ), .ZN(new_n5221_));
  NOR3_X1    g04965(.A1(new_n5221_), .A2(\a[47] ), .A3(\a[48] ), .ZN(new_n5222_));
  INV_X1     g04966(.I(\a[48] ), .ZN(new_n5223_));
  NOR3_X1    g04967(.A1(new_n4701_), .A2(new_n5223_), .A3(\a[49] ), .ZN(new_n5224_));
  NOR2_X1    g04968(.A1(new_n5224_), .A2(new_n5222_), .ZN(new_n5225_));
  NOR2_X1    g04969(.A1(new_n5225_), .A2(new_n258_), .ZN(new_n5226_));
  XOR2_X1    g04970(.A1(\a[49] ), .A2(\a[50] ), .Z(new_n5227_));
  NAND2_X1   g04971(.A1(new_n5025_), .A2(new_n5227_), .ZN(new_n5228_));
  NOR2_X1    g04972(.A1(new_n5228_), .A2(new_n267_), .ZN(new_n5229_));
  XOR2_X1    g04973(.A1(\a[47] ), .A2(\a[48] ), .Z(new_n5230_));
  NAND2_X1   g04974(.A1(new_n5230_), .A2(new_n5227_), .ZN(new_n5231_));
  NOR4_X1    g04975(.A1(new_n5229_), .A2(new_n261_), .A3(new_n5226_), .A4(new_n5231_), .ZN(new_n5232_));
  XOR2_X1    g04976(.A1(new_n5232_), .A2(new_n5220_), .Z(new_n5233_));
  NOR2_X1    g04977(.A1(new_n5026_), .A2(new_n5220_), .ZN(new_n5234_));
  XNOR2_X1   g04978(.A1(new_n5233_), .A2(new_n5234_), .ZN(new_n5235_));
  XOR2_X1    g04979(.A1(new_n5219_), .A2(new_n5235_), .Z(new_n5236_));
  NOR2_X1    g04980(.A1(new_n5215_), .A2(new_n5236_), .ZN(new_n5237_));
  INV_X1     g04981(.I(new_n5215_), .ZN(new_n5238_));
  XNOR2_X1   g04982(.A1(new_n5219_), .A2(new_n5235_), .ZN(new_n5239_));
  NOR2_X1    g04983(.A1(new_n5238_), .A2(new_n5239_), .ZN(new_n5240_));
  NOR2_X1    g04984(.A1(new_n5240_), .A2(new_n5237_), .ZN(new_n5241_));
  INV_X1     g04985(.I(new_n5241_), .ZN(new_n5242_));
  OAI22_X1   g04986(.A1(new_n4208_), .A2(new_n450_), .B1(new_n403_), .B2(new_n4203_), .ZN(new_n5243_));
  INV_X1     g04987(.I(new_n4362_), .ZN(new_n5244_));
  NAND2_X1   g04988(.A1(new_n5244_), .A2(\b[5] ), .ZN(new_n5245_));
  AOI21_X1   g04989(.A1(new_n5243_), .A2(new_n5245_), .B(new_n4211_), .ZN(new_n5246_));
  NAND2_X1   g04990(.A1(new_n454_), .A2(new_n5246_), .ZN(new_n5247_));
  XOR2_X1    g04991(.A1(new_n5247_), .A2(\a[44] ), .Z(new_n5248_));
  NOR2_X1    g04992(.A1(new_n5242_), .A2(new_n5248_), .ZN(new_n5249_));
  INV_X1     g04993(.I(new_n5249_), .ZN(new_n5250_));
  NAND2_X1   g04994(.A1(new_n5242_), .A2(new_n5248_), .ZN(new_n5251_));
  NAND2_X1   g04995(.A1(new_n5250_), .A2(new_n5251_), .ZN(new_n5252_));
  OAI22_X1   g04996(.A1(new_n3736_), .A2(new_n617_), .B1(new_n510_), .B2(new_n3731_), .ZN(new_n5253_));
  NAND2_X1   g04997(.A1(new_n4730_), .A2(\b[8] ), .ZN(new_n5254_));
  AOI21_X1   g04998(.A1(new_n5253_), .A2(new_n5254_), .B(new_n3739_), .ZN(new_n5255_));
  NAND2_X1   g04999(.A1(new_n616_), .A2(new_n5255_), .ZN(new_n5256_));
  XOR2_X1    g05000(.A1(new_n5256_), .A2(\a[41] ), .Z(new_n5257_));
  XNOR2_X1   g05001(.A1(new_n5252_), .A2(new_n5257_), .ZN(new_n5258_));
  OAI22_X1   g05002(.A1(new_n3298_), .A2(new_n795_), .B1(new_n717_), .B2(new_n3293_), .ZN(new_n5259_));
  NAND2_X1   g05003(.A1(new_n4227_), .A2(\b[11] ), .ZN(new_n5260_));
  AOI21_X1   g05004(.A1(new_n5259_), .A2(new_n5260_), .B(new_n3301_), .ZN(new_n5261_));
  NAND2_X1   g05005(.A1(new_n799_), .A2(new_n5261_), .ZN(new_n5262_));
  XOR2_X1    g05006(.A1(new_n5262_), .A2(\a[38] ), .Z(new_n5263_));
  NOR2_X1    g05007(.A1(new_n5258_), .A2(new_n5263_), .ZN(new_n5264_));
  INV_X1     g05008(.I(new_n5264_), .ZN(new_n5265_));
  NAND2_X1   g05009(.A1(new_n5258_), .A2(new_n5263_), .ZN(new_n5266_));
  NAND2_X1   g05010(.A1(new_n5265_), .A2(new_n5266_), .ZN(new_n5267_));
  OAI22_X1   g05011(.A1(new_n2846_), .A2(new_n992_), .B1(new_n904_), .B2(new_n2841_), .ZN(new_n5268_));
  NAND2_X1   g05012(.A1(new_n3755_), .A2(\b[14] ), .ZN(new_n5269_));
  AOI21_X1   g05013(.A1(new_n5268_), .A2(new_n5269_), .B(new_n2849_), .ZN(new_n5270_));
  NAND2_X1   g05014(.A1(new_n991_), .A2(new_n5270_), .ZN(new_n5271_));
  XOR2_X1    g05015(.A1(new_n5271_), .A2(\a[35] ), .Z(new_n5272_));
  XOR2_X1    g05016(.A1(new_n5267_), .A2(new_n5272_), .Z(new_n5273_));
  INV_X1     g05017(.I(new_n5273_), .ZN(new_n5274_));
  OAI22_X1   g05018(.A1(new_n2452_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n2447_), .ZN(new_n5275_));
  NAND2_X1   g05019(.A1(new_n3312_), .A2(\b[17] ), .ZN(new_n5276_));
  AOI21_X1   g05020(.A1(new_n5275_), .A2(new_n5276_), .B(new_n2455_), .ZN(new_n5277_));
  NAND2_X1   g05021(.A1(new_n1225_), .A2(new_n5277_), .ZN(new_n5278_));
  XOR2_X1    g05022(.A1(new_n5278_), .A2(\a[32] ), .Z(new_n5279_));
  NOR2_X1    g05023(.A1(new_n5274_), .A2(new_n5279_), .ZN(new_n5280_));
  INV_X1     g05024(.I(new_n5279_), .ZN(new_n5281_));
  NOR2_X1    g05025(.A1(new_n5273_), .A2(new_n5281_), .ZN(new_n5282_));
  NOR2_X1    g05026(.A1(new_n5280_), .A2(new_n5282_), .ZN(new_n5283_));
  OAI22_X1   g05027(.A1(new_n2084_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n2079_), .ZN(new_n5284_));
  NAND2_X1   g05028(.A1(new_n2864_), .A2(\b[20] ), .ZN(new_n5285_));
  AOI21_X1   g05029(.A1(new_n5284_), .A2(new_n5285_), .B(new_n2087_), .ZN(new_n5286_));
  NAND2_X1   g05030(.A1(new_n1517_), .A2(new_n5286_), .ZN(new_n5287_));
  XOR2_X1    g05031(.A1(new_n5287_), .A2(\a[29] ), .Z(new_n5288_));
  XOR2_X1    g05032(.A1(new_n5283_), .A2(new_n5288_), .Z(new_n5289_));
  OAI22_X1   g05033(.A1(new_n1760_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n1755_), .ZN(new_n5290_));
  NAND2_X1   g05034(.A1(new_n2470_), .A2(\b[23] ), .ZN(new_n5291_));
  AOI21_X1   g05035(.A1(new_n5290_), .A2(new_n5291_), .B(new_n1763_), .ZN(new_n5292_));
  NAND2_X1   g05036(.A1(new_n1828_), .A2(new_n5292_), .ZN(new_n5293_));
  XOR2_X1    g05037(.A1(new_n5293_), .A2(\a[26] ), .Z(new_n5294_));
  XOR2_X1    g05038(.A1(new_n5289_), .A2(new_n5294_), .Z(new_n5295_));
  OAI22_X1   g05039(.A1(new_n1444_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n1439_), .ZN(new_n5296_));
  NAND2_X1   g05040(.A1(new_n2098_), .A2(\b[26] ), .ZN(new_n5297_));
  AOI21_X1   g05041(.A1(new_n5296_), .A2(new_n5297_), .B(new_n1447_), .ZN(new_n5298_));
  NAND2_X1   g05042(.A1(new_n2174_), .A2(new_n5298_), .ZN(new_n5299_));
  XOR2_X1    g05043(.A1(new_n5299_), .A2(\a[23] ), .Z(new_n5300_));
  XOR2_X1    g05044(.A1(new_n5295_), .A2(new_n5300_), .Z(new_n5301_));
  OAI22_X1   g05045(.A1(new_n1168_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n1163_), .ZN(new_n5302_));
  NAND2_X1   g05046(.A1(new_n1774_), .A2(\b[29] ), .ZN(new_n5303_));
  AOI21_X1   g05047(.A1(new_n5302_), .A2(new_n5303_), .B(new_n1171_), .ZN(new_n5304_));
  NAND2_X1   g05048(.A1(new_n2546_), .A2(new_n5304_), .ZN(new_n5305_));
  XOR2_X1    g05049(.A1(new_n5305_), .A2(\a[20] ), .Z(new_n5306_));
  XOR2_X1    g05050(.A1(new_n5301_), .A2(new_n5306_), .Z(new_n5307_));
  XOR2_X1    g05051(.A1(new_n5111_), .A2(new_n5116_), .Z(new_n5308_));
  AOI21_X1   g05052(.A1(new_n5116_), .A2(new_n5120_), .B(new_n5308_), .ZN(new_n5309_));
  XOR2_X1    g05053(.A1(new_n5309_), .A2(new_n5307_), .Z(new_n5310_));
  OAI22_X1   g05054(.A1(new_n940_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n935_), .ZN(new_n5311_));
  NAND2_X1   g05055(.A1(new_n1458_), .A2(\b[32] ), .ZN(new_n5312_));
  AOI21_X1   g05056(.A1(new_n5311_), .A2(new_n5312_), .B(new_n943_), .ZN(new_n5313_));
  NAND2_X1   g05057(.A1(new_n2963_), .A2(new_n5313_), .ZN(new_n5314_));
  XOR2_X1    g05058(.A1(new_n5314_), .A2(\a[17] ), .Z(new_n5315_));
  XOR2_X1    g05059(.A1(new_n5310_), .A2(new_n5315_), .Z(new_n5316_));
  OAI22_X1   g05060(.A1(new_n757_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n752_), .ZN(new_n5317_));
  NAND2_X1   g05061(.A1(new_n1182_), .A2(\b[35] ), .ZN(new_n5318_));
  AOI21_X1   g05062(.A1(new_n5317_), .A2(new_n5318_), .B(new_n760_), .ZN(new_n5319_));
  NAND2_X1   g05063(.A1(new_n3411_), .A2(new_n5319_), .ZN(new_n5320_));
  XOR2_X1    g05064(.A1(new_n5320_), .A2(\a[14] ), .Z(new_n5321_));
  XOR2_X1    g05065(.A1(new_n5316_), .A2(new_n5321_), .Z(new_n5322_));
  XOR2_X1    g05066(.A1(new_n5133_), .A2(new_n5138_), .Z(new_n5323_));
  OAI21_X1   g05067(.A1(new_n5138_), .A2(new_n5142_), .B(new_n5323_), .ZN(new_n5324_));
  XNOR2_X1   g05068(.A1(new_n5324_), .A2(new_n5322_), .ZN(new_n5325_));
  OAI22_X1   g05069(.A1(new_n582_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n577_), .ZN(new_n5326_));
  NAND2_X1   g05070(.A1(new_n960_), .A2(\b[38] ), .ZN(new_n5327_));
  AOI21_X1   g05071(.A1(new_n5326_), .A2(new_n5327_), .B(new_n585_), .ZN(new_n5328_));
  NAND2_X1   g05072(.A1(new_n3844_), .A2(new_n5328_), .ZN(new_n5329_));
  XOR2_X1    g05073(.A1(new_n5329_), .A2(\a[11] ), .Z(new_n5330_));
  INV_X1     g05074(.I(new_n5330_), .ZN(new_n5331_));
  XOR2_X1    g05075(.A1(new_n5325_), .A2(new_n5331_), .Z(new_n5332_));
  OAI22_X1   g05076(.A1(new_n437_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n431_), .ZN(new_n5333_));
  NAND2_X1   g05077(.A1(new_n775_), .A2(\b[41] ), .ZN(new_n5334_));
  AOI21_X1   g05078(.A1(new_n5333_), .A2(new_n5334_), .B(new_n440_), .ZN(new_n5335_));
  NAND2_X1   g05079(.A1(new_n4320_), .A2(new_n5335_), .ZN(new_n5336_));
  XOR2_X1    g05080(.A1(new_n5336_), .A2(\a[8] ), .Z(new_n5337_));
  XNOR2_X1   g05081(.A1(new_n5332_), .A2(new_n5337_), .ZN(new_n5338_));
  XOR2_X1    g05082(.A1(new_n5211_), .A2(new_n5338_), .Z(new_n5339_));
  XOR2_X1    g05083(.A1(new_n5339_), .A2(new_n5208_), .Z(new_n5340_));
  XOR2_X1    g05084(.A1(new_n5340_), .A2(new_n5202_), .Z(new_n5341_));
  INV_X1     g05085(.I(new_n5183_), .ZN(new_n5342_));
  NAND2_X1   g05086(.A1(new_n5189_), .A2(new_n5187_), .ZN(new_n5343_));
  XOR2_X1    g05087(.A1(new_n5018_), .A2(new_n5168_), .Z(new_n5344_));
  OAI21_X1   g05088(.A1(new_n5342_), .A2(new_n5344_), .B(new_n5343_), .ZN(new_n5345_));
  XOR2_X1    g05089(.A1(new_n5341_), .A2(new_n5345_), .Z(\f[49] ));
  XOR2_X1    g05090(.A1(new_n5338_), .A2(new_n5208_), .Z(new_n5347_));
  INV_X1     g05091(.I(new_n5347_), .ZN(new_n5348_));
  XOR2_X1    g05092(.A1(new_n5211_), .A2(new_n5348_), .Z(new_n5349_));
  NAND2_X1   g05093(.A1(new_n5349_), .A2(new_n5202_), .ZN(new_n5350_));
  NAND2_X1   g05094(.A1(new_n5341_), .A2(new_n5345_), .ZN(new_n5351_));
  NAND2_X1   g05095(.A1(new_n5351_), .A2(new_n5350_), .ZN(new_n5352_));
  INV_X1     g05096(.I(new_n5332_), .ZN(new_n5353_));
  NOR2_X1    g05097(.A1(new_n5353_), .A2(new_n5337_), .ZN(new_n5354_));
  OAI22_X1   g05098(.A1(new_n1760_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n1755_), .ZN(new_n5355_));
  NAND2_X1   g05099(.A1(new_n2470_), .A2(\b[24] ), .ZN(new_n5356_));
  AOI21_X1   g05100(.A1(new_n5355_), .A2(new_n5356_), .B(new_n1763_), .ZN(new_n5357_));
  NAND2_X1   g05101(.A1(new_n1926_), .A2(new_n5357_), .ZN(new_n5358_));
  XOR2_X1    g05102(.A1(new_n5358_), .A2(\a[26] ), .Z(new_n5359_));
  OAI22_X1   g05103(.A1(new_n2084_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n2079_), .ZN(new_n5360_));
  NAND2_X1   g05104(.A1(new_n2864_), .A2(\b[21] ), .ZN(new_n5361_));
  AOI21_X1   g05105(.A1(new_n5360_), .A2(new_n5361_), .B(new_n2087_), .ZN(new_n5362_));
  NAND2_X1   g05106(.A1(new_n1604_), .A2(new_n5362_), .ZN(new_n5363_));
  XOR2_X1    g05107(.A1(new_n5363_), .A2(\a[29] ), .Z(new_n5364_));
  NOR3_X1    g05108(.A1(new_n5280_), .A2(new_n5282_), .A3(new_n5288_), .ZN(new_n5365_));
  NOR2_X1    g05109(.A1(new_n5252_), .A2(new_n5257_), .ZN(new_n5366_));
  OAI22_X1   g05110(.A1(new_n4711_), .A2(new_n347_), .B1(new_n393_), .B2(new_n4706_), .ZN(new_n5367_));
  OAI21_X1   g05111(.A1(new_n290_), .A2(new_n4873_), .B(new_n5367_), .ZN(new_n5368_));
  AOI21_X1   g05112(.A1(new_n352_), .A2(new_n4713_), .B(new_n5368_), .ZN(new_n5369_));
  INV_X1     g05113(.I(new_n5232_), .ZN(new_n5370_));
  NOR3_X1    g05114(.A1(new_n5370_), .A2(new_n5220_), .A3(new_n5026_), .ZN(new_n5371_));
  XNOR2_X1   g05115(.A1(\a[49] ), .A2(\a[50] ), .ZN(new_n5372_));
  NOR3_X1    g05116(.A1(new_n5372_), .A2(new_n5230_), .A3(new_n292_), .ZN(new_n5373_));
  OAI21_X1   g05117(.A1(new_n5224_), .A2(new_n5222_), .B(\b[1] ), .ZN(new_n5374_));
  INV_X1     g05118(.I(new_n5374_), .ZN(new_n5375_));
  XOR2_X1    g05119(.A1(\a[47] ), .A2(\a[49] ), .Z(new_n5376_));
  XNOR2_X1   g05120(.A1(\a[47] ), .A2(\a[50] ), .ZN(new_n5377_));
  OAI21_X1   g05121(.A1(new_n5230_), .A2(new_n5376_), .B(new_n5377_), .ZN(new_n5378_));
  OAI22_X1   g05122(.A1(new_n258_), .A2(new_n5378_), .B1(new_n5375_), .B2(new_n5373_), .ZN(new_n5379_));
  NOR2_X1    g05123(.A1(new_n5231_), .A2(new_n278_), .ZN(new_n5380_));
  NAND3_X1   g05124(.A1(new_n5379_), .A2(new_n5220_), .A3(new_n5380_), .ZN(new_n5381_));
  NAND3_X1   g05125(.A1(new_n5025_), .A2(new_n5227_), .A3(\b[2] ), .ZN(new_n5382_));
  NOR2_X1    g05126(.A1(new_n5221_), .A2(\a[47] ), .ZN(new_n5383_));
  NOR2_X1    g05127(.A1(new_n4701_), .A2(\a[49] ), .ZN(new_n5384_));
  NOR2_X1    g05128(.A1(new_n5383_), .A2(new_n5384_), .ZN(new_n5385_));
  XOR2_X1    g05129(.A1(\a[47] ), .A2(\a[50] ), .Z(new_n5386_));
  AOI21_X1   g05130(.A1(new_n5385_), .A2(new_n5025_), .B(new_n5386_), .ZN(new_n5387_));
  AOI22_X1   g05131(.A1(new_n5387_), .A2(\b[0] ), .B1(new_n5382_), .B2(new_n5374_), .ZN(new_n5388_));
  INV_X1     g05132(.I(new_n278_), .ZN(new_n5389_));
  NAND2_X1   g05133(.A1(new_n4701_), .A2(\a[48] ), .ZN(new_n5390_));
  NAND2_X1   g05134(.A1(new_n5223_), .A2(\a[47] ), .ZN(new_n5391_));
  NAND2_X1   g05135(.A1(new_n5221_), .A2(\a[50] ), .ZN(new_n5392_));
  NAND2_X1   g05136(.A1(new_n5220_), .A2(\a[49] ), .ZN(new_n5393_));
  AOI22_X1   g05137(.A1(new_n5390_), .A2(new_n5391_), .B1(new_n5392_), .B2(new_n5393_), .ZN(new_n5394_));
  NAND2_X1   g05138(.A1(new_n5389_), .A2(new_n5394_), .ZN(new_n5395_));
  OAI21_X1   g05139(.A1(new_n5388_), .A2(new_n5395_), .B(\a[50] ), .ZN(new_n5396_));
  NAND2_X1   g05140(.A1(new_n5381_), .A2(new_n5396_), .ZN(new_n5397_));
  XOR2_X1    g05141(.A1(new_n5371_), .A2(new_n5397_), .Z(new_n5398_));
  XOR2_X1    g05142(.A1(new_n5398_), .A2(new_n4701_), .Z(new_n5399_));
  XOR2_X1    g05143(.A1(new_n5399_), .A2(new_n5369_), .Z(new_n5400_));
  INV_X1     g05144(.I(new_n5219_), .ZN(new_n5401_));
  OAI21_X1   g05145(.A1(new_n5238_), .A2(new_n5235_), .B(new_n5401_), .ZN(new_n5402_));
  XNOR2_X1   g05146(.A1(new_n5402_), .A2(new_n5400_), .ZN(new_n5403_));
  OAI22_X1   g05147(.A1(new_n4208_), .A2(new_n495_), .B1(new_n450_), .B2(new_n4203_), .ZN(new_n5404_));
  NAND2_X1   g05148(.A1(new_n5244_), .A2(\b[6] ), .ZN(new_n5405_));
  AOI21_X1   g05149(.A1(new_n5404_), .A2(new_n5405_), .B(new_n4211_), .ZN(new_n5406_));
  NAND2_X1   g05150(.A1(new_n494_), .A2(new_n5406_), .ZN(new_n5407_));
  XOR2_X1    g05151(.A1(new_n5407_), .A2(\a[44] ), .Z(new_n5408_));
  XNOR2_X1   g05152(.A1(new_n5403_), .A2(new_n5408_), .ZN(new_n5409_));
  XOR2_X1    g05153(.A1(new_n5409_), .A2(new_n5249_), .Z(new_n5410_));
  OAI22_X1   g05154(.A1(new_n3736_), .A2(new_n659_), .B1(new_n617_), .B2(new_n3731_), .ZN(new_n5411_));
  NAND2_X1   g05155(.A1(new_n4730_), .A2(\b[9] ), .ZN(new_n5412_));
  AOI21_X1   g05156(.A1(new_n5411_), .A2(new_n5412_), .B(new_n3739_), .ZN(new_n5413_));
  NAND2_X1   g05157(.A1(new_n663_), .A2(new_n5413_), .ZN(new_n5414_));
  XOR2_X1    g05158(.A1(new_n5414_), .A2(\a[41] ), .Z(new_n5415_));
  XNOR2_X1   g05159(.A1(new_n5410_), .A2(new_n5415_), .ZN(new_n5416_));
  OAI22_X1   g05160(.A1(new_n3298_), .A2(new_n848_), .B1(new_n795_), .B2(new_n3293_), .ZN(new_n5417_));
  NAND2_X1   g05161(.A1(new_n4227_), .A2(\b[12] ), .ZN(new_n5418_));
  AOI21_X1   g05162(.A1(new_n5417_), .A2(new_n5418_), .B(new_n3301_), .ZN(new_n5419_));
  NAND2_X1   g05163(.A1(new_n847_), .A2(new_n5419_), .ZN(new_n5420_));
  XOR2_X1    g05164(.A1(new_n5420_), .A2(\a[38] ), .Z(new_n5421_));
  XOR2_X1    g05165(.A1(new_n5416_), .A2(new_n5421_), .Z(new_n5422_));
  NAND2_X1   g05166(.A1(new_n5422_), .A2(new_n5366_), .ZN(new_n5423_));
  XOR2_X1    g05167(.A1(new_n5416_), .A2(new_n5421_), .Z(new_n5424_));
  OAI21_X1   g05168(.A1(new_n5366_), .A2(new_n5424_), .B(new_n5423_), .ZN(new_n5425_));
  XOR2_X1    g05169(.A1(new_n5425_), .A2(new_n5265_), .Z(new_n5426_));
  OAI22_X1   g05170(.A1(new_n2846_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n2841_), .ZN(new_n5427_));
  NAND2_X1   g05171(.A1(new_n3755_), .A2(\b[15] ), .ZN(new_n5428_));
  AOI21_X1   g05172(.A1(new_n5427_), .A2(new_n5428_), .B(new_n2849_), .ZN(new_n5429_));
  NAND2_X1   g05173(.A1(new_n1047_), .A2(new_n5429_), .ZN(new_n5430_));
  XOR2_X1    g05174(.A1(new_n5430_), .A2(\a[35] ), .Z(new_n5431_));
  XNOR2_X1   g05175(.A1(new_n5426_), .A2(new_n5431_), .ZN(new_n5432_));
  OR2_X2     g05176(.A1(new_n5267_), .A2(new_n5272_), .Z(new_n5433_));
  XNOR2_X1   g05177(.A1(new_n5432_), .A2(new_n5433_), .ZN(new_n5434_));
  OAI22_X1   g05178(.A1(new_n2452_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n2447_), .ZN(new_n5435_));
  NAND2_X1   g05179(.A1(new_n3312_), .A2(\b[18] ), .ZN(new_n5436_));
  AOI21_X1   g05180(.A1(new_n5435_), .A2(new_n5436_), .B(new_n2455_), .ZN(new_n5437_));
  NAND2_X1   g05181(.A1(new_n1304_), .A2(new_n5437_), .ZN(new_n5438_));
  XOR2_X1    g05182(.A1(new_n5438_), .A2(\a[32] ), .Z(new_n5439_));
  INV_X1     g05183(.I(new_n5439_), .ZN(new_n5440_));
  XOR2_X1    g05184(.A1(new_n5434_), .A2(new_n5440_), .Z(new_n5441_));
  NOR2_X1    g05185(.A1(new_n5274_), .A2(new_n5279_), .ZN(new_n5442_));
  XNOR2_X1   g05186(.A1(new_n5441_), .A2(new_n5442_), .ZN(new_n5443_));
  XOR2_X1    g05187(.A1(new_n5443_), .A2(new_n5365_), .Z(new_n5444_));
  XOR2_X1    g05188(.A1(new_n5444_), .A2(new_n5364_), .Z(new_n5445_));
  XOR2_X1    g05189(.A1(new_n5445_), .A2(new_n5359_), .Z(new_n5446_));
  NOR2_X1    g05190(.A1(new_n5289_), .A2(new_n5294_), .ZN(new_n5447_));
  XOR2_X1    g05191(.A1(new_n5446_), .A2(new_n5447_), .Z(new_n5448_));
  OAI22_X1   g05192(.A1(new_n1444_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n1439_), .ZN(new_n5449_));
  NAND2_X1   g05193(.A1(new_n2098_), .A2(\b[27] ), .ZN(new_n5450_));
  AOI21_X1   g05194(.A1(new_n5449_), .A2(new_n5450_), .B(new_n1447_), .ZN(new_n5451_));
  NAND2_X1   g05195(.A1(new_n2276_), .A2(new_n5451_), .ZN(new_n5452_));
  XOR2_X1    g05196(.A1(new_n5452_), .A2(\a[23] ), .Z(new_n5453_));
  XOR2_X1    g05197(.A1(new_n5448_), .A2(new_n5453_), .Z(new_n5454_));
  INV_X1     g05198(.I(new_n5295_), .ZN(new_n5455_));
  NOR2_X1    g05199(.A1(new_n5455_), .A2(new_n5300_), .ZN(new_n5456_));
  NAND2_X1   g05200(.A1(new_n5454_), .A2(new_n5456_), .ZN(new_n5457_));
  INV_X1     g05201(.I(new_n5457_), .ZN(new_n5458_));
  NOR2_X1    g05202(.A1(new_n5454_), .A2(new_n5456_), .ZN(new_n5459_));
  NOR2_X1    g05203(.A1(new_n5458_), .A2(new_n5459_), .ZN(new_n5460_));
  OAI22_X1   g05204(.A1(new_n1168_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n1163_), .ZN(new_n5461_));
  NAND2_X1   g05205(.A1(new_n1774_), .A2(\b[30] ), .ZN(new_n5462_));
  AOI21_X1   g05206(.A1(new_n5461_), .A2(new_n5462_), .B(new_n1171_), .ZN(new_n5463_));
  NAND2_X1   g05207(.A1(new_n2659_), .A2(new_n5463_), .ZN(new_n5464_));
  XOR2_X1    g05208(.A1(new_n5464_), .A2(\a[20] ), .Z(new_n5465_));
  XNOR2_X1   g05209(.A1(new_n5460_), .A2(new_n5465_), .ZN(new_n5466_));
  NAND2_X1   g05210(.A1(new_n5301_), .A2(new_n5306_), .ZN(new_n5467_));
  INV_X1     g05211(.I(new_n5307_), .ZN(new_n5468_));
  OAI21_X1   g05212(.A1(new_n5309_), .A2(new_n5468_), .B(new_n5467_), .ZN(new_n5469_));
  XOR2_X1    g05213(.A1(new_n5469_), .A2(new_n5466_), .Z(new_n5470_));
  INV_X1     g05214(.I(new_n5470_), .ZN(new_n5471_));
  OAI22_X1   g05215(.A1(new_n940_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n935_), .ZN(new_n5472_));
  NAND2_X1   g05216(.A1(new_n1458_), .A2(\b[33] ), .ZN(new_n5473_));
  AOI21_X1   g05217(.A1(new_n5472_), .A2(new_n5473_), .B(new_n943_), .ZN(new_n5474_));
  NAND2_X1   g05218(.A1(new_n3101_), .A2(new_n5474_), .ZN(new_n5475_));
  XOR2_X1    g05219(.A1(new_n5475_), .A2(\a[17] ), .Z(new_n5476_));
  NOR2_X1    g05220(.A1(new_n5471_), .A2(new_n5476_), .ZN(new_n5477_));
  NAND2_X1   g05221(.A1(new_n5471_), .A2(new_n5476_), .ZN(new_n5478_));
  INV_X1     g05222(.I(new_n5478_), .ZN(new_n5479_));
  NOR2_X1    g05223(.A1(new_n5479_), .A2(new_n5477_), .ZN(new_n5480_));
  INV_X1     g05224(.I(new_n5310_), .ZN(new_n5481_));
  NOR2_X1    g05225(.A1(new_n5481_), .A2(new_n5315_), .ZN(new_n5482_));
  XOR2_X1    g05226(.A1(new_n5480_), .A2(new_n5482_), .Z(new_n5483_));
  OAI22_X1   g05227(.A1(new_n757_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n752_), .ZN(new_n5484_));
  NAND2_X1   g05228(.A1(new_n1182_), .A2(\b[36] ), .ZN(new_n5485_));
  AOI21_X1   g05229(.A1(new_n5484_), .A2(new_n5485_), .B(new_n760_), .ZN(new_n5486_));
  NAND2_X1   g05230(.A1(new_n3565_), .A2(new_n5486_), .ZN(new_n5487_));
  XOR2_X1    g05231(.A1(new_n5487_), .A2(\a[14] ), .Z(new_n5488_));
  INV_X1     g05232(.I(new_n5488_), .ZN(new_n5489_));
  XOR2_X1    g05233(.A1(new_n5483_), .A2(new_n5489_), .Z(new_n5490_));
  INV_X1     g05234(.I(new_n5490_), .ZN(new_n5491_));
  NAND2_X1   g05235(.A1(new_n5316_), .A2(new_n5321_), .ZN(new_n5492_));
  NAND2_X1   g05236(.A1(new_n5324_), .A2(new_n5322_), .ZN(new_n5493_));
  NAND2_X1   g05237(.A1(new_n5493_), .A2(new_n5492_), .ZN(new_n5494_));
  XOR2_X1    g05238(.A1(new_n5494_), .A2(new_n5491_), .Z(new_n5495_));
  OAI22_X1   g05239(.A1(new_n582_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n577_), .ZN(new_n5496_));
  NAND2_X1   g05240(.A1(new_n960_), .A2(\b[39] ), .ZN(new_n5497_));
  AOI21_X1   g05241(.A1(new_n5496_), .A2(new_n5497_), .B(new_n585_), .ZN(new_n5498_));
  NAND2_X1   g05242(.A1(new_n3996_), .A2(new_n5498_), .ZN(new_n5499_));
  XOR2_X1    g05243(.A1(new_n5499_), .A2(\a[11] ), .Z(new_n5500_));
  XNOR2_X1   g05244(.A1(new_n5495_), .A2(new_n5500_), .ZN(new_n5501_));
  NAND2_X1   g05245(.A1(new_n5325_), .A2(new_n5331_), .ZN(new_n5502_));
  XNOR2_X1   g05246(.A1(new_n5501_), .A2(new_n5502_), .ZN(new_n5503_));
  INV_X1     g05247(.I(new_n5503_), .ZN(new_n5504_));
  OAI22_X1   g05248(.A1(new_n437_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n431_), .ZN(new_n5505_));
  NAND2_X1   g05249(.A1(new_n775_), .A2(\b[42] ), .ZN(new_n5506_));
  AOI21_X1   g05250(.A1(new_n5505_), .A2(new_n5506_), .B(new_n440_), .ZN(new_n5507_));
  NAND2_X1   g05251(.A1(new_n4500_), .A2(new_n5507_), .ZN(new_n5508_));
  XOR2_X1    g05252(.A1(new_n5508_), .A2(\a[8] ), .Z(new_n5509_));
  NOR2_X1    g05253(.A1(new_n5504_), .A2(new_n5509_), .ZN(new_n5510_));
  INV_X1     g05254(.I(new_n5510_), .ZN(new_n5511_));
  NAND2_X1   g05255(.A1(new_n5504_), .A2(new_n5509_), .ZN(new_n5512_));
  NAND2_X1   g05256(.A1(new_n5511_), .A2(new_n5512_), .ZN(new_n5513_));
  XOR2_X1    g05257(.A1(new_n5503_), .A2(new_n5509_), .Z(new_n5514_));
  NOR2_X1    g05258(.A1(new_n5514_), .A2(new_n5354_), .ZN(new_n5515_));
  AOI21_X1   g05259(.A1(new_n5354_), .A2(new_n5513_), .B(new_n5515_), .ZN(new_n5516_));
  OAI22_X1   g05260(.A1(new_n364_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n320_), .ZN(new_n5517_));
  NAND2_X1   g05261(.A1(new_n594_), .A2(\b[45] ), .ZN(new_n5518_));
  AOI21_X1   g05262(.A1(new_n5517_), .A2(new_n5518_), .B(new_n312_), .ZN(new_n5519_));
  NAND2_X1   g05263(.A1(new_n5004_), .A2(new_n5519_), .ZN(new_n5520_));
  XOR2_X1    g05264(.A1(new_n5520_), .A2(\a[5] ), .Z(new_n5521_));
  NOR2_X1    g05265(.A1(new_n5338_), .A2(new_n5208_), .ZN(new_n5522_));
  NOR2_X1    g05266(.A1(new_n5162_), .A2(new_n5167_), .ZN(new_n5523_));
  NOR2_X1    g05267(.A1(new_n5523_), .A2(new_n5348_), .ZN(new_n5524_));
  NAND2_X1   g05268(.A1(new_n5210_), .A2(new_n5524_), .ZN(new_n5525_));
  NOR2_X1    g05269(.A1(new_n5525_), .A2(new_n5522_), .ZN(new_n5526_));
  XOR2_X1    g05270(.A1(new_n5526_), .A2(new_n5521_), .Z(new_n5527_));
  XOR2_X1    g05271(.A1(new_n5527_), .A2(new_n5516_), .Z(new_n5528_));
  OAI21_X1   g05272(.A1(new_n4997_), .A2(new_n5197_), .B(new_n5178_), .ZN(new_n5529_));
  NAND3_X1   g05273(.A1(new_n5170_), .A2(new_n5171_), .A3(new_n5529_), .ZN(new_n5530_));
  OAI21_X1   g05274(.A1(\b[47] ), .A2(\b[49] ), .B(\b[48] ), .ZN(new_n5531_));
  NAND2_X1   g05275(.A1(new_n5530_), .A2(new_n5531_), .ZN(new_n5532_));
  XNOR2_X1   g05276(.A1(\b[49] ), .A2(\b[50] ), .ZN(new_n5533_));
  INV_X1     g05277(.I(new_n5533_), .ZN(new_n5534_));
  NAND2_X1   g05278(.A1(new_n5532_), .A2(new_n5534_), .ZN(new_n5535_));
  XOR2_X1    g05279(.A1(\b[49] ), .A2(\b[50] ), .Z(new_n5536_));
  OAI21_X1   g05280(.A1(new_n5532_), .A2(new_n5536_), .B(new_n5535_), .ZN(new_n5537_));
  INV_X1     g05281(.I(\b[50] ), .ZN(new_n5538_));
  OAI22_X1   g05282(.A1(new_n405_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n404_), .ZN(new_n5539_));
  NAND2_X1   g05283(.A1(new_n279_), .A2(\b[48] ), .ZN(new_n5540_));
  AOI21_X1   g05284(.A1(new_n5539_), .A2(new_n5540_), .B(new_n264_), .ZN(new_n5541_));
  NAND2_X1   g05285(.A1(new_n5537_), .A2(new_n5541_), .ZN(new_n5542_));
  XOR2_X1    g05286(.A1(new_n5542_), .A2(\a[2] ), .Z(new_n5543_));
  INV_X1     g05287(.I(new_n5543_), .ZN(new_n5544_));
  XOR2_X1    g05288(.A1(new_n5528_), .A2(new_n5544_), .Z(new_n5545_));
  NAND2_X1   g05289(.A1(new_n5352_), .A2(new_n5545_), .ZN(new_n5546_));
  XOR2_X1    g05290(.A1(new_n5528_), .A2(new_n5544_), .Z(new_n5547_));
  OAI21_X1   g05291(.A1(new_n5352_), .A2(new_n5547_), .B(new_n5546_), .ZN(\f[50] ));
  INV_X1     g05292(.I(new_n5521_), .ZN(new_n5549_));
  NOR2_X1    g05293(.A1(new_n5516_), .A2(new_n5549_), .ZN(new_n5550_));
  XOR2_X1    g05294(.A1(new_n5516_), .A2(new_n5549_), .Z(new_n5551_));
  NOR3_X1    g05295(.A1(new_n5525_), .A2(new_n5522_), .A3(new_n5551_), .ZN(new_n5552_));
  NOR2_X1    g05296(.A1(new_n5552_), .A2(new_n5550_), .ZN(new_n5553_));
  NAND2_X1   g05297(.A1(new_n5514_), .A2(new_n5354_), .ZN(new_n5554_));
  NAND2_X1   g05298(.A1(new_n5554_), .A2(new_n5512_), .ZN(new_n5555_));
  INV_X1     g05299(.I(new_n5371_), .ZN(new_n5556_));
  NOR2_X1    g05300(.A1(new_n5556_), .A2(new_n5397_), .ZN(new_n5557_));
  NOR2_X1    g05301(.A1(new_n5223_), .A2(\a[47] ), .ZN(new_n5558_));
  NOR2_X1    g05302(.A1(new_n4701_), .A2(\a[48] ), .ZN(new_n5559_));
  NOR4_X1    g05303(.A1(new_n5558_), .A2(new_n5559_), .A3(new_n5383_), .A4(new_n5384_), .ZN(new_n5560_));
  NOR3_X1    g05304(.A1(new_n5560_), .A2(new_n267_), .A3(new_n5386_), .ZN(new_n5561_));
  NOR2_X1    g05305(.A1(new_n295_), .A2(new_n296_), .ZN(new_n5562_));
  AOI21_X1   g05306(.A1(new_n289_), .A2(new_n291_), .B(new_n293_), .ZN(new_n5563_));
  OAI21_X1   g05307(.A1(new_n5563_), .A2(new_n5562_), .B(new_n5394_), .ZN(new_n5564_));
  NAND3_X1   g05308(.A1(new_n5025_), .A2(new_n5227_), .A3(\b[3] ), .ZN(new_n5565_));
  OAI21_X1   g05309(.A1(new_n5224_), .A2(new_n5222_), .B(\b[2] ), .ZN(new_n5566_));
  NAND2_X1   g05310(.A1(new_n5565_), .A2(new_n5566_), .ZN(new_n5567_));
  NOR3_X1    g05311(.A1(new_n5564_), .A2(new_n5567_), .A3(new_n5561_), .ZN(new_n5568_));
  NOR2_X1    g05312(.A1(new_n5568_), .A2(new_n5220_), .ZN(new_n5569_));
  NOR4_X1    g05313(.A1(new_n5564_), .A2(new_n5567_), .A3(new_n5561_), .A4(\a[50] ), .ZN(new_n5570_));
  XNOR2_X1   g05314(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n5571_));
  NOR2_X1    g05315(.A1(new_n5571_), .A2(new_n258_), .ZN(new_n5572_));
  INV_X1     g05316(.I(new_n5572_), .ZN(new_n5573_));
  NOR3_X1    g05317(.A1(new_n5569_), .A2(new_n5570_), .A3(new_n5573_), .ZN(new_n5574_));
  NAND4_X1   g05318(.A1(new_n298_), .A2(new_n5394_), .A3(new_n5565_), .A4(new_n5566_), .ZN(new_n5575_));
  OAI21_X1   g05319(.A1(new_n5575_), .A2(new_n5561_), .B(\a[50] ), .ZN(new_n5576_));
  NAND2_X1   g05320(.A1(new_n5387_), .A2(\b[1] ), .ZN(new_n5577_));
  AOI21_X1   g05321(.A1(new_n294_), .A2(new_n297_), .B(new_n5231_), .ZN(new_n5578_));
  NAND3_X1   g05322(.A1(new_n4701_), .A2(new_n5223_), .A3(\a[49] ), .ZN(new_n5579_));
  NAND3_X1   g05323(.A1(new_n5221_), .A2(\a[47] ), .A3(\a[48] ), .ZN(new_n5580_));
  NAND2_X1   g05324(.A1(new_n5579_), .A2(new_n5580_), .ZN(new_n5581_));
  NOR2_X1    g05325(.A1(new_n5372_), .A2(new_n5230_), .ZN(new_n5582_));
  AOI22_X1   g05326(.A1(new_n5582_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n5581_), .ZN(new_n5583_));
  NAND4_X1   g05327(.A1(new_n5578_), .A2(new_n5583_), .A3(new_n5577_), .A4(new_n5220_), .ZN(new_n5584_));
  AOI21_X1   g05328(.A1(new_n5576_), .A2(new_n5584_), .B(new_n5572_), .ZN(new_n5585_));
  NOR2_X1    g05329(.A1(new_n5574_), .A2(new_n5585_), .ZN(new_n5586_));
  XOR2_X1    g05330(.A1(new_n5557_), .A2(new_n5586_), .Z(new_n5587_));
  INV_X1     g05331(.I(new_n4706_), .ZN(new_n5588_));
  AOI22_X1   g05332(.A1(\b[6] ), .A2(new_n4710_), .B1(new_n5588_), .B2(\b[5] ), .ZN(new_n5589_));
  NOR2_X1    g05333(.A1(new_n4873_), .A2(new_n393_), .ZN(new_n5590_));
  OAI21_X1   g05334(.A1(new_n5589_), .A2(new_n5590_), .B(new_n4713_), .ZN(new_n5591_));
  NOR2_X1    g05335(.A1(new_n524_), .A2(new_n5591_), .ZN(new_n5592_));
  XOR2_X1    g05336(.A1(new_n5592_), .A2(new_n4701_), .Z(new_n5593_));
  NOR2_X1    g05337(.A1(new_n5401_), .A2(new_n5235_), .ZN(new_n5594_));
  NAND2_X1   g05338(.A1(new_n5215_), .A2(new_n5594_), .ZN(new_n5595_));
  NAND2_X1   g05339(.A1(new_n5369_), .A2(new_n4701_), .ZN(new_n5596_));
  NOR2_X1    g05340(.A1(new_n5369_), .A2(new_n4701_), .ZN(new_n5597_));
  NOR3_X1    g05341(.A1(new_n5594_), .A2(new_n5398_), .A3(new_n5597_), .ZN(new_n5598_));
  NAND4_X1   g05342(.A1(new_n5595_), .A2(new_n5400_), .A3(new_n5596_), .A4(new_n5598_), .ZN(new_n5599_));
  XOR2_X1    g05343(.A1(new_n5599_), .A2(new_n5593_), .Z(new_n5600_));
  XNOR2_X1   g05344(.A1(new_n5600_), .A2(new_n5587_), .ZN(new_n5601_));
  OAI22_X1   g05345(.A1(new_n4208_), .A2(new_n510_), .B1(new_n495_), .B2(new_n4203_), .ZN(new_n5602_));
  NAND2_X1   g05346(.A1(new_n5244_), .A2(\b[7] ), .ZN(new_n5603_));
  AOI21_X1   g05347(.A1(new_n5602_), .A2(new_n5603_), .B(new_n4211_), .ZN(new_n5604_));
  NAND2_X1   g05348(.A1(new_n518_), .A2(new_n5604_), .ZN(new_n5605_));
  XOR2_X1    g05349(.A1(new_n5605_), .A2(\a[44] ), .Z(new_n5606_));
  INV_X1     g05350(.I(new_n5403_), .ZN(new_n5607_));
  NAND2_X1   g05351(.A1(new_n5607_), .A2(new_n5408_), .ZN(new_n5608_));
  NAND3_X1   g05352(.A1(new_n5409_), .A2(new_n5251_), .A3(new_n5608_), .ZN(new_n5609_));
  XOR2_X1    g05353(.A1(new_n5609_), .A2(new_n5606_), .Z(new_n5610_));
  XNOR2_X1   g05354(.A1(new_n5610_), .A2(new_n5601_), .ZN(new_n5611_));
  OAI22_X1   g05355(.A1(new_n3736_), .A2(new_n717_), .B1(new_n659_), .B2(new_n3731_), .ZN(new_n5612_));
  NAND2_X1   g05356(.A1(new_n4730_), .A2(\b[10] ), .ZN(new_n5613_));
  AOI21_X1   g05357(.A1(new_n5612_), .A2(new_n5613_), .B(new_n3739_), .ZN(new_n5614_));
  NAND2_X1   g05358(.A1(new_n716_), .A2(new_n5614_), .ZN(new_n5615_));
  XOR2_X1    g05359(.A1(new_n5615_), .A2(\a[41] ), .Z(new_n5616_));
  NAND2_X1   g05360(.A1(new_n5410_), .A2(new_n5415_), .ZN(new_n5617_));
  OAI21_X1   g05361(.A1(new_n5416_), .A2(new_n5366_), .B(new_n5617_), .ZN(new_n5618_));
  XOR2_X1    g05362(.A1(new_n5618_), .A2(new_n5616_), .Z(new_n5619_));
  XNOR2_X1   g05363(.A1(new_n5619_), .A2(new_n5611_), .ZN(new_n5620_));
  OAI22_X1   g05364(.A1(new_n3298_), .A2(new_n904_), .B1(new_n848_), .B2(new_n3293_), .ZN(new_n5621_));
  NAND2_X1   g05365(.A1(new_n4227_), .A2(\b[13] ), .ZN(new_n5622_));
  AOI21_X1   g05366(.A1(new_n5621_), .A2(new_n5622_), .B(new_n3301_), .ZN(new_n5623_));
  NAND2_X1   g05367(.A1(new_n907_), .A2(new_n5623_), .ZN(new_n5624_));
  XOR2_X1    g05368(.A1(new_n5624_), .A2(new_n3288_), .Z(new_n5625_));
  XOR2_X1    g05369(.A1(new_n5416_), .A2(new_n5366_), .Z(new_n5626_));
  NAND2_X1   g05370(.A1(new_n5626_), .A2(new_n5421_), .ZN(new_n5627_));
  NAND2_X1   g05371(.A1(new_n5627_), .A2(new_n5265_), .ZN(new_n5628_));
  NOR2_X1    g05372(.A1(new_n5425_), .A2(new_n5628_), .ZN(new_n5629_));
  XOR2_X1    g05373(.A1(new_n5629_), .A2(new_n5625_), .Z(new_n5630_));
  XNOR2_X1   g05374(.A1(new_n5630_), .A2(new_n5620_), .ZN(new_n5631_));
  OAI22_X1   g05375(.A1(new_n2846_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n2841_), .ZN(new_n5632_));
  NAND2_X1   g05376(.A1(new_n3755_), .A2(\b[16] ), .ZN(new_n5633_));
  AOI21_X1   g05377(.A1(new_n5632_), .A2(new_n5633_), .B(new_n2849_), .ZN(new_n5634_));
  NAND2_X1   g05378(.A1(new_n1123_), .A2(new_n5634_), .ZN(new_n5635_));
  XOR2_X1    g05379(.A1(new_n5635_), .A2(\a[35] ), .Z(new_n5636_));
  INV_X1     g05380(.I(new_n5426_), .ZN(new_n5637_));
  NAND2_X1   g05381(.A1(new_n5637_), .A2(new_n5431_), .ZN(new_n5638_));
  NAND3_X1   g05382(.A1(new_n5432_), .A2(new_n5638_), .A3(new_n5433_), .ZN(new_n5639_));
  XOR2_X1    g05383(.A1(new_n5639_), .A2(new_n5636_), .Z(new_n5640_));
  XNOR2_X1   g05384(.A1(new_n5640_), .A2(new_n5631_), .ZN(new_n5641_));
  OAI22_X1   g05385(.A1(new_n2452_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n2447_), .ZN(new_n5642_));
  NAND2_X1   g05386(.A1(new_n3312_), .A2(\b[19] ), .ZN(new_n5643_));
  AOI21_X1   g05387(.A1(new_n5642_), .A2(new_n5643_), .B(new_n2455_), .ZN(new_n5644_));
  NAND2_X1   g05388(.A1(new_n1396_), .A2(new_n5644_), .ZN(new_n5645_));
  XOR2_X1    g05389(.A1(new_n5645_), .A2(new_n2442_), .Z(new_n5646_));
  INV_X1     g05390(.I(new_n5434_), .ZN(new_n5647_));
  NOR2_X1    g05391(.A1(new_n5647_), .A2(new_n5440_), .ZN(new_n5648_));
  NOR3_X1    g05392(.A1(new_n5441_), .A2(new_n5648_), .A3(new_n5442_), .ZN(new_n5649_));
  XOR2_X1    g05393(.A1(new_n5649_), .A2(new_n5646_), .Z(new_n5650_));
  XNOR2_X1   g05394(.A1(new_n5650_), .A2(new_n5641_), .ZN(new_n5651_));
  OAI22_X1   g05395(.A1(new_n2084_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n2079_), .ZN(new_n5652_));
  NAND2_X1   g05396(.A1(new_n2864_), .A2(\b[22] ), .ZN(new_n5653_));
  AOI21_X1   g05397(.A1(new_n5652_), .A2(new_n5653_), .B(new_n2087_), .ZN(new_n5654_));
  NAND2_X1   g05398(.A1(new_n1708_), .A2(new_n5654_), .ZN(new_n5655_));
  XOR2_X1    g05399(.A1(new_n5655_), .A2(\a[29] ), .Z(new_n5656_));
  INV_X1     g05400(.I(new_n5364_), .ZN(new_n5657_));
  NAND2_X1   g05401(.A1(new_n5443_), .A2(new_n5364_), .ZN(new_n5658_));
  OR2_X2     g05402(.A1(new_n5443_), .A2(new_n5364_), .Z(new_n5659_));
  NAND3_X1   g05403(.A1(new_n5659_), .A2(new_n5365_), .A3(new_n5658_), .ZN(new_n5660_));
  OAI21_X1   g05404(.A1(new_n5657_), .A2(new_n5443_), .B(new_n5660_), .ZN(new_n5661_));
  XOR2_X1    g05405(.A1(new_n5661_), .A2(new_n5656_), .Z(new_n5662_));
  XNOR2_X1   g05406(.A1(new_n5662_), .A2(new_n5651_), .ZN(new_n5663_));
  OAI22_X1   g05407(.A1(new_n1760_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n1755_), .ZN(new_n5664_));
  NAND2_X1   g05408(.A1(new_n2470_), .A2(\b[25] ), .ZN(new_n5665_));
  AOI21_X1   g05409(.A1(new_n5664_), .A2(new_n5665_), .B(new_n1763_), .ZN(new_n5666_));
  NAND2_X1   g05410(.A1(new_n2042_), .A2(new_n5666_), .ZN(new_n5667_));
  XOR2_X1    g05411(.A1(new_n5667_), .A2(new_n1750_), .Z(new_n5668_));
  XOR2_X1    g05412(.A1(new_n5443_), .A2(new_n5364_), .Z(new_n5669_));
  XOR2_X1    g05413(.A1(new_n5669_), .A2(new_n5365_), .Z(new_n5670_));
  AOI22_X1   g05414(.A1(new_n5446_), .A2(new_n5447_), .B1(new_n5359_), .B2(new_n5670_), .ZN(new_n5671_));
  XOR2_X1    g05415(.A1(new_n5671_), .A2(new_n5668_), .Z(new_n5672_));
  XNOR2_X1   g05416(.A1(new_n5672_), .A2(new_n5663_), .ZN(new_n5673_));
  OAI22_X1   g05417(.A1(new_n1444_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n1439_), .ZN(new_n5674_));
  NAND2_X1   g05418(.A1(new_n2098_), .A2(\b[28] ), .ZN(new_n5675_));
  AOI21_X1   g05419(.A1(new_n5674_), .A2(new_n5675_), .B(new_n1447_), .ZN(new_n5676_));
  NAND2_X1   g05420(.A1(new_n2404_), .A2(new_n5676_), .ZN(new_n5677_));
  XOR2_X1    g05421(.A1(new_n5677_), .A2(\a[23] ), .Z(new_n5678_));
  INV_X1     g05422(.I(new_n5453_), .ZN(new_n5679_));
  OAI21_X1   g05423(.A1(new_n5448_), .A2(new_n5679_), .B(new_n5457_), .ZN(new_n5680_));
  XNOR2_X1   g05424(.A1(new_n5680_), .A2(new_n5678_), .ZN(new_n5681_));
  XOR2_X1    g05425(.A1(new_n5681_), .A2(new_n5673_), .Z(new_n5682_));
  OAI22_X1   g05426(.A1(new_n1168_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n1163_), .ZN(new_n5683_));
  NAND2_X1   g05427(.A1(new_n1774_), .A2(\b[31] ), .ZN(new_n5684_));
  AOI21_X1   g05428(.A1(new_n5683_), .A2(new_n5684_), .B(new_n1171_), .ZN(new_n5685_));
  NAND2_X1   g05429(.A1(new_n2797_), .A2(new_n5685_), .ZN(new_n5686_));
  XOR2_X1    g05430(.A1(new_n5686_), .A2(\a[20] ), .Z(new_n5687_));
  OAI21_X1   g05431(.A1(new_n5458_), .A2(new_n5459_), .B(new_n5465_), .ZN(new_n5688_));
  OAI21_X1   g05432(.A1(new_n5469_), .A2(new_n5466_), .B(new_n5688_), .ZN(new_n5689_));
  XOR2_X1    g05433(.A1(new_n5689_), .A2(new_n5687_), .Z(new_n5690_));
  XNOR2_X1   g05434(.A1(new_n5690_), .A2(new_n5682_), .ZN(new_n5691_));
  OAI22_X1   g05435(.A1(new_n940_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n935_), .ZN(new_n5692_));
  NAND2_X1   g05436(.A1(new_n1458_), .A2(\b[34] ), .ZN(new_n5693_));
  AOI21_X1   g05437(.A1(new_n5692_), .A2(new_n5693_), .B(new_n943_), .ZN(new_n5694_));
  NAND2_X1   g05438(.A1(new_n3246_), .A2(new_n5694_), .ZN(new_n5695_));
  XOR2_X1    g05439(.A1(new_n5695_), .A2(\a[17] ), .Z(new_n5696_));
  NOR3_X1    g05440(.A1(new_n5479_), .A2(new_n5477_), .A3(new_n5482_), .ZN(new_n5697_));
  XOR2_X1    g05441(.A1(new_n5697_), .A2(new_n5696_), .Z(new_n5698_));
  XOR2_X1    g05442(.A1(new_n5698_), .A2(new_n5691_), .Z(new_n5699_));
  OAI22_X1   g05443(.A1(new_n757_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n752_), .ZN(new_n5700_));
  NAND2_X1   g05444(.A1(new_n1182_), .A2(\b[37] ), .ZN(new_n5701_));
  AOI21_X1   g05445(.A1(new_n5700_), .A2(new_n5701_), .B(new_n760_), .ZN(new_n5702_));
  NAND2_X1   g05446(.A1(new_n3700_), .A2(new_n5702_), .ZN(new_n5703_));
  XOR2_X1    g05447(.A1(new_n5703_), .A2(\a[14] ), .Z(new_n5704_));
  NOR2_X1    g05448(.A1(new_n5483_), .A2(new_n5489_), .ZN(new_n5705_));
  NOR2_X1    g05449(.A1(new_n5491_), .A2(new_n5705_), .ZN(new_n5706_));
  NAND2_X1   g05450(.A1(new_n5494_), .A2(new_n5706_), .ZN(new_n5707_));
  XOR2_X1    g05451(.A1(new_n5707_), .A2(new_n5704_), .Z(new_n5708_));
  XNOR2_X1   g05452(.A1(new_n5708_), .A2(new_n5699_), .ZN(new_n5709_));
  OAI22_X1   g05453(.A1(new_n582_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n577_), .ZN(new_n5710_));
  NAND2_X1   g05454(.A1(new_n960_), .A2(\b[40] ), .ZN(new_n5711_));
  AOI21_X1   g05455(.A1(new_n5710_), .A2(new_n5711_), .B(new_n585_), .ZN(new_n5712_));
  NAND2_X1   g05456(.A1(new_n4017_), .A2(new_n5712_), .ZN(new_n5713_));
  XOR2_X1    g05457(.A1(new_n5713_), .A2(\a[11] ), .Z(new_n5714_));
  INV_X1     g05458(.I(new_n5495_), .ZN(new_n5715_));
  NAND2_X1   g05459(.A1(new_n5715_), .A2(new_n5500_), .ZN(new_n5716_));
  NAND3_X1   g05460(.A1(new_n5501_), .A2(new_n5716_), .A3(new_n5502_), .ZN(new_n5717_));
  XOR2_X1    g05461(.A1(new_n5717_), .A2(new_n5714_), .Z(new_n5718_));
  XNOR2_X1   g05462(.A1(new_n5718_), .A2(new_n5709_), .ZN(new_n5719_));
  OAI22_X1   g05463(.A1(new_n437_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n431_), .ZN(new_n5720_));
  NAND2_X1   g05464(.A1(new_n775_), .A2(\b[43] ), .ZN(new_n5721_));
  AOI21_X1   g05465(.A1(new_n5720_), .A2(new_n5721_), .B(new_n440_), .ZN(new_n5722_));
  NAND2_X1   g05466(.A1(new_n4513_), .A2(new_n5722_), .ZN(new_n5723_));
  XOR2_X1    g05467(.A1(new_n5723_), .A2(\a[8] ), .Z(new_n5724_));
  XNOR2_X1   g05468(.A1(new_n5719_), .A2(new_n5724_), .ZN(new_n5725_));
  OAI22_X1   g05469(.A1(new_n364_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n320_), .ZN(new_n5726_));
  NAND2_X1   g05470(.A1(new_n594_), .A2(\b[46] ), .ZN(new_n5727_));
  AOI21_X1   g05471(.A1(new_n5726_), .A2(new_n5727_), .B(new_n312_), .ZN(new_n5728_));
  NAND2_X1   g05472(.A1(new_n5177_), .A2(new_n5728_), .ZN(new_n5729_));
  XOR2_X1    g05473(.A1(new_n5729_), .A2(\a[5] ), .Z(new_n5730_));
  INV_X1     g05474(.I(new_n5730_), .ZN(new_n5731_));
  XOR2_X1    g05475(.A1(new_n5725_), .A2(new_n5731_), .Z(new_n5732_));
  NOR2_X1    g05476(.A1(new_n5732_), .A2(new_n5555_), .ZN(new_n5733_));
  INV_X1     g05477(.I(new_n5555_), .ZN(new_n5734_));
  XOR2_X1    g05478(.A1(new_n5725_), .A2(new_n5730_), .Z(new_n5735_));
  NOR2_X1    g05479(.A1(new_n5735_), .A2(new_n5734_), .ZN(new_n5736_));
  NOR2_X1    g05480(.A1(new_n5733_), .A2(new_n5736_), .ZN(new_n5737_));
  INV_X1     g05481(.I(\b[51] ), .ZN(new_n5738_));
  XOR2_X1    g05482(.A1(new_n5532_), .A2(\b[49] ), .Z(new_n5739_));
  NAND2_X1   g05483(.A1(new_n5739_), .A2(new_n5534_), .ZN(new_n5740_));
  XOR2_X1    g05484(.A1(new_n5740_), .A2(new_n5738_), .Z(new_n5741_));
  NAND2_X1   g05485(.A1(new_n283_), .A2(\b[51] ), .ZN(new_n5742_));
  NAND2_X1   g05486(.A1(new_n279_), .A2(\b[49] ), .ZN(new_n5743_));
  AOI21_X1   g05487(.A1(\b[50] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n5744_));
  NAND4_X1   g05488(.A1(new_n5741_), .A2(new_n5742_), .A3(new_n5743_), .A4(new_n5744_), .ZN(new_n5745_));
  XOR2_X1    g05489(.A1(new_n5745_), .A2(\a[2] ), .Z(new_n5746_));
  XOR2_X1    g05490(.A1(new_n5737_), .A2(new_n5746_), .Z(new_n5747_));
  XOR2_X1    g05491(.A1(new_n5737_), .A2(new_n5746_), .Z(new_n5748_));
  NAND2_X1   g05492(.A1(new_n5553_), .A2(new_n5748_), .ZN(new_n5749_));
  OAI21_X1   g05493(.A1(new_n5553_), .A2(new_n5747_), .B(new_n5749_), .ZN(new_n5750_));
  XOR2_X1    g05494(.A1(new_n5352_), .A2(new_n5544_), .Z(new_n5751_));
  NAND2_X1   g05495(.A1(new_n5751_), .A2(new_n5528_), .ZN(new_n5752_));
  XOR2_X1    g05496(.A1(new_n5752_), .A2(new_n5750_), .Z(new_n5753_));
  NAND2_X1   g05497(.A1(new_n5352_), .A2(new_n5544_), .ZN(new_n5754_));
  XOR2_X1    g05498(.A1(new_n5753_), .A2(new_n5754_), .Z(\f[51] ));
  INV_X1     g05499(.I(new_n5553_), .ZN(new_n5756_));
  XOR2_X1    g05500(.A1(new_n5725_), .A2(new_n5734_), .Z(new_n5757_));
  NOR3_X1    g05501(.A1(new_n5756_), .A2(new_n5731_), .A3(new_n5757_), .ZN(new_n5758_));
  AOI21_X1   g05502(.A1(new_n5756_), .A2(new_n5731_), .B(new_n5758_), .ZN(new_n5759_));
  XOR2_X1    g05503(.A1(new_n5691_), .A2(new_n5696_), .Z(new_n5760_));
  NAND2_X1   g05504(.A1(new_n5760_), .A2(new_n5696_), .ZN(new_n5761_));
  NAND2_X1   g05505(.A1(new_n5760_), .A2(new_n5697_), .ZN(new_n5762_));
  XOR2_X1    g05506(.A1(new_n5673_), .A2(new_n5678_), .Z(new_n5763_));
  NAND2_X1   g05507(.A1(new_n5763_), .A2(new_n5678_), .ZN(new_n5764_));
  INV_X1     g05508(.I(new_n5680_), .ZN(new_n5765_));
  NAND2_X1   g05509(.A1(new_n5763_), .A2(new_n5765_), .ZN(new_n5766_));
  NAND2_X1   g05510(.A1(new_n5582_), .A2(\b[4] ), .ZN(new_n5767_));
  NAND2_X1   g05511(.A1(new_n5581_), .A2(\b[3] ), .ZN(new_n5768_));
  AOI22_X1   g05512(.A1(new_n5767_), .A2(new_n5768_), .B1(\b[2] ), .B2(new_n5387_), .ZN(new_n5769_));
  OAI21_X1   g05513(.A1(new_n424_), .A2(new_n5231_), .B(new_n5769_), .ZN(new_n5770_));
  INV_X1     g05514(.I(new_n5770_), .ZN(new_n5771_));
  NOR3_X1    g05515(.A1(new_n5388_), .A2(\a[50] ), .A3(new_n5395_), .ZN(new_n5772_));
  AOI21_X1   g05516(.A1(new_n5379_), .A2(new_n5380_), .B(new_n5220_), .ZN(new_n5773_));
  NOR2_X1    g05517(.A1(new_n5773_), .A2(new_n5772_), .ZN(new_n5774_));
  NAND3_X1   g05518(.A1(new_n5576_), .A2(new_n5584_), .A3(new_n5572_), .ZN(new_n5775_));
  OAI21_X1   g05519(.A1(new_n5569_), .A2(new_n5570_), .B(new_n5573_), .ZN(new_n5776_));
  NAND3_X1   g05520(.A1(new_n5776_), .A2(new_n5775_), .A3(new_n5774_), .ZN(new_n5777_));
  NOR3_X1    g05521(.A1(new_n5569_), .A2(new_n5570_), .A3(new_n5573_), .ZN(new_n5778_));
  INV_X1     g05522(.I(new_n5778_), .ZN(new_n5779_));
  AOI21_X1   g05523(.A1(new_n5777_), .A2(new_n5556_), .B(new_n5779_), .ZN(new_n5780_));
  NOR3_X1    g05524(.A1(new_n5574_), .A2(new_n5585_), .A3(new_n5397_), .ZN(new_n5781_));
  NOR3_X1    g05525(.A1(new_n5781_), .A2(new_n5371_), .A3(new_n5778_), .ZN(new_n5782_));
  INV_X1     g05526(.I(\a[53] ), .ZN(new_n5783_));
  XOR2_X1    g05527(.A1(\a[50] ), .A2(\a[51] ), .Z(new_n5784_));
  XNOR2_X1   g05528(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n5785_));
  NAND2_X1   g05529(.A1(new_n5785_), .A2(new_n5784_), .ZN(new_n5786_));
  NOR2_X1    g05530(.A1(new_n5786_), .A2(new_n267_), .ZN(new_n5787_));
  INV_X1     g05531(.I(\a[52] ), .ZN(new_n5788_));
  NOR3_X1    g05532(.A1(new_n5788_), .A2(\a[50] ), .A3(\a[51] ), .ZN(new_n5789_));
  NAND2_X1   g05533(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n5790_));
  NOR2_X1    g05534(.A1(new_n5790_), .A2(\a[52] ), .ZN(new_n5791_));
  NOR2_X1    g05535(.A1(new_n5791_), .A2(new_n5789_), .ZN(new_n5792_));
  NOR2_X1    g05536(.A1(new_n5792_), .A2(new_n258_), .ZN(new_n5793_));
  XNOR2_X1   g05537(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n5794_));
  NOR2_X1    g05538(.A1(new_n5571_), .A2(new_n5794_), .ZN(new_n5795_));
  INV_X1     g05539(.I(new_n5795_), .ZN(new_n5796_));
  NOR4_X1    g05540(.A1(new_n5787_), .A2(new_n5796_), .A3(new_n261_), .A4(new_n5793_), .ZN(new_n5797_));
  XOR2_X1    g05541(.A1(new_n5797_), .A2(new_n5783_), .Z(new_n5798_));
  NAND2_X1   g05542(.A1(new_n5573_), .A2(\a[53] ), .ZN(new_n5799_));
  XOR2_X1    g05543(.A1(new_n5798_), .A2(new_n5799_), .Z(new_n5800_));
  NOR3_X1    g05544(.A1(new_n5800_), .A2(new_n5780_), .A3(new_n5782_), .ZN(new_n5801_));
  NOR2_X1    g05545(.A1(new_n5782_), .A2(new_n5780_), .ZN(new_n5802_));
  XNOR2_X1   g05546(.A1(new_n5798_), .A2(new_n5799_), .ZN(new_n5803_));
  NOR2_X1    g05547(.A1(new_n5802_), .A2(new_n5803_), .ZN(new_n5804_));
  OAI21_X1   g05548(.A1(new_n5804_), .A2(new_n5801_), .B(new_n5220_), .ZN(new_n5805_));
  NAND2_X1   g05549(.A1(new_n5802_), .A2(new_n5803_), .ZN(new_n5806_));
  OAI21_X1   g05550(.A1(new_n5780_), .A2(new_n5782_), .B(new_n5800_), .ZN(new_n5807_));
  NAND3_X1   g05551(.A1(new_n5806_), .A2(new_n5807_), .A3(\a[50] ), .ZN(new_n5808_));
  AOI21_X1   g05552(.A1(new_n5805_), .A2(new_n5808_), .B(new_n5771_), .ZN(new_n5809_));
  AOI21_X1   g05553(.A1(new_n5806_), .A2(new_n5807_), .B(\a[50] ), .ZN(new_n5810_));
  NOR3_X1    g05554(.A1(new_n5804_), .A2(new_n5801_), .A3(new_n5220_), .ZN(new_n5811_));
  NOR3_X1    g05555(.A1(new_n5811_), .A2(new_n5810_), .A3(new_n5770_), .ZN(new_n5812_));
  OAI22_X1   g05556(.A1(new_n4711_), .A2(new_n450_), .B1(new_n403_), .B2(new_n4706_), .ZN(new_n5813_));
  INV_X1     g05557(.I(new_n4873_), .ZN(new_n5814_));
  NAND2_X1   g05558(.A1(new_n5814_), .A2(\b[5] ), .ZN(new_n5815_));
  AOI21_X1   g05559(.A1(new_n5813_), .A2(new_n5815_), .B(new_n4714_), .ZN(new_n5816_));
  NAND2_X1   g05560(.A1(new_n454_), .A2(new_n5816_), .ZN(new_n5817_));
  XOR2_X1    g05561(.A1(new_n5817_), .A2(\a[47] ), .Z(new_n5818_));
  NOR3_X1    g05562(.A1(new_n5812_), .A2(new_n5809_), .A3(new_n5818_), .ZN(new_n5819_));
  OAI21_X1   g05563(.A1(new_n5811_), .A2(new_n5810_), .B(new_n5770_), .ZN(new_n5820_));
  NAND3_X1   g05564(.A1(new_n5805_), .A2(new_n5808_), .A3(new_n5771_), .ZN(new_n5821_));
  INV_X1     g05565(.I(new_n5818_), .ZN(new_n5822_));
  AOI21_X1   g05566(.A1(new_n5820_), .A2(new_n5821_), .B(new_n5822_), .ZN(new_n5823_));
  NOR2_X1    g05567(.A1(new_n5823_), .A2(new_n5819_), .ZN(new_n5824_));
  OAI22_X1   g05568(.A1(new_n4208_), .A2(new_n617_), .B1(new_n510_), .B2(new_n4203_), .ZN(new_n5825_));
  NAND2_X1   g05569(.A1(new_n5244_), .A2(\b[8] ), .ZN(new_n5826_));
  AOI21_X1   g05570(.A1(new_n5825_), .A2(new_n5826_), .B(new_n4211_), .ZN(new_n5827_));
  NAND2_X1   g05571(.A1(new_n616_), .A2(new_n5827_), .ZN(new_n5828_));
  XOR2_X1    g05572(.A1(new_n5828_), .A2(\a[44] ), .Z(new_n5829_));
  NOR2_X1    g05573(.A1(new_n5824_), .A2(new_n5829_), .ZN(new_n5830_));
  INV_X1     g05574(.I(new_n5824_), .ZN(new_n5831_));
  INV_X1     g05575(.I(new_n5829_), .ZN(new_n5832_));
  NOR2_X1    g05576(.A1(new_n5831_), .A2(new_n5832_), .ZN(new_n5833_));
  NOR2_X1    g05577(.A1(new_n5833_), .A2(new_n5830_), .ZN(new_n5834_));
  INV_X1     g05578(.I(new_n5834_), .ZN(new_n5835_));
  OAI22_X1   g05579(.A1(new_n3736_), .A2(new_n795_), .B1(new_n717_), .B2(new_n3731_), .ZN(new_n5836_));
  NAND2_X1   g05580(.A1(new_n4730_), .A2(\b[11] ), .ZN(new_n5837_));
  AOI21_X1   g05581(.A1(new_n5836_), .A2(new_n5837_), .B(new_n3739_), .ZN(new_n5838_));
  AND3_X2    g05582(.A1(new_n799_), .A2(new_n3726_), .A3(new_n5838_), .Z(new_n5839_));
  AOI21_X1   g05583(.A1(new_n799_), .A2(new_n5838_), .B(new_n3726_), .ZN(new_n5840_));
  NOR2_X1    g05584(.A1(new_n5839_), .A2(new_n5840_), .ZN(new_n5841_));
  NOR2_X1    g05585(.A1(new_n5835_), .A2(new_n5841_), .ZN(new_n5842_));
  INV_X1     g05586(.I(new_n5841_), .ZN(new_n5843_));
  NOR2_X1    g05587(.A1(new_n5843_), .A2(new_n5834_), .ZN(new_n5844_));
  NOR2_X1    g05588(.A1(new_n5842_), .A2(new_n5844_), .ZN(new_n5845_));
  INV_X1     g05589(.I(new_n5845_), .ZN(new_n5846_));
  OAI22_X1   g05590(.A1(new_n3298_), .A2(new_n992_), .B1(new_n904_), .B2(new_n3293_), .ZN(new_n5847_));
  NAND2_X1   g05591(.A1(new_n4227_), .A2(\b[14] ), .ZN(new_n5848_));
  AOI21_X1   g05592(.A1(new_n5847_), .A2(new_n5848_), .B(new_n3301_), .ZN(new_n5849_));
  NAND2_X1   g05593(.A1(new_n991_), .A2(new_n5849_), .ZN(new_n5850_));
  XOR2_X1    g05594(.A1(new_n5850_), .A2(\a[38] ), .Z(new_n5851_));
  INV_X1     g05595(.I(new_n5851_), .ZN(new_n5852_));
  NAND2_X1   g05596(.A1(new_n5846_), .A2(new_n5852_), .ZN(new_n5853_));
  NOR2_X1    g05597(.A1(new_n5846_), .A2(new_n5852_), .ZN(new_n5854_));
  INV_X1     g05598(.I(new_n5854_), .ZN(new_n5855_));
  AND2_X2    g05599(.A1(new_n5855_), .A2(new_n5853_), .Z(new_n5856_));
  OAI22_X1   g05600(.A1(new_n2846_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n2841_), .ZN(new_n5857_));
  NAND2_X1   g05601(.A1(new_n3755_), .A2(\b[17] ), .ZN(new_n5858_));
  AOI21_X1   g05602(.A1(new_n5857_), .A2(new_n5858_), .B(new_n2849_), .ZN(new_n5859_));
  NAND2_X1   g05603(.A1(new_n1225_), .A2(new_n5859_), .ZN(new_n5860_));
  XOR2_X1    g05604(.A1(new_n5860_), .A2(\a[35] ), .Z(new_n5861_));
  XOR2_X1    g05605(.A1(new_n5856_), .A2(new_n5861_), .Z(new_n5862_));
  OAI22_X1   g05606(.A1(new_n2452_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n2447_), .ZN(new_n5863_));
  NAND2_X1   g05607(.A1(new_n3312_), .A2(\b[20] ), .ZN(new_n5864_));
  AOI21_X1   g05608(.A1(new_n5863_), .A2(new_n5864_), .B(new_n2455_), .ZN(new_n5865_));
  NAND2_X1   g05609(.A1(new_n1517_), .A2(new_n5865_), .ZN(new_n5866_));
  XOR2_X1    g05610(.A1(new_n5866_), .A2(\a[32] ), .Z(new_n5867_));
  NOR2_X1    g05611(.A1(new_n5862_), .A2(new_n5867_), .ZN(new_n5868_));
  INV_X1     g05612(.I(new_n5868_), .ZN(new_n5869_));
  NAND2_X1   g05613(.A1(new_n5862_), .A2(new_n5867_), .ZN(new_n5870_));
  NAND2_X1   g05614(.A1(new_n5869_), .A2(new_n5870_), .ZN(new_n5871_));
  OAI22_X1   g05615(.A1(new_n2084_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n2079_), .ZN(new_n5872_));
  NAND2_X1   g05616(.A1(new_n2864_), .A2(\b[23] ), .ZN(new_n5873_));
  AOI21_X1   g05617(.A1(new_n5872_), .A2(new_n5873_), .B(new_n2087_), .ZN(new_n5874_));
  NAND2_X1   g05618(.A1(new_n1828_), .A2(new_n5874_), .ZN(new_n5875_));
  XOR2_X1    g05619(.A1(new_n5875_), .A2(\a[29] ), .Z(new_n5876_));
  AND2_X2    g05620(.A1(new_n5871_), .A2(new_n5876_), .Z(new_n5877_));
  NOR2_X1    g05621(.A1(new_n5871_), .A2(new_n5876_), .ZN(new_n5878_));
  NOR2_X1    g05622(.A1(new_n5877_), .A2(new_n5878_), .ZN(new_n5879_));
  OAI22_X1   g05623(.A1(new_n1760_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n1755_), .ZN(new_n5880_));
  NAND2_X1   g05624(.A1(new_n2470_), .A2(\b[26] ), .ZN(new_n5881_));
  AOI21_X1   g05625(.A1(new_n5880_), .A2(new_n5881_), .B(new_n1763_), .ZN(new_n5882_));
  NAND2_X1   g05626(.A1(new_n2174_), .A2(new_n5882_), .ZN(new_n5883_));
  XOR2_X1    g05627(.A1(new_n5883_), .A2(\a[26] ), .Z(new_n5884_));
  XOR2_X1    g05628(.A1(new_n5879_), .A2(new_n5884_), .Z(new_n5885_));
  OAI22_X1   g05629(.A1(new_n1444_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n1439_), .ZN(new_n5886_));
  NAND2_X1   g05630(.A1(new_n2098_), .A2(\b[29] ), .ZN(new_n5887_));
  AOI21_X1   g05631(.A1(new_n5886_), .A2(new_n5887_), .B(new_n1447_), .ZN(new_n5888_));
  NAND2_X1   g05632(.A1(new_n2546_), .A2(new_n5888_), .ZN(new_n5889_));
  XOR2_X1    g05633(.A1(new_n5889_), .A2(\a[23] ), .Z(new_n5890_));
  XNOR2_X1   g05634(.A1(new_n5890_), .A2(new_n5885_), .ZN(new_n5891_));
  OAI22_X1   g05635(.A1(new_n1168_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n1163_), .ZN(new_n5892_));
  NAND2_X1   g05636(.A1(new_n1774_), .A2(\b[32] ), .ZN(new_n5893_));
  AOI21_X1   g05637(.A1(new_n5892_), .A2(new_n5893_), .B(new_n1171_), .ZN(new_n5894_));
  NAND2_X1   g05638(.A1(new_n2963_), .A2(new_n5894_), .ZN(new_n5895_));
  XOR2_X1    g05639(.A1(new_n5895_), .A2(\a[20] ), .Z(new_n5896_));
  INV_X1     g05640(.I(new_n5896_), .ZN(new_n5897_));
  XOR2_X1    g05641(.A1(new_n5891_), .A2(new_n5897_), .Z(new_n5898_));
  AOI21_X1   g05642(.A1(new_n5764_), .A2(new_n5766_), .B(new_n5898_), .ZN(new_n5899_));
  NAND2_X1   g05643(.A1(new_n5766_), .A2(new_n5764_), .ZN(new_n5900_));
  XOR2_X1    g05644(.A1(new_n5891_), .A2(new_n5896_), .Z(new_n5901_));
  NOR2_X1    g05645(.A1(new_n5900_), .A2(new_n5901_), .ZN(new_n5902_));
  NOR2_X1    g05646(.A1(new_n5902_), .A2(new_n5899_), .ZN(new_n5903_));
  OAI22_X1   g05647(.A1(new_n940_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n935_), .ZN(new_n5904_));
  NAND2_X1   g05648(.A1(new_n1458_), .A2(\b[35] ), .ZN(new_n5905_));
  AOI21_X1   g05649(.A1(new_n5904_), .A2(new_n5905_), .B(new_n943_), .ZN(new_n5906_));
  NAND2_X1   g05650(.A1(new_n3411_), .A2(new_n5906_), .ZN(new_n5907_));
  XOR2_X1    g05651(.A1(new_n5907_), .A2(\a[17] ), .Z(new_n5908_));
  XOR2_X1    g05652(.A1(new_n5903_), .A2(new_n5908_), .Z(new_n5909_));
  OAI22_X1   g05653(.A1(new_n757_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n752_), .ZN(new_n5910_));
  NAND2_X1   g05654(.A1(new_n1182_), .A2(\b[38] ), .ZN(new_n5911_));
  AOI21_X1   g05655(.A1(new_n5910_), .A2(new_n5911_), .B(new_n760_), .ZN(new_n5912_));
  NAND2_X1   g05656(.A1(new_n3844_), .A2(new_n5912_), .ZN(new_n5913_));
  XOR2_X1    g05657(.A1(new_n5913_), .A2(\a[14] ), .Z(new_n5914_));
  XNOR2_X1   g05658(.A1(new_n5909_), .A2(new_n5914_), .ZN(new_n5915_));
  AOI21_X1   g05659(.A1(new_n5762_), .A2(new_n5761_), .B(new_n5915_), .ZN(new_n5916_));
  NAND2_X1   g05660(.A1(new_n5762_), .A2(new_n5761_), .ZN(new_n5917_));
  XOR2_X1    g05661(.A1(new_n5909_), .A2(new_n5914_), .Z(new_n5918_));
  NOR2_X1    g05662(.A1(new_n5917_), .A2(new_n5918_), .ZN(new_n5919_));
  NOR2_X1    g05663(.A1(new_n5919_), .A2(new_n5916_), .ZN(new_n5920_));
  OAI22_X1   g05664(.A1(new_n582_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n577_), .ZN(new_n5921_));
  NAND2_X1   g05665(.A1(new_n960_), .A2(\b[41] ), .ZN(new_n5922_));
  AOI21_X1   g05666(.A1(new_n5921_), .A2(new_n5922_), .B(new_n585_), .ZN(new_n5923_));
  NAND2_X1   g05667(.A1(new_n4320_), .A2(new_n5923_), .ZN(new_n5924_));
  XOR2_X1    g05668(.A1(new_n5924_), .A2(\a[11] ), .Z(new_n5925_));
  XOR2_X1    g05669(.A1(new_n5920_), .A2(new_n5925_), .Z(new_n5926_));
  OAI22_X1   g05670(.A1(new_n437_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n431_), .ZN(new_n5927_));
  NAND2_X1   g05671(.A1(new_n775_), .A2(\b[44] ), .ZN(new_n5928_));
  AOI21_X1   g05672(.A1(new_n5927_), .A2(new_n5928_), .B(new_n440_), .ZN(new_n5929_));
  NAND2_X1   g05673(.A1(new_n4833_), .A2(new_n5929_), .ZN(new_n5930_));
  XOR2_X1    g05674(.A1(new_n5930_), .A2(\a[8] ), .Z(new_n5931_));
  NOR2_X1    g05675(.A1(new_n5926_), .A2(new_n5931_), .ZN(new_n5932_));
  INV_X1     g05676(.I(new_n5932_), .ZN(new_n5933_));
  NAND2_X1   g05677(.A1(new_n5926_), .A2(new_n5931_), .ZN(new_n5934_));
  NAND2_X1   g05678(.A1(new_n5933_), .A2(new_n5934_), .ZN(new_n5935_));
  INV_X1     g05679(.I(new_n5935_), .ZN(new_n5936_));
  OAI22_X1   g05680(.A1(new_n364_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n320_), .ZN(new_n5937_));
  NAND2_X1   g05681(.A1(new_n594_), .A2(\b[47] ), .ZN(new_n5938_));
  AOI21_X1   g05682(.A1(new_n5937_), .A2(new_n5938_), .B(new_n312_), .ZN(new_n5939_));
  NAND2_X1   g05683(.A1(new_n5196_), .A2(new_n5939_), .ZN(new_n5940_));
  XOR2_X1    g05684(.A1(new_n5940_), .A2(\a[5] ), .Z(new_n5941_));
  INV_X1     g05685(.I(new_n5941_), .ZN(new_n5942_));
  NOR2_X1    g05686(.A1(new_n5936_), .A2(new_n5942_), .ZN(new_n5943_));
  NOR2_X1    g05687(.A1(new_n5935_), .A2(new_n5941_), .ZN(new_n5944_));
  NOR2_X1    g05688(.A1(new_n5943_), .A2(new_n5944_), .ZN(new_n5945_));
  OAI21_X1   g05689(.A1(new_n5197_), .A2(new_n5738_), .B(new_n5538_), .ZN(new_n5946_));
  NAND3_X1   g05690(.A1(new_n5530_), .A2(new_n5531_), .A3(new_n5946_), .ZN(new_n5947_));
  OAI21_X1   g05691(.A1(\b[49] ), .A2(\b[51] ), .B(\b[50] ), .ZN(new_n5948_));
  NAND2_X1   g05692(.A1(new_n5947_), .A2(new_n5948_), .ZN(new_n5949_));
  XNOR2_X1   g05693(.A1(\b[51] ), .A2(\b[52] ), .ZN(new_n5950_));
  INV_X1     g05694(.I(new_n5950_), .ZN(new_n5951_));
  NAND2_X1   g05695(.A1(new_n5949_), .A2(new_n5951_), .ZN(new_n5952_));
  XOR2_X1    g05696(.A1(\b[51] ), .A2(\b[52] ), .Z(new_n5953_));
  OAI21_X1   g05697(.A1(new_n5949_), .A2(new_n5953_), .B(new_n5952_), .ZN(new_n5954_));
  INV_X1     g05698(.I(\b[52] ), .ZN(new_n5955_));
  OAI22_X1   g05699(.A1(new_n405_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n404_), .ZN(new_n5956_));
  NAND2_X1   g05700(.A1(new_n279_), .A2(\b[50] ), .ZN(new_n5957_));
  AOI21_X1   g05701(.A1(new_n5956_), .A2(new_n5957_), .B(new_n264_), .ZN(new_n5958_));
  NAND2_X1   g05702(.A1(new_n5954_), .A2(new_n5958_), .ZN(new_n5959_));
  XOR2_X1    g05703(.A1(new_n5959_), .A2(\a[2] ), .Z(new_n5960_));
  INV_X1     g05704(.I(new_n5960_), .ZN(new_n5961_));
  XOR2_X1    g05705(.A1(new_n5945_), .A2(new_n5961_), .Z(new_n5962_));
  XOR2_X1    g05706(.A1(new_n5945_), .A2(new_n5961_), .Z(new_n5963_));
  NAND2_X1   g05707(.A1(new_n5759_), .A2(new_n5963_), .ZN(new_n5964_));
  OAI21_X1   g05708(.A1(new_n5759_), .A2(new_n5962_), .B(new_n5964_), .ZN(new_n5965_));
  NOR2_X1    g05709(.A1(new_n5754_), .A2(new_n5750_), .ZN(new_n5966_));
  NOR2_X1    g05710(.A1(new_n5752_), .A2(new_n5966_), .ZN(new_n5967_));
  INV_X1     g05711(.I(new_n5746_), .ZN(new_n5968_));
  XOR2_X1    g05712(.A1(new_n5553_), .A2(new_n5737_), .Z(new_n5969_));
  NOR2_X1    g05713(.A1(new_n5969_), .A2(new_n5968_), .ZN(new_n5970_));
  NOR2_X1    g05714(.A1(new_n5967_), .A2(new_n5970_), .ZN(new_n5971_));
  OAI21_X1   g05715(.A1(new_n5968_), .A2(new_n5969_), .B(new_n5965_), .ZN(new_n5972_));
  OAI22_X1   g05716(.A1(new_n5971_), .A2(new_n5965_), .B1(new_n5967_), .B2(new_n5972_), .ZN(\f[52] ));
  XNOR2_X1   g05717(.A1(new_n5759_), .A2(new_n5945_), .ZN(new_n5974_));
  OAI21_X1   g05718(.A1(new_n5967_), .A2(new_n5970_), .B(new_n5965_), .ZN(new_n5975_));
  OAI21_X1   g05719(.A1(new_n5961_), .A2(new_n5974_), .B(new_n5975_), .ZN(new_n5976_));
  OAI22_X1   g05720(.A1(new_n437_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n431_), .ZN(new_n5977_));
  NAND2_X1   g05721(.A1(new_n775_), .A2(\b[45] ), .ZN(new_n5978_));
  AOI21_X1   g05722(.A1(new_n5977_), .A2(new_n5978_), .B(new_n440_), .ZN(new_n5979_));
  NAND2_X1   g05723(.A1(new_n5004_), .A2(new_n5979_), .ZN(new_n5980_));
  XOR2_X1    g05724(.A1(new_n5980_), .A2(\a[8] ), .Z(new_n5981_));
  INV_X1     g05725(.I(new_n5981_), .ZN(new_n5982_));
  OAI22_X1   g05726(.A1(new_n582_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n577_), .ZN(new_n5983_));
  NAND2_X1   g05727(.A1(new_n960_), .A2(\b[42] ), .ZN(new_n5984_));
  AOI21_X1   g05728(.A1(new_n5983_), .A2(new_n5984_), .B(new_n585_), .ZN(new_n5985_));
  NAND2_X1   g05729(.A1(new_n4500_), .A2(new_n5985_), .ZN(new_n5986_));
  XOR2_X1    g05730(.A1(new_n5986_), .A2(\a[11] ), .Z(new_n5987_));
  NOR3_X1    g05731(.A1(new_n5919_), .A2(new_n5916_), .A3(new_n5925_), .ZN(new_n5988_));
  INV_X1     g05732(.I(new_n5856_), .ZN(new_n5989_));
  NOR2_X1    g05733(.A1(new_n5989_), .A2(new_n5861_), .ZN(new_n5990_));
  NOR2_X1    g05734(.A1(new_n5845_), .A2(new_n5851_), .ZN(new_n5991_));
  INV_X1     g05735(.I(new_n5991_), .ZN(new_n5992_));
  NAND2_X1   g05736(.A1(new_n5824_), .A2(new_n5832_), .ZN(new_n5993_));
  INV_X1     g05737(.I(new_n5993_), .ZN(new_n5994_));
  XOR2_X1    g05738(.A1(new_n5770_), .A2(new_n5220_), .Z(new_n5995_));
  OAI21_X1   g05739(.A1(new_n5781_), .A2(new_n5371_), .B(new_n5778_), .ZN(new_n5996_));
  NAND3_X1   g05740(.A1(new_n5777_), .A2(new_n5556_), .A3(new_n5779_), .ZN(new_n5997_));
  NAND3_X1   g05741(.A1(new_n5996_), .A2(new_n5997_), .A3(new_n5995_), .ZN(new_n5998_));
  XOR2_X1    g05742(.A1(new_n5770_), .A2(\a[50] ), .Z(new_n5999_));
  OAI21_X1   g05743(.A1(new_n5782_), .A2(new_n5780_), .B(new_n5999_), .ZN(new_n6000_));
  AOI22_X1   g05744(.A1(new_n6000_), .A2(new_n5998_), .B1(new_n5803_), .B2(new_n5995_), .ZN(new_n6001_));
  INV_X1     g05745(.I(new_n5797_), .ZN(new_n6002_));
  NOR3_X1    g05746(.A1(new_n6002_), .A2(new_n5783_), .A3(new_n5572_), .ZN(new_n6003_));
  XOR2_X1    g05747(.A1(\a[52] ), .A2(\a[53] ), .Z(new_n6004_));
  NOR2_X1    g05748(.A1(new_n5571_), .A2(new_n6004_), .ZN(new_n6005_));
  NOR2_X1    g05749(.A1(new_n5792_), .A2(new_n267_), .ZN(new_n6006_));
  AOI21_X1   g05750(.A1(\b[2] ), .A2(new_n6005_), .B(new_n6006_), .ZN(new_n6007_));
  XNOR2_X1   g05751(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n6008_));
  XNOR2_X1   g05752(.A1(\a[50] ), .A2(\a[52] ), .ZN(new_n6009_));
  NAND2_X1   g05753(.A1(new_n6008_), .A2(new_n6009_), .ZN(new_n6010_));
  XNOR2_X1   g05754(.A1(\a[50] ), .A2(\a[53] ), .ZN(new_n6011_));
  NAND2_X1   g05755(.A1(new_n6010_), .A2(new_n6011_), .ZN(new_n6012_));
  NOR2_X1    g05756(.A1(new_n6012_), .A2(new_n258_), .ZN(new_n6013_));
  NOR2_X1    g05757(.A1(new_n5796_), .A2(new_n278_), .ZN(new_n6014_));
  OAI21_X1   g05758(.A1(new_n6013_), .A2(new_n6007_), .B(new_n6014_), .ZN(new_n6015_));
  NOR2_X1    g05759(.A1(new_n6015_), .A2(\a[53] ), .ZN(new_n6016_));
  NAND2_X1   g05760(.A1(new_n6015_), .A2(\a[53] ), .ZN(new_n6017_));
  INV_X1     g05761(.I(new_n6017_), .ZN(new_n6018_));
  OAI21_X1   g05762(.A1(new_n6018_), .A2(new_n6016_), .B(new_n6003_), .ZN(new_n6019_));
  INV_X1     g05763(.I(new_n6003_), .ZN(new_n6020_));
  INV_X1     g05764(.I(new_n6016_), .ZN(new_n6021_));
  NAND3_X1   g05765(.A1(new_n6020_), .A2(new_n6021_), .A3(new_n6017_), .ZN(new_n6022_));
  NAND2_X1   g05766(.A1(new_n6022_), .A2(new_n6019_), .ZN(new_n6023_));
  OAI22_X1   g05767(.A1(new_n5228_), .A2(new_n347_), .B1(new_n393_), .B2(new_n5225_), .ZN(new_n6024_));
  NAND2_X1   g05768(.A1(new_n5387_), .A2(\b[3] ), .ZN(new_n6025_));
  AOI21_X1   g05769(.A1(new_n6024_), .A2(new_n6025_), .B(new_n5231_), .ZN(new_n6026_));
  NAND3_X1   g05770(.A1(new_n352_), .A2(new_n5220_), .A3(new_n6026_), .ZN(new_n6027_));
  AOI21_X1   g05771(.A1(new_n352_), .A2(new_n6026_), .B(new_n5220_), .ZN(new_n6028_));
  INV_X1     g05772(.I(new_n6028_), .ZN(new_n6029_));
  AOI21_X1   g05773(.A1(new_n6027_), .A2(new_n6029_), .B(new_n6023_), .ZN(new_n6030_));
  NAND3_X1   g05774(.A1(new_n6029_), .A2(new_n6023_), .A3(new_n6027_), .ZN(new_n6031_));
  INV_X1     g05775(.I(new_n6031_), .ZN(new_n6032_));
  OAI21_X1   g05776(.A1(new_n6030_), .A2(new_n6032_), .B(new_n6001_), .ZN(new_n6033_));
  NOR3_X1    g05777(.A1(new_n5782_), .A2(new_n5780_), .A3(new_n5999_), .ZN(new_n6034_));
  AOI21_X1   g05778(.A1(new_n5996_), .A2(new_n5997_), .B(new_n5995_), .ZN(new_n6035_));
  OAI22_X1   g05779(.A1(new_n6034_), .A2(new_n6035_), .B1(new_n5800_), .B2(new_n5999_), .ZN(new_n6036_));
  INV_X1     g05780(.I(new_n6027_), .ZN(new_n6037_));
  OAI21_X1   g05781(.A1(new_n6037_), .A2(new_n6028_), .B(new_n6023_), .ZN(new_n6038_));
  AOI21_X1   g05782(.A1(new_n6021_), .A2(new_n6017_), .B(new_n6020_), .ZN(new_n6039_));
  NOR3_X1    g05783(.A1(new_n6018_), .A2(new_n6016_), .A3(new_n6003_), .ZN(new_n6040_));
  NOR2_X1    g05784(.A1(new_n6039_), .A2(new_n6040_), .ZN(new_n6041_));
  NAND3_X1   g05785(.A1(new_n6041_), .A2(new_n6029_), .A3(new_n6027_), .ZN(new_n6042_));
  NAND2_X1   g05786(.A1(new_n6038_), .A2(new_n6042_), .ZN(new_n6043_));
  NAND2_X1   g05787(.A1(new_n6043_), .A2(new_n6036_), .ZN(new_n6044_));
  NAND2_X1   g05788(.A1(new_n6033_), .A2(new_n6044_), .ZN(new_n6045_));
  OAI22_X1   g05789(.A1(new_n4711_), .A2(new_n495_), .B1(new_n450_), .B2(new_n4706_), .ZN(new_n6046_));
  NAND2_X1   g05790(.A1(new_n5814_), .A2(\b[6] ), .ZN(new_n6047_));
  AOI21_X1   g05791(.A1(new_n6046_), .A2(new_n6047_), .B(new_n4714_), .ZN(new_n6048_));
  NAND2_X1   g05792(.A1(new_n494_), .A2(new_n6048_), .ZN(new_n6049_));
  XOR2_X1    g05793(.A1(new_n6049_), .A2(\a[47] ), .Z(new_n6050_));
  NOR2_X1    g05794(.A1(new_n6045_), .A2(new_n6050_), .ZN(new_n6051_));
  OAI21_X1   g05795(.A1(new_n6037_), .A2(new_n6028_), .B(new_n6041_), .ZN(new_n6052_));
  AOI21_X1   g05796(.A1(new_n6052_), .A2(new_n6031_), .B(new_n6036_), .ZN(new_n6053_));
  AOI21_X1   g05797(.A1(new_n6038_), .A2(new_n6042_), .B(new_n6001_), .ZN(new_n6054_));
  NOR2_X1    g05798(.A1(new_n6053_), .A2(new_n6054_), .ZN(new_n6055_));
  XOR2_X1    g05799(.A1(new_n6049_), .A2(new_n4701_), .Z(new_n6056_));
  NOR2_X1    g05800(.A1(new_n6055_), .A2(new_n6056_), .ZN(new_n6057_));
  OAI21_X1   g05801(.A1(new_n6057_), .A2(new_n6051_), .B(new_n5819_), .ZN(new_n6058_));
  NAND3_X1   g05802(.A1(new_n5820_), .A2(new_n5821_), .A3(new_n5822_), .ZN(new_n6059_));
  AOI21_X1   g05803(.A1(new_n6033_), .A2(new_n6044_), .B(new_n6050_), .ZN(new_n6060_));
  NOR3_X1    g05804(.A1(new_n6053_), .A2(new_n6054_), .A3(new_n6056_), .ZN(new_n6061_));
  OAI21_X1   g05805(.A1(new_n6060_), .A2(new_n6061_), .B(new_n6059_), .ZN(new_n6062_));
  OAI22_X1   g05806(.A1(new_n4208_), .A2(new_n659_), .B1(new_n617_), .B2(new_n4203_), .ZN(new_n6063_));
  NAND2_X1   g05807(.A1(new_n5244_), .A2(\b[9] ), .ZN(new_n6064_));
  AOI21_X1   g05808(.A1(new_n6063_), .A2(new_n6064_), .B(new_n4211_), .ZN(new_n6065_));
  NAND3_X1   g05809(.A1(new_n663_), .A2(new_n4198_), .A3(new_n6065_), .ZN(new_n6066_));
  INV_X1     g05810(.I(new_n6066_), .ZN(new_n6067_));
  AOI21_X1   g05811(.A1(new_n663_), .A2(new_n6065_), .B(new_n4198_), .ZN(new_n6068_));
  NOR2_X1    g05812(.A1(new_n6067_), .A2(new_n6068_), .ZN(new_n6069_));
  AOI21_X1   g05813(.A1(new_n6058_), .A2(new_n6062_), .B(new_n6069_), .ZN(new_n6070_));
  NAND2_X1   g05814(.A1(new_n6055_), .A2(new_n6056_), .ZN(new_n6071_));
  NAND2_X1   g05815(.A1(new_n6045_), .A2(new_n6050_), .ZN(new_n6072_));
  AOI21_X1   g05816(.A1(new_n6071_), .A2(new_n6072_), .B(new_n6059_), .ZN(new_n6073_));
  OAI21_X1   g05817(.A1(new_n6053_), .A2(new_n6054_), .B(new_n6056_), .ZN(new_n6074_));
  NAND3_X1   g05818(.A1(new_n6033_), .A2(new_n6044_), .A3(new_n6050_), .ZN(new_n6075_));
  AOI21_X1   g05819(.A1(new_n6074_), .A2(new_n6075_), .B(new_n5819_), .ZN(new_n6076_));
  INV_X1     g05820(.I(new_n6068_), .ZN(new_n6077_));
  NAND2_X1   g05821(.A1(new_n6077_), .A2(new_n6066_), .ZN(new_n6078_));
  NOR3_X1    g05822(.A1(new_n6078_), .A2(new_n6073_), .A3(new_n6076_), .ZN(new_n6079_));
  OAI22_X1   g05823(.A1(new_n3736_), .A2(new_n848_), .B1(new_n795_), .B2(new_n3731_), .ZN(new_n6080_));
  NAND2_X1   g05824(.A1(new_n4730_), .A2(\b[12] ), .ZN(new_n6081_));
  AOI21_X1   g05825(.A1(new_n6080_), .A2(new_n6081_), .B(new_n3739_), .ZN(new_n6082_));
  AND3_X2    g05826(.A1(new_n847_), .A2(new_n3726_), .A3(new_n6082_), .Z(new_n6083_));
  AOI21_X1   g05827(.A1(new_n847_), .A2(new_n6082_), .B(new_n3726_), .ZN(new_n6084_));
  NOR2_X1    g05828(.A1(new_n6083_), .A2(new_n6084_), .ZN(new_n6085_));
  NOR3_X1    g05829(.A1(new_n6070_), .A2(new_n6079_), .A3(new_n6085_), .ZN(new_n6086_));
  NAND2_X1   g05830(.A1(new_n6058_), .A2(new_n6062_), .ZN(new_n6087_));
  NAND2_X1   g05831(.A1(new_n6087_), .A2(new_n6078_), .ZN(new_n6088_));
  NAND3_X1   g05832(.A1(new_n6069_), .A2(new_n6058_), .A3(new_n6062_), .ZN(new_n6089_));
  INV_X1     g05833(.I(new_n6085_), .ZN(new_n6090_));
  AOI21_X1   g05834(.A1(new_n6088_), .A2(new_n6089_), .B(new_n6090_), .ZN(new_n6091_));
  OAI21_X1   g05835(.A1(new_n6091_), .A2(new_n6086_), .B(new_n5994_), .ZN(new_n6092_));
  AOI21_X1   g05836(.A1(new_n6088_), .A2(new_n6089_), .B(new_n6085_), .ZN(new_n6093_));
  NOR3_X1    g05837(.A1(new_n6070_), .A2(new_n6079_), .A3(new_n6090_), .ZN(new_n6094_));
  OAI21_X1   g05838(.A1(new_n6093_), .A2(new_n6094_), .B(new_n5993_), .ZN(new_n6095_));
  NAND2_X1   g05839(.A1(new_n6092_), .A2(new_n6095_), .ZN(new_n6096_));
  NOR2_X1    g05840(.A1(new_n5834_), .A2(new_n5841_), .ZN(new_n6097_));
  INV_X1     g05841(.I(new_n6097_), .ZN(new_n6098_));
  NOR2_X1    g05842(.A1(new_n6096_), .A2(new_n6098_), .ZN(new_n6099_));
  NAND3_X1   g05843(.A1(new_n6088_), .A2(new_n6090_), .A3(new_n6089_), .ZN(new_n6100_));
  OAI21_X1   g05844(.A1(new_n6070_), .A2(new_n6079_), .B(new_n6085_), .ZN(new_n6101_));
  AOI21_X1   g05845(.A1(new_n6100_), .A2(new_n6101_), .B(new_n5993_), .ZN(new_n6102_));
  OAI21_X1   g05846(.A1(new_n6070_), .A2(new_n6079_), .B(new_n6090_), .ZN(new_n6103_));
  NAND3_X1   g05847(.A1(new_n6088_), .A2(new_n6085_), .A3(new_n6089_), .ZN(new_n6104_));
  AOI21_X1   g05848(.A1(new_n6104_), .A2(new_n6103_), .B(new_n5994_), .ZN(new_n6105_));
  NOR2_X1    g05849(.A1(new_n6102_), .A2(new_n6105_), .ZN(new_n6106_));
  NOR2_X1    g05850(.A1(new_n6106_), .A2(new_n6097_), .ZN(new_n6107_));
  OAI22_X1   g05851(.A1(new_n3298_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n3293_), .ZN(new_n6108_));
  NAND2_X1   g05852(.A1(new_n4227_), .A2(\b[15] ), .ZN(new_n6109_));
  AOI21_X1   g05853(.A1(new_n6108_), .A2(new_n6109_), .B(new_n3301_), .ZN(new_n6110_));
  AND3_X2    g05854(.A1(new_n1047_), .A2(new_n3288_), .A3(new_n6110_), .Z(new_n6111_));
  AOI21_X1   g05855(.A1(new_n1047_), .A2(new_n6110_), .B(new_n3288_), .ZN(new_n6112_));
  NOR2_X1    g05856(.A1(new_n6111_), .A2(new_n6112_), .ZN(new_n6113_));
  NOR3_X1    g05857(.A1(new_n6107_), .A2(new_n6099_), .A3(new_n6113_), .ZN(new_n6114_));
  INV_X1     g05858(.I(new_n6114_), .ZN(new_n6115_));
  OAI21_X1   g05859(.A1(new_n6107_), .A2(new_n6099_), .B(new_n6113_), .ZN(new_n6116_));
  AOI21_X1   g05860(.A1(new_n6115_), .A2(new_n6116_), .B(new_n5992_), .ZN(new_n6117_));
  NOR2_X1    g05861(.A1(new_n6107_), .A2(new_n6099_), .ZN(new_n6118_));
  XOR2_X1    g05862(.A1(new_n6118_), .A2(new_n6113_), .Z(new_n6119_));
  NOR2_X1    g05863(.A1(new_n6119_), .A2(new_n5991_), .ZN(new_n6120_));
  NOR2_X1    g05864(.A1(new_n6120_), .A2(new_n6117_), .ZN(new_n6121_));
  OAI22_X1   g05865(.A1(new_n2846_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n2841_), .ZN(new_n6122_));
  NAND2_X1   g05866(.A1(new_n3755_), .A2(\b[18] ), .ZN(new_n6123_));
  AOI21_X1   g05867(.A1(new_n6122_), .A2(new_n6123_), .B(new_n2849_), .ZN(new_n6124_));
  NAND2_X1   g05868(.A1(new_n1304_), .A2(new_n6124_), .ZN(new_n6125_));
  XOR2_X1    g05869(.A1(new_n6125_), .A2(\a[35] ), .Z(new_n6126_));
  XNOR2_X1   g05870(.A1(new_n6121_), .A2(new_n6126_), .ZN(new_n6127_));
  OAI22_X1   g05871(.A1(new_n2452_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n2447_), .ZN(new_n6128_));
  NAND2_X1   g05872(.A1(new_n3312_), .A2(\b[21] ), .ZN(new_n6129_));
  AOI21_X1   g05873(.A1(new_n6128_), .A2(new_n6129_), .B(new_n2455_), .ZN(new_n6130_));
  NAND2_X1   g05874(.A1(new_n1604_), .A2(new_n6130_), .ZN(new_n6131_));
  XOR2_X1    g05875(.A1(new_n6131_), .A2(\a[32] ), .Z(new_n6132_));
  XOR2_X1    g05876(.A1(new_n6127_), .A2(new_n6132_), .Z(new_n6133_));
  NAND2_X1   g05877(.A1(new_n6133_), .A2(new_n5990_), .ZN(new_n6134_));
  XOR2_X1    g05878(.A1(new_n6127_), .A2(new_n6132_), .Z(new_n6135_));
  OAI21_X1   g05879(.A1(new_n5990_), .A2(new_n6135_), .B(new_n6134_), .ZN(new_n6136_));
  XOR2_X1    g05880(.A1(new_n6136_), .A2(new_n5869_), .Z(new_n6137_));
  OAI22_X1   g05881(.A1(new_n2084_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n2079_), .ZN(new_n6138_));
  NAND2_X1   g05882(.A1(new_n2864_), .A2(\b[24] ), .ZN(new_n6139_));
  AOI21_X1   g05883(.A1(new_n6138_), .A2(new_n6139_), .B(new_n2087_), .ZN(new_n6140_));
  NAND2_X1   g05884(.A1(new_n1926_), .A2(new_n6140_), .ZN(new_n6141_));
  XOR2_X1    g05885(.A1(new_n6141_), .A2(\a[29] ), .Z(new_n6142_));
  XNOR2_X1   g05886(.A1(new_n6137_), .A2(new_n6142_), .ZN(new_n6143_));
  NOR2_X1    g05887(.A1(new_n5871_), .A2(new_n5876_), .ZN(new_n6144_));
  XNOR2_X1   g05888(.A1(new_n6143_), .A2(new_n6144_), .ZN(new_n6145_));
  OAI22_X1   g05889(.A1(new_n1760_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n1755_), .ZN(new_n6146_));
  NAND2_X1   g05890(.A1(new_n2470_), .A2(\b[27] ), .ZN(new_n6147_));
  AOI21_X1   g05891(.A1(new_n6146_), .A2(new_n6147_), .B(new_n1763_), .ZN(new_n6148_));
  NAND2_X1   g05892(.A1(new_n2276_), .A2(new_n6148_), .ZN(new_n6149_));
  XOR2_X1    g05893(.A1(new_n6149_), .A2(\a[26] ), .Z(new_n6150_));
  XOR2_X1    g05894(.A1(new_n6145_), .A2(new_n6150_), .Z(new_n6151_));
  NOR3_X1    g05895(.A1(new_n5877_), .A2(new_n5878_), .A3(new_n5884_), .ZN(new_n6152_));
  XNOR2_X1   g05896(.A1(new_n6151_), .A2(new_n6152_), .ZN(new_n6153_));
  OAI22_X1   g05897(.A1(new_n1444_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n1439_), .ZN(new_n6154_));
  NAND2_X1   g05898(.A1(new_n2098_), .A2(\b[30] ), .ZN(new_n6155_));
  AOI21_X1   g05899(.A1(new_n6154_), .A2(new_n6155_), .B(new_n1447_), .ZN(new_n6156_));
  NAND2_X1   g05900(.A1(new_n2659_), .A2(new_n6156_), .ZN(new_n6157_));
  XOR2_X1    g05901(.A1(new_n6157_), .A2(\a[23] ), .Z(new_n6158_));
  XOR2_X1    g05902(.A1(new_n6153_), .A2(new_n6158_), .Z(new_n6159_));
  INV_X1     g05903(.I(new_n6159_), .ZN(new_n6160_));
  NAND2_X1   g05904(.A1(new_n5890_), .A2(new_n5885_), .ZN(new_n6161_));
  OAI21_X1   g05905(.A1(new_n5900_), .A2(new_n5891_), .B(new_n6161_), .ZN(new_n6162_));
  XOR2_X1    g05906(.A1(new_n6162_), .A2(new_n6160_), .Z(new_n6163_));
  INV_X1     g05907(.I(new_n6163_), .ZN(new_n6164_));
  OAI22_X1   g05908(.A1(new_n1168_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n1163_), .ZN(new_n6165_));
  NAND2_X1   g05909(.A1(new_n1774_), .A2(\b[33] ), .ZN(new_n6166_));
  AOI21_X1   g05910(.A1(new_n6165_), .A2(new_n6166_), .B(new_n1171_), .ZN(new_n6167_));
  NAND2_X1   g05911(.A1(new_n3101_), .A2(new_n6167_), .ZN(new_n6168_));
  XOR2_X1    g05912(.A1(new_n6168_), .A2(\a[20] ), .Z(new_n6169_));
  NOR2_X1    g05913(.A1(new_n6164_), .A2(new_n6169_), .ZN(new_n6170_));
  NAND2_X1   g05914(.A1(new_n6164_), .A2(new_n6169_), .ZN(new_n6171_));
  INV_X1     g05915(.I(new_n6171_), .ZN(new_n6172_));
  NOR2_X1    g05916(.A1(new_n6172_), .A2(new_n6170_), .ZN(new_n6173_));
  INV_X1     g05917(.I(new_n5903_), .ZN(new_n6174_));
  XNOR2_X1   g05918(.A1(new_n5900_), .A2(new_n5891_), .ZN(new_n6175_));
  OAI21_X1   g05919(.A1(new_n5897_), .A2(new_n6175_), .B(new_n6174_), .ZN(new_n6176_));
  INV_X1     g05920(.I(new_n6176_), .ZN(new_n6177_));
  XOR2_X1    g05921(.A1(new_n6173_), .A2(new_n6177_), .Z(new_n6178_));
  OAI22_X1   g05922(.A1(new_n940_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n935_), .ZN(new_n6179_));
  NAND2_X1   g05923(.A1(new_n1458_), .A2(\b[36] ), .ZN(new_n6180_));
  AOI21_X1   g05924(.A1(new_n6179_), .A2(new_n6180_), .B(new_n943_), .ZN(new_n6181_));
  NAND2_X1   g05925(.A1(new_n3565_), .A2(new_n6181_), .ZN(new_n6182_));
  XOR2_X1    g05926(.A1(new_n6182_), .A2(\a[17] ), .Z(new_n6183_));
  INV_X1     g05927(.I(new_n6183_), .ZN(new_n6184_));
  XOR2_X1    g05928(.A1(new_n6178_), .A2(new_n6184_), .Z(new_n6185_));
  INV_X1     g05929(.I(new_n6185_), .ZN(new_n6186_));
  NAND2_X1   g05930(.A1(new_n6174_), .A2(new_n5908_), .ZN(new_n6187_));
  OAI21_X1   g05931(.A1(new_n5917_), .A2(new_n5909_), .B(new_n6187_), .ZN(new_n6188_));
  XOR2_X1    g05932(.A1(new_n6188_), .A2(new_n6186_), .Z(new_n6189_));
  OAI22_X1   g05933(.A1(new_n757_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n752_), .ZN(new_n6190_));
  NAND2_X1   g05934(.A1(new_n1182_), .A2(\b[39] ), .ZN(new_n6191_));
  AOI21_X1   g05935(.A1(new_n6190_), .A2(new_n6191_), .B(new_n760_), .ZN(new_n6192_));
  NAND2_X1   g05936(.A1(new_n3996_), .A2(new_n6192_), .ZN(new_n6193_));
  XOR2_X1    g05937(.A1(new_n6193_), .A2(\a[14] ), .Z(new_n6194_));
  XOR2_X1    g05938(.A1(new_n6189_), .A2(new_n6194_), .Z(new_n6195_));
  XOR2_X1    g05939(.A1(new_n5917_), .A2(new_n5909_), .Z(new_n6196_));
  AOI21_X1   g05940(.A1(new_n6196_), .A2(new_n5914_), .B(new_n5920_), .ZN(new_n6197_));
  XOR2_X1    g05941(.A1(new_n6195_), .A2(new_n6197_), .Z(new_n6198_));
  XOR2_X1    g05942(.A1(new_n6198_), .A2(new_n5988_), .Z(new_n6199_));
  XOR2_X1    g05943(.A1(new_n6199_), .A2(new_n5987_), .Z(new_n6200_));
  XOR2_X1    g05944(.A1(new_n6200_), .A2(new_n5982_), .Z(new_n6201_));
  XOR2_X1    g05945(.A1(new_n6201_), .A2(new_n5932_), .Z(new_n6202_));
  OAI22_X1   g05946(.A1(new_n364_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n320_), .ZN(new_n6203_));
  NAND2_X1   g05947(.A1(new_n594_), .A2(\b[48] ), .ZN(new_n6204_));
  AOI21_X1   g05948(.A1(new_n6203_), .A2(new_n6204_), .B(new_n312_), .ZN(new_n6205_));
  NAND2_X1   g05949(.A1(new_n5537_), .A2(new_n6205_), .ZN(new_n6206_));
  XOR2_X1    g05950(.A1(new_n6206_), .A2(\a[5] ), .Z(new_n6207_));
  INV_X1     g05951(.I(new_n5943_), .ZN(new_n6208_));
  XOR2_X1    g05952(.A1(new_n5725_), .A2(new_n5734_), .Z(new_n6209_));
  OAI21_X1   g05953(.A1(new_n5731_), .A2(new_n6209_), .B(new_n5756_), .ZN(new_n6210_));
  NAND2_X1   g05954(.A1(new_n6209_), .A2(new_n5731_), .ZN(new_n6211_));
  NAND4_X1   g05955(.A1(new_n6210_), .A2(new_n6208_), .A3(new_n5945_), .A4(new_n6211_), .ZN(new_n6212_));
  XOR2_X1    g05956(.A1(new_n6212_), .A2(new_n6207_), .Z(new_n6213_));
  XNOR2_X1   g05957(.A1(new_n6213_), .A2(new_n6202_), .ZN(new_n6214_));
  INV_X1     g05958(.I(\b[53] ), .ZN(new_n6215_));
  XOR2_X1    g05959(.A1(new_n5949_), .A2(\b[51] ), .Z(new_n6216_));
  AND3_X2    g05960(.A1(new_n6216_), .A2(new_n6215_), .A3(new_n5951_), .Z(new_n6217_));
  AOI21_X1   g05961(.A1(new_n6216_), .A2(new_n5951_), .B(new_n6215_), .ZN(new_n6218_));
  OR2_X2     g05962(.A1(new_n6217_), .A2(new_n6218_), .Z(new_n6219_));
  OAI22_X1   g05963(.A1(new_n405_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n404_), .ZN(new_n6220_));
  NAND2_X1   g05964(.A1(new_n279_), .A2(\b[51] ), .ZN(new_n6221_));
  AOI21_X1   g05965(.A1(new_n6220_), .A2(new_n6221_), .B(new_n264_), .ZN(new_n6222_));
  NAND2_X1   g05966(.A1(new_n6219_), .A2(new_n6222_), .ZN(new_n6223_));
  XOR2_X1    g05967(.A1(new_n6223_), .A2(\a[2] ), .Z(new_n6224_));
  XOR2_X1    g05968(.A1(new_n6214_), .A2(new_n6224_), .Z(new_n6225_));
  NAND2_X1   g05969(.A1(new_n5976_), .A2(new_n6225_), .ZN(new_n6226_));
  XOR2_X1    g05970(.A1(new_n6214_), .A2(new_n6224_), .Z(new_n6227_));
  OAI21_X1   g05971(.A1(new_n5976_), .A2(new_n6227_), .B(new_n6226_), .ZN(\f[53] ));
  OAI21_X1   g05972(.A1(new_n5738_), .A2(new_n6215_), .B(new_n5955_), .ZN(new_n6229_));
  NAND3_X1   g05973(.A1(new_n5947_), .A2(new_n5948_), .A3(new_n6229_), .ZN(new_n6230_));
  OAI21_X1   g05974(.A1(\b[51] ), .A2(\b[53] ), .B(\b[52] ), .ZN(new_n6231_));
  NAND2_X1   g05975(.A1(new_n6230_), .A2(new_n6231_), .ZN(new_n6232_));
  XNOR2_X1   g05976(.A1(\b[53] ), .A2(\b[54] ), .ZN(new_n6233_));
  INV_X1     g05977(.I(new_n6233_), .ZN(new_n6234_));
  NAND2_X1   g05978(.A1(new_n6232_), .A2(new_n6234_), .ZN(new_n6235_));
  XOR2_X1    g05979(.A1(\b[53] ), .A2(\b[54] ), .Z(new_n6236_));
  OAI21_X1   g05980(.A1(new_n6232_), .A2(new_n6236_), .B(new_n6235_), .ZN(new_n6237_));
  INV_X1     g05981(.I(\b[54] ), .ZN(new_n6238_));
  OAI22_X1   g05982(.A1(new_n405_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n404_), .ZN(new_n6239_));
  NAND2_X1   g05983(.A1(new_n279_), .A2(\b[52] ), .ZN(new_n6240_));
  AOI21_X1   g05984(.A1(new_n6239_), .A2(new_n6240_), .B(new_n264_), .ZN(new_n6241_));
  NAND2_X1   g05985(.A1(new_n6237_), .A2(new_n6241_), .ZN(new_n6242_));
  XOR2_X1    g05986(.A1(new_n6242_), .A2(\a[2] ), .Z(new_n6243_));
  OAI22_X1   g05987(.A1(new_n364_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n320_), .ZN(new_n6244_));
  NAND2_X1   g05988(.A1(new_n594_), .A2(\b[49] ), .ZN(new_n6245_));
  AOI21_X1   g05989(.A1(new_n6244_), .A2(new_n6245_), .B(new_n312_), .ZN(new_n6246_));
  NAND2_X1   g05990(.A1(new_n5741_), .A2(new_n6246_), .ZN(new_n6247_));
  XOR2_X1    g05991(.A1(new_n6247_), .A2(\a[5] ), .Z(new_n6248_));
  INV_X1     g05992(.I(new_n6248_), .ZN(new_n6249_));
  AOI21_X1   g05993(.A1(new_n5991_), .A2(new_n6116_), .B(new_n6114_), .ZN(new_n6250_));
  AOI21_X1   g05994(.A1(new_n5819_), .A2(new_n6075_), .B(new_n6060_), .ZN(new_n6251_));
  OAI21_X1   g05995(.A1(new_n6036_), .A2(new_n6032_), .B(new_n6052_), .ZN(new_n6252_));
  NAND2_X1   g05996(.A1(\a[53] ), .A2(\a[54] ), .ZN(new_n6253_));
  OR2_X2     g05997(.A1(\a[53] ), .A2(\a[54] ), .Z(new_n6254_));
  NAND2_X1   g05998(.A1(new_n6254_), .A2(new_n6253_), .ZN(new_n6255_));
  NOR2_X1    g05999(.A1(new_n6255_), .A2(new_n258_), .ZN(new_n6256_));
  NOR4_X1    g06000(.A1(new_n6015_), .A2(new_n6002_), .A3(new_n5783_), .A4(new_n5572_), .ZN(new_n6257_));
  OAI22_X1   g06001(.A1(new_n5786_), .A2(new_n290_), .B1(new_n292_), .B2(new_n5792_), .ZN(new_n6258_));
  OAI21_X1   g06002(.A1(new_n267_), .A2(new_n6012_), .B(new_n6258_), .ZN(new_n6259_));
  NOR2_X1    g06003(.A1(new_n677_), .A2(new_n5796_), .ZN(new_n6260_));
  AND3_X2    g06004(.A1(new_n6259_), .A2(new_n5783_), .A3(new_n6260_), .Z(new_n6261_));
  AOI21_X1   g06005(.A1(new_n6259_), .A2(new_n6260_), .B(new_n5783_), .ZN(new_n6262_));
  NOR2_X1    g06006(.A1(new_n6261_), .A2(new_n6262_), .ZN(new_n6263_));
  NOR2_X1    g06007(.A1(new_n6263_), .A2(new_n6257_), .ZN(new_n6264_));
  INV_X1     g06008(.I(new_n6264_), .ZN(new_n6265_));
  NAND2_X1   g06009(.A1(new_n6263_), .A2(new_n6257_), .ZN(new_n6266_));
  AOI21_X1   g06010(.A1(new_n6265_), .A2(new_n6266_), .B(new_n6256_), .ZN(new_n6267_));
  NAND3_X1   g06011(.A1(new_n6265_), .A2(new_n6266_), .A3(new_n6256_), .ZN(new_n6268_));
  INV_X1     g06012(.I(new_n6268_), .ZN(new_n6269_));
  OAI22_X1   g06013(.A1(new_n5228_), .A2(new_n403_), .B1(new_n347_), .B2(new_n5225_), .ZN(new_n6270_));
  OAI21_X1   g06014(.A1(new_n393_), .A2(new_n5378_), .B(new_n6270_), .ZN(new_n6271_));
  AND3_X2    g06015(.A1(new_n402_), .A2(new_n5394_), .A3(new_n6271_), .Z(new_n6272_));
  XOR2_X1    g06016(.A1(new_n6272_), .A2(\a[50] ), .Z(new_n6273_));
  OAI21_X1   g06017(.A1(new_n6269_), .A2(new_n6267_), .B(new_n6273_), .ZN(new_n6274_));
  INV_X1     g06018(.I(new_n6256_), .ZN(new_n6275_));
  INV_X1     g06019(.I(new_n6266_), .ZN(new_n6276_));
  OAI21_X1   g06020(.A1(new_n6276_), .A2(new_n6264_), .B(new_n6275_), .ZN(new_n6277_));
  XOR2_X1    g06021(.A1(new_n6272_), .A2(new_n5220_), .Z(new_n6278_));
  NAND3_X1   g06022(.A1(new_n6278_), .A2(new_n6277_), .A3(new_n6268_), .ZN(new_n6279_));
  NAND2_X1   g06023(.A1(new_n6274_), .A2(new_n6279_), .ZN(new_n6280_));
  NAND2_X1   g06024(.A1(new_n6280_), .A2(new_n6252_), .ZN(new_n6281_));
  AOI21_X1   g06025(.A1(new_n6001_), .A2(new_n6031_), .B(new_n6030_), .ZN(new_n6282_));
  NOR3_X1    g06026(.A1(new_n6269_), .A2(new_n6267_), .A3(new_n6278_), .ZN(new_n6283_));
  AOI21_X1   g06027(.A1(new_n6277_), .A2(new_n6268_), .B(new_n6273_), .ZN(new_n6284_));
  OAI21_X1   g06028(.A1(new_n6283_), .A2(new_n6284_), .B(new_n6282_), .ZN(new_n6285_));
  NAND2_X1   g06029(.A1(new_n6281_), .A2(new_n6285_), .ZN(new_n6286_));
  OAI22_X1   g06030(.A1(new_n4711_), .A2(new_n510_), .B1(new_n495_), .B2(new_n4706_), .ZN(new_n6287_));
  NAND2_X1   g06031(.A1(new_n5814_), .A2(\b[7] ), .ZN(new_n6288_));
  AOI21_X1   g06032(.A1(new_n6287_), .A2(new_n6288_), .B(new_n4714_), .ZN(new_n6289_));
  NAND2_X1   g06033(.A1(new_n518_), .A2(new_n6289_), .ZN(new_n6290_));
  XOR2_X1    g06034(.A1(new_n6290_), .A2(new_n4701_), .Z(new_n6291_));
  XOR2_X1    g06035(.A1(new_n6286_), .A2(new_n6291_), .Z(new_n6292_));
  NAND3_X1   g06036(.A1(new_n6281_), .A2(new_n6285_), .A3(new_n6291_), .ZN(new_n6293_));
  AOI21_X1   g06037(.A1(new_n6274_), .A2(new_n6279_), .B(new_n6282_), .ZN(new_n6294_));
  NAND3_X1   g06038(.A1(new_n6273_), .A2(new_n6277_), .A3(new_n6268_), .ZN(new_n6295_));
  OAI21_X1   g06039(.A1(new_n6269_), .A2(new_n6267_), .B(new_n6278_), .ZN(new_n6296_));
  AOI21_X1   g06040(.A1(new_n6295_), .A2(new_n6296_), .B(new_n6252_), .ZN(new_n6297_));
  XOR2_X1    g06041(.A1(new_n6290_), .A2(\a[47] ), .Z(new_n6298_));
  OAI21_X1   g06042(.A1(new_n6297_), .A2(new_n6294_), .B(new_n6298_), .ZN(new_n6299_));
  NAND2_X1   g06043(.A1(new_n6299_), .A2(new_n6293_), .ZN(new_n6300_));
  NAND2_X1   g06044(.A1(new_n6300_), .A2(new_n6251_), .ZN(new_n6301_));
  OAI21_X1   g06045(.A1(new_n6292_), .A2(new_n6251_), .B(new_n6301_), .ZN(new_n6302_));
  INV_X1     g06046(.I(new_n6302_), .ZN(new_n6303_));
  OAI22_X1   g06047(.A1(new_n4208_), .A2(new_n717_), .B1(new_n659_), .B2(new_n4203_), .ZN(new_n6304_));
  NAND2_X1   g06048(.A1(new_n5244_), .A2(\b[10] ), .ZN(new_n6305_));
  AOI21_X1   g06049(.A1(new_n6304_), .A2(new_n6305_), .B(new_n4211_), .ZN(new_n6306_));
  NAND2_X1   g06050(.A1(new_n716_), .A2(new_n6306_), .ZN(new_n6307_));
  XOR2_X1    g06051(.A1(new_n6307_), .A2(\a[44] ), .Z(new_n6308_));
  INV_X1     g06052(.I(new_n6308_), .ZN(new_n6309_));
  OAI21_X1   g06053(.A1(new_n6070_), .A2(new_n6079_), .B(new_n5993_), .ZN(new_n6310_));
  NAND2_X1   g06054(.A1(new_n6087_), .A2(new_n6069_), .ZN(new_n6311_));
  AOI21_X1   g06055(.A1(new_n6310_), .A2(new_n6311_), .B(new_n6309_), .ZN(new_n6312_));
  AOI21_X1   g06056(.A1(new_n6088_), .A2(new_n6089_), .B(new_n5994_), .ZN(new_n6313_));
  INV_X1     g06057(.I(new_n6311_), .ZN(new_n6314_));
  NOR3_X1    g06058(.A1(new_n6313_), .A2(new_n6308_), .A3(new_n6314_), .ZN(new_n6315_));
  OAI21_X1   g06059(.A1(new_n6315_), .A2(new_n6312_), .B(new_n6303_), .ZN(new_n6316_));
  OAI21_X1   g06060(.A1(new_n6313_), .A2(new_n6314_), .B(new_n6308_), .ZN(new_n6317_));
  NAND3_X1   g06061(.A1(new_n6310_), .A2(new_n6309_), .A3(new_n6311_), .ZN(new_n6318_));
  NAND3_X1   g06062(.A1(new_n6317_), .A2(new_n6318_), .A3(new_n6302_), .ZN(new_n6319_));
  NAND2_X1   g06063(.A1(new_n6316_), .A2(new_n6319_), .ZN(new_n6320_));
  OAI22_X1   g06064(.A1(new_n3736_), .A2(new_n904_), .B1(new_n848_), .B2(new_n3731_), .ZN(new_n6321_));
  NAND2_X1   g06065(.A1(new_n4730_), .A2(\b[13] ), .ZN(new_n6322_));
  AOI21_X1   g06066(.A1(new_n6321_), .A2(new_n6322_), .B(new_n3739_), .ZN(new_n6323_));
  NAND2_X1   g06067(.A1(new_n907_), .A2(new_n6323_), .ZN(new_n6324_));
  XOR2_X1    g06068(.A1(new_n6324_), .A2(\a[41] ), .Z(new_n6325_));
  AOI21_X1   g06069(.A1(new_n6088_), .A2(new_n6089_), .B(new_n5993_), .ZN(new_n6326_));
  NOR3_X1    g06070(.A1(new_n6070_), .A2(new_n6079_), .A3(new_n5994_), .ZN(new_n6327_));
  OAI21_X1   g06071(.A1(new_n6326_), .A2(new_n6327_), .B(new_n6085_), .ZN(new_n6328_));
  NAND2_X1   g06072(.A1(new_n6328_), .A2(new_n6098_), .ZN(new_n6329_));
  OAI21_X1   g06073(.A1(new_n6096_), .A2(new_n6329_), .B(new_n6325_), .ZN(new_n6330_));
  INV_X1     g06074(.I(new_n6325_), .ZN(new_n6331_));
  OAI21_X1   g06075(.A1(new_n6070_), .A2(new_n6079_), .B(new_n5994_), .ZN(new_n6332_));
  NAND3_X1   g06076(.A1(new_n6088_), .A2(new_n6089_), .A3(new_n5993_), .ZN(new_n6333_));
  NAND2_X1   g06077(.A1(new_n6333_), .A2(new_n6332_), .ZN(new_n6334_));
  AOI21_X1   g06078(.A1(new_n6334_), .A2(new_n6085_), .B(new_n6097_), .ZN(new_n6335_));
  NAND3_X1   g06079(.A1(new_n6106_), .A2(new_n6331_), .A3(new_n6335_), .ZN(new_n6336_));
  AOI21_X1   g06080(.A1(new_n6336_), .A2(new_n6330_), .B(new_n6320_), .ZN(new_n6337_));
  INV_X1     g06081(.I(new_n6320_), .ZN(new_n6338_));
  AOI21_X1   g06082(.A1(new_n6106_), .A2(new_n6335_), .B(new_n6331_), .ZN(new_n6339_));
  NOR3_X1    g06083(.A1(new_n6096_), .A2(new_n6329_), .A3(new_n6325_), .ZN(new_n6340_));
  NOR3_X1    g06084(.A1(new_n6338_), .A2(new_n6340_), .A3(new_n6339_), .ZN(new_n6341_));
  NOR2_X1    g06085(.A1(new_n6341_), .A2(new_n6337_), .ZN(new_n6342_));
  OAI22_X1   g06086(.A1(new_n3298_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n3293_), .ZN(new_n6343_));
  NAND2_X1   g06087(.A1(new_n4227_), .A2(\b[16] ), .ZN(new_n6344_));
  AOI21_X1   g06088(.A1(new_n6343_), .A2(new_n6344_), .B(new_n3301_), .ZN(new_n6345_));
  NAND2_X1   g06089(.A1(new_n1123_), .A2(new_n6345_), .ZN(new_n6346_));
  XOR2_X1    g06090(.A1(new_n6346_), .A2(\a[38] ), .Z(new_n6347_));
  XOR2_X1    g06091(.A1(new_n6342_), .A2(new_n6347_), .Z(new_n6348_));
  NOR3_X1    g06092(.A1(new_n6341_), .A2(new_n6337_), .A3(new_n6347_), .ZN(new_n6349_));
  OAI21_X1   g06093(.A1(new_n6340_), .A2(new_n6339_), .B(new_n6338_), .ZN(new_n6350_));
  NAND3_X1   g06094(.A1(new_n6336_), .A2(new_n6330_), .A3(new_n6320_), .ZN(new_n6351_));
  INV_X1     g06095(.I(new_n6347_), .ZN(new_n6352_));
  AOI21_X1   g06096(.A1(new_n6350_), .A2(new_n6351_), .B(new_n6352_), .ZN(new_n6353_));
  OAI21_X1   g06097(.A1(new_n6353_), .A2(new_n6349_), .B(new_n6250_), .ZN(new_n6354_));
  OAI21_X1   g06098(.A1(new_n6348_), .A2(new_n6250_), .B(new_n6354_), .ZN(new_n6355_));
  OAI22_X1   g06099(.A1(new_n2846_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n2841_), .ZN(new_n6356_));
  NAND2_X1   g06100(.A1(new_n3755_), .A2(\b[19] ), .ZN(new_n6357_));
  AOI21_X1   g06101(.A1(new_n6356_), .A2(new_n6357_), .B(new_n2849_), .ZN(new_n6358_));
  NAND2_X1   g06102(.A1(new_n1396_), .A2(new_n6358_), .ZN(new_n6359_));
  XOR2_X1    g06103(.A1(new_n6359_), .A2(new_n2836_), .Z(new_n6360_));
  NAND2_X1   g06104(.A1(new_n6121_), .A2(new_n6126_), .ZN(new_n6361_));
  OAI21_X1   g06105(.A1(new_n6127_), .A2(new_n5990_), .B(new_n6361_), .ZN(new_n6362_));
  XOR2_X1    g06106(.A1(new_n6362_), .A2(new_n6360_), .Z(new_n6363_));
  XOR2_X1    g06107(.A1(new_n6363_), .A2(new_n6355_), .Z(new_n6364_));
  OAI22_X1   g06108(.A1(new_n2452_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n2447_), .ZN(new_n6365_));
  NAND2_X1   g06109(.A1(new_n3312_), .A2(\b[22] ), .ZN(new_n6366_));
  AOI21_X1   g06110(.A1(new_n6365_), .A2(new_n6366_), .B(new_n2455_), .ZN(new_n6367_));
  NAND2_X1   g06111(.A1(new_n1708_), .A2(new_n6367_), .ZN(new_n6368_));
  XOR2_X1    g06112(.A1(new_n6368_), .A2(new_n2442_), .Z(new_n6369_));
  XOR2_X1    g06113(.A1(new_n6127_), .A2(new_n5990_), .Z(new_n6370_));
  NAND2_X1   g06114(.A1(new_n6370_), .A2(new_n6132_), .ZN(new_n6371_));
  NAND2_X1   g06115(.A1(new_n6371_), .A2(new_n5869_), .ZN(new_n6372_));
  NOR2_X1    g06116(.A1(new_n6136_), .A2(new_n6372_), .ZN(new_n6373_));
  XOR2_X1    g06117(.A1(new_n6373_), .A2(new_n6369_), .Z(new_n6374_));
  XOR2_X1    g06118(.A1(new_n6374_), .A2(new_n6364_), .Z(new_n6375_));
  OAI22_X1   g06119(.A1(new_n2084_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n2079_), .ZN(new_n6376_));
  NAND2_X1   g06120(.A1(new_n2864_), .A2(\b[25] ), .ZN(new_n6377_));
  AOI21_X1   g06121(.A1(new_n6376_), .A2(new_n6377_), .B(new_n2087_), .ZN(new_n6378_));
  NAND2_X1   g06122(.A1(new_n2042_), .A2(new_n6378_), .ZN(new_n6379_));
  XOR2_X1    g06123(.A1(new_n6379_), .A2(\a[29] ), .Z(new_n6380_));
  NAND2_X1   g06124(.A1(new_n6143_), .A2(new_n6144_), .ZN(new_n6381_));
  NAND2_X1   g06125(.A1(new_n6137_), .A2(new_n6142_), .ZN(new_n6382_));
  NAND2_X1   g06126(.A1(new_n6381_), .A2(new_n6382_), .ZN(new_n6383_));
  XOR2_X1    g06127(.A1(new_n6383_), .A2(new_n6380_), .Z(new_n6384_));
  XOR2_X1    g06128(.A1(new_n6384_), .A2(new_n6375_), .Z(new_n6385_));
  OAI22_X1   g06129(.A1(new_n1760_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n1755_), .ZN(new_n6386_));
  NAND2_X1   g06130(.A1(new_n2470_), .A2(\b[28] ), .ZN(new_n6387_));
  AOI21_X1   g06131(.A1(new_n6386_), .A2(new_n6387_), .B(new_n1763_), .ZN(new_n6388_));
  NAND2_X1   g06132(.A1(new_n2404_), .A2(new_n6388_), .ZN(new_n6389_));
  XOR2_X1    g06133(.A1(new_n6389_), .A2(\a[26] ), .Z(new_n6390_));
  NAND2_X1   g06134(.A1(new_n6145_), .A2(new_n6150_), .ZN(new_n6391_));
  XNOR2_X1   g06135(.A1(new_n6391_), .A2(new_n6390_), .ZN(new_n6392_));
  XOR2_X1    g06136(.A1(new_n6385_), .A2(new_n6392_), .Z(new_n6393_));
  OAI22_X1   g06137(.A1(new_n1444_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n1439_), .ZN(new_n6394_));
  NAND2_X1   g06138(.A1(new_n2098_), .A2(\b[31] ), .ZN(new_n6395_));
  AOI21_X1   g06139(.A1(new_n6394_), .A2(new_n6395_), .B(new_n1447_), .ZN(new_n6396_));
  NAND2_X1   g06140(.A1(new_n2797_), .A2(new_n6396_), .ZN(new_n6397_));
  XOR2_X1    g06141(.A1(new_n6397_), .A2(\a[23] ), .Z(new_n6398_));
  INV_X1     g06142(.I(new_n6153_), .ZN(new_n6399_));
  NAND2_X1   g06143(.A1(new_n6399_), .A2(new_n6158_), .ZN(new_n6400_));
  OAI21_X1   g06144(.A1(new_n6162_), .A2(new_n6160_), .B(new_n6400_), .ZN(new_n6401_));
  XOR2_X1    g06145(.A1(new_n6401_), .A2(new_n6398_), .Z(new_n6402_));
  XNOR2_X1   g06146(.A1(new_n6402_), .A2(new_n6393_), .ZN(new_n6403_));
  OAI22_X1   g06147(.A1(new_n1168_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n1163_), .ZN(new_n6404_));
  NAND2_X1   g06148(.A1(new_n1774_), .A2(\b[34] ), .ZN(new_n6405_));
  AOI21_X1   g06149(.A1(new_n6404_), .A2(new_n6405_), .B(new_n1171_), .ZN(new_n6406_));
  NAND2_X1   g06150(.A1(new_n3246_), .A2(new_n6406_), .ZN(new_n6407_));
  XOR2_X1    g06151(.A1(new_n6407_), .A2(\a[20] ), .Z(new_n6408_));
  NOR3_X1    g06152(.A1(new_n6172_), .A2(new_n6170_), .A3(new_n6177_), .ZN(new_n6409_));
  XOR2_X1    g06153(.A1(new_n6409_), .A2(new_n6408_), .Z(new_n6410_));
  XOR2_X1    g06154(.A1(new_n6410_), .A2(new_n6403_), .Z(new_n6411_));
  OAI22_X1   g06155(.A1(new_n940_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n935_), .ZN(new_n6412_));
  NAND2_X1   g06156(.A1(new_n1458_), .A2(\b[37] ), .ZN(new_n6413_));
  AOI21_X1   g06157(.A1(new_n6412_), .A2(new_n6413_), .B(new_n943_), .ZN(new_n6414_));
  NAND2_X1   g06158(.A1(new_n3700_), .A2(new_n6414_), .ZN(new_n6415_));
  XOR2_X1    g06159(.A1(new_n6415_), .A2(\a[17] ), .Z(new_n6416_));
  NOR2_X1    g06160(.A1(new_n6178_), .A2(new_n6184_), .ZN(new_n6417_));
  NOR2_X1    g06161(.A1(new_n6186_), .A2(new_n6417_), .ZN(new_n6418_));
  NAND2_X1   g06162(.A1(new_n6418_), .A2(new_n6188_), .ZN(new_n6419_));
  XOR2_X1    g06163(.A1(new_n6419_), .A2(new_n6416_), .Z(new_n6420_));
  XNOR2_X1   g06164(.A1(new_n6420_), .A2(new_n6411_), .ZN(new_n6421_));
  OAI22_X1   g06165(.A1(new_n757_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n752_), .ZN(new_n6422_));
  NAND2_X1   g06166(.A1(new_n1182_), .A2(\b[40] ), .ZN(new_n6423_));
  AOI21_X1   g06167(.A1(new_n6422_), .A2(new_n6423_), .B(new_n760_), .ZN(new_n6424_));
  NAND2_X1   g06168(.A1(new_n4017_), .A2(new_n6424_), .ZN(new_n6425_));
  XOR2_X1    g06169(.A1(new_n6425_), .A2(new_n747_), .Z(new_n6426_));
  INV_X1     g06170(.I(new_n6194_), .ZN(new_n6427_));
  NOR2_X1    g06171(.A1(new_n6189_), .A2(new_n6427_), .ZN(new_n6428_));
  NOR3_X1    g06172(.A1(new_n6195_), .A2(new_n6428_), .A3(new_n6197_), .ZN(new_n6429_));
  XOR2_X1    g06173(.A1(new_n6429_), .A2(new_n6426_), .Z(new_n6430_));
  XNOR2_X1   g06174(.A1(new_n6430_), .A2(new_n6421_), .ZN(new_n6431_));
  OAI22_X1   g06175(.A1(new_n582_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n577_), .ZN(new_n6432_));
  NAND2_X1   g06176(.A1(new_n960_), .A2(\b[43] ), .ZN(new_n6433_));
  AOI21_X1   g06177(.A1(new_n6432_), .A2(new_n6433_), .B(new_n585_), .ZN(new_n6434_));
  NAND2_X1   g06178(.A1(new_n4513_), .A2(new_n6434_), .ZN(new_n6435_));
  XOR2_X1    g06179(.A1(new_n6435_), .A2(\a[11] ), .Z(new_n6436_));
  AOI21_X1   g06180(.A1(new_n6198_), .A2(new_n5987_), .B(new_n5988_), .ZN(new_n6437_));
  XOR2_X1    g06181(.A1(new_n6437_), .A2(new_n6436_), .Z(new_n6438_));
  XOR2_X1    g06182(.A1(new_n6431_), .A2(new_n6438_), .Z(new_n6439_));
  OAI22_X1   g06183(.A1(new_n437_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n431_), .ZN(new_n6440_));
  NAND2_X1   g06184(.A1(new_n775_), .A2(\b[46] ), .ZN(new_n6441_));
  AOI21_X1   g06185(.A1(new_n6440_), .A2(new_n6441_), .B(new_n440_), .ZN(new_n6442_));
  NAND2_X1   g06186(.A1(new_n5177_), .A2(new_n6442_), .ZN(new_n6443_));
  XOR2_X1    g06187(.A1(new_n6443_), .A2(\a[8] ), .Z(new_n6444_));
  NAND2_X1   g06188(.A1(new_n6201_), .A2(new_n5933_), .ZN(new_n6445_));
  XOR2_X1    g06189(.A1(new_n6198_), .A2(new_n5987_), .Z(new_n6446_));
  XOR2_X1    g06190(.A1(new_n6446_), .A2(new_n5988_), .Z(new_n6447_));
  NOR2_X1    g06191(.A1(new_n6447_), .A2(new_n5982_), .ZN(new_n6448_));
  NOR2_X1    g06192(.A1(new_n6445_), .A2(new_n6448_), .ZN(new_n6449_));
  XOR2_X1    g06193(.A1(new_n6449_), .A2(new_n6444_), .Z(new_n6450_));
  XOR2_X1    g06194(.A1(new_n6450_), .A2(new_n6439_), .Z(new_n6451_));
  NOR2_X1    g06195(.A1(new_n6451_), .A2(new_n6249_), .ZN(new_n6452_));
  INV_X1     g06196(.I(new_n6452_), .ZN(new_n6453_));
  NAND2_X1   g06197(.A1(new_n6451_), .A2(new_n6249_), .ZN(new_n6454_));
  NAND2_X1   g06198(.A1(new_n6453_), .A2(new_n6454_), .ZN(new_n6455_));
  AND2_X2    g06199(.A1(new_n6455_), .A2(new_n6243_), .Z(new_n6456_));
  NOR2_X1    g06200(.A1(new_n6455_), .A2(new_n6243_), .ZN(new_n6457_));
  NOR2_X1    g06201(.A1(new_n6456_), .A2(new_n6457_), .ZN(new_n6458_));
  INV_X1     g06202(.I(new_n6458_), .ZN(new_n6459_));
  INV_X1     g06203(.I(new_n6214_), .ZN(new_n6460_));
  NAND2_X1   g06204(.A1(new_n5976_), .A2(new_n6460_), .ZN(new_n6461_));
  XOR2_X1    g06205(.A1(new_n6461_), .A2(new_n6459_), .Z(new_n6462_));
  INV_X1     g06206(.I(new_n6224_), .ZN(new_n6463_));
  XOR2_X1    g06207(.A1(new_n5976_), .A2(new_n6460_), .Z(new_n6464_));
  NAND2_X1   g06208(.A1(new_n6464_), .A2(new_n6463_), .ZN(new_n6465_));
  XOR2_X1    g06209(.A1(new_n6462_), .A2(new_n6465_), .Z(\f[54] ));
  INV_X1     g06210(.I(\b[55] ), .ZN(new_n6467_));
  XOR2_X1    g06211(.A1(new_n6232_), .A2(\b[53] ), .Z(new_n6468_));
  AND3_X2    g06212(.A1(new_n6468_), .A2(new_n6467_), .A3(new_n6234_), .Z(new_n6469_));
  AOI21_X1   g06213(.A1(new_n6468_), .A2(new_n6234_), .B(new_n6467_), .ZN(new_n6470_));
  OR2_X2     g06214(.A1(new_n6469_), .A2(new_n6470_), .Z(new_n6471_));
  NOR2_X1    g06215(.A1(new_n405_), .A2(new_n6467_), .ZN(new_n6472_));
  NOR2_X1    g06216(.A1(new_n280_), .A2(new_n6215_), .ZN(new_n6473_));
  NOR2_X1    g06217(.A1(new_n404_), .A2(new_n6238_), .ZN(new_n6474_));
  NOR4_X1    g06218(.A1(new_n6472_), .A2(new_n264_), .A3(new_n6473_), .A4(new_n6474_), .ZN(new_n6475_));
  NAND2_X1   g06219(.A1(new_n6471_), .A2(new_n6475_), .ZN(new_n6476_));
  XOR2_X1    g06220(.A1(new_n6439_), .A2(new_n6444_), .Z(new_n6477_));
  NAND2_X1   g06221(.A1(new_n6477_), .A2(new_n6444_), .ZN(new_n6478_));
  NAND2_X1   g06222(.A1(new_n6449_), .A2(new_n6477_), .ZN(new_n6479_));
  NAND2_X1   g06223(.A1(new_n6479_), .A2(new_n6478_), .ZN(new_n6480_));
  INV_X1     g06224(.I(new_n6480_), .ZN(new_n6481_));
  XOR2_X1    g06225(.A1(new_n6403_), .A2(new_n6408_), .Z(new_n6482_));
  NAND2_X1   g06226(.A1(new_n6482_), .A2(new_n6408_), .ZN(new_n6483_));
  NAND2_X1   g06227(.A1(new_n6482_), .A2(new_n6409_), .ZN(new_n6484_));
  OAI22_X1   g06228(.A1(new_n2452_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n2447_), .ZN(new_n6485_));
  NAND2_X1   g06229(.A1(new_n3312_), .A2(\b[23] ), .ZN(new_n6486_));
  AOI21_X1   g06230(.A1(new_n6485_), .A2(new_n6486_), .B(new_n2455_), .ZN(new_n6487_));
  AND3_X2    g06231(.A1(new_n1828_), .A2(new_n2442_), .A3(new_n6487_), .Z(new_n6488_));
  AOI21_X1   g06232(.A1(new_n1828_), .A2(new_n6487_), .B(new_n2442_), .ZN(new_n6489_));
  NOR2_X1    g06233(.A1(new_n6488_), .A2(new_n6489_), .ZN(new_n6490_));
  NAND3_X1   g06234(.A1(new_n6350_), .A2(new_n6351_), .A3(new_n6352_), .ZN(new_n6491_));
  OAI21_X1   g06235(.A1(new_n6250_), .A2(new_n6353_), .B(new_n6491_), .ZN(new_n6492_));
  AOI21_X1   g06236(.A1(new_n6281_), .A2(new_n6285_), .B(new_n6291_), .ZN(new_n6493_));
  OAI21_X1   g06237(.A1(new_n6251_), .A2(new_n6493_), .B(new_n6293_), .ZN(new_n6494_));
  INV_X1     g06238(.I(new_n6494_), .ZN(new_n6495_));
  OAI21_X1   g06239(.A1(new_n6282_), .A2(new_n6284_), .B(new_n6295_), .ZN(new_n6496_));
  OAI21_X1   g06240(.A1(new_n6263_), .A2(new_n6257_), .B(new_n6275_), .ZN(new_n6497_));
  OAI22_X1   g06241(.A1(new_n5786_), .A2(new_n393_), .B1(new_n290_), .B2(new_n5792_), .ZN(new_n6498_));
  OAI21_X1   g06242(.A1(new_n292_), .A2(new_n6012_), .B(new_n6498_), .ZN(new_n6499_));
  NAND4_X1   g06243(.A1(new_n6499_), .A2(new_n5783_), .A3(new_n334_), .A4(new_n5795_), .ZN(new_n6500_));
  NAND3_X1   g06244(.A1(new_n6499_), .A2(new_n334_), .A3(new_n5795_), .ZN(new_n6501_));
  NAND2_X1   g06245(.A1(new_n6501_), .A2(\a[53] ), .ZN(new_n6502_));
  NAND2_X1   g06246(.A1(new_n6502_), .A2(new_n6500_), .ZN(new_n6503_));
  XOR2_X1    g06247(.A1(\a[53] ), .A2(\a[54] ), .Z(new_n6504_));
  XNOR2_X1   g06248(.A1(\a[55] ), .A2(\a[56] ), .ZN(new_n6505_));
  AND2_X2    g06249(.A1(new_n6505_), .A2(new_n6504_), .Z(new_n6506_));
  INV_X1     g06250(.I(\a[55] ), .ZN(new_n6507_));
  NAND3_X1   g06251(.A1(new_n6507_), .A2(\a[53] ), .A3(\a[54] ), .ZN(new_n6508_));
  OAI21_X1   g06252(.A1(new_n6507_), .A2(new_n6254_), .B(new_n6508_), .ZN(new_n6509_));
  NAND2_X1   g06253(.A1(new_n6509_), .A2(\b[0] ), .ZN(new_n6510_));
  XNOR2_X1   g06254(.A1(\a[55] ), .A2(\a[56] ), .ZN(new_n6511_));
  NOR2_X1    g06255(.A1(new_n6255_), .A2(new_n6511_), .ZN(new_n6512_));
  NAND3_X1   g06256(.A1(new_n6510_), .A2(new_n6512_), .A3(new_n260_), .ZN(new_n6513_));
  AOI21_X1   g06257(.A1(\b[1] ), .A2(new_n6506_), .B(new_n6513_), .ZN(new_n6514_));
  NOR3_X1    g06258(.A1(new_n6514_), .A2(\a[56] ), .A3(new_n6275_), .ZN(new_n6515_));
  INV_X1     g06259(.I(\a[56] ), .ZN(new_n6516_));
  NAND2_X1   g06260(.A1(new_n6514_), .A2(new_n6516_), .ZN(new_n6517_));
  NAND2_X1   g06261(.A1(new_n6506_), .A2(\b[1] ), .ZN(new_n6518_));
  NAND4_X1   g06262(.A1(new_n6518_), .A2(new_n260_), .A3(new_n6510_), .A4(new_n6512_), .ZN(new_n6519_));
  NAND2_X1   g06263(.A1(new_n6519_), .A2(\a[56] ), .ZN(new_n6520_));
  AOI22_X1   g06264(.A1(new_n6517_), .A2(new_n6520_), .B1(new_n6516_), .B2(new_n6256_), .ZN(new_n6521_));
  NOR2_X1    g06265(.A1(new_n6521_), .A2(new_n6515_), .ZN(new_n6522_));
  XOR2_X1    g06266(.A1(new_n6522_), .A2(new_n6503_), .Z(new_n6523_));
  NAND2_X1   g06267(.A1(new_n6523_), .A2(new_n6497_), .ZN(new_n6524_));
  INV_X1     g06268(.I(new_n6497_), .ZN(new_n6525_));
  NOR2_X1    g06269(.A1(new_n6522_), .A2(new_n6503_), .ZN(new_n6526_));
  INV_X1     g06270(.I(new_n6503_), .ZN(new_n6527_));
  INV_X1     g06271(.I(new_n6515_), .ZN(new_n6528_));
  NOR2_X1    g06272(.A1(new_n6519_), .A2(\a[56] ), .ZN(new_n6529_));
  NOR2_X1    g06273(.A1(new_n6514_), .A2(new_n6516_), .ZN(new_n6530_));
  OAI22_X1   g06274(.A1(new_n6530_), .A2(new_n6529_), .B1(\a[56] ), .B2(new_n6275_), .ZN(new_n6531_));
  NAND2_X1   g06275(.A1(new_n6531_), .A2(new_n6528_), .ZN(new_n6532_));
  NOR2_X1    g06276(.A1(new_n6527_), .A2(new_n6532_), .ZN(new_n6533_));
  OAI21_X1   g06277(.A1(new_n6526_), .A2(new_n6533_), .B(new_n6525_), .ZN(new_n6534_));
  NAND2_X1   g06278(.A1(new_n6524_), .A2(new_n6534_), .ZN(new_n6535_));
  OAI22_X1   g06279(.A1(new_n5228_), .A2(new_n450_), .B1(new_n403_), .B2(new_n5225_), .ZN(new_n6536_));
  NAND2_X1   g06280(.A1(new_n5387_), .A2(\b[5] ), .ZN(new_n6537_));
  AOI21_X1   g06281(.A1(new_n6536_), .A2(new_n6537_), .B(new_n5231_), .ZN(new_n6538_));
  NAND2_X1   g06282(.A1(new_n454_), .A2(new_n6538_), .ZN(new_n6539_));
  XOR2_X1    g06283(.A1(new_n6539_), .A2(\a[50] ), .Z(new_n6540_));
  XOR2_X1    g06284(.A1(new_n6535_), .A2(new_n6540_), .Z(new_n6541_));
  NAND2_X1   g06285(.A1(new_n6541_), .A2(new_n6496_), .ZN(new_n6542_));
  AOI21_X1   g06286(.A1(new_n6252_), .A2(new_n6296_), .B(new_n6283_), .ZN(new_n6543_));
  XOR2_X1    g06287(.A1(new_n6539_), .A2(new_n5220_), .Z(new_n6544_));
  XOR2_X1    g06288(.A1(new_n6535_), .A2(new_n6544_), .Z(new_n6545_));
  NAND2_X1   g06289(.A1(new_n6545_), .A2(new_n6543_), .ZN(new_n6546_));
  NAND2_X1   g06290(.A1(new_n6542_), .A2(new_n6546_), .ZN(new_n6547_));
  OAI22_X1   g06291(.A1(new_n4711_), .A2(new_n617_), .B1(new_n510_), .B2(new_n4706_), .ZN(new_n6548_));
  NAND2_X1   g06292(.A1(new_n5814_), .A2(\b[8] ), .ZN(new_n6549_));
  AOI21_X1   g06293(.A1(new_n6548_), .A2(new_n6549_), .B(new_n4714_), .ZN(new_n6550_));
  NAND2_X1   g06294(.A1(new_n616_), .A2(new_n6550_), .ZN(new_n6551_));
  XOR2_X1    g06295(.A1(new_n6551_), .A2(\a[47] ), .Z(new_n6552_));
  INV_X1     g06296(.I(new_n6552_), .ZN(new_n6553_));
  XOR2_X1    g06297(.A1(new_n6547_), .A2(new_n6553_), .Z(new_n6554_));
  NOR2_X1    g06298(.A1(new_n6554_), .A2(new_n6495_), .ZN(new_n6555_));
  XOR2_X1    g06299(.A1(new_n6547_), .A2(new_n6553_), .Z(new_n6556_));
  NAND2_X1   g06300(.A1(new_n6556_), .A2(new_n6495_), .ZN(new_n6557_));
  INV_X1     g06301(.I(new_n6557_), .ZN(new_n6558_));
  OAI22_X1   g06302(.A1(new_n4208_), .A2(new_n795_), .B1(new_n717_), .B2(new_n4203_), .ZN(new_n6559_));
  NAND2_X1   g06303(.A1(new_n5244_), .A2(\b[11] ), .ZN(new_n6560_));
  AOI21_X1   g06304(.A1(new_n6559_), .A2(new_n6560_), .B(new_n4211_), .ZN(new_n6561_));
  NAND2_X1   g06305(.A1(new_n799_), .A2(new_n6561_), .ZN(new_n6562_));
  XOR2_X1    g06306(.A1(new_n6562_), .A2(\a[44] ), .Z(new_n6563_));
  INV_X1     g06307(.I(new_n6563_), .ZN(new_n6564_));
  OAI21_X1   g06308(.A1(new_n6558_), .A2(new_n6555_), .B(new_n6564_), .ZN(new_n6565_));
  INV_X1     g06309(.I(new_n6555_), .ZN(new_n6566_));
  NAND3_X1   g06310(.A1(new_n6566_), .A2(new_n6557_), .A3(new_n6563_), .ZN(new_n6567_));
  OAI22_X1   g06311(.A1(new_n3736_), .A2(new_n992_), .B1(new_n904_), .B2(new_n3731_), .ZN(new_n6568_));
  NAND2_X1   g06312(.A1(new_n4730_), .A2(\b[14] ), .ZN(new_n6569_));
  AOI21_X1   g06313(.A1(new_n6568_), .A2(new_n6569_), .B(new_n3739_), .ZN(new_n6570_));
  NAND2_X1   g06314(.A1(new_n991_), .A2(new_n6570_), .ZN(new_n6571_));
  XOR2_X1    g06315(.A1(new_n6571_), .A2(\a[41] ), .Z(new_n6572_));
  INV_X1     g06316(.I(new_n6572_), .ZN(new_n6573_));
  NAND3_X1   g06317(.A1(new_n6565_), .A2(new_n6567_), .A3(new_n6573_), .ZN(new_n6574_));
  INV_X1     g06318(.I(new_n6574_), .ZN(new_n6575_));
  AOI21_X1   g06319(.A1(new_n6565_), .A2(new_n6567_), .B(new_n6573_), .ZN(new_n6576_));
  OAI22_X1   g06320(.A1(new_n3298_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n3293_), .ZN(new_n6577_));
  NAND2_X1   g06321(.A1(new_n4227_), .A2(\b[17] ), .ZN(new_n6578_));
  AOI21_X1   g06322(.A1(new_n6577_), .A2(new_n6578_), .B(new_n3301_), .ZN(new_n6579_));
  NAND2_X1   g06323(.A1(new_n1225_), .A2(new_n6579_), .ZN(new_n6580_));
  XOR2_X1    g06324(.A1(new_n6580_), .A2(\a[38] ), .Z(new_n6581_));
  NOR3_X1    g06325(.A1(new_n6581_), .A2(new_n6575_), .A3(new_n6576_), .ZN(new_n6582_));
  INV_X1     g06326(.I(new_n6576_), .ZN(new_n6583_));
  XOR2_X1    g06327(.A1(new_n6580_), .A2(new_n3288_), .Z(new_n6584_));
  AOI21_X1   g06328(.A1(new_n6583_), .A2(new_n6574_), .B(new_n6584_), .ZN(new_n6585_));
  OAI21_X1   g06329(.A1(new_n6582_), .A2(new_n6585_), .B(new_n6492_), .ZN(new_n6586_));
  NAND2_X1   g06330(.A1(new_n6116_), .A2(new_n5991_), .ZN(new_n6587_));
  NAND2_X1   g06331(.A1(new_n6587_), .A2(new_n6115_), .ZN(new_n6588_));
  OAI21_X1   g06332(.A1(new_n6341_), .A2(new_n6337_), .B(new_n6347_), .ZN(new_n6589_));
  AOI21_X1   g06333(.A1(new_n6588_), .A2(new_n6589_), .B(new_n6349_), .ZN(new_n6590_));
  NOR2_X1    g06334(.A1(new_n6575_), .A2(new_n6576_), .ZN(new_n6591_));
  XOR2_X1    g06335(.A1(new_n6591_), .A2(new_n6584_), .Z(new_n6592_));
  NAND2_X1   g06336(.A1(new_n6592_), .A2(new_n6590_), .ZN(new_n6593_));
  OAI22_X1   g06337(.A1(new_n2846_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n2841_), .ZN(new_n6594_));
  NAND2_X1   g06338(.A1(new_n3755_), .A2(\b[20] ), .ZN(new_n6595_));
  AOI21_X1   g06339(.A1(new_n6594_), .A2(new_n6595_), .B(new_n2849_), .ZN(new_n6596_));
  NAND2_X1   g06340(.A1(new_n1517_), .A2(new_n6596_), .ZN(new_n6597_));
  XOR2_X1    g06341(.A1(new_n6597_), .A2(\a[35] ), .Z(new_n6598_));
  AOI21_X1   g06342(.A1(new_n6586_), .A2(new_n6593_), .B(new_n6598_), .ZN(new_n6599_));
  NAND3_X1   g06343(.A1(new_n6586_), .A2(new_n6593_), .A3(new_n6598_), .ZN(new_n6600_));
  INV_X1     g06344(.I(new_n6600_), .ZN(new_n6601_));
  OAI21_X1   g06345(.A1(new_n6601_), .A2(new_n6599_), .B(new_n6490_), .ZN(new_n6602_));
  INV_X1     g06346(.I(new_n6490_), .ZN(new_n6603_));
  INV_X1     g06347(.I(new_n6599_), .ZN(new_n6604_));
  NAND3_X1   g06348(.A1(new_n6604_), .A2(new_n6603_), .A3(new_n6600_), .ZN(new_n6605_));
  NAND2_X1   g06349(.A1(new_n6605_), .A2(new_n6602_), .ZN(new_n6606_));
  OAI22_X1   g06350(.A1(new_n2084_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n2079_), .ZN(new_n6607_));
  NAND2_X1   g06351(.A1(new_n2864_), .A2(\b[26] ), .ZN(new_n6608_));
  AOI21_X1   g06352(.A1(new_n6607_), .A2(new_n6608_), .B(new_n2087_), .ZN(new_n6609_));
  NAND2_X1   g06353(.A1(new_n2174_), .A2(new_n6609_), .ZN(new_n6610_));
  XOR2_X1    g06354(.A1(new_n6610_), .A2(\a[29] ), .Z(new_n6611_));
  XOR2_X1    g06355(.A1(new_n6606_), .A2(new_n6611_), .Z(new_n6612_));
  OAI22_X1   g06356(.A1(new_n1760_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n1755_), .ZN(new_n6613_));
  NAND2_X1   g06357(.A1(new_n2470_), .A2(\b[29] ), .ZN(new_n6614_));
  AOI21_X1   g06358(.A1(new_n6613_), .A2(new_n6614_), .B(new_n1763_), .ZN(new_n6615_));
  NAND2_X1   g06359(.A1(new_n2546_), .A2(new_n6615_), .ZN(new_n6616_));
  XOR2_X1    g06360(.A1(new_n6616_), .A2(\a[26] ), .Z(new_n6617_));
  XOR2_X1    g06361(.A1(new_n6617_), .A2(new_n6612_), .Z(new_n6618_));
  OAI22_X1   g06362(.A1(new_n1444_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n1439_), .ZN(new_n6619_));
  NAND2_X1   g06363(.A1(new_n2098_), .A2(\b[32] ), .ZN(new_n6620_));
  AOI21_X1   g06364(.A1(new_n6619_), .A2(new_n6620_), .B(new_n1447_), .ZN(new_n6621_));
  NAND2_X1   g06365(.A1(new_n2963_), .A2(new_n6621_), .ZN(new_n6622_));
  XOR2_X1    g06366(.A1(new_n6622_), .A2(\a[23] ), .Z(new_n6623_));
  XOR2_X1    g06367(.A1(new_n6618_), .A2(new_n6623_), .Z(new_n6624_));
  INV_X1     g06368(.I(new_n6624_), .ZN(new_n6625_));
  OAI22_X1   g06369(.A1(new_n1168_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n1163_), .ZN(new_n6626_));
  NAND2_X1   g06370(.A1(new_n1774_), .A2(\b[35] ), .ZN(new_n6627_));
  AOI21_X1   g06371(.A1(new_n6626_), .A2(new_n6627_), .B(new_n1171_), .ZN(new_n6628_));
  NAND2_X1   g06372(.A1(new_n3411_), .A2(new_n6628_), .ZN(new_n6629_));
  XOR2_X1    g06373(.A1(new_n6629_), .A2(\a[20] ), .Z(new_n6630_));
  NOR2_X1    g06374(.A1(new_n6625_), .A2(new_n6630_), .ZN(new_n6631_));
  NAND2_X1   g06375(.A1(new_n6625_), .A2(new_n6630_), .ZN(new_n6632_));
  INV_X1     g06376(.I(new_n6632_), .ZN(new_n6633_));
  NOR2_X1    g06377(.A1(new_n6633_), .A2(new_n6631_), .ZN(new_n6634_));
  OAI22_X1   g06378(.A1(new_n940_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n935_), .ZN(new_n6635_));
  NAND2_X1   g06379(.A1(new_n1458_), .A2(\b[38] ), .ZN(new_n6636_));
  AOI21_X1   g06380(.A1(new_n6635_), .A2(new_n6636_), .B(new_n943_), .ZN(new_n6637_));
  NAND2_X1   g06381(.A1(new_n3844_), .A2(new_n6637_), .ZN(new_n6638_));
  XOR2_X1    g06382(.A1(new_n6638_), .A2(\a[17] ), .Z(new_n6639_));
  XOR2_X1    g06383(.A1(new_n6634_), .A2(new_n6639_), .Z(new_n6640_));
  AOI21_X1   g06384(.A1(new_n6483_), .A2(new_n6484_), .B(new_n6640_), .ZN(new_n6641_));
  NAND2_X1   g06385(.A1(new_n6483_), .A2(new_n6484_), .ZN(new_n6642_));
  INV_X1     g06386(.I(new_n6639_), .ZN(new_n6643_));
  XOR2_X1    g06387(.A1(new_n6634_), .A2(new_n6643_), .Z(new_n6644_));
  NOR2_X1    g06388(.A1(new_n6642_), .A2(new_n6644_), .ZN(new_n6645_));
  NOR2_X1    g06389(.A1(new_n6645_), .A2(new_n6641_), .ZN(new_n6646_));
  OAI22_X1   g06390(.A1(new_n757_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n752_), .ZN(new_n6647_));
  NAND2_X1   g06391(.A1(new_n1182_), .A2(\b[41] ), .ZN(new_n6648_));
  AOI21_X1   g06392(.A1(new_n6647_), .A2(new_n6648_), .B(new_n760_), .ZN(new_n6649_));
  NAND2_X1   g06393(.A1(new_n4320_), .A2(new_n6649_), .ZN(new_n6650_));
  XOR2_X1    g06394(.A1(new_n6650_), .A2(\a[14] ), .Z(new_n6651_));
  XOR2_X1    g06395(.A1(new_n6646_), .A2(new_n6651_), .Z(new_n6652_));
  OAI22_X1   g06396(.A1(new_n582_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n577_), .ZN(new_n6653_));
  NAND2_X1   g06397(.A1(new_n960_), .A2(\b[44] ), .ZN(new_n6654_));
  AOI21_X1   g06398(.A1(new_n6653_), .A2(new_n6654_), .B(new_n585_), .ZN(new_n6655_));
  NAND2_X1   g06399(.A1(new_n4833_), .A2(new_n6655_), .ZN(new_n6656_));
  XOR2_X1    g06400(.A1(new_n6656_), .A2(\a[11] ), .Z(new_n6657_));
  XOR2_X1    g06401(.A1(new_n6652_), .A2(new_n6657_), .Z(new_n6658_));
  OAI22_X1   g06402(.A1(new_n437_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n431_), .ZN(new_n6659_));
  NAND2_X1   g06403(.A1(new_n775_), .A2(\b[47] ), .ZN(new_n6660_));
  AOI21_X1   g06404(.A1(new_n6659_), .A2(new_n6660_), .B(new_n440_), .ZN(new_n6661_));
  NAND2_X1   g06405(.A1(new_n5196_), .A2(new_n6661_), .ZN(new_n6662_));
  XOR2_X1    g06406(.A1(new_n6662_), .A2(\a[8] ), .Z(new_n6663_));
  XOR2_X1    g06407(.A1(new_n6658_), .A2(new_n6663_), .Z(new_n6664_));
  OAI22_X1   g06408(.A1(new_n364_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n320_), .ZN(new_n6665_));
  NAND2_X1   g06409(.A1(new_n594_), .A2(\b[50] ), .ZN(new_n6666_));
  AOI21_X1   g06410(.A1(new_n6665_), .A2(new_n6666_), .B(new_n312_), .ZN(new_n6667_));
  NAND2_X1   g06411(.A1(new_n5954_), .A2(new_n6667_), .ZN(new_n6668_));
  XOR2_X1    g06412(.A1(new_n6668_), .A2(\a[5] ), .Z(new_n6669_));
  INV_X1     g06413(.I(new_n6669_), .ZN(new_n6670_));
  XOR2_X1    g06414(.A1(new_n6664_), .A2(new_n6670_), .Z(new_n6671_));
  NOR2_X1    g06415(.A1(new_n6481_), .A2(new_n6671_), .ZN(new_n6672_));
  XOR2_X1    g06416(.A1(new_n6664_), .A2(new_n6669_), .Z(new_n6673_));
  NOR2_X1    g06417(.A1(new_n6480_), .A2(new_n6673_), .ZN(new_n6674_));
  NOR2_X1    g06418(.A1(new_n6672_), .A2(new_n6674_), .ZN(new_n6675_));
  INV_X1     g06419(.I(new_n6675_), .ZN(new_n6676_));
  XOR2_X1    g06420(.A1(new_n6454_), .A2(new_n6676_), .Z(new_n6677_));
  XOR2_X1    g06421(.A1(new_n6677_), .A2(\a[2] ), .Z(new_n6678_));
  XNOR2_X1   g06422(.A1(new_n6678_), .A2(new_n6476_), .ZN(new_n6679_));
  INV_X1     g06423(.I(new_n6679_), .ZN(new_n6680_));
  INV_X1     g06424(.I(new_n5976_), .ZN(new_n6681_));
  NOR2_X1    g06425(.A1(new_n6459_), .A2(new_n6224_), .ZN(new_n6682_));
  NOR3_X1    g06426(.A1(new_n6681_), .A2(new_n6214_), .A3(new_n6682_), .ZN(new_n6683_));
  NOR2_X1    g06427(.A1(new_n6683_), .A2(new_n6456_), .ZN(new_n6684_));
  OR2_X2     g06428(.A1(new_n6679_), .A2(new_n6456_), .Z(new_n6685_));
  OAI22_X1   g06429(.A1(new_n6684_), .A2(new_n6680_), .B1(new_n6683_), .B2(new_n6685_), .ZN(\f[55] ));
  XOR2_X1    g06430(.A1(new_n6476_), .A2(new_n271_), .Z(new_n6687_));
  NOR2_X1    g06431(.A1(new_n6684_), .A2(new_n6679_), .ZN(new_n6688_));
  AOI21_X1   g06432(.A1(new_n6677_), .A2(new_n6687_), .B(new_n6688_), .ZN(new_n6689_));
  NOR2_X1    g06433(.A1(new_n6652_), .A2(new_n6657_), .ZN(new_n6690_));
  OAI22_X1   g06434(.A1(new_n582_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n577_), .ZN(new_n6691_));
  NAND2_X1   g06435(.A1(new_n960_), .A2(\b[45] ), .ZN(new_n6692_));
  AOI21_X1   g06436(.A1(new_n6691_), .A2(new_n6692_), .B(new_n585_), .ZN(new_n6693_));
  NAND2_X1   g06437(.A1(new_n5004_), .A2(new_n6693_), .ZN(new_n6694_));
  XOR2_X1    g06438(.A1(new_n6694_), .A2(\a[11] ), .Z(new_n6695_));
  OAI22_X1   g06439(.A1(new_n757_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n752_), .ZN(new_n6696_));
  NAND2_X1   g06440(.A1(new_n1182_), .A2(\b[42] ), .ZN(new_n6697_));
  AOI21_X1   g06441(.A1(new_n6696_), .A2(new_n6697_), .B(new_n760_), .ZN(new_n6698_));
  NAND2_X1   g06442(.A1(new_n4500_), .A2(new_n6698_), .ZN(new_n6699_));
  XOR2_X1    g06443(.A1(new_n6699_), .A2(\a[14] ), .Z(new_n6700_));
  INV_X1     g06444(.I(new_n6651_), .ZN(new_n6701_));
  NAND2_X1   g06445(.A1(new_n6646_), .A2(new_n6701_), .ZN(new_n6702_));
  OAI22_X1   g06446(.A1(new_n2084_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n2079_), .ZN(new_n6703_));
  NAND2_X1   g06447(.A1(new_n2864_), .A2(\b[27] ), .ZN(new_n6704_));
  AOI21_X1   g06448(.A1(new_n6703_), .A2(new_n6704_), .B(new_n2087_), .ZN(new_n6705_));
  NAND2_X1   g06449(.A1(new_n2276_), .A2(new_n6705_), .ZN(new_n6706_));
  XOR2_X1    g06450(.A1(new_n6706_), .A2(\a[29] ), .Z(new_n6707_));
  OAI22_X1   g06451(.A1(new_n2452_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n2447_), .ZN(new_n6708_));
  NAND2_X1   g06452(.A1(new_n3312_), .A2(\b[24] ), .ZN(new_n6709_));
  AOI21_X1   g06453(.A1(new_n6708_), .A2(new_n6709_), .B(new_n2455_), .ZN(new_n6710_));
  NAND2_X1   g06454(.A1(new_n1926_), .A2(new_n6710_), .ZN(new_n6711_));
  XOR2_X1    g06455(.A1(new_n6711_), .A2(\a[32] ), .Z(new_n6712_));
  INV_X1     g06456(.I(new_n6712_), .ZN(new_n6713_));
  INV_X1     g06457(.I(new_n6582_), .ZN(new_n6714_));
  OAI21_X1   g06458(.A1(new_n6590_), .A2(new_n6585_), .B(new_n6714_), .ZN(new_n6715_));
  AOI21_X1   g06459(.A1(new_n6565_), .A2(new_n6567_), .B(new_n6572_), .ZN(new_n6716_));
  INV_X1     g06460(.I(new_n6535_), .ZN(new_n6717_));
  NAND2_X1   g06461(.A1(new_n6527_), .A2(new_n6532_), .ZN(new_n6718_));
  AOI21_X1   g06462(.A1(new_n6497_), .A2(new_n6718_), .B(new_n6533_), .ZN(new_n6719_));
  NAND4_X1   g06463(.A1(new_n6519_), .A2(new_n6516_), .A3(new_n258_), .A4(new_n6255_), .ZN(new_n6720_));
  INV_X1     g06464(.I(new_n6509_), .ZN(new_n6721_));
  NOR2_X1    g06465(.A1(new_n6721_), .A2(new_n267_), .ZN(new_n6722_));
  NAND2_X1   g06466(.A1(new_n6505_), .A2(new_n6504_), .ZN(new_n6723_));
  NOR2_X1    g06467(.A1(new_n6723_), .A2(new_n292_), .ZN(new_n6724_));
  XNOR2_X1   g06468(.A1(\a[53] ), .A2(\a[54] ), .ZN(new_n6725_));
  XNOR2_X1   g06469(.A1(\a[53] ), .A2(\a[55] ), .ZN(new_n6726_));
  NAND2_X1   g06470(.A1(new_n6725_), .A2(new_n6726_), .ZN(new_n6727_));
  XNOR2_X1   g06471(.A1(\a[53] ), .A2(\a[56] ), .ZN(new_n6728_));
  NAND2_X1   g06472(.A1(new_n6727_), .A2(new_n6728_), .ZN(new_n6729_));
  OAI22_X1   g06473(.A1(new_n6722_), .A2(new_n6724_), .B1(new_n6729_), .B2(new_n258_), .ZN(new_n6730_));
  INV_X1     g06474(.I(new_n6512_), .ZN(new_n6731_));
  NOR2_X1    g06475(.A1(new_n6731_), .A2(new_n278_), .ZN(new_n6732_));
  NAND3_X1   g06476(.A1(new_n6730_), .A2(new_n6516_), .A3(new_n6732_), .ZN(new_n6733_));
  AOI21_X1   g06477(.A1(new_n6730_), .A2(new_n6732_), .B(new_n6516_), .ZN(new_n6734_));
  INV_X1     g06478(.I(new_n6734_), .ZN(new_n6735_));
  AOI21_X1   g06479(.A1(new_n6735_), .A2(new_n6733_), .B(new_n6720_), .ZN(new_n6736_));
  NOR4_X1    g06480(.A1(new_n6514_), .A2(\a[56] ), .A3(\b[0] ), .A4(new_n6504_), .ZN(new_n6737_));
  INV_X1     g06481(.I(new_n6733_), .ZN(new_n6738_));
  NOR3_X1    g06482(.A1(new_n6738_), .A2(new_n6737_), .A3(new_n6734_), .ZN(new_n6739_));
  NOR2_X1    g06483(.A1(new_n6736_), .A2(new_n6739_), .ZN(new_n6740_));
  NOR2_X1    g06484(.A1(new_n351_), .A2(\b[5] ), .ZN(new_n6741_));
  XOR2_X1    g06485(.A1(new_n330_), .A2(new_n290_), .Z(new_n6742_));
  AOI21_X1   g06486(.A1(new_n6742_), .A2(new_n348_), .B(new_n347_), .ZN(new_n6743_));
  OAI22_X1   g06487(.A1(new_n5786_), .A2(new_n347_), .B1(new_n393_), .B2(new_n5792_), .ZN(new_n6744_));
  INV_X1     g06488(.I(new_n6012_), .ZN(new_n6745_));
  NAND2_X1   g06489(.A1(new_n6745_), .A2(\b[3] ), .ZN(new_n6746_));
  AOI21_X1   g06490(.A1(new_n6746_), .A2(new_n6744_), .B(new_n5796_), .ZN(new_n6747_));
  OAI21_X1   g06491(.A1(new_n6741_), .A2(new_n6743_), .B(new_n6747_), .ZN(new_n6748_));
  XOR2_X1    g06492(.A1(new_n6748_), .A2(new_n5783_), .Z(new_n6749_));
  NAND2_X1   g06493(.A1(new_n6749_), .A2(new_n6740_), .ZN(new_n6750_));
  OR2_X2     g06494(.A1(new_n6736_), .A2(new_n6739_), .Z(new_n6751_));
  NOR2_X1    g06495(.A1(new_n6748_), .A2(\a[53] ), .ZN(new_n6752_));
  AOI21_X1   g06496(.A1(new_n352_), .A2(new_n6747_), .B(new_n5783_), .ZN(new_n6753_));
  NOR2_X1    g06497(.A1(new_n6753_), .A2(new_n6752_), .ZN(new_n6754_));
  NAND2_X1   g06498(.A1(new_n6754_), .A2(new_n6751_), .ZN(new_n6755_));
  AOI21_X1   g06499(.A1(new_n6750_), .A2(new_n6755_), .B(new_n6719_), .ZN(new_n6756_));
  NAND2_X1   g06500(.A1(new_n6522_), .A2(new_n6503_), .ZN(new_n6757_));
  OAI21_X1   g06501(.A1(new_n6525_), .A2(new_n6526_), .B(new_n6757_), .ZN(new_n6758_));
  NAND2_X1   g06502(.A1(new_n6749_), .A2(new_n6751_), .ZN(new_n6759_));
  NAND2_X1   g06503(.A1(new_n6754_), .A2(new_n6740_), .ZN(new_n6760_));
  AOI21_X1   g06504(.A1(new_n6759_), .A2(new_n6760_), .B(new_n6758_), .ZN(new_n6761_));
  OAI22_X1   g06505(.A1(new_n5228_), .A2(new_n495_), .B1(new_n450_), .B2(new_n5225_), .ZN(new_n6762_));
  NAND2_X1   g06506(.A1(new_n5387_), .A2(\b[6] ), .ZN(new_n6763_));
  AOI21_X1   g06507(.A1(new_n6762_), .A2(new_n6763_), .B(new_n5231_), .ZN(new_n6764_));
  OAI21_X1   g06508(.A1(new_n493_), .A2(new_n490_), .B(new_n6764_), .ZN(new_n6765_));
  XOR2_X1    g06509(.A1(new_n6765_), .A2(\a[50] ), .Z(new_n6766_));
  NOR3_X1    g06510(.A1(new_n6756_), .A2(new_n6761_), .A3(new_n6766_), .ZN(new_n6767_));
  NOR2_X1    g06511(.A1(new_n6754_), .A2(new_n6751_), .ZN(new_n6768_));
  NOR3_X1    g06512(.A1(new_n6740_), .A2(new_n6753_), .A3(new_n6752_), .ZN(new_n6769_));
  OAI21_X1   g06513(.A1(new_n6768_), .A2(new_n6769_), .B(new_n6758_), .ZN(new_n6770_));
  NAND2_X1   g06514(.A1(new_n6759_), .A2(new_n6760_), .ZN(new_n6771_));
  NAND2_X1   g06515(.A1(new_n6771_), .A2(new_n6719_), .ZN(new_n6772_));
  INV_X1     g06516(.I(new_n6766_), .ZN(new_n6773_));
  AOI21_X1   g06517(.A1(new_n6772_), .A2(new_n6770_), .B(new_n6773_), .ZN(new_n6774_));
  NOR2_X1    g06518(.A1(new_n6774_), .A2(new_n6767_), .ZN(new_n6775_));
  NAND2_X1   g06519(.A1(new_n6543_), .A2(new_n6544_), .ZN(new_n6776_));
  NAND2_X1   g06520(.A1(new_n6496_), .A2(new_n6540_), .ZN(new_n6777_));
  NAND2_X1   g06521(.A1(new_n6776_), .A2(new_n6777_), .ZN(new_n6778_));
  NAND3_X1   g06522(.A1(new_n6778_), .A2(new_n6717_), .A3(new_n6775_), .ZN(new_n6779_));
  NAND3_X1   g06523(.A1(new_n6772_), .A2(new_n6770_), .A3(new_n6773_), .ZN(new_n6780_));
  OAI21_X1   g06524(.A1(new_n6756_), .A2(new_n6761_), .B(new_n6766_), .ZN(new_n6781_));
  NAND2_X1   g06525(.A1(new_n6780_), .A2(new_n6781_), .ZN(new_n6782_));
  NOR2_X1    g06526(.A1(new_n6496_), .A2(new_n6540_), .ZN(new_n6783_));
  NOR2_X1    g06527(.A1(new_n6543_), .A2(new_n6544_), .ZN(new_n6784_));
  OAI21_X1   g06528(.A1(new_n6784_), .A2(new_n6783_), .B(new_n6717_), .ZN(new_n6785_));
  NAND2_X1   g06529(.A1(new_n6785_), .A2(new_n6782_), .ZN(new_n6786_));
  NOR2_X1    g06530(.A1(new_n6543_), .A2(new_n6540_), .ZN(new_n6787_));
  NAND3_X1   g06531(.A1(new_n6786_), .A2(new_n6779_), .A3(new_n6787_), .ZN(new_n6788_));
  NOR2_X1    g06532(.A1(new_n6785_), .A2(new_n6782_), .ZN(new_n6789_));
  AOI21_X1   g06533(.A1(new_n6776_), .A2(new_n6777_), .B(new_n6535_), .ZN(new_n6790_));
  NOR2_X1    g06534(.A1(new_n6790_), .A2(new_n6775_), .ZN(new_n6791_));
  NAND2_X1   g06535(.A1(new_n6496_), .A2(new_n6544_), .ZN(new_n6792_));
  OAI21_X1   g06536(.A1(new_n6789_), .A2(new_n6791_), .B(new_n6792_), .ZN(new_n6793_));
  OAI22_X1   g06537(.A1(new_n4711_), .A2(new_n659_), .B1(new_n617_), .B2(new_n4706_), .ZN(new_n6794_));
  NAND2_X1   g06538(.A1(new_n5814_), .A2(\b[9] ), .ZN(new_n6795_));
  AOI21_X1   g06539(.A1(new_n6794_), .A2(new_n6795_), .B(new_n4714_), .ZN(new_n6796_));
  NAND2_X1   g06540(.A1(new_n663_), .A2(new_n6796_), .ZN(new_n6797_));
  XOR2_X1    g06541(.A1(new_n6797_), .A2(\a[47] ), .Z(new_n6798_));
  AOI21_X1   g06542(.A1(new_n6793_), .A2(new_n6788_), .B(new_n6798_), .ZN(new_n6799_));
  NOR3_X1    g06543(.A1(new_n6789_), .A2(new_n6791_), .A3(new_n6792_), .ZN(new_n6800_));
  AOI21_X1   g06544(.A1(new_n6786_), .A2(new_n6779_), .B(new_n6787_), .ZN(new_n6801_));
  INV_X1     g06545(.I(new_n6798_), .ZN(new_n6802_));
  NOR3_X1    g06546(.A1(new_n6800_), .A2(new_n6801_), .A3(new_n6802_), .ZN(new_n6803_));
  INV_X1     g06547(.I(new_n6547_), .ZN(new_n6804_));
  NOR2_X1    g06548(.A1(new_n6494_), .A2(new_n6552_), .ZN(new_n6805_));
  OAI21_X1   g06549(.A1(new_n6059_), .A2(new_n6061_), .B(new_n6074_), .ZN(new_n6806_));
  NAND2_X1   g06550(.A1(new_n6806_), .A2(new_n6299_), .ZN(new_n6807_));
  AOI21_X1   g06551(.A1(new_n6807_), .A2(new_n6293_), .B(new_n6553_), .ZN(new_n6808_));
  OAI21_X1   g06552(.A1(new_n6805_), .A2(new_n6808_), .B(new_n6804_), .ZN(new_n6809_));
  NOR3_X1    g06553(.A1(new_n6803_), .A2(new_n6799_), .A3(new_n6809_), .ZN(new_n6810_));
  OAI21_X1   g06554(.A1(new_n6800_), .A2(new_n6801_), .B(new_n6802_), .ZN(new_n6811_));
  NAND3_X1   g06555(.A1(new_n6793_), .A2(new_n6788_), .A3(new_n6798_), .ZN(new_n6812_));
  NAND3_X1   g06556(.A1(new_n6807_), .A2(new_n6293_), .A3(new_n6553_), .ZN(new_n6813_));
  NAND2_X1   g06557(.A1(new_n6494_), .A2(new_n6552_), .ZN(new_n6814_));
  AOI21_X1   g06558(.A1(new_n6814_), .A2(new_n6813_), .B(new_n6547_), .ZN(new_n6815_));
  AOI21_X1   g06559(.A1(new_n6811_), .A2(new_n6812_), .B(new_n6815_), .ZN(new_n6816_));
  NOR2_X1    g06560(.A1(new_n6495_), .A2(new_n6552_), .ZN(new_n6817_));
  INV_X1     g06561(.I(new_n6817_), .ZN(new_n6818_));
  NOR3_X1    g06562(.A1(new_n6810_), .A2(new_n6816_), .A3(new_n6818_), .ZN(new_n6819_));
  NAND3_X1   g06563(.A1(new_n6811_), .A2(new_n6812_), .A3(new_n6815_), .ZN(new_n6820_));
  OAI21_X1   g06564(.A1(new_n6803_), .A2(new_n6799_), .B(new_n6809_), .ZN(new_n6821_));
  AOI21_X1   g06565(.A1(new_n6821_), .A2(new_n6820_), .B(new_n6817_), .ZN(new_n6822_));
  OAI22_X1   g06566(.A1(new_n4208_), .A2(new_n848_), .B1(new_n795_), .B2(new_n4203_), .ZN(new_n6823_));
  NAND2_X1   g06567(.A1(new_n5244_), .A2(\b[12] ), .ZN(new_n6824_));
  AOI21_X1   g06568(.A1(new_n6823_), .A2(new_n6824_), .B(new_n4211_), .ZN(new_n6825_));
  NAND2_X1   g06569(.A1(new_n847_), .A2(new_n6825_), .ZN(new_n6826_));
  XOR2_X1    g06570(.A1(new_n6826_), .A2(\a[44] ), .Z(new_n6827_));
  NOR3_X1    g06571(.A1(new_n6819_), .A2(new_n6822_), .A3(new_n6827_), .ZN(new_n6828_));
  NAND3_X1   g06572(.A1(new_n6821_), .A2(new_n6820_), .A3(new_n6817_), .ZN(new_n6829_));
  OAI21_X1   g06573(.A1(new_n6810_), .A2(new_n6816_), .B(new_n6818_), .ZN(new_n6830_));
  INV_X1     g06574(.I(new_n6827_), .ZN(new_n6831_));
  AOI21_X1   g06575(.A1(new_n6830_), .A2(new_n6829_), .B(new_n6831_), .ZN(new_n6832_));
  NOR3_X1    g06576(.A1(new_n6558_), .A2(new_n6555_), .A3(new_n6563_), .ZN(new_n6833_));
  INV_X1     g06577(.I(new_n6833_), .ZN(new_n6834_));
  NOR3_X1    g06578(.A1(new_n6828_), .A2(new_n6832_), .A3(new_n6834_), .ZN(new_n6835_));
  NAND3_X1   g06579(.A1(new_n6830_), .A2(new_n6829_), .A3(new_n6831_), .ZN(new_n6836_));
  OAI21_X1   g06580(.A1(new_n6819_), .A2(new_n6822_), .B(new_n6827_), .ZN(new_n6837_));
  AOI21_X1   g06581(.A1(new_n6837_), .A2(new_n6836_), .B(new_n6833_), .ZN(new_n6838_));
  OAI22_X1   g06582(.A1(new_n3736_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n3731_), .ZN(new_n6839_));
  NAND2_X1   g06583(.A1(new_n4730_), .A2(\b[15] ), .ZN(new_n6840_));
  AOI21_X1   g06584(.A1(new_n6839_), .A2(new_n6840_), .B(new_n3739_), .ZN(new_n6841_));
  NAND2_X1   g06585(.A1(new_n1047_), .A2(new_n6841_), .ZN(new_n6842_));
  XOR2_X1    g06586(.A1(new_n6842_), .A2(\a[41] ), .Z(new_n6843_));
  NOR3_X1    g06587(.A1(new_n6835_), .A2(new_n6838_), .A3(new_n6843_), .ZN(new_n6844_));
  NAND3_X1   g06588(.A1(new_n6837_), .A2(new_n6836_), .A3(new_n6833_), .ZN(new_n6845_));
  OAI21_X1   g06589(.A1(new_n6828_), .A2(new_n6832_), .B(new_n6834_), .ZN(new_n6846_));
  INV_X1     g06590(.I(new_n6843_), .ZN(new_n6847_));
  AOI21_X1   g06591(.A1(new_n6846_), .A2(new_n6845_), .B(new_n6847_), .ZN(new_n6848_));
  OAI21_X1   g06592(.A1(new_n6844_), .A2(new_n6848_), .B(new_n6716_), .ZN(new_n6849_));
  INV_X1     g06593(.I(new_n6716_), .ZN(new_n6850_));
  AOI21_X1   g06594(.A1(new_n6846_), .A2(new_n6845_), .B(new_n6843_), .ZN(new_n6851_));
  NOR3_X1    g06595(.A1(new_n6835_), .A2(new_n6838_), .A3(new_n6847_), .ZN(new_n6852_));
  OAI21_X1   g06596(.A1(new_n6852_), .A2(new_n6851_), .B(new_n6850_), .ZN(new_n6853_));
  OAI22_X1   g06597(.A1(new_n3298_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n3293_), .ZN(new_n6854_));
  NAND2_X1   g06598(.A1(new_n4227_), .A2(\b[18] ), .ZN(new_n6855_));
  AOI21_X1   g06599(.A1(new_n6854_), .A2(new_n6855_), .B(new_n3301_), .ZN(new_n6856_));
  NAND2_X1   g06600(.A1(new_n1304_), .A2(new_n6856_), .ZN(new_n6857_));
  XOR2_X1    g06601(.A1(new_n6857_), .A2(\a[38] ), .Z(new_n6858_));
  AOI21_X1   g06602(.A1(new_n6853_), .A2(new_n6849_), .B(new_n6858_), .ZN(new_n6859_));
  NAND3_X1   g06603(.A1(new_n6846_), .A2(new_n6845_), .A3(new_n6847_), .ZN(new_n6860_));
  OAI21_X1   g06604(.A1(new_n6835_), .A2(new_n6838_), .B(new_n6843_), .ZN(new_n6861_));
  AOI21_X1   g06605(.A1(new_n6861_), .A2(new_n6860_), .B(new_n6850_), .ZN(new_n6862_));
  OAI21_X1   g06606(.A1(new_n6835_), .A2(new_n6838_), .B(new_n6847_), .ZN(new_n6863_));
  NAND3_X1   g06607(.A1(new_n6846_), .A2(new_n6845_), .A3(new_n6843_), .ZN(new_n6864_));
  AOI21_X1   g06608(.A1(new_n6863_), .A2(new_n6864_), .B(new_n6716_), .ZN(new_n6865_));
  INV_X1     g06609(.I(new_n6858_), .ZN(new_n6866_));
  NOR3_X1    g06610(.A1(new_n6862_), .A2(new_n6865_), .A3(new_n6866_), .ZN(new_n6867_));
  OAI21_X1   g06611(.A1(new_n6859_), .A2(new_n6867_), .B(new_n6715_), .ZN(new_n6868_));
  INV_X1     g06612(.I(new_n6585_), .ZN(new_n6869_));
  AOI21_X1   g06613(.A1(new_n6492_), .A2(new_n6869_), .B(new_n6582_), .ZN(new_n6870_));
  NOR3_X1    g06614(.A1(new_n6862_), .A2(new_n6865_), .A3(new_n6858_), .ZN(new_n6871_));
  AOI21_X1   g06615(.A1(new_n6853_), .A2(new_n6849_), .B(new_n6866_), .ZN(new_n6872_));
  OAI21_X1   g06616(.A1(new_n6872_), .A2(new_n6871_), .B(new_n6870_), .ZN(new_n6873_));
  OAI22_X1   g06617(.A1(new_n2846_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n2841_), .ZN(new_n6874_));
  NAND2_X1   g06618(.A1(new_n3755_), .A2(\b[21] ), .ZN(new_n6875_));
  AOI21_X1   g06619(.A1(new_n6874_), .A2(new_n6875_), .B(new_n2849_), .ZN(new_n6876_));
  NAND2_X1   g06620(.A1(new_n1604_), .A2(new_n6876_), .ZN(new_n6877_));
  XOR2_X1    g06621(.A1(new_n6877_), .A2(\a[35] ), .Z(new_n6878_));
  INV_X1     g06622(.I(new_n6878_), .ZN(new_n6879_));
  NAND3_X1   g06623(.A1(new_n6873_), .A2(new_n6868_), .A3(new_n6879_), .ZN(new_n6880_));
  OAI21_X1   g06624(.A1(new_n6862_), .A2(new_n6865_), .B(new_n6866_), .ZN(new_n6881_));
  NAND3_X1   g06625(.A1(new_n6853_), .A2(new_n6849_), .A3(new_n6858_), .ZN(new_n6882_));
  AOI21_X1   g06626(.A1(new_n6881_), .A2(new_n6882_), .B(new_n6870_), .ZN(new_n6883_));
  NAND3_X1   g06627(.A1(new_n6853_), .A2(new_n6849_), .A3(new_n6866_), .ZN(new_n6884_));
  OAI21_X1   g06628(.A1(new_n6862_), .A2(new_n6865_), .B(new_n6858_), .ZN(new_n6885_));
  AOI21_X1   g06629(.A1(new_n6885_), .A2(new_n6884_), .B(new_n6715_), .ZN(new_n6886_));
  OAI21_X1   g06630(.A1(new_n6883_), .A2(new_n6886_), .B(new_n6878_), .ZN(new_n6887_));
  AOI21_X1   g06631(.A1(new_n6887_), .A2(new_n6880_), .B(new_n6604_), .ZN(new_n6888_));
  NOR3_X1    g06632(.A1(new_n6883_), .A2(new_n6886_), .A3(new_n6878_), .ZN(new_n6889_));
  AOI21_X1   g06633(.A1(new_n6873_), .A2(new_n6868_), .B(new_n6879_), .ZN(new_n6890_));
  NOR3_X1    g06634(.A1(new_n6889_), .A2(new_n6890_), .A3(new_n6599_), .ZN(new_n6891_));
  OAI21_X1   g06635(.A1(new_n6891_), .A2(new_n6888_), .B(new_n6602_), .ZN(new_n6892_));
  AOI21_X1   g06636(.A1(new_n6604_), .A2(new_n6600_), .B(new_n6603_), .ZN(new_n6893_));
  OAI21_X1   g06637(.A1(new_n6889_), .A2(new_n6890_), .B(new_n6599_), .ZN(new_n6894_));
  NAND3_X1   g06638(.A1(new_n6887_), .A2(new_n6880_), .A3(new_n6604_), .ZN(new_n6895_));
  NAND3_X1   g06639(.A1(new_n6894_), .A2(new_n6895_), .A3(new_n6893_), .ZN(new_n6896_));
  AOI21_X1   g06640(.A1(new_n6892_), .A2(new_n6896_), .B(new_n6713_), .ZN(new_n6897_));
  AOI21_X1   g06641(.A1(new_n6894_), .A2(new_n6895_), .B(new_n6893_), .ZN(new_n6898_));
  NOR3_X1    g06642(.A1(new_n6891_), .A2(new_n6888_), .A3(new_n6602_), .ZN(new_n6899_));
  NOR3_X1    g06643(.A1(new_n6899_), .A2(new_n6898_), .A3(new_n6712_), .ZN(new_n6900_));
  OAI21_X1   g06644(.A1(new_n6900_), .A2(new_n6897_), .B(new_n6707_), .ZN(new_n6901_));
  XOR2_X1    g06645(.A1(new_n6706_), .A2(new_n2074_), .Z(new_n6902_));
  OAI21_X1   g06646(.A1(new_n6899_), .A2(new_n6898_), .B(new_n6712_), .ZN(new_n6903_));
  NAND3_X1   g06647(.A1(new_n6892_), .A2(new_n6896_), .A3(new_n6713_), .ZN(new_n6904_));
  NAND3_X1   g06648(.A1(new_n6903_), .A2(new_n6904_), .A3(new_n6902_), .ZN(new_n6905_));
  NOR2_X1    g06649(.A1(new_n6606_), .A2(new_n6611_), .ZN(new_n6906_));
  NAND3_X1   g06650(.A1(new_n6901_), .A2(new_n6905_), .A3(new_n6906_), .ZN(new_n6907_));
  AOI21_X1   g06651(.A1(new_n6903_), .A2(new_n6904_), .B(new_n6902_), .ZN(new_n6908_));
  NOR3_X1    g06652(.A1(new_n6900_), .A2(new_n6897_), .A3(new_n6707_), .ZN(new_n6909_));
  INV_X1     g06653(.I(new_n6906_), .ZN(new_n6910_));
  OAI21_X1   g06654(.A1(new_n6909_), .A2(new_n6908_), .B(new_n6910_), .ZN(new_n6911_));
  OAI22_X1   g06655(.A1(new_n1760_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n1755_), .ZN(new_n6912_));
  NAND2_X1   g06656(.A1(new_n2470_), .A2(\b[30] ), .ZN(new_n6913_));
  AOI21_X1   g06657(.A1(new_n6912_), .A2(new_n6913_), .B(new_n1763_), .ZN(new_n6914_));
  NAND2_X1   g06658(.A1(new_n2659_), .A2(new_n6914_), .ZN(new_n6915_));
  XOR2_X1    g06659(.A1(new_n6915_), .A2(\a[26] ), .Z(new_n6916_));
  AOI21_X1   g06660(.A1(new_n6911_), .A2(new_n6907_), .B(new_n6916_), .ZN(new_n6917_));
  NOR3_X1    g06661(.A1(new_n6909_), .A2(new_n6908_), .A3(new_n6910_), .ZN(new_n6918_));
  AOI21_X1   g06662(.A1(new_n6901_), .A2(new_n6905_), .B(new_n6906_), .ZN(new_n6919_));
  INV_X1     g06663(.I(new_n6916_), .ZN(new_n6920_));
  NOR3_X1    g06664(.A1(new_n6918_), .A2(new_n6919_), .A3(new_n6920_), .ZN(new_n6921_));
  INV_X1     g06665(.I(new_n6612_), .ZN(new_n6922_));
  NOR2_X1    g06666(.A1(new_n6617_), .A2(new_n6922_), .ZN(new_n6923_));
  INV_X1     g06667(.I(new_n6923_), .ZN(new_n6924_));
  NOR3_X1    g06668(.A1(new_n6921_), .A2(new_n6917_), .A3(new_n6924_), .ZN(new_n6925_));
  OAI21_X1   g06669(.A1(new_n6918_), .A2(new_n6919_), .B(new_n6920_), .ZN(new_n6926_));
  NAND3_X1   g06670(.A1(new_n6911_), .A2(new_n6907_), .A3(new_n6916_), .ZN(new_n6927_));
  AOI21_X1   g06671(.A1(new_n6926_), .A2(new_n6927_), .B(new_n6923_), .ZN(new_n6928_));
  OAI22_X1   g06672(.A1(new_n1444_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n1439_), .ZN(new_n6929_));
  NAND2_X1   g06673(.A1(new_n2098_), .A2(\b[33] ), .ZN(new_n6930_));
  AOI21_X1   g06674(.A1(new_n6929_), .A2(new_n6930_), .B(new_n1447_), .ZN(new_n6931_));
  NAND2_X1   g06675(.A1(new_n3101_), .A2(new_n6931_), .ZN(new_n6932_));
  XOR2_X1    g06676(.A1(new_n6932_), .A2(\a[23] ), .Z(new_n6933_));
  NOR3_X1    g06677(.A1(new_n6925_), .A2(new_n6928_), .A3(new_n6933_), .ZN(new_n6934_));
  OAI21_X1   g06678(.A1(new_n6925_), .A2(new_n6928_), .B(new_n6933_), .ZN(new_n6935_));
  INV_X1     g06679(.I(new_n6935_), .ZN(new_n6936_));
  NOR2_X1    g06680(.A1(new_n6936_), .A2(new_n6934_), .ZN(new_n6937_));
  NOR2_X1    g06681(.A1(new_n6618_), .A2(new_n6623_), .ZN(new_n6938_));
  XOR2_X1    g06682(.A1(new_n6937_), .A2(new_n6938_), .Z(new_n6939_));
  OAI22_X1   g06683(.A1(new_n1168_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n1163_), .ZN(new_n6940_));
  NAND2_X1   g06684(.A1(new_n1774_), .A2(\b[36] ), .ZN(new_n6941_));
  AOI21_X1   g06685(.A1(new_n6940_), .A2(new_n6941_), .B(new_n1171_), .ZN(new_n6942_));
  NAND2_X1   g06686(.A1(new_n3565_), .A2(new_n6942_), .ZN(new_n6943_));
  XOR2_X1    g06687(.A1(new_n6943_), .A2(\a[20] ), .Z(new_n6944_));
  XNOR2_X1   g06688(.A1(new_n6939_), .A2(new_n6944_), .ZN(new_n6945_));
  OAI21_X1   g06689(.A1(new_n6642_), .A2(new_n6631_), .B(new_n6632_), .ZN(new_n6946_));
  XNOR2_X1   g06690(.A1(new_n6946_), .A2(new_n6945_), .ZN(new_n6947_));
  OAI22_X1   g06691(.A1(new_n940_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n935_), .ZN(new_n6948_));
  NAND2_X1   g06692(.A1(new_n1458_), .A2(\b[39] ), .ZN(new_n6949_));
  AOI21_X1   g06693(.A1(new_n6948_), .A2(new_n6949_), .B(new_n943_), .ZN(new_n6950_));
  NAND2_X1   g06694(.A1(new_n3996_), .A2(new_n6950_), .ZN(new_n6951_));
  XOR2_X1    g06695(.A1(new_n6951_), .A2(\a[17] ), .Z(new_n6952_));
  XNOR2_X1   g06696(.A1(new_n6947_), .A2(new_n6952_), .ZN(new_n6953_));
  XOR2_X1    g06697(.A1(new_n6642_), .A2(new_n6634_), .Z(new_n6954_));
  OAI22_X1   g06698(.A1(new_n6954_), .A2(new_n6643_), .B1(new_n6641_), .B2(new_n6645_), .ZN(new_n6955_));
  XOR2_X1    g06699(.A1(new_n6953_), .A2(new_n6955_), .Z(new_n6956_));
  XOR2_X1    g06700(.A1(new_n6956_), .A2(new_n6702_), .Z(new_n6957_));
  XNOR2_X1   g06701(.A1(new_n6957_), .A2(new_n6700_), .ZN(new_n6958_));
  XNOR2_X1   g06702(.A1(new_n6958_), .A2(new_n6695_), .ZN(new_n6959_));
  XOR2_X1    g06703(.A1(new_n6959_), .A2(new_n6690_), .Z(new_n6960_));
  OAI22_X1   g06704(.A1(new_n437_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n431_), .ZN(new_n6961_));
  NAND2_X1   g06705(.A1(new_n775_), .A2(\b[48] ), .ZN(new_n6962_));
  AOI21_X1   g06706(.A1(new_n6961_), .A2(new_n6962_), .B(new_n440_), .ZN(new_n6963_));
  NAND2_X1   g06707(.A1(new_n5537_), .A2(new_n6963_), .ZN(new_n6964_));
  XOR2_X1    g06708(.A1(new_n6964_), .A2(\a[8] ), .Z(new_n6965_));
  INV_X1     g06709(.I(new_n6965_), .ZN(new_n6966_));
  XOR2_X1    g06710(.A1(new_n6960_), .A2(new_n6966_), .Z(new_n6967_));
  INV_X1     g06711(.I(new_n6663_), .ZN(new_n6968_));
  XOR2_X1    g06712(.A1(new_n6480_), .A2(new_n6968_), .Z(new_n6969_));
  NAND2_X1   g06713(.A1(new_n6969_), .A2(new_n6658_), .ZN(new_n6970_));
  XNOR2_X1   g06714(.A1(new_n6970_), .A2(new_n6967_), .ZN(new_n6971_));
  NOR2_X1    g06715(.A1(new_n6481_), .A2(new_n6663_), .ZN(new_n6972_));
  XNOR2_X1   g06716(.A1(new_n6971_), .A2(new_n6972_), .ZN(new_n6973_));
  OAI22_X1   g06717(.A1(new_n364_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n320_), .ZN(new_n6974_));
  NAND2_X1   g06718(.A1(new_n594_), .A2(\b[51] ), .ZN(new_n6975_));
  AOI21_X1   g06719(.A1(new_n6974_), .A2(new_n6975_), .B(new_n312_), .ZN(new_n6976_));
  NAND2_X1   g06720(.A1(new_n6219_), .A2(new_n6976_), .ZN(new_n6977_));
  XOR2_X1    g06721(.A1(new_n6977_), .A2(\a[5] ), .Z(new_n6978_));
  INV_X1     g06722(.I(new_n6978_), .ZN(new_n6979_));
  XNOR2_X1   g06723(.A1(new_n6480_), .A2(new_n6664_), .ZN(new_n6980_));
  NOR2_X1    g06724(.A1(new_n6980_), .A2(new_n6670_), .ZN(new_n6981_));
  NOR3_X1    g06725(.A1(new_n6452_), .A2(new_n6676_), .A3(new_n6981_), .ZN(new_n6982_));
  XOR2_X1    g06726(.A1(new_n6982_), .A2(new_n6979_), .Z(new_n6983_));
  XOR2_X1    g06727(.A1(new_n6973_), .A2(new_n6983_), .Z(new_n6984_));
  OAI21_X1   g06728(.A1(new_n6215_), .A2(new_n6467_), .B(new_n6238_), .ZN(new_n6985_));
  NAND3_X1   g06729(.A1(new_n6230_), .A2(new_n6231_), .A3(new_n6985_), .ZN(new_n6986_));
  OAI21_X1   g06730(.A1(\b[53] ), .A2(\b[55] ), .B(\b[54] ), .ZN(new_n6987_));
  NAND2_X1   g06731(.A1(new_n6986_), .A2(new_n6987_), .ZN(new_n6988_));
  XNOR2_X1   g06732(.A1(\b[55] ), .A2(\b[56] ), .ZN(new_n6989_));
  INV_X1     g06733(.I(new_n6989_), .ZN(new_n6990_));
  XOR2_X1    g06734(.A1(\b[55] ), .A2(\b[56] ), .Z(new_n6991_));
  NOR2_X1    g06735(.A1(new_n6988_), .A2(new_n6991_), .ZN(new_n6992_));
  AOI21_X1   g06736(.A1(new_n6988_), .A2(new_n6990_), .B(new_n6992_), .ZN(new_n6993_));
  INV_X1     g06737(.I(new_n6993_), .ZN(new_n6994_));
  INV_X1     g06738(.I(\b[56] ), .ZN(new_n6995_));
  OAI22_X1   g06739(.A1(new_n405_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n404_), .ZN(new_n6996_));
  NAND2_X1   g06740(.A1(new_n279_), .A2(\b[54] ), .ZN(new_n6997_));
  AOI21_X1   g06741(.A1(new_n6996_), .A2(new_n6997_), .B(new_n264_), .ZN(new_n6998_));
  NAND2_X1   g06742(.A1(new_n6994_), .A2(new_n6998_), .ZN(new_n6999_));
  XOR2_X1    g06743(.A1(new_n6999_), .A2(\a[2] ), .Z(new_n7000_));
  XOR2_X1    g06744(.A1(new_n6984_), .A2(new_n7000_), .Z(new_n7001_));
  INV_X1     g06745(.I(new_n6984_), .ZN(new_n7002_));
  NOR2_X1    g06746(.A1(new_n7002_), .A2(new_n7000_), .ZN(new_n7003_));
  INV_X1     g06747(.I(new_n7000_), .ZN(new_n7004_));
  NOR2_X1    g06748(.A1(new_n6984_), .A2(new_n7004_), .ZN(new_n7005_));
  OAI21_X1   g06749(.A1(new_n7003_), .A2(new_n7005_), .B(new_n6689_), .ZN(new_n7006_));
  OAI21_X1   g06750(.A1(new_n6689_), .A2(new_n7001_), .B(new_n7006_), .ZN(\f[56] ));
  INV_X1     g06751(.I(new_n6982_), .ZN(new_n7008_));
  XOR2_X1    g06752(.A1(new_n6973_), .A2(new_n6978_), .Z(new_n7009_));
  AOI21_X1   g06753(.A1(new_n6979_), .A2(new_n7008_), .B(new_n7009_), .ZN(new_n7010_));
  OAI21_X1   g06754(.A1(new_n6870_), .A2(new_n6867_), .B(new_n6881_), .ZN(new_n7011_));
  AOI21_X1   g06755(.A1(new_n6758_), .A2(new_n6755_), .B(new_n6768_), .ZN(new_n7012_));
  NAND2_X1   g06756(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n7013_));
  OR2_X2     g06757(.A1(\a[56] ), .A2(\a[57] ), .Z(new_n7014_));
  NAND2_X1   g06758(.A1(new_n7014_), .A2(new_n7013_), .ZN(new_n7015_));
  NOR2_X1    g06759(.A1(new_n7015_), .A2(new_n258_), .ZN(new_n7016_));
  INV_X1     g06760(.I(new_n7016_), .ZN(new_n7017_));
  NOR3_X1    g06761(.A1(new_n6738_), .A2(new_n6720_), .A3(new_n6734_), .ZN(new_n7018_));
  NOR2_X1    g06762(.A1(new_n6721_), .A2(new_n292_), .ZN(new_n7019_));
  NOR2_X1    g06763(.A1(new_n6723_), .A2(new_n290_), .ZN(new_n7020_));
  OAI22_X1   g06764(.A1(new_n7019_), .A2(new_n7020_), .B1(new_n6729_), .B2(new_n267_), .ZN(new_n7021_));
  NOR2_X1    g06765(.A1(new_n677_), .A2(new_n6731_), .ZN(new_n7022_));
  AND3_X2    g06766(.A1(new_n7021_), .A2(new_n6516_), .A3(new_n7022_), .Z(new_n7023_));
  AOI21_X1   g06767(.A1(new_n7021_), .A2(new_n7022_), .B(new_n6516_), .ZN(new_n7024_));
  NOR2_X1    g06768(.A1(new_n7023_), .A2(new_n7024_), .ZN(new_n7025_));
  NOR2_X1    g06769(.A1(new_n7018_), .A2(new_n7025_), .ZN(new_n7026_));
  NAND2_X1   g06770(.A1(new_n7018_), .A2(new_n7025_), .ZN(new_n7027_));
  INV_X1     g06771(.I(new_n7027_), .ZN(new_n7028_));
  OAI21_X1   g06772(.A1(new_n7028_), .A2(new_n7026_), .B(new_n7017_), .ZN(new_n7029_));
  NAND3_X1   g06773(.A1(new_n6735_), .A2(new_n6737_), .A3(new_n6733_), .ZN(new_n7030_));
  INV_X1     g06774(.I(new_n7025_), .ZN(new_n7031_));
  NAND2_X1   g06775(.A1(new_n7031_), .A2(new_n7030_), .ZN(new_n7032_));
  NAND3_X1   g06776(.A1(new_n7032_), .A2(new_n7027_), .A3(new_n7016_), .ZN(new_n7033_));
  OAI22_X1   g06777(.A1(new_n5786_), .A2(new_n403_), .B1(new_n347_), .B2(new_n5792_), .ZN(new_n7034_));
  OAI21_X1   g06778(.A1(new_n393_), .A2(new_n6012_), .B(new_n7034_), .ZN(new_n7035_));
  NAND3_X1   g06779(.A1(new_n402_), .A2(new_n5795_), .A3(new_n7035_), .ZN(new_n7036_));
  XOR2_X1    g06780(.A1(new_n7036_), .A2(new_n5783_), .Z(new_n7037_));
  NAND3_X1   g06781(.A1(new_n7029_), .A2(new_n7033_), .A3(new_n7037_), .ZN(new_n7038_));
  AOI21_X1   g06782(.A1(new_n7032_), .A2(new_n7027_), .B(new_n7016_), .ZN(new_n7039_));
  NOR3_X1    g06783(.A1(new_n7028_), .A2(new_n7017_), .A3(new_n7026_), .ZN(new_n7040_));
  XOR2_X1    g06784(.A1(new_n7036_), .A2(\a[53] ), .Z(new_n7041_));
  OAI21_X1   g06785(.A1(new_n7040_), .A2(new_n7039_), .B(new_n7041_), .ZN(new_n7042_));
  AOI21_X1   g06786(.A1(new_n7038_), .A2(new_n7042_), .B(new_n7012_), .ZN(new_n7043_));
  OAI21_X1   g06787(.A1(new_n6719_), .A2(new_n6769_), .B(new_n6750_), .ZN(new_n7044_));
  AOI21_X1   g06788(.A1(new_n7029_), .A2(new_n7033_), .B(new_n7041_), .ZN(new_n7045_));
  INV_X1     g06789(.I(new_n7045_), .ZN(new_n7046_));
  NAND3_X1   g06790(.A1(new_n7029_), .A2(new_n7033_), .A3(new_n7041_), .ZN(new_n7047_));
  AOI21_X1   g06791(.A1(new_n7046_), .A2(new_n7047_), .B(new_n7044_), .ZN(new_n7048_));
  NOR2_X1    g06792(.A1(new_n7048_), .A2(new_n7043_), .ZN(new_n7049_));
  INV_X1     g06793(.I(new_n7049_), .ZN(new_n7050_));
  OAI22_X1   g06794(.A1(new_n5228_), .A2(new_n510_), .B1(new_n495_), .B2(new_n5225_), .ZN(new_n7051_));
  NAND2_X1   g06795(.A1(new_n5387_), .A2(\b[7] ), .ZN(new_n7052_));
  AOI21_X1   g06796(.A1(new_n7051_), .A2(new_n7052_), .B(new_n5231_), .ZN(new_n7053_));
  NAND3_X1   g06797(.A1(new_n518_), .A2(new_n5220_), .A3(new_n7053_), .ZN(new_n7054_));
  NOR2_X1    g06798(.A1(new_n516_), .A2(\b[9] ), .ZN(new_n7055_));
  AOI21_X1   g06799(.A1(new_n512_), .A2(new_n511_), .B(new_n510_), .ZN(new_n7056_));
  OAI21_X1   g06800(.A1(new_n7055_), .A2(new_n7056_), .B(new_n7053_), .ZN(new_n7057_));
  NAND2_X1   g06801(.A1(new_n7057_), .A2(\a[50] ), .ZN(new_n7058_));
  NAND2_X1   g06802(.A1(new_n7058_), .A2(new_n7054_), .ZN(new_n7059_));
  NAND2_X1   g06803(.A1(new_n6787_), .A2(new_n6775_), .ZN(new_n7060_));
  NAND2_X1   g06804(.A1(new_n6790_), .A2(new_n7060_), .ZN(new_n7061_));
  NOR3_X1    g06805(.A1(new_n6756_), .A2(new_n6761_), .A3(new_n6773_), .ZN(new_n7062_));
  INV_X1     g06806(.I(new_n7062_), .ZN(new_n7063_));
  AOI21_X1   g06807(.A1(new_n7061_), .A2(new_n7063_), .B(new_n7059_), .ZN(new_n7064_));
  NAND3_X1   g06808(.A1(new_n7061_), .A2(new_n7059_), .A3(new_n7063_), .ZN(new_n7065_));
  INV_X1     g06809(.I(new_n7065_), .ZN(new_n7066_));
  NOR2_X1    g06810(.A1(new_n7066_), .A2(new_n7064_), .ZN(new_n7067_));
  NOR2_X1    g06811(.A1(new_n7067_), .A2(new_n7050_), .ZN(new_n7068_));
  NOR3_X1    g06812(.A1(new_n7066_), .A2(new_n7049_), .A3(new_n7064_), .ZN(new_n7069_));
  NOR2_X1    g06813(.A1(new_n7068_), .A2(new_n7069_), .ZN(new_n7070_));
  INV_X1     g06814(.I(new_n7070_), .ZN(new_n7071_));
  OAI22_X1   g06815(.A1(new_n4711_), .A2(new_n717_), .B1(new_n659_), .B2(new_n4706_), .ZN(new_n7072_));
  NAND2_X1   g06816(.A1(new_n5814_), .A2(\b[10] ), .ZN(new_n7073_));
  AOI21_X1   g06817(.A1(new_n7072_), .A2(new_n7073_), .B(new_n4714_), .ZN(new_n7074_));
  NAND2_X1   g06818(.A1(new_n716_), .A2(new_n7074_), .ZN(new_n7075_));
  XOR2_X1    g06819(.A1(new_n7075_), .A2(\a[47] ), .Z(new_n7076_));
  NOR3_X1    g06820(.A1(new_n6803_), .A2(new_n6799_), .A3(new_n6818_), .ZN(new_n7077_));
  OAI21_X1   g06821(.A1(new_n6800_), .A2(new_n6801_), .B(new_n6798_), .ZN(new_n7078_));
  OAI21_X1   g06822(.A1(new_n7077_), .A2(new_n6809_), .B(new_n7078_), .ZN(new_n7079_));
  NAND2_X1   g06823(.A1(new_n7079_), .A2(new_n7076_), .ZN(new_n7080_));
  INV_X1     g06824(.I(new_n7076_), .ZN(new_n7081_));
  NAND3_X1   g06825(.A1(new_n6811_), .A2(new_n6812_), .A3(new_n6817_), .ZN(new_n7082_));
  NAND2_X1   g06826(.A1(new_n7082_), .A2(new_n6815_), .ZN(new_n7083_));
  NAND3_X1   g06827(.A1(new_n7083_), .A2(new_n7081_), .A3(new_n7078_), .ZN(new_n7084_));
  AOI21_X1   g06828(.A1(new_n7080_), .A2(new_n7084_), .B(new_n7071_), .ZN(new_n7085_));
  AOI21_X1   g06829(.A1(new_n7083_), .A2(new_n7078_), .B(new_n7081_), .ZN(new_n7086_));
  NOR2_X1    g06830(.A1(new_n7079_), .A2(new_n7076_), .ZN(new_n7087_));
  NOR3_X1    g06831(.A1(new_n7087_), .A2(new_n7086_), .A3(new_n7070_), .ZN(new_n7088_));
  NOR2_X1    g06832(.A1(new_n7088_), .A2(new_n7085_), .ZN(new_n7089_));
  OAI22_X1   g06833(.A1(new_n4208_), .A2(new_n904_), .B1(new_n848_), .B2(new_n4203_), .ZN(new_n7090_));
  NAND2_X1   g06834(.A1(new_n5244_), .A2(\b[13] ), .ZN(new_n7091_));
  AOI21_X1   g06835(.A1(new_n7090_), .A2(new_n7091_), .B(new_n4211_), .ZN(new_n7092_));
  NAND2_X1   g06836(.A1(new_n907_), .A2(new_n7092_), .ZN(new_n7093_));
  XOR2_X1    g06837(.A1(new_n7093_), .A2(\a[44] ), .Z(new_n7094_));
  INV_X1     g06838(.I(new_n7094_), .ZN(new_n7095_));
  OAI21_X1   g06839(.A1(new_n6558_), .A2(new_n6555_), .B(new_n6563_), .ZN(new_n7096_));
  INV_X1     g06840(.I(new_n7096_), .ZN(new_n7097_));
  NOR3_X1    g06841(.A1(new_n6828_), .A2(new_n6832_), .A3(new_n7097_), .ZN(new_n7098_));
  NOR2_X1    g06842(.A1(new_n7098_), .A2(new_n7095_), .ZN(new_n7099_));
  NOR4_X1    g06843(.A1(new_n6828_), .A2(new_n6832_), .A3(new_n7097_), .A4(new_n7094_), .ZN(new_n7100_));
  OAI21_X1   g06844(.A1(new_n7099_), .A2(new_n7100_), .B(new_n7089_), .ZN(new_n7101_));
  OAI21_X1   g06845(.A1(new_n7087_), .A2(new_n7086_), .B(new_n7070_), .ZN(new_n7102_));
  NAND3_X1   g06846(.A1(new_n7080_), .A2(new_n7084_), .A3(new_n7071_), .ZN(new_n7103_));
  NAND2_X1   g06847(.A1(new_n7102_), .A2(new_n7103_), .ZN(new_n7104_));
  NAND3_X1   g06848(.A1(new_n6837_), .A2(new_n6836_), .A3(new_n7096_), .ZN(new_n7105_));
  NAND2_X1   g06849(.A1(new_n7105_), .A2(new_n7094_), .ZN(new_n7106_));
  NAND4_X1   g06850(.A1(new_n6837_), .A2(new_n6836_), .A3(new_n7095_), .A4(new_n7096_), .ZN(new_n7107_));
  NAND3_X1   g06851(.A1(new_n7106_), .A2(new_n7104_), .A3(new_n7107_), .ZN(new_n7108_));
  OAI22_X1   g06852(.A1(new_n3736_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n3731_), .ZN(new_n7109_));
  NAND2_X1   g06853(.A1(new_n4730_), .A2(\b[16] ), .ZN(new_n7110_));
  AOI21_X1   g06854(.A1(new_n7109_), .A2(new_n7110_), .B(new_n3739_), .ZN(new_n7111_));
  NAND2_X1   g06855(.A1(new_n1123_), .A2(new_n7111_), .ZN(new_n7112_));
  XOR2_X1    g06856(.A1(new_n7112_), .A2(\a[41] ), .Z(new_n7113_));
  INV_X1     g06857(.I(new_n7113_), .ZN(new_n7114_));
  NAND3_X1   g06858(.A1(new_n7101_), .A2(new_n7108_), .A3(new_n7114_), .ZN(new_n7115_));
  AOI21_X1   g06859(.A1(new_n7106_), .A2(new_n7107_), .B(new_n7104_), .ZN(new_n7116_));
  NOR3_X1    g06860(.A1(new_n7099_), .A2(new_n7089_), .A3(new_n7100_), .ZN(new_n7117_));
  OAI21_X1   g06861(.A1(new_n7117_), .A2(new_n7116_), .B(new_n7113_), .ZN(new_n7118_));
  OAI21_X1   g06862(.A1(new_n6850_), .A2(new_n6848_), .B(new_n6860_), .ZN(new_n7119_));
  NAND3_X1   g06863(.A1(new_n7118_), .A2(new_n7115_), .A3(new_n7119_), .ZN(new_n7120_));
  NOR3_X1    g06864(.A1(new_n7117_), .A2(new_n7116_), .A3(new_n7113_), .ZN(new_n7121_));
  AOI21_X1   g06865(.A1(new_n7101_), .A2(new_n7108_), .B(new_n7114_), .ZN(new_n7122_));
  AOI21_X1   g06866(.A1(new_n6716_), .A2(new_n6861_), .B(new_n6844_), .ZN(new_n7123_));
  OAI21_X1   g06867(.A1(new_n7121_), .A2(new_n7122_), .B(new_n7123_), .ZN(new_n7124_));
  OAI22_X1   g06868(.A1(new_n3298_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n3293_), .ZN(new_n7125_));
  NAND2_X1   g06869(.A1(new_n4227_), .A2(\b[19] ), .ZN(new_n7126_));
  AOI21_X1   g06870(.A1(new_n7125_), .A2(new_n7126_), .B(new_n3301_), .ZN(new_n7127_));
  NAND2_X1   g06871(.A1(new_n1396_), .A2(new_n7127_), .ZN(new_n7128_));
  XOR2_X1    g06872(.A1(new_n7128_), .A2(\a[38] ), .Z(new_n7129_));
  AOI21_X1   g06873(.A1(new_n7124_), .A2(new_n7120_), .B(new_n7129_), .ZN(new_n7130_));
  INV_X1     g06874(.I(new_n7130_), .ZN(new_n7131_));
  NAND3_X1   g06875(.A1(new_n7124_), .A2(new_n7120_), .A3(new_n7129_), .ZN(new_n7132_));
  NAND2_X1   g06876(.A1(new_n7131_), .A2(new_n7132_), .ZN(new_n7133_));
  INV_X1     g06877(.I(new_n7129_), .ZN(new_n7134_));
  NAND3_X1   g06878(.A1(new_n7124_), .A2(new_n7120_), .A3(new_n7134_), .ZN(new_n7135_));
  NOR3_X1    g06879(.A1(new_n7121_), .A2(new_n7122_), .A3(new_n7123_), .ZN(new_n7136_));
  AOI21_X1   g06880(.A1(new_n7118_), .A2(new_n7115_), .B(new_n7119_), .ZN(new_n7137_));
  OAI21_X1   g06881(.A1(new_n7136_), .A2(new_n7137_), .B(new_n7129_), .ZN(new_n7138_));
  AOI21_X1   g06882(.A1(new_n7138_), .A2(new_n7135_), .B(new_n7011_), .ZN(new_n7139_));
  AOI21_X1   g06883(.A1(new_n7133_), .A2(new_n7011_), .B(new_n7139_), .ZN(new_n7140_));
  OAI22_X1   g06884(.A1(new_n2846_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n2841_), .ZN(new_n7141_));
  NAND2_X1   g06885(.A1(new_n3755_), .A2(\b[22] ), .ZN(new_n7142_));
  AOI21_X1   g06886(.A1(new_n7141_), .A2(new_n7142_), .B(new_n2849_), .ZN(new_n7143_));
  NAND2_X1   g06887(.A1(new_n1708_), .A2(new_n7143_), .ZN(new_n7144_));
  XOR2_X1    g06888(.A1(new_n7144_), .A2(\a[35] ), .Z(new_n7145_));
  INV_X1     g06889(.I(new_n7145_), .ZN(new_n7146_));
  OAI21_X1   g06890(.A1(new_n6889_), .A2(new_n6890_), .B(new_n6604_), .ZN(new_n7147_));
  NOR3_X1    g06891(.A1(new_n6883_), .A2(new_n6886_), .A3(new_n6879_), .ZN(new_n7148_));
  INV_X1     g06892(.I(new_n7148_), .ZN(new_n7149_));
  AOI21_X1   g06893(.A1(new_n7147_), .A2(new_n7149_), .B(new_n7146_), .ZN(new_n7150_));
  AOI21_X1   g06894(.A1(new_n6887_), .A2(new_n6880_), .B(new_n6599_), .ZN(new_n7151_));
  NOR3_X1    g06895(.A1(new_n7151_), .A2(new_n7145_), .A3(new_n7148_), .ZN(new_n7152_));
  OAI21_X1   g06896(.A1(new_n7150_), .A2(new_n7152_), .B(new_n7140_), .ZN(new_n7153_));
  INV_X1     g06897(.I(new_n7132_), .ZN(new_n7154_));
  OAI21_X1   g06898(.A1(new_n7154_), .A2(new_n7130_), .B(new_n7011_), .ZN(new_n7155_));
  AOI21_X1   g06899(.A1(new_n6715_), .A2(new_n6882_), .B(new_n6859_), .ZN(new_n7156_));
  NOR3_X1    g06900(.A1(new_n7136_), .A2(new_n7137_), .A3(new_n7129_), .ZN(new_n7157_));
  AOI21_X1   g06901(.A1(new_n7124_), .A2(new_n7120_), .B(new_n7134_), .ZN(new_n7158_));
  OAI21_X1   g06902(.A1(new_n7157_), .A2(new_n7158_), .B(new_n7156_), .ZN(new_n7159_));
  NAND2_X1   g06903(.A1(new_n7155_), .A2(new_n7159_), .ZN(new_n7160_));
  OAI21_X1   g06904(.A1(new_n7151_), .A2(new_n7148_), .B(new_n7145_), .ZN(new_n7161_));
  NAND3_X1   g06905(.A1(new_n7147_), .A2(new_n7146_), .A3(new_n7149_), .ZN(new_n7162_));
  NAND3_X1   g06906(.A1(new_n7161_), .A2(new_n7162_), .A3(new_n7160_), .ZN(new_n7163_));
  NAND2_X1   g06907(.A1(new_n7153_), .A2(new_n7163_), .ZN(new_n7164_));
  OAI22_X1   g06908(.A1(new_n2452_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n2447_), .ZN(new_n7165_));
  NAND2_X1   g06909(.A1(new_n3312_), .A2(\b[25] ), .ZN(new_n7166_));
  AOI21_X1   g06910(.A1(new_n7165_), .A2(new_n7166_), .B(new_n2455_), .ZN(new_n7167_));
  NAND2_X1   g06911(.A1(new_n2042_), .A2(new_n7167_), .ZN(new_n7168_));
  XOR2_X1    g06912(.A1(new_n7168_), .A2(\a[32] ), .Z(new_n7169_));
  AOI21_X1   g06913(.A1(new_n6894_), .A2(new_n6895_), .B(new_n6713_), .ZN(new_n7170_));
  OAI21_X1   g06914(.A1(new_n6891_), .A2(new_n6888_), .B(new_n6713_), .ZN(new_n7171_));
  NAND3_X1   g06915(.A1(new_n6894_), .A2(new_n6895_), .A3(new_n6712_), .ZN(new_n7172_));
  AOI21_X1   g06916(.A1(new_n7171_), .A2(new_n7172_), .B(new_n6893_), .ZN(new_n7173_));
  OAI21_X1   g06917(.A1(new_n7173_), .A2(new_n7170_), .B(new_n7169_), .ZN(new_n7174_));
  INV_X1     g06918(.I(new_n7169_), .ZN(new_n7175_));
  INV_X1     g06919(.I(new_n7170_), .ZN(new_n7176_));
  AOI21_X1   g06920(.A1(new_n6894_), .A2(new_n6895_), .B(new_n6712_), .ZN(new_n7177_));
  NOR3_X1    g06921(.A1(new_n6891_), .A2(new_n6888_), .A3(new_n6713_), .ZN(new_n7178_));
  OAI21_X1   g06922(.A1(new_n7178_), .A2(new_n7177_), .B(new_n6602_), .ZN(new_n7179_));
  NAND3_X1   g06923(.A1(new_n7179_), .A2(new_n7175_), .A3(new_n7176_), .ZN(new_n7180_));
  AOI21_X1   g06924(.A1(new_n7180_), .A2(new_n7174_), .B(new_n7164_), .ZN(new_n7181_));
  AOI21_X1   g06925(.A1(new_n7161_), .A2(new_n7162_), .B(new_n7160_), .ZN(new_n7182_));
  NOR3_X1    g06926(.A1(new_n7150_), .A2(new_n7152_), .A3(new_n7140_), .ZN(new_n7183_));
  NOR2_X1    g06927(.A1(new_n7182_), .A2(new_n7183_), .ZN(new_n7184_));
  AOI21_X1   g06928(.A1(new_n7179_), .A2(new_n7176_), .B(new_n7175_), .ZN(new_n7185_));
  NOR3_X1    g06929(.A1(new_n7173_), .A2(new_n7169_), .A3(new_n7170_), .ZN(new_n7186_));
  NOR3_X1    g06930(.A1(new_n7185_), .A2(new_n7186_), .A3(new_n7184_), .ZN(new_n7187_));
  NOR2_X1    g06931(.A1(new_n7187_), .A2(new_n7181_), .ZN(new_n7188_));
  OAI22_X1   g06932(.A1(new_n2084_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n2079_), .ZN(new_n7189_));
  NAND2_X1   g06933(.A1(new_n2864_), .A2(\b[28] ), .ZN(new_n7190_));
  AOI21_X1   g06934(.A1(new_n7189_), .A2(new_n7190_), .B(new_n2087_), .ZN(new_n7191_));
  NAND2_X1   g06935(.A1(new_n2404_), .A2(new_n7191_), .ZN(new_n7192_));
  XOR2_X1    g06936(.A1(new_n7192_), .A2(\a[29] ), .Z(new_n7193_));
  INV_X1     g06937(.I(new_n7193_), .ZN(new_n7194_));
  NOR3_X1    g06938(.A1(new_n6891_), .A2(new_n6888_), .A3(new_n6712_), .ZN(new_n7195_));
  OAI21_X1   g06939(.A1(new_n7195_), .A2(new_n7170_), .B(new_n6602_), .ZN(new_n7196_));
  INV_X1     g06940(.I(new_n7196_), .ZN(new_n7197_));
  NOR3_X1    g06941(.A1(new_n7195_), .A2(new_n7170_), .A3(new_n6602_), .ZN(new_n7198_));
  OAI21_X1   g06942(.A1(new_n7197_), .A2(new_n7198_), .B(new_n6707_), .ZN(new_n7199_));
  AOI21_X1   g06943(.A1(new_n6907_), .A2(new_n7199_), .B(new_n7194_), .ZN(new_n7200_));
  INV_X1     g06944(.I(new_n7198_), .ZN(new_n7201_));
  AOI21_X1   g06945(.A1(new_n7201_), .A2(new_n7196_), .B(new_n6902_), .ZN(new_n7202_));
  NOR3_X1    g06946(.A1(new_n6918_), .A2(new_n7193_), .A3(new_n7202_), .ZN(new_n7203_));
  OAI21_X1   g06947(.A1(new_n7203_), .A2(new_n7200_), .B(new_n7188_), .ZN(new_n7204_));
  OAI21_X1   g06948(.A1(new_n7185_), .A2(new_n7186_), .B(new_n7184_), .ZN(new_n7205_));
  NAND3_X1   g06949(.A1(new_n7180_), .A2(new_n7174_), .A3(new_n7164_), .ZN(new_n7206_));
  NAND2_X1   g06950(.A1(new_n7205_), .A2(new_n7206_), .ZN(new_n7207_));
  OAI21_X1   g06951(.A1(new_n6918_), .A2(new_n7202_), .B(new_n7193_), .ZN(new_n7208_));
  NAND3_X1   g06952(.A1(new_n6907_), .A2(new_n7194_), .A3(new_n7199_), .ZN(new_n7209_));
  NAND3_X1   g06953(.A1(new_n7208_), .A2(new_n7207_), .A3(new_n7209_), .ZN(new_n7210_));
  NAND2_X1   g06954(.A1(new_n7204_), .A2(new_n7210_), .ZN(new_n7211_));
  OAI22_X1   g06955(.A1(new_n1760_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n1755_), .ZN(new_n7212_));
  NAND2_X1   g06956(.A1(new_n2470_), .A2(\b[31] ), .ZN(new_n7213_));
  AOI21_X1   g06957(.A1(new_n7212_), .A2(new_n7213_), .B(new_n1763_), .ZN(new_n7214_));
  NAND3_X1   g06958(.A1(new_n2797_), .A2(new_n1750_), .A3(new_n7214_), .ZN(new_n7215_));
  INV_X1     g06959(.I(new_n7215_), .ZN(new_n7216_));
  AOI21_X1   g06960(.A1(new_n2797_), .A2(new_n7214_), .B(new_n1750_), .ZN(new_n7217_));
  NOR2_X1    g06961(.A1(new_n7216_), .A2(new_n7217_), .ZN(new_n7218_));
  AOI21_X1   g06962(.A1(new_n6911_), .A2(new_n6907_), .B(new_n6920_), .ZN(new_n7219_));
  OAI21_X1   g06963(.A1(new_n6925_), .A2(new_n7219_), .B(new_n7218_), .ZN(new_n7220_));
  NAND3_X1   g06964(.A1(new_n6926_), .A2(new_n6927_), .A3(new_n6923_), .ZN(new_n7221_));
  INV_X1     g06965(.I(new_n7218_), .ZN(new_n7222_));
  INV_X1     g06966(.I(new_n7219_), .ZN(new_n7223_));
  NAND3_X1   g06967(.A1(new_n7221_), .A2(new_n7222_), .A3(new_n7223_), .ZN(new_n7224_));
  AOI21_X1   g06968(.A1(new_n7220_), .A2(new_n7224_), .B(new_n7211_), .ZN(new_n7225_));
  AOI21_X1   g06969(.A1(new_n7208_), .A2(new_n7209_), .B(new_n7207_), .ZN(new_n7226_));
  NOR3_X1    g06970(.A1(new_n7203_), .A2(new_n7188_), .A3(new_n7200_), .ZN(new_n7227_));
  NOR2_X1    g06971(.A1(new_n7227_), .A2(new_n7226_), .ZN(new_n7228_));
  AOI21_X1   g06972(.A1(new_n7221_), .A2(new_n7223_), .B(new_n7222_), .ZN(new_n7229_));
  NOR3_X1    g06973(.A1(new_n6925_), .A2(new_n7218_), .A3(new_n7219_), .ZN(new_n7230_));
  NOR3_X1    g06974(.A1(new_n7228_), .A2(new_n7230_), .A3(new_n7229_), .ZN(new_n7231_));
  NOR2_X1    g06975(.A1(new_n7231_), .A2(new_n7225_), .ZN(new_n7232_));
  OAI22_X1   g06976(.A1(new_n1444_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n1439_), .ZN(new_n7233_));
  NAND2_X1   g06977(.A1(new_n2098_), .A2(\b[34] ), .ZN(new_n7234_));
  AOI21_X1   g06978(.A1(new_n7233_), .A2(new_n7234_), .B(new_n1447_), .ZN(new_n7235_));
  NAND2_X1   g06979(.A1(new_n3246_), .A2(new_n7235_), .ZN(new_n7236_));
  XOR2_X1    g06980(.A1(new_n7236_), .A2(\a[23] ), .Z(new_n7237_));
  INV_X1     g06981(.I(new_n6934_), .ZN(new_n7238_));
  INV_X1     g06982(.I(new_n6938_), .ZN(new_n7239_));
  NAND3_X1   g06983(.A1(new_n7238_), .A2(new_n6935_), .A3(new_n7239_), .ZN(new_n7240_));
  XOR2_X1    g06984(.A1(new_n7240_), .A2(new_n7237_), .Z(new_n7241_));
  XOR2_X1    g06985(.A1(new_n7241_), .A2(new_n7232_), .Z(new_n7242_));
  OAI22_X1   g06986(.A1(new_n1168_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n1163_), .ZN(new_n7243_));
  NAND2_X1   g06987(.A1(new_n1774_), .A2(\b[37] ), .ZN(new_n7244_));
  AOI21_X1   g06988(.A1(new_n7243_), .A2(new_n7244_), .B(new_n1171_), .ZN(new_n7245_));
  NAND2_X1   g06989(.A1(new_n3700_), .A2(new_n7245_), .ZN(new_n7246_));
  XOR2_X1    g06990(.A1(new_n7246_), .A2(\a[20] ), .Z(new_n7247_));
  INV_X1     g06991(.I(new_n6939_), .ZN(new_n7248_));
  NAND2_X1   g06992(.A1(new_n7248_), .A2(new_n6944_), .ZN(new_n7249_));
  NAND3_X1   g06993(.A1(new_n6946_), .A2(new_n7249_), .A3(new_n6945_), .ZN(new_n7250_));
  XOR2_X1    g06994(.A1(new_n7250_), .A2(new_n7247_), .Z(new_n7251_));
  XOR2_X1    g06995(.A1(new_n7251_), .A2(new_n7242_), .Z(new_n7252_));
  OAI22_X1   g06996(.A1(new_n940_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n935_), .ZN(new_n7253_));
  NAND2_X1   g06997(.A1(new_n1458_), .A2(\b[40] ), .ZN(new_n7254_));
  AOI21_X1   g06998(.A1(new_n7253_), .A2(new_n7254_), .B(new_n943_), .ZN(new_n7255_));
  NAND2_X1   g06999(.A1(new_n4017_), .A2(new_n7255_), .ZN(new_n7256_));
  XOR2_X1    g07000(.A1(new_n7256_), .A2(\a[17] ), .Z(new_n7257_));
  INV_X1     g07001(.I(new_n6947_), .ZN(new_n7258_));
  NAND2_X1   g07002(.A1(new_n7258_), .A2(new_n6952_), .ZN(new_n7259_));
  NAND3_X1   g07003(.A1(new_n6953_), .A2(new_n7259_), .A3(new_n6955_), .ZN(new_n7260_));
  XOR2_X1    g07004(.A1(new_n7260_), .A2(new_n7257_), .Z(new_n7261_));
  XOR2_X1    g07005(.A1(new_n7261_), .A2(new_n7252_), .Z(new_n7262_));
  OAI22_X1   g07006(.A1(new_n757_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n752_), .ZN(new_n7263_));
  NAND2_X1   g07007(.A1(new_n1182_), .A2(\b[43] ), .ZN(new_n7264_));
  AOI21_X1   g07008(.A1(new_n7263_), .A2(new_n7264_), .B(new_n760_), .ZN(new_n7265_));
  NAND2_X1   g07009(.A1(new_n4513_), .A2(new_n7265_), .ZN(new_n7266_));
  XOR2_X1    g07010(.A1(new_n7266_), .A2(\a[14] ), .Z(new_n7267_));
  XOR2_X1    g07011(.A1(new_n6956_), .A2(new_n6700_), .Z(new_n7268_));
  NAND2_X1   g07012(.A1(new_n7268_), .A2(new_n6702_), .ZN(new_n7269_));
  NAND2_X1   g07013(.A1(new_n6956_), .A2(new_n6700_), .ZN(new_n7270_));
  NAND2_X1   g07014(.A1(new_n7269_), .A2(new_n7270_), .ZN(new_n7271_));
  XOR2_X1    g07015(.A1(new_n7271_), .A2(new_n7267_), .Z(new_n7272_));
  XOR2_X1    g07016(.A1(new_n7272_), .A2(new_n7262_), .Z(new_n7273_));
  OAI22_X1   g07017(.A1(new_n582_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n577_), .ZN(new_n7274_));
  NAND2_X1   g07018(.A1(new_n960_), .A2(\b[46] ), .ZN(new_n7275_));
  AOI21_X1   g07019(.A1(new_n7274_), .A2(new_n7275_), .B(new_n585_), .ZN(new_n7276_));
  NAND2_X1   g07020(.A1(new_n5177_), .A2(new_n7276_), .ZN(new_n7277_));
  XOR2_X1    g07021(.A1(new_n7277_), .A2(\a[11] ), .Z(new_n7278_));
  XOR2_X1    g07022(.A1(new_n6956_), .A2(new_n6700_), .Z(new_n7279_));
  XOR2_X1    g07023(.A1(new_n7279_), .A2(new_n6702_), .Z(new_n7280_));
  AOI21_X1   g07024(.A1(new_n7280_), .A2(new_n6695_), .B(new_n6690_), .ZN(new_n7281_));
  NAND2_X1   g07025(.A1(new_n6959_), .A2(new_n7281_), .ZN(new_n7282_));
  XOR2_X1    g07026(.A1(new_n7282_), .A2(new_n7278_), .Z(new_n7283_));
  XOR2_X1    g07027(.A1(new_n7283_), .A2(new_n7273_), .Z(new_n7284_));
  OAI22_X1   g07028(.A1(new_n437_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n431_), .ZN(new_n7285_));
  NAND2_X1   g07029(.A1(new_n775_), .A2(\b[49] ), .ZN(new_n7286_));
  AOI21_X1   g07030(.A1(new_n7285_), .A2(new_n7286_), .B(new_n440_), .ZN(new_n7287_));
  NAND2_X1   g07031(.A1(new_n5741_), .A2(new_n7287_), .ZN(new_n7288_));
  XOR2_X1    g07032(.A1(new_n7288_), .A2(\a[8] ), .Z(new_n7289_));
  NOR2_X1    g07033(.A1(new_n6658_), .A2(new_n6968_), .ZN(new_n7290_));
  NAND2_X1   g07034(.A1(new_n6481_), .A2(new_n7290_), .ZN(new_n7291_));
  NOR2_X1    g07035(.A1(new_n6960_), .A2(new_n6966_), .ZN(new_n7292_));
  NOR2_X1    g07036(.A1(new_n7292_), .A2(new_n7290_), .ZN(new_n7293_));
  NAND3_X1   g07037(.A1(new_n7291_), .A2(new_n6967_), .A3(new_n7293_), .ZN(new_n7294_));
  XOR2_X1    g07038(.A1(new_n7294_), .A2(new_n7289_), .Z(new_n7295_));
  XOR2_X1    g07039(.A1(new_n7295_), .A2(new_n7284_), .Z(new_n7296_));
  OAI22_X1   g07040(.A1(new_n364_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n320_), .ZN(new_n7297_));
  NAND2_X1   g07041(.A1(new_n594_), .A2(\b[52] ), .ZN(new_n7298_));
  AOI21_X1   g07042(.A1(new_n7297_), .A2(new_n7298_), .B(new_n312_), .ZN(new_n7299_));
  NAND2_X1   g07043(.A1(new_n6237_), .A2(new_n7299_), .ZN(new_n7300_));
  XOR2_X1    g07044(.A1(new_n7300_), .A2(new_n308_), .Z(new_n7301_));
  NAND2_X1   g07045(.A1(new_n7296_), .A2(new_n7301_), .ZN(new_n7302_));
  OR2_X2     g07046(.A1(new_n7296_), .A2(new_n7301_), .Z(new_n7303_));
  NAND2_X1   g07047(.A1(new_n7303_), .A2(new_n7302_), .ZN(new_n7304_));
  INV_X1     g07048(.I(\b[57] ), .ZN(new_n7305_));
  XOR2_X1    g07049(.A1(new_n6988_), .A2(\b[55] ), .Z(new_n7306_));
  NAND2_X1   g07050(.A1(new_n7306_), .A2(new_n6990_), .ZN(new_n7307_));
  XOR2_X1    g07051(.A1(new_n7307_), .A2(new_n7305_), .Z(new_n7308_));
  NAND2_X1   g07052(.A1(new_n283_), .A2(\b[57] ), .ZN(new_n7309_));
  NAND2_X1   g07053(.A1(new_n279_), .A2(\b[55] ), .ZN(new_n7310_));
  AOI21_X1   g07054(.A1(\b[56] ), .A2(new_n266_), .B(new_n264_), .ZN(new_n7311_));
  NAND4_X1   g07055(.A1(new_n7308_), .A2(new_n7309_), .A3(new_n7310_), .A4(new_n7311_), .ZN(new_n7312_));
  XOR2_X1    g07056(.A1(new_n7312_), .A2(\a[2] ), .Z(new_n7313_));
  XOR2_X1    g07057(.A1(new_n7304_), .A2(new_n7313_), .Z(new_n7314_));
  XOR2_X1    g07058(.A1(new_n7304_), .A2(new_n7313_), .Z(new_n7315_));
  NOR2_X1    g07059(.A1(new_n7315_), .A2(new_n7010_), .ZN(new_n7316_));
  AOI21_X1   g07060(.A1(new_n7010_), .A2(new_n7314_), .B(new_n7316_), .ZN(new_n7317_));
  AOI21_X1   g07061(.A1(new_n6689_), .A2(new_n7002_), .B(new_n7000_), .ZN(new_n7318_));
  XNOR2_X1   g07062(.A1(new_n7318_), .A2(new_n7317_), .ZN(\f[57] ));
  NOR2_X1    g07063(.A1(new_n7049_), .A2(new_n7059_), .ZN(new_n7320_));
  INV_X1     g07064(.I(new_n7320_), .ZN(new_n7321_));
  NOR2_X1    g07065(.A1(new_n6792_), .A2(new_n6782_), .ZN(new_n7322_));
  NAND2_X1   g07066(.A1(new_n6718_), .A2(new_n6497_), .ZN(new_n7323_));
  AOI21_X1   g07067(.A1(new_n7323_), .A2(new_n6757_), .B(new_n6769_), .ZN(new_n7324_));
  NOR3_X1    g07068(.A1(new_n7040_), .A2(new_n7039_), .A3(new_n7041_), .ZN(new_n7325_));
  AOI21_X1   g07069(.A1(new_n7029_), .A2(new_n7033_), .B(new_n7037_), .ZN(new_n7326_));
  OAI22_X1   g07070(.A1(new_n7325_), .A2(new_n7326_), .B1(new_n7324_), .B2(new_n6768_), .ZN(new_n7327_));
  NOR3_X1    g07071(.A1(new_n7040_), .A2(new_n7039_), .A3(new_n7037_), .ZN(new_n7328_));
  OAI21_X1   g07072(.A1(new_n7045_), .A2(new_n7328_), .B(new_n7012_), .ZN(new_n7329_));
  NAND3_X1   g07073(.A1(new_n7329_), .A2(new_n7327_), .A3(new_n7059_), .ZN(new_n7330_));
  XOR2_X1    g07074(.A1(new_n7057_), .A2(\a[50] ), .Z(new_n7331_));
  OAI21_X1   g07075(.A1(new_n7048_), .A2(new_n7043_), .B(new_n7331_), .ZN(new_n7332_));
  AOI21_X1   g07076(.A1(new_n7332_), .A2(new_n7330_), .B(new_n7062_), .ZN(new_n7333_));
  OAI21_X1   g07077(.A1(new_n6785_), .A2(new_n7322_), .B(new_n7333_), .ZN(new_n7334_));
  NAND2_X1   g07078(.A1(new_n7334_), .A2(new_n7321_), .ZN(new_n7335_));
  AOI21_X1   g07079(.A1(new_n7044_), .A2(new_n7042_), .B(new_n7325_), .ZN(new_n7336_));
  NOR2_X1    g07080(.A1(new_n7026_), .A2(new_n7016_), .ZN(new_n7337_));
  INV_X1     g07081(.I(new_n7337_), .ZN(new_n7338_));
  OAI22_X1   g07082(.A1(new_n6721_), .A2(new_n290_), .B1(new_n6723_), .B2(new_n393_), .ZN(new_n7339_));
  OAI21_X1   g07083(.A1(new_n292_), .A2(new_n6729_), .B(new_n7339_), .ZN(new_n7340_));
  NAND3_X1   g07084(.A1(new_n7340_), .A2(new_n334_), .A3(new_n6512_), .ZN(new_n7341_));
  XOR2_X1    g07085(.A1(new_n7341_), .A2(new_n6516_), .Z(new_n7342_));
  INV_X1     g07086(.I(\a[59] ), .ZN(new_n7343_));
  XOR2_X1    g07087(.A1(\a[56] ), .A2(\a[57] ), .Z(new_n7344_));
  XNOR2_X1   g07088(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n7345_));
  NAND2_X1   g07089(.A1(new_n7345_), .A2(new_n7344_), .ZN(new_n7346_));
  NOR2_X1    g07090(.A1(new_n7346_), .A2(new_n267_), .ZN(new_n7347_));
  INV_X1     g07091(.I(\a[58] ), .ZN(new_n7348_));
  NOR2_X1    g07092(.A1(new_n7014_), .A2(new_n7348_), .ZN(new_n7349_));
  NOR2_X1    g07093(.A1(new_n7013_), .A2(\a[58] ), .ZN(new_n7350_));
  NOR2_X1    g07094(.A1(new_n7349_), .A2(new_n7350_), .ZN(new_n7351_));
  NOR2_X1    g07095(.A1(new_n7351_), .A2(new_n258_), .ZN(new_n7352_));
  XNOR2_X1   g07096(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n7353_));
  OR2_X2     g07097(.A1(new_n7015_), .A2(new_n7353_), .Z(new_n7354_));
  NOR4_X1    g07098(.A1(new_n7347_), .A2(new_n7352_), .A3(new_n7354_), .A4(new_n261_), .ZN(new_n7355_));
  XOR2_X1    g07099(.A1(new_n7355_), .A2(new_n7343_), .Z(new_n7356_));
  NOR2_X1    g07100(.A1(new_n7017_), .A2(\a[59] ), .ZN(new_n7357_));
  XOR2_X1    g07101(.A1(new_n7356_), .A2(new_n7357_), .Z(new_n7358_));
  XOR2_X1    g07102(.A1(new_n7358_), .A2(new_n7342_), .Z(new_n7359_));
  NAND2_X1   g07103(.A1(new_n7359_), .A2(new_n7338_), .ZN(new_n7360_));
  NOR2_X1    g07104(.A1(new_n7358_), .A2(new_n7342_), .ZN(new_n7361_));
  XOR2_X1    g07105(.A1(new_n7341_), .A2(\a[56] ), .Z(new_n7362_));
  XNOR2_X1   g07106(.A1(new_n7356_), .A2(new_n7357_), .ZN(new_n7363_));
  NOR2_X1    g07107(.A1(new_n7363_), .A2(new_n7362_), .ZN(new_n7364_));
  OAI21_X1   g07108(.A1(new_n7364_), .A2(new_n7361_), .B(new_n7337_), .ZN(new_n7365_));
  NAND2_X1   g07109(.A1(new_n7360_), .A2(new_n7365_), .ZN(new_n7366_));
  OAI22_X1   g07110(.A1(new_n5786_), .A2(new_n450_), .B1(new_n403_), .B2(new_n5792_), .ZN(new_n7367_));
  NAND2_X1   g07111(.A1(new_n6745_), .A2(\b[5] ), .ZN(new_n7368_));
  AOI21_X1   g07112(.A1(new_n7368_), .A2(new_n7367_), .B(new_n5796_), .ZN(new_n7369_));
  NAND2_X1   g07113(.A1(new_n454_), .A2(new_n7369_), .ZN(new_n7370_));
  XOR2_X1    g07114(.A1(new_n7370_), .A2(new_n5783_), .Z(new_n7371_));
  XOR2_X1    g07115(.A1(new_n7366_), .A2(new_n7371_), .Z(new_n7372_));
  NOR2_X1    g07116(.A1(new_n7372_), .A2(new_n7336_), .ZN(new_n7373_));
  INV_X1     g07117(.I(new_n7336_), .ZN(new_n7374_));
  NAND3_X1   g07118(.A1(new_n7360_), .A2(new_n7371_), .A3(new_n7365_), .ZN(new_n7375_));
  XOR2_X1    g07119(.A1(new_n7358_), .A2(new_n7362_), .Z(new_n7376_));
  NOR2_X1    g07120(.A1(new_n7376_), .A2(new_n7337_), .ZN(new_n7377_));
  INV_X1     g07121(.I(new_n7365_), .ZN(new_n7378_));
  XOR2_X1    g07122(.A1(new_n7370_), .A2(\a[53] ), .Z(new_n7379_));
  OAI21_X1   g07123(.A1(new_n7377_), .A2(new_n7378_), .B(new_n7379_), .ZN(new_n7380_));
  AOI21_X1   g07124(.A1(new_n7380_), .A2(new_n7375_), .B(new_n7374_), .ZN(new_n7381_));
  NOR2_X1    g07125(.A1(new_n7373_), .A2(new_n7381_), .ZN(new_n7382_));
  OAI22_X1   g07126(.A1(new_n5228_), .A2(new_n617_), .B1(new_n510_), .B2(new_n5225_), .ZN(new_n7383_));
  NAND2_X1   g07127(.A1(new_n5387_), .A2(\b[8] ), .ZN(new_n7384_));
  AOI21_X1   g07128(.A1(new_n7383_), .A2(new_n7384_), .B(new_n5231_), .ZN(new_n7385_));
  NAND2_X1   g07129(.A1(new_n616_), .A2(new_n7385_), .ZN(new_n7386_));
  XOR2_X1    g07130(.A1(new_n7386_), .A2(\a[50] ), .Z(new_n7387_));
  NOR2_X1    g07131(.A1(new_n7382_), .A2(new_n7387_), .ZN(new_n7388_));
  INV_X1     g07132(.I(new_n7382_), .ZN(new_n7389_));
  INV_X1     g07133(.I(new_n7387_), .ZN(new_n7390_));
  NOR2_X1    g07134(.A1(new_n7389_), .A2(new_n7390_), .ZN(new_n7391_));
  OAI21_X1   g07135(.A1(new_n7391_), .A2(new_n7388_), .B(new_n7335_), .ZN(new_n7392_));
  NOR3_X1    g07136(.A1(new_n7048_), .A2(new_n7043_), .A3(new_n7331_), .ZN(new_n7393_));
  AOI21_X1   g07137(.A1(new_n7329_), .A2(new_n7327_), .B(new_n7059_), .ZN(new_n7394_));
  OAI21_X1   g07138(.A1(new_n7393_), .A2(new_n7394_), .B(new_n7063_), .ZN(new_n7395_));
  AOI21_X1   g07139(.A1(new_n6790_), .A2(new_n7060_), .B(new_n7395_), .ZN(new_n7396_));
  NOR2_X1    g07140(.A1(new_n7396_), .A2(new_n7320_), .ZN(new_n7397_));
  NOR2_X1    g07141(.A1(new_n7389_), .A2(new_n7387_), .ZN(new_n7398_));
  NOR2_X1    g07142(.A1(new_n7382_), .A2(new_n7390_), .ZN(new_n7399_));
  OAI21_X1   g07143(.A1(new_n7398_), .A2(new_n7399_), .B(new_n7397_), .ZN(new_n7400_));
  NAND2_X1   g07144(.A1(new_n7392_), .A2(new_n7400_), .ZN(new_n7401_));
  OAI22_X1   g07145(.A1(new_n4711_), .A2(new_n795_), .B1(new_n717_), .B2(new_n4706_), .ZN(new_n7402_));
  NAND2_X1   g07146(.A1(new_n5814_), .A2(\b[11] ), .ZN(new_n7403_));
  AOI21_X1   g07147(.A1(new_n7402_), .A2(new_n7403_), .B(new_n4714_), .ZN(new_n7404_));
  NAND2_X1   g07148(.A1(new_n799_), .A2(new_n7404_), .ZN(new_n7405_));
  XOR2_X1    g07149(.A1(new_n7405_), .A2(\a[47] ), .Z(new_n7406_));
  INV_X1     g07150(.I(new_n7406_), .ZN(new_n7407_));
  NAND2_X1   g07151(.A1(new_n7401_), .A2(new_n7407_), .ZN(new_n7408_));
  NAND3_X1   g07152(.A1(new_n7400_), .A2(new_n7392_), .A3(new_n7406_), .ZN(new_n7409_));
  NAND2_X1   g07153(.A1(new_n7408_), .A2(new_n7409_), .ZN(new_n7410_));
  OAI22_X1   g07154(.A1(new_n4208_), .A2(new_n992_), .B1(new_n904_), .B2(new_n4203_), .ZN(new_n7411_));
  NAND2_X1   g07155(.A1(new_n5244_), .A2(\b[14] ), .ZN(new_n7412_));
  AOI21_X1   g07156(.A1(new_n7411_), .A2(new_n7412_), .B(new_n4211_), .ZN(new_n7413_));
  NAND2_X1   g07157(.A1(new_n991_), .A2(new_n7413_), .ZN(new_n7414_));
  XOR2_X1    g07158(.A1(new_n7414_), .A2(\a[44] ), .Z(new_n7415_));
  INV_X1     g07159(.I(new_n7415_), .ZN(new_n7416_));
  NAND2_X1   g07160(.A1(new_n7410_), .A2(new_n7416_), .ZN(new_n7417_));
  NAND3_X1   g07161(.A1(new_n7408_), .A2(new_n7409_), .A3(new_n7415_), .ZN(new_n7418_));
  NAND2_X1   g07162(.A1(new_n7417_), .A2(new_n7418_), .ZN(new_n7419_));
  OAI22_X1   g07163(.A1(new_n3736_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n3731_), .ZN(new_n7420_));
  NAND2_X1   g07164(.A1(new_n4730_), .A2(\b[17] ), .ZN(new_n7421_));
  AOI21_X1   g07165(.A1(new_n7420_), .A2(new_n7421_), .B(new_n3739_), .ZN(new_n7422_));
  NAND2_X1   g07166(.A1(new_n1225_), .A2(new_n7422_), .ZN(new_n7423_));
  XOR2_X1    g07167(.A1(new_n7423_), .A2(\a[41] ), .Z(new_n7424_));
  OAI21_X1   g07168(.A1(new_n7121_), .A2(new_n7119_), .B(new_n7118_), .ZN(new_n7425_));
  NAND2_X1   g07169(.A1(new_n7425_), .A2(new_n7424_), .ZN(new_n7426_));
  INV_X1     g07170(.I(new_n7424_), .ZN(new_n7427_));
  NAND3_X1   g07171(.A1(new_n7118_), .A2(new_n7115_), .A3(new_n7123_), .ZN(new_n7428_));
  NAND3_X1   g07172(.A1(new_n7428_), .A2(new_n7118_), .A3(new_n7427_), .ZN(new_n7429_));
  AOI21_X1   g07173(.A1(new_n7426_), .A2(new_n7429_), .B(new_n7419_), .ZN(new_n7430_));
  INV_X1     g07174(.I(new_n7419_), .ZN(new_n7431_));
  AOI21_X1   g07175(.A1(new_n7428_), .A2(new_n7118_), .B(new_n7427_), .ZN(new_n7432_));
  NOR2_X1    g07176(.A1(new_n7425_), .A2(new_n7424_), .ZN(new_n7433_));
  NOR3_X1    g07177(.A1(new_n7433_), .A2(new_n7432_), .A3(new_n7431_), .ZN(new_n7434_));
  OAI22_X1   g07178(.A1(new_n3298_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n3293_), .ZN(new_n7435_));
  NAND2_X1   g07179(.A1(new_n4227_), .A2(\b[20] ), .ZN(new_n7436_));
  AOI21_X1   g07180(.A1(new_n7435_), .A2(new_n7436_), .B(new_n3301_), .ZN(new_n7437_));
  NAND2_X1   g07181(.A1(new_n1517_), .A2(new_n7437_), .ZN(new_n7438_));
  XOR2_X1    g07182(.A1(new_n7438_), .A2(\a[38] ), .Z(new_n7439_));
  INV_X1     g07183(.I(new_n7439_), .ZN(new_n7440_));
  OAI21_X1   g07184(.A1(new_n7434_), .A2(new_n7430_), .B(new_n7440_), .ZN(new_n7441_));
  OAI21_X1   g07185(.A1(new_n7433_), .A2(new_n7432_), .B(new_n7431_), .ZN(new_n7442_));
  NAND3_X1   g07186(.A1(new_n7426_), .A2(new_n7429_), .A3(new_n7419_), .ZN(new_n7443_));
  NAND3_X1   g07187(.A1(new_n7442_), .A2(new_n7443_), .A3(new_n7439_), .ZN(new_n7444_));
  NAND2_X1   g07188(.A1(new_n7441_), .A2(new_n7444_), .ZN(new_n7445_));
  OAI21_X1   g07189(.A1(new_n7156_), .A2(new_n7158_), .B(new_n7135_), .ZN(new_n7446_));
  OAI22_X1   g07190(.A1(new_n2846_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n2841_), .ZN(new_n7447_));
  NAND2_X1   g07191(.A1(new_n3755_), .A2(\b[23] ), .ZN(new_n7448_));
  AOI21_X1   g07192(.A1(new_n7447_), .A2(new_n7448_), .B(new_n2849_), .ZN(new_n7449_));
  NAND2_X1   g07193(.A1(new_n1828_), .A2(new_n7449_), .ZN(new_n7450_));
  XOR2_X1    g07194(.A1(new_n7450_), .A2(\a[35] ), .Z(new_n7451_));
  INV_X1     g07195(.I(new_n7451_), .ZN(new_n7452_));
  NAND2_X1   g07196(.A1(new_n7446_), .A2(new_n7452_), .ZN(new_n7453_));
  AOI21_X1   g07197(.A1(new_n7011_), .A2(new_n7138_), .B(new_n7157_), .ZN(new_n7454_));
  NAND2_X1   g07198(.A1(new_n7454_), .A2(new_n7451_), .ZN(new_n7455_));
  NAND2_X1   g07199(.A1(new_n7455_), .A2(new_n7453_), .ZN(new_n7456_));
  NAND2_X1   g07200(.A1(new_n7445_), .A2(new_n7456_), .ZN(new_n7457_));
  XOR2_X1    g07201(.A1(new_n7446_), .A2(new_n7452_), .Z(new_n7458_));
  NAND3_X1   g07202(.A1(new_n7458_), .A2(new_n7441_), .A3(new_n7444_), .ZN(new_n7459_));
  OAI22_X1   g07203(.A1(new_n2452_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n2447_), .ZN(new_n7460_));
  NAND2_X1   g07204(.A1(new_n3312_), .A2(\b[26] ), .ZN(new_n7461_));
  AOI21_X1   g07205(.A1(new_n7460_), .A2(new_n7461_), .B(new_n2455_), .ZN(new_n7462_));
  NAND2_X1   g07206(.A1(new_n2174_), .A2(new_n7462_), .ZN(new_n7463_));
  XOR2_X1    g07207(.A1(new_n7463_), .A2(\a[32] ), .Z(new_n7464_));
  INV_X1     g07208(.I(new_n7464_), .ZN(new_n7465_));
  AOI21_X1   g07209(.A1(new_n7459_), .A2(new_n7457_), .B(new_n7465_), .ZN(new_n7466_));
  INV_X1     g07210(.I(new_n7457_), .ZN(new_n7467_));
  XOR2_X1    g07211(.A1(new_n7446_), .A2(new_n7451_), .Z(new_n7468_));
  NOR2_X1    g07212(.A1(new_n7468_), .A2(new_n7445_), .ZN(new_n7469_));
  NOR3_X1    g07213(.A1(new_n7467_), .A2(new_n7469_), .A3(new_n7464_), .ZN(new_n7470_));
  NOR2_X1    g07214(.A1(new_n7470_), .A2(new_n7466_), .ZN(new_n7471_));
  OAI22_X1   g07215(.A1(new_n2084_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n2079_), .ZN(new_n7472_));
  NAND2_X1   g07216(.A1(new_n2864_), .A2(\b[29] ), .ZN(new_n7473_));
  AOI21_X1   g07217(.A1(new_n7472_), .A2(new_n7473_), .B(new_n2087_), .ZN(new_n7474_));
  NAND2_X1   g07218(.A1(new_n2546_), .A2(new_n7474_), .ZN(new_n7475_));
  XOR2_X1    g07219(.A1(new_n7475_), .A2(\a[29] ), .Z(new_n7476_));
  NOR2_X1    g07220(.A1(new_n7471_), .A2(new_n7476_), .ZN(new_n7477_));
  INV_X1     g07221(.I(new_n7471_), .ZN(new_n7478_));
  INV_X1     g07222(.I(new_n7476_), .ZN(new_n7479_));
  NOR2_X1    g07223(.A1(new_n7478_), .A2(new_n7479_), .ZN(new_n7480_));
  NOR2_X1    g07224(.A1(new_n7480_), .A2(new_n7477_), .ZN(new_n7481_));
  OAI22_X1   g07225(.A1(new_n1760_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n1755_), .ZN(new_n7482_));
  NAND2_X1   g07226(.A1(new_n2470_), .A2(\b[32] ), .ZN(new_n7483_));
  AOI21_X1   g07227(.A1(new_n7482_), .A2(new_n7483_), .B(new_n1763_), .ZN(new_n7484_));
  NAND2_X1   g07228(.A1(new_n2963_), .A2(new_n7484_), .ZN(new_n7485_));
  XOR2_X1    g07229(.A1(new_n7485_), .A2(\a[26] ), .Z(new_n7486_));
  NOR2_X1    g07230(.A1(new_n7481_), .A2(new_n7486_), .ZN(new_n7487_));
  INV_X1     g07231(.I(new_n7487_), .ZN(new_n7488_));
  NAND2_X1   g07232(.A1(new_n7481_), .A2(new_n7486_), .ZN(new_n7489_));
  OAI22_X1   g07233(.A1(new_n1444_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n1439_), .ZN(new_n7490_));
  NAND2_X1   g07234(.A1(new_n2098_), .A2(\b[35] ), .ZN(new_n7491_));
  AOI21_X1   g07235(.A1(new_n7490_), .A2(new_n7491_), .B(new_n1447_), .ZN(new_n7492_));
  NAND2_X1   g07236(.A1(new_n3411_), .A2(new_n7492_), .ZN(new_n7493_));
  XOR2_X1    g07237(.A1(new_n7493_), .A2(\a[23] ), .Z(new_n7494_));
  INV_X1     g07238(.I(new_n7494_), .ZN(new_n7495_));
  AOI21_X1   g07239(.A1(new_n7488_), .A2(new_n7489_), .B(new_n7495_), .ZN(new_n7496_));
  INV_X1     g07240(.I(new_n7489_), .ZN(new_n7497_));
  NOR3_X1    g07241(.A1(new_n7497_), .A2(new_n7487_), .A3(new_n7494_), .ZN(new_n7498_));
  NOR2_X1    g07242(.A1(new_n7496_), .A2(new_n7498_), .ZN(new_n7499_));
  OAI22_X1   g07243(.A1(new_n1168_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n1163_), .ZN(new_n7500_));
  NAND2_X1   g07244(.A1(new_n1774_), .A2(\b[38] ), .ZN(new_n7501_));
  AOI21_X1   g07245(.A1(new_n7500_), .A2(new_n7501_), .B(new_n1171_), .ZN(new_n7502_));
  NAND2_X1   g07246(.A1(new_n3844_), .A2(new_n7502_), .ZN(new_n7503_));
  XOR2_X1    g07247(.A1(new_n7503_), .A2(\a[20] ), .Z(new_n7504_));
  INV_X1     g07248(.I(new_n7237_), .ZN(new_n7505_));
  OAI21_X1   g07249(.A1(new_n7230_), .A2(new_n7229_), .B(new_n7228_), .ZN(new_n7506_));
  NAND3_X1   g07250(.A1(new_n7220_), .A2(new_n7211_), .A3(new_n7224_), .ZN(new_n7507_));
  NAND3_X1   g07251(.A1(new_n7506_), .A2(new_n7507_), .A3(new_n7505_), .ZN(new_n7508_));
  OAI21_X1   g07252(.A1(new_n7231_), .A2(new_n7225_), .B(new_n7237_), .ZN(new_n7509_));
  AOI22_X1   g07253(.A1(new_n7509_), .A2(new_n7508_), .B1(new_n7505_), .B2(new_n7240_), .ZN(new_n7510_));
  XOR2_X1    g07254(.A1(new_n7510_), .A2(new_n7504_), .Z(new_n7511_));
  XOR2_X1    g07255(.A1(new_n7511_), .A2(new_n7499_), .Z(new_n7512_));
  OAI22_X1   g07256(.A1(new_n940_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n935_), .ZN(new_n7513_));
  NAND2_X1   g07257(.A1(new_n1458_), .A2(\b[41] ), .ZN(new_n7514_));
  AOI21_X1   g07258(.A1(new_n7513_), .A2(new_n7514_), .B(new_n943_), .ZN(new_n7515_));
  NAND2_X1   g07259(.A1(new_n4320_), .A2(new_n7515_), .ZN(new_n7516_));
  XOR2_X1    g07260(.A1(new_n7516_), .A2(\a[17] ), .Z(new_n7517_));
  XNOR2_X1   g07261(.A1(new_n7512_), .A2(new_n7517_), .ZN(new_n7518_));
  OAI22_X1   g07262(.A1(new_n757_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n752_), .ZN(new_n7519_));
  NAND2_X1   g07263(.A1(new_n1182_), .A2(\b[44] ), .ZN(new_n7520_));
  AOI21_X1   g07264(.A1(new_n7519_), .A2(new_n7520_), .B(new_n760_), .ZN(new_n7521_));
  NAND2_X1   g07265(.A1(new_n4833_), .A2(new_n7521_), .ZN(new_n7522_));
  XOR2_X1    g07266(.A1(new_n7522_), .A2(\a[14] ), .Z(new_n7523_));
  NOR2_X1    g07267(.A1(new_n7518_), .A2(new_n7523_), .ZN(new_n7524_));
  AND2_X2    g07268(.A1(new_n7518_), .A2(new_n7523_), .Z(new_n7525_));
  NOR2_X1    g07269(.A1(new_n7525_), .A2(new_n7524_), .ZN(new_n7526_));
  OAI22_X1   g07270(.A1(new_n582_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n577_), .ZN(new_n7527_));
  NAND2_X1   g07271(.A1(new_n960_), .A2(\b[47] ), .ZN(new_n7528_));
  AOI21_X1   g07272(.A1(new_n7527_), .A2(new_n7528_), .B(new_n585_), .ZN(new_n7529_));
  NAND2_X1   g07273(.A1(new_n5196_), .A2(new_n7529_), .ZN(new_n7530_));
  XOR2_X1    g07274(.A1(new_n7530_), .A2(\a[11] ), .Z(new_n7531_));
  XOR2_X1    g07275(.A1(new_n7526_), .A2(new_n7531_), .Z(new_n7532_));
  OAI22_X1   g07276(.A1(new_n437_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n431_), .ZN(new_n7533_));
  NAND2_X1   g07277(.A1(new_n775_), .A2(\b[50] ), .ZN(new_n7534_));
  AOI21_X1   g07278(.A1(new_n7533_), .A2(new_n7534_), .B(new_n440_), .ZN(new_n7535_));
  NAND2_X1   g07279(.A1(new_n5954_), .A2(new_n7535_), .ZN(new_n7536_));
  XOR2_X1    g07280(.A1(new_n7536_), .A2(\a[8] ), .Z(new_n7537_));
  XNOR2_X1   g07281(.A1(new_n7532_), .A2(new_n7537_), .ZN(new_n7538_));
  OAI22_X1   g07282(.A1(new_n364_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n320_), .ZN(new_n7539_));
  NAND2_X1   g07283(.A1(new_n594_), .A2(\b[53] ), .ZN(new_n7540_));
  AOI21_X1   g07284(.A1(new_n7539_), .A2(new_n7540_), .B(new_n312_), .ZN(new_n7541_));
  NAND2_X1   g07285(.A1(new_n6471_), .A2(new_n7541_), .ZN(new_n7542_));
  XOR2_X1    g07286(.A1(new_n7542_), .A2(\a[5] ), .Z(new_n7543_));
  XOR2_X1    g07287(.A1(new_n7538_), .A2(new_n7543_), .Z(new_n7544_));
  XOR2_X1    g07288(.A1(new_n7010_), .A2(new_n7301_), .Z(new_n7545_));
  NAND2_X1   g07289(.A1(new_n7545_), .A2(new_n7296_), .ZN(new_n7546_));
  XOR2_X1    g07290(.A1(new_n7546_), .A2(new_n7544_), .Z(new_n7547_));
  NAND2_X1   g07291(.A1(new_n7010_), .A2(new_n7301_), .ZN(new_n7548_));
  XOR2_X1    g07292(.A1(new_n7547_), .A2(new_n7548_), .Z(new_n7549_));
  OAI21_X1   g07293(.A1(new_n6467_), .A2(new_n7305_), .B(new_n6995_), .ZN(new_n7550_));
  NAND3_X1   g07294(.A1(new_n6986_), .A2(new_n6987_), .A3(new_n7550_), .ZN(new_n7551_));
  OAI21_X1   g07295(.A1(\b[55] ), .A2(\b[57] ), .B(\b[56] ), .ZN(new_n7552_));
  NAND2_X1   g07296(.A1(new_n7551_), .A2(new_n7552_), .ZN(new_n7553_));
  XNOR2_X1   g07297(.A1(\b[57] ), .A2(\b[58] ), .ZN(new_n7554_));
  INV_X1     g07298(.I(new_n7554_), .ZN(new_n7555_));
  XOR2_X1    g07299(.A1(\b[57] ), .A2(\b[58] ), .Z(new_n7556_));
  NOR2_X1    g07300(.A1(new_n7553_), .A2(new_n7556_), .ZN(new_n7557_));
  AOI21_X1   g07301(.A1(new_n7553_), .A2(new_n7555_), .B(new_n7557_), .ZN(new_n7558_));
  INV_X1     g07302(.I(new_n7558_), .ZN(new_n7559_));
  INV_X1     g07303(.I(\b[58] ), .ZN(new_n7560_));
  OAI22_X1   g07304(.A1(new_n405_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n404_), .ZN(new_n7561_));
  NAND2_X1   g07305(.A1(new_n279_), .A2(\b[56] ), .ZN(new_n7562_));
  AOI21_X1   g07306(.A1(new_n7561_), .A2(new_n7562_), .B(new_n264_), .ZN(new_n7563_));
  NAND2_X1   g07307(.A1(new_n7559_), .A2(new_n7563_), .ZN(new_n7564_));
  XOR2_X1    g07308(.A1(new_n7564_), .A2(\a[2] ), .Z(new_n7565_));
  XOR2_X1    g07309(.A1(new_n7549_), .A2(new_n7565_), .Z(new_n7566_));
  INV_X1     g07310(.I(new_n7005_), .ZN(new_n7567_));
  NAND2_X1   g07311(.A1(new_n7317_), .A2(new_n7567_), .ZN(new_n7568_));
  AOI21_X1   g07312(.A1(new_n6689_), .A2(new_n7005_), .B(new_n7568_), .ZN(new_n7569_));
  INV_X1     g07313(.I(new_n7313_), .ZN(new_n7570_));
  XNOR2_X1   g07314(.A1(new_n7010_), .A2(new_n7304_), .ZN(new_n7571_));
  NOR2_X1    g07315(.A1(new_n7571_), .A2(new_n7570_), .ZN(new_n7572_));
  INV_X1     g07316(.I(new_n7572_), .ZN(new_n7573_));
  AND2_X2    g07317(.A1(new_n7569_), .A2(new_n7573_), .Z(new_n7574_));
  NAND3_X1   g07318(.A1(new_n7569_), .A2(new_n7566_), .A3(new_n7573_), .ZN(new_n7575_));
  OAI21_X1   g07319(.A1(new_n7574_), .A2(new_n7566_), .B(new_n7575_), .ZN(\f[58] ));
  NOR3_X1    g07320(.A1(new_n7525_), .A2(new_n7524_), .A3(new_n7531_), .ZN(new_n7577_));
  INV_X1     g07321(.I(new_n7577_), .ZN(new_n7578_));
  INV_X1     g07322(.I(new_n7524_), .ZN(new_n7579_));
  NOR2_X1    g07323(.A1(new_n7512_), .A2(new_n7517_), .ZN(new_n7580_));
  INV_X1     g07324(.I(new_n7580_), .ZN(new_n7581_));
  INV_X1     g07325(.I(new_n7504_), .ZN(new_n7582_));
  XOR2_X1    g07326(.A1(new_n7510_), .A2(new_n7499_), .Z(new_n7583_));
  NOR2_X1    g07327(.A1(new_n7583_), .A2(new_n7582_), .ZN(new_n7584_));
  NOR2_X1    g07328(.A1(new_n7478_), .A2(new_n7476_), .ZN(new_n7585_));
  INV_X1     g07329(.I(new_n7585_), .ZN(new_n7586_));
  OAI22_X1   g07330(.A1(new_n2084_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n2079_), .ZN(new_n7587_));
  NAND2_X1   g07331(.A1(new_n2864_), .A2(\b[30] ), .ZN(new_n7588_));
  AOI21_X1   g07332(.A1(new_n7587_), .A2(new_n7588_), .B(new_n2087_), .ZN(new_n7589_));
  NAND2_X1   g07333(.A1(new_n2659_), .A2(new_n7589_), .ZN(new_n7590_));
  XOR2_X1    g07334(.A1(new_n7590_), .A2(\a[29] ), .Z(new_n7591_));
  OAI22_X1   g07335(.A1(new_n2452_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n2447_), .ZN(new_n7592_));
  NAND2_X1   g07336(.A1(new_n3312_), .A2(\b[27] ), .ZN(new_n7593_));
  AOI21_X1   g07337(.A1(new_n7592_), .A2(new_n7593_), .B(new_n2455_), .ZN(new_n7594_));
  NAND2_X1   g07338(.A1(new_n2276_), .A2(new_n7594_), .ZN(new_n7595_));
  XOR2_X1    g07339(.A1(new_n7595_), .A2(\a[32] ), .Z(new_n7596_));
  INV_X1     g07340(.I(new_n7596_), .ZN(new_n7597_));
  OAI21_X1   g07341(.A1(new_n7467_), .A2(new_n7469_), .B(new_n7464_), .ZN(new_n7598_));
  AOI21_X1   g07342(.A1(new_n7360_), .A2(new_n7365_), .B(new_n7371_), .ZN(new_n7599_));
  OAI21_X1   g07343(.A1(new_n7599_), .A2(new_n7336_), .B(new_n7375_), .ZN(new_n7600_));
  NAND2_X1   g07344(.A1(new_n7358_), .A2(new_n7342_), .ZN(new_n7601_));
  OAI21_X1   g07345(.A1(new_n7337_), .A2(new_n7361_), .B(new_n7601_), .ZN(new_n7602_));
  NOR4_X1    g07346(.A1(new_n7355_), .A2(\a[59] ), .A3(\b[0] ), .A4(new_n7344_), .ZN(new_n7603_));
  INV_X1     g07347(.I(new_n7354_), .ZN(new_n7604_));
  NOR2_X1    g07348(.A1(new_n7351_), .A2(new_n267_), .ZN(new_n7605_));
  NOR2_X1    g07349(.A1(new_n7346_), .A2(new_n292_), .ZN(new_n7606_));
  XNOR2_X1   g07350(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n7607_));
  XNOR2_X1   g07351(.A1(\a[56] ), .A2(\a[58] ), .ZN(new_n7608_));
  NAND2_X1   g07352(.A1(new_n7607_), .A2(new_n7608_), .ZN(new_n7609_));
  XNOR2_X1   g07353(.A1(\a[56] ), .A2(\a[59] ), .ZN(new_n7610_));
  NAND2_X1   g07354(.A1(new_n7609_), .A2(new_n7610_), .ZN(new_n7611_));
  OAI22_X1   g07355(.A1(new_n7605_), .A2(new_n7606_), .B1(new_n7611_), .B2(new_n258_), .ZN(new_n7612_));
  NAND3_X1   g07356(.A1(new_n7612_), .A2(new_n5389_), .A3(new_n7604_), .ZN(new_n7613_));
  XOR2_X1    g07357(.A1(new_n7613_), .A2(\a[59] ), .Z(new_n7614_));
  XOR2_X1    g07358(.A1(new_n7614_), .A2(new_n7603_), .Z(new_n7615_));
  OAI22_X1   g07359(.A1(new_n6721_), .A2(new_n393_), .B1(new_n6723_), .B2(new_n347_), .ZN(new_n7616_));
  INV_X1     g07360(.I(new_n6729_), .ZN(new_n7617_));
  NAND2_X1   g07361(.A1(new_n7617_), .A2(\b[3] ), .ZN(new_n7618_));
  AOI21_X1   g07362(.A1(new_n7618_), .A2(new_n7616_), .B(new_n6731_), .ZN(new_n7619_));
  NAND2_X1   g07363(.A1(new_n352_), .A2(new_n7619_), .ZN(new_n7620_));
  XOR2_X1    g07364(.A1(new_n7620_), .A2(\a[56] ), .Z(new_n7621_));
  NOR2_X1    g07365(.A1(new_n7621_), .A2(new_n7615_), .ZN(new_n7622_));
  XOR2_X1    g07366(.A1(new_n7613_), .A2(new_n7343_), .Z(new_n7623_));
  XOR2_X1    g07367(.A1(new_n7623_), .A2(new_n7603_), .Z(new_n7624_));
  XOR2_X1    g07368(.A1(new_n7620_), .A2(new_n6516_), .Z(new_n7625_));
  NOR2_X1    g07369(.A1(new_n7625_), .A2(new_n7624_), .ZN(new_n7626_));
  OAI21_X1   g07370(.A1(new_n7622_), .A2(new_n7626_), .B(new_n7602_), .ZN(new_n7627_));
  NAND2_X1   g07371(.A1(new_n7363_), .A2(new_n7362_), .ZN(new_n7628_));
  AOI21_X1   g07372(.A1(new_n7338_), .A2(new_n7628_), .B(new_n7364_), .ZN(new_n7629_));
  NOR2_X1    g07373(.A1(new_n7621_), .A2(new_n7624_), .ZN(new_n7630_));
  NOR2_X1    g07374(.A1(new_n7625_), .A2(new_n7615_), .ZN(new_n7631_));
  OAI21_X1   g07375(.A1(new_n7630_), .A2(new_n7631_), .B(new_n7629_), .ZN(new_n7632_));
  OAI22_X1   g07376(.A1(new_n5786_), .A2(new_n495_), .B1(new_n450_), .B2(new_n5792_), .ZN(new_n7633_));
  NAND2_X1   g07377(.A1(new_n6745_), .A2(\b[6] ), .ZN(new_n7634_));
  AOI21_X1   g07378(.A1(new_n7634_), .A2(new_n7633_), .B(new_n5796_), .ZN(new_n7635_));
  NAND2_X1   g07379(.A1(new_n494_), .A2(new_n7635_), .ZN(new_n7636_));
  XOR2_X1    g07380(.A1(new_n7636_), .A2(new_n5783_), .Z(new_n7637_));
  NAND3_X1   g07381(.A1(new_n7632_), .A2(new_n7627_), .A3(new_n7637_), .ZN(new_n7638_));
  NAND2_X1   g07382(.A1(new_n7625_), .A2(new_n7624_), .ZN(new_n7639_));
  NAND2_X1   g07383(.A1(new_n7621_), .A2(new_n7615_), .ZN(new_n7640_));
  AOI21_X1   g07384(.A1(new_n7639_), .A2(new_n7640_), .B(new_n7629_), .ZN(new_n7641_));
  NAND2_X1   g07385(.A1(new_n7625_), .A2(new_n7615_), .ZN(new_n7642_));
  NAND2_X1   g07386(.A1(new_n7621_), .A2(new_n7624_), .ZN(new_n7643_));
  AOI21_X1   g07387(.A1(new_n7642_), .A2(new_n7643_), .B(new_n7602_), .ZN(new_n7644_));
  XOR2_X1    g07388(.A1(new_n7636_), .A2(\a[53] ), .Z(new_n7645_));
  OAI21_X1   g07389(.A1(new_n7641_), .A2(new_n7644_), .B(new_n7645_), .ZN(new_n7646_));
  NAND2_X1   g07390(.A1(new_n7646_), .A2(new_n7638_), .ZN(new_n7647_));
  NAND2_X1   g07391(.A1(new_n7647_), .A2(new_n7600_), .ZN(new_n7648_));
  NOR3_X1    g07392(.A1(new_n7377_), .A2(new_n7379_), .A3(new_n7378_), .ZN(new_n7649_));
  AOI21_X1   g07393(.A1(new_n7374_), .A2(new_n7380_), .B(new_n7649_), .ZN(new_n7650_));
  NOR3_X1    g07394(.A1(new_n7641_), .A2(new_n7644_), .A3(new_n7645_), .ZN(new_n7651_));
  AOI21_X1   g07395(.A1(new_n7632_), .A2(new_n7627_), .B(new_n7637_), .ZN(new_n7652_));
  NOR2_X1    g07396(.A1(new_n7652_), .A2(new_n7651_), .ZN(new_n7653_));
  NAND2_X1   g07397(.A1(new_n7653_), .A2(new_n7650_), .ZN(new_n7654_));
  OAI22_X1   g07398(.A1(new_n5228_), .A2(new_n659_), .B1(new_n617_), .B2(new_n5225_), .ZN(new_n7655_));
  NAND2_X1   g07399(.A1(new_n5387_), .A2(\b[9] ), .ZN(new_n7656_));
  AOI21_X1   g07400(.A1(new_n7655_), .A2(new_n7656_), .B(new_n5231_), .ZN(new_n7657_));
  OAI21_X1   g07401(.A1(new_n661_), .A2(new_n662_), .B(new_n7657_), .ZN(new_n7658_));
  XOR2_X1    g07402(.A1(new_n7658_), .A2(\a[50] ), .Z(new_n7659_));
  AOI21_X1   g07403(.A1(new_n7654_), .A2(new_n7648_), .B(new_n7659_), .ZN(new_n7660_));
  NOR2_X1    g07404(.A1(new_n7653_), .A2(new_n7650_), .ZN(new_n7661_));
  NOR2_X1    g07405(.A1(new_n7647_), .A2(new_n7600_), .ZN(new_n7662_));
  INV_X1     g07406(.I(new_n7659_), .ZN(new_n7663_));
  NOR3_X1    g07407(.A1(new_n7661_), .A2(new_n7662_), .A3(new_n7663_), .ZN(new_n7664_));
  NOR2_X1    g07408(.A1(new_n7664_), .A2(new_n7660_), .ZN(new_n7665_));
  NAND3_X1   g07409(.A1(new_n7334_), .A2(new_n7321_), .A3(new_n7390_), .ZN(new_n7666_));
  OAI21_X1   g07410(.A1(new_n7396_), .A2(new_n7320_), .B(new_n7387_), .ZN(new_n7667_));
  NAND2_X1   g07411(.A1(new_n7667_), .A2(new_n7666_), .ZN(new_n7668_));
  NAND3_X1   g07412(.A1(new_n7668_), .A2(new_n7382_), .A3(new_n7665_), .ZN(new_n7669_));
  OR2_X2     g07413(.A1(new_n7664_), .A2(new_n7660_), .Z(new_n7670_));
  NOR3_X1    g07414(.A1(new_n7396_), .A2(new_n7320_), .A3(new_n7387_), .ZN(new_n7671_));
  AOI21_X1   g07415(.A1(new_n7334_), .A2(new_n7321_), .B(new_n7390_), .ZN(new_n7672_));
  OAI21_X1   g07416(.A1(new_n7671_), .A2(new_n7672_), .B(new_n7382_), .ZN(new_n7673_));
  NAND2_X1   g07417(.A1(new_n7673_), .A2(new_n7670_), .ZN(new_n7674_));
  NOR2_X1    g07418(.A1(new_n7397_), .A2(new_n7387_), .ZN(new_n7675_));
  NAND3_X1   g07419(.A1(new_n7674_), .A2(new_n7669_), .A3(new_n7675_), .ZN(new_n7676_));
  NOR2_X1    g07420(.A1(new_n7673_), .A2(new_n7670_), .ZN(new_n7677_));
  AOI21_X1   g07421(.A1(new_n7668_), .A2(new_n7382_), .B(new_n7665_), .ZN(new_n7678_));
  NAND2_X1   g07422(.A1(new_n7335_), .A2(new_n7390_), .ZN(new_n7679_));
  OAI21_X1   g07423(.A1(new_n7677_), .A2(new_n7678_), .B(new_n7679_), .ZN(new_n7680_));
  OAI22_X1   g07424(.A1(new_n4711_), .A2(new_n848_), .B1(new_n795_), .B2(new_n4706_), .ZN(new_n7681_));
  NAND2_X1   g07425(.A1(new_n5814_), .A2(\b[12] ), .ZN(new_n7682_));
  AOI21_X1   g07426(.A1(new_n7681_), .A2(new_n7682_), .B(new_n4714_), .ZN(new_n7683_));
  NAND2_X1   g07427(.A1(new_n847_), .A2(new_n7683_), .ZN(new_n7684_));
  XOR2_X1    g07428(.A1(new_n7684_), .A2(\a[47] ), .Z(new_n7685_));
  INV_X1     g07429(.I(new_n7685_), .ZN(new_n7686_));
  NAND3_X1   g07430(.A1(new_n7680_), .A2(new_n7676_), .A3(new_n7686_), .ZN(new_n7687_));
  NOR3_X1    g07431(.A1(new_n7677_), .A2(new_n7678_), .A3(new_n7679_), .ZN(new_n7688_));
  AOI21_X1   g07432(.A1(new_n7674_), .A2(new_n7669_), .B(new_n7675_), .ZN(new_n7689_));
  OAI21_X1   g07433(.A1(new_n7688_), .A2(new_n7689_), .B(new_n7685_), .ZN(new_n7690_));
  NAND2_X1   g07434(.A1(new_n7690_), .A2(new_n7687_), .ZN(new_n7691_));
  OAI22_X1   g07435(.A1(new_n4208_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n4203_), .ZN(new_n7692_));
  NAND2_X1   g07436(.A1(new_n5244_), .A2(\b[15] ), .ZN(new_n7693_));
  AOI21_X1   g07437(.A1(new_n7692_), .A2(new_n7693_), .B(new_n4211_), .ZN(new_n7694_));
  NAND2_X1   g07438(.A1(new_n1047_), .A2(new_n7694_), .ZN(new_n7695_));
  XOR2_X1    g07439(.A1(new_n7695_), .A2(\a[44] ), .Z(new_n7696_));
  INV_X1     g07440(.I(new_n7696_), .ZN(new_n7697_));
  NAND3_X1   g07441(.A1(new_n7392_), .A2(new_n7400_), .A3(new_n7407_), .ZN(new_n7698_));
  NAND3_X1   g07442(.A1(new_n7400_), .A2(new_n7392_), .A3(new_n7407_), .ZN(new_n7699_));
  NAND3_X1   g07443(.A1(new_n7410_), .A2(new_n7416_), .A3(new_n7699_), .ZN(new_n7700_));
  AOI21_X1   g07444(.A1(new_n7700_), .A2(new_n7698_), .B(new_n7697_), .ZN(new_n7701_));
  NAND3_X1   g07445(.A1(new_n7700_), .A2(new_n7697_), .A3(new_n7698_), .ZN(new_n7702_));
  INV_X1     g07446(.I(new_n7702_), .ZN(new_n7703_));
  NOR2_X1    g07447(.A1(new_n7703_), .A2(new_n7701_), .ZN(new_n7704_));
  NOR2_X1    g07448(.A1(new_n7704_), .A2(new_n7691_), .ZN(new_n7705_));
  INV_X1     g07449(.I(new_n7691_), .ZN(new_n7706_));
  INV_X1     g07450(.I(new_n7701_), .ZN(new_n7707_));
  NAND2_X1   g07451(.A1(new_n7707_), .A2(new_n7702_), .ZN(new_n7708_));
  NOR2_X1    g07452(.A1(new_n7708_), .A2(new_n7706_), .ZN(new_n7709_));
  NOR2_X1    g07453(.A1(new_n7709_), .A2(new_n7705_), .ZN(new_n7710_));
  OAI22_X1   g07454(.A1(new_n3736_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n3731_), .ZN(new_n7711_));
  NAND2_X1   g07455(.A1(new_n4730_), .A2(\b[18] ), .ZN(new_n7712_));
  AOI21_X1   g07456(.A1(new_n7711_), .A2(new_n7712_), .B(new_n3739_), .ZN(new_n7713_));
  NAND2_X1   g07457(.A1(new_n1304_), .A2(new_n7713_), .ZN(new_n7714_));
  XOR2_X1    g07458(.A1(new_n7714_), .A2(\a[41] ), .Z(new_n7715_));
  INV_X1     g07459(.I(new_n7715_), .ZN(new_n7716_));
  NAND2_X1   g07460(.A1(new_n7710_), .A2(new_n7716_), .ZN(new_n7717_));
  NAND2_X1   g07461(.A1(new_n7708_), .A2(new_n7706_), .ZN(new_n7718_));
  NAND2_X1   g07462(.A1(new_n7704_), .A2(new_n7691_), .ZN(new_n7719_));
  NAND2_X1   g07463(.A1(new_n7718_), .A2(new_n7719_), .ZN(new_n7720_));
  NAND2_X1   g07464(.A1(new_n7720_), .A2(new_n7715_), .ZN(new_n7721_));
  NAND2_X1   g07465(.A1(new_n7717_), .A2(new_n7721_), .ZN(new_n7722_));
  OAI22_X1   g07466(.A1(new_n3298_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n3293_), .ZN(new_n7723_));
  NAND2_X1   g07467(.A1(new_n4227_), .A2(\b[21] ), .ZN(new_n7724_));
  AOI21_X1   g07468(.A1(new_n7723_), .A2(new_n7724_), .B(new_n3301_), .ZN(new_n7725_));
  NAND2_X1   g07469(.A1(new_n1604_), .A2(new_n7725_), .ZN(new_n7726_));
  XOR2_X1    g07470(.A1(new_n7726_), .A2(\a[38] ), .Z(new_n7727_));
  XOR2_X1    g07471(.A1(new_n7722_), .A2(new_n7727_), .Z(new_n7728_));
  NOR2_X1    g07472(.A1(new_n7158_), .A2(new_n7156_), .ZN(new_n7729_));
  OAI21_X1   g07473(.A1(new_n7729_), .A2(new_n7157_), .B(new_n7440_), .ZN(new_n7730_));
  OAI22_X1   g07474(.A1(new_n7440_), .A2(new_n7446_), .B1(new_n7434_), .B2(new_n7430_), .ZN(new_n7731_));
  OAI22_X1   g07475(.A1(new_n2846_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n2841_), .ZN(new_n7732_));
  NAND2_X1   g07476(.A1(new_n3755_), .A2(\b[24] ), .ZN(new_n7733_));
  AOI21_X1   g07477(.A1(new_n7732_), .A2(new_n7733_), .B(new_n2849_), .ZN(new_n7734_));
  NAND2_X1   g07478(.A1(new_n1926_), .A2(new_n7734_), .ZN(new_n7735_));
  XOR2_X1    g07479(.A1(new_n7735_), .A2(\a[35] ), .Z(new_n7736_));
  INV_X1     g07480(.I(new_n7736_), .ZN(new_n7737_));
  NAND3_X1   g07481(.A1(new_n7731_), .A2(new_n7730_), .A3(new_n7737_), .ZN(new_n7738_));
  NAND2_X1   g07482(.A1(new_n7138_), .A2(new_n7011_), .ZN(new_n7739_));
  AOI21_X1   g07483(.A1(new_n7739_), .A2(new_n7135_), .B(new_n7439_), .ZN(new_n7740_));
  AOI22_X1   g07484(.A1(new_n7454_), .A2(new_n7439_), .B1(new_n7442_), .B2(new_n7443_), .ZN(new_n7741_));
  OAI21_X1   g07485(.A1(new_n7741_), .A2(new_n7740_), .B(new_n7736_), .ZN(new_n7742_));
  AOI21_X1   g07486(.A1(new_n7742_), .A2(new_n7738_), .B(new_n7728_), .ZN(new_n7743_));
  INV_X1     g07487(.I(new_n7727_), .ZN(new_n7744_));
  XOR2_X1    g07488(.A1(new_n7722_), .A2(new_n7744_), .Z(new_n7745_));
  OAI21_X1   g07489(.A1(new_n7741_), .A2(new_n7740_), .B(new_n7737_), .ZN(new_n7746_));
  NAND3_X1   g07490(.A1(new_n7731_), .A2(new_n7730_), .A3(new_n7736_), .ZN(new_n7747_));
  AOI21_X1   g07491(.A1(new_n7746_), .A2(new_n7747_), .B(new_n7745_), .ZN(new_n7748_));
  AOI21_X1   g07492(.A1(new_n7441_), .A2(new_n7444_), .B(new_n7446_), .ZN(new_n7749_));
  AOI21_X1   g07493(.A1(new_n7442_), .A2(new_n7443_), .B(new_n7439_), .ZN(new_n7750_));
  NOR3_X1    g07494(.A1(new_n7434_), .A2(new_n7430_), .A3(new_n7440_), .ZN(new_n7751_));
  NOR3_X1    g07495(.A1(new_n7751_), .A2(new_n7750_), .A3(new_n7454_), .ZN(new_n7752_));
  OAI21_X1   g07496(.A1(new_n7752_), .A2(new_n7749_), .B(new_n7451_), .ZN(new_n7753_));
  NOR3_X1    g07497(.A1(new_n7743_), .A2(new_n7748_), .A3(new_n7753_), .ZN(new_n7754_));
  NOR3_X1    g07498(.A1(new_n7741_), .A2(new_n7740_), .A3(new_n7736_), .ZN(new_n7755_));
  AOI21_X1   g07499(.A1(new_n7731_), .A2(new_n7730_), .B(new_n7737_), .ZN(new_n7756_));
  OAI21_X1   g07500(.A1(new_n7755_), .A2(new_n7756_), .B(new_n7745_), .ZN(new_n7757_));
  AOI21_X1   g07501(.A1(new_n7731_), .A2(new_n7730_), .B(new_n7736_), .ZN(new_n7758_));
  NOR3_X1    g07502(.A1(new_n7741_), .A2(new_n7740_), .A3(new_n7737_), .ZN(new_n7759_));
  OAI21_X1   g07503(.A1(new_n7759_), .A2(new_n7758_), .B(new_n7728_), .ZN(new_n7760_));
  OAI21_X1   g07504(.A1(new_n7751_), .A2(new_n7750_), .B(new_n7454_), .ZN(new_n7761_));
  NAND3_X1   g07505(.A1(new_n7441_), .A2(new_n7444_), .A3(new_n7446_), .ZN(new_n7762_));
  AOI21_X1   g07506(.A1(new_n7761_), .A2(new_n7762_), .B(new_n7452_), .ZN(new_n7763_));
  AOI21_X1   g07507(.A1(new_n7757_), .A2(new_n7760_), .B(new_n7763_), .ZN(new_n7764_));
  OAI21_X1   g07508(.A1(new_n7764_), .A2(new_n7754_), .B(new_n7598_), .ZN(new_n7765_));
  NAND3_X1   g07509(.A1(new_n7757_), .A2(new_n7760_), .A3(new_n7763_), .ZN(new_n7766_));
  OAI21_X1   g07510(.A1(new_n7743_), .A2(new_n7748_), .B(new_n7753_), .ZN(new_n7767_));
  NAND3_X1   g07511(.A1(new_n7767_), .A2(new_n7766_), .A3(new_n7466_), .ZN(new_n7768_));
  AOI21_X1   g07512(.A1(new_n7765_), .A2(new_n7768_), .B(new_n7597_), .ZN(new_n7769_));
  AOI21_X1   g07513(.A1(new_n7767_), .A2(new_n7766_), .B(new_n7466_), .ZN(new_n7770_));
  NOR3_X1    g07514(.A1(new_n7764_), .A2(new_n7754_), .A3(new_n7598_), .ZN(new_n7771_));
  NOR3_X1    g07515(.A1(new_n7770_), .A2(new_n7771_), .A3(new_n7596_), .ZN(new_n7772_));
  OAI21_X1   g07516(.A1(new_n7772_), .A2(new_n7769_), .B(new_n7591_), .ZN(new_n7773_));
  INV_X1     g07517(.I(new_n7591_), .ZN(new_n7774_));
  OAI21_X1   g07518(.A1(new_n7770_), .A2(new_n7771_), .B(new_n7596_), .ZN(new_n7775_));
  NAND3_X1   g07519(.A1(new_n7765_), .A2(new_n7768_), .A3(new_n7597_), .ZN(new_n7776_));
  NAND3_X1   g07520(.A1(new_n7775_), .A2(new_n7776_), .A3(new_n7774_), .ZN(new_n7777_));
  AOI21_X1   g07521(.A1(new_n7773_), .A2(new_n7777_), .B(new_n7586_), .ZN(new_n7778_));
  AOI21_X1   g07522(.A1(new_n7775_), .A2(new_n7776_), .B(new_n7774_), .ZN(new_n7779_));
  NOR3_X1    g07523(.A1(new_n7772_), .A2(new_n7769_), .A3(new_n7591_), .ZN(new_n7780_));
  NOR3_X1    g07524(.A1(new_n7780_), .A2(new_n7779_), .A3(new_n7585_), .ZN(new_n7781_));
  OAI22_X1   g07525(.A1(new_n1760_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n1755_), .ZN(new_n7782_));
  NAND2_X1   g07526(.A1(new_n2470_), .A2(\b[33] ), .ZN(new_n7783_));
  AOI21_X1   g07527(.A1(new_n7782_), .A2(new_n7783_), .B(new_n1763_), .ZN(new_n7784_));
  NAND2_X1   g07528(.A1(new_n3101_), .A2(new_n7784_), .ZN(new_n7785_));
  XOR2_X1    g07529(.A1(new_n7785_), .A2(\a[26] ), .Z(new_n7786_));
  NOR3_X1    g07530(.A1(new_n7781_), .A2(new_n7778_), .A3(new_n7786_), .ZN(new_n7787_));
  OAI21_X1   g07531(.A1(new_n7780_), .A2(new_n7779_), .B(new_n7585_), .ZN(new_n7788_));
  NAND3_X1   g07532(.A1(new_n7773_), .A2(new_n7777_), .A3(new_n7586_), .ZN(new_n7789_));
  INV_X1     g07533(.I(new_n7786_), .ZN(new_n7790_));
  AOI21_X1   g07534(.A1(new_n7788_), .A2(new_n7789_), .B(new_n7790_), .ZN(new_n7791_));
  NOR2_X1    g07535(.A1(new_n7481_), .A2(new_n7486_), .ZN(new_n7792_));
  INV_X1     g07536(.I(new_n7792_), .ZN(new_n7793_));
  NOR3_X1    g07537(.A1(new_n7787_), .A2(new_n7791_), .A3(new_n7793_), .ZN(new_n7794_));
  NAND3_X1   g07538(.A1(new_n7788_), .A2(new_n7789_), .A3(new_n7790_), .ZN(new_n7795_));
  OAI21_X1   g07539(.A1(new_n7781_), .A2(new_n7778_), .B(new_n7786_), .ZN(new_n7796_));
  AOI21_X1   g07540(.A1(new_n7796_), .A2(new_n7795_), .B(new_n7792_), .ZN(new_n7797_));
  OAI22_X1   g07541(.A1(new_n1444_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n1439_), .ZN(new_n7798_));
  NAND2_X1   g07542(.A1(new_n2098_), .A2(\b[36] ), .ZN(new_n7799_));
  AOI21_X1   g07543(.A1(new_n7798_), .A2(new_n7799_), .B(new_n1447_), .ZN(new_n7800_));
  NAND2_X1   g07544(.A1(new_n3565_), .A2(new_n7800_), .ZN(new_n7801_));
  XOR2_X1    g07545(.A1(new_n7801_), .A2(\a[23] ), .Z(new_n7802_));
  NOR3_X1    g07546(.A1(new_n7794_), .A2(new_n7797_), .A3(new_n7802_), .ZN(new_n7803_));
  NAND3_X1   g07547(.A1(new_n7796_), .A2(new_n7795_), .A3(new_n7792_), .ZN(new_n7804_));
  OAI21_X1   g07548(.A1(new_n7787_), .A2(new_n7791_), .B(new_n7793_), .ZN(new_n7805_));
  INV_X1     g07549(.I(new_n7802_), .ZN(new_n7806_));
  AOI21_X1   g07550(.A1(new_n7805_), .A2(new_n7804_), .B(new_n7806_), .ZN(new_n7807_));
  OAI21_X1   g07551(.A1(new_n7497_), .A2(new_n7487_), .B(new_n7494_), .ZN(new_n7808_));
  NAND3_X1   g07552(.A1(new_n7488_), .A2(new_n7489_), .A3(new_n7495_), .ZN(new_n7809_));
  NAND2_X1   g07553(.A1(new_n7808_), .A2(new_n7809_), .ZN(new_n7810_));
  OAI21_X1   g07554(.A1(new_n7510_), .A2(new_n7810_), .B(new_n7808_), .ZN(new_n7811_));
  NOR3_X1    g07555(.A1(new_n7811_), .A2(new_n7803_), .A3(new_n7807_), .ZN(new_n7812_));
  NAND3_X1   g07556(.A1(new_n7805_), .A2(new_n7804_), .A3(new_n7806_), .ZN(new_n7813_));
  OAI21_X1   g07557(.A1(new_n7794_), .A2(new_n7797_), .B(new_n7802_), .ZN(new_n7814_));
  NOR3_X1    g07558(.A1(new_n6936_), .A2(new_n6934_), .A3(new_n6938_), .ZN(new_n7815_));
  NOR3_X1    g07559(.A1(new_n7231_), .A2(new_n7225_), .A3(new_n7237_), .ZN(new_n7816_));
  AOI21_X1   g07560(.A1(new_n7506_), .A2(new_n7507_), .B(new_n7505_), .ZN(new_n7817_));
  OAI22_X1   g07561(.A1(new_n7816_), .A2(new_n7817_), .B1(new_n7237_), .B2(new_n7815_), .ZN(new_n7818_));
  NAND2_X1   g07562(.A1(new_n7818_), .A2(new_n7499_), .ZN(new_n7819_));
  AOI22_X1   g07563(.A1(new_n7819_), .A2(new_n7808_), .B1(new_n7814_), .B2(new_n7813_), .ZN(new_n7820_));
  OAI22_X1   g07564(.A1(new_n1168_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n1163_), .ZN(new_n7821_));
  NAND2_X1   g07565(.A1(new_n1774_), .A2(\b[39] ), .ZN(new_n7822_));
  AOI21_X1   g07566(.A1(new_n7821_), .A2(new_n7822_), .B(new_n1171_), .ZN(new_n7823_));
  NAND2_X1   g07567(.A1(new_n3996_), .A2(new_n7823_), .ZN(new_n7824_));
  XOR2_X1    g07568(.A1(new_n7824_), .A2(\a[20] ), .Z(new_n7825_));
  NOR3_X1    g07569(.A1(new_n7820_), .A2(new_n7812_), .A3(new_n7825_), .ZN(new_n7826_));
  AOI21_X1   g07570(.A1(new_n7818_), .A2(new_n7499_), .B(new_n7496_), .ZN(new_n7827_));
  NAND3_X1   g07571(.A1(new_n7827_), .A2(new_n7813_), .A3(new_n7814_), .ZN(new_n7828_));
  OAI21_X1   g07572(.A1(new_n7803_), .A2(new_n7807_), .B(new_n7811_), .ZN(new_n7829_));
  INV_X1     g07573(.I(new_n7825_), .ZN(new_n7830_));
  AOI21_X1   g07574(.A1(new_n7829_), .A2(new_n7828_), .B(new_n7830_), .ZN(new_n7831_));
  OAI21_X1   g07575(.A1(new_n7831_), .A2(new_n7826_), .B(new_n7584_), .ZN(new_n7832_));
  XOR2_X1    g07576(.A1(new_n7510_), .A2(new_n7810_), .Z(new_n7833_));
  NAND2_X1   g07577(.A1(new_n7833_), .A2(new_n7504_), .ZN(new_n7834_));
  AOI21_X1   g07578(.A1(new_n7829_), .A2(new_n7828_), .B(new_n7825_), .ZN(new_n7835_));
  NOR3_X1    g07579(.A1(new_n7820_), .A2(new_n7812_), .A3(new_n7830_), .ZN(new_n7836_));
  OAI21_X1   g07580(.A1(new_n7835_), .A2(new_n7836_), .B(new_n7834_), .ZN(new_n7837_));
  OAI22_X1   g07581(.A1(new_n940_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n935_), .ZN(new_n7838_));
  NAND2_X1   g07582(.A1(new_n1458_), .A2(\b[42] ), .ZN(new_n7839_));
  AOI21_X1   g07583(.A1(new_n7838_), .A2(new_n7839_), .B(new_n943_), .ZN(new_n7840_));
  NAND2_X1   g07584(.A1(new_n4500_), .A2(new_n7840_), .ZN(new_n7841_));
  XOR2_X1    g07585(.A1(new_n7841_), .A2(\a[17] ), .Z(new_n7842_));
  AOI21_X1   g07586(.A1(new_n7832_), .A2(new_n7837_), .B(new_n7842_), .ZN(new_n7843_));
  NAND3_X1   g07587(.A1(new_n7832_), .A2(new_n7837_), .A3(new_n7842_), .ZN(new_n7844_));
  INV_X1     g07588(.I(new_n7844_), .ZN(new_n7845_));
  NOR2_X1    g07589(.A1(new_n7845_), .A2(new_n7843_), .ZN(new_n7846_));
  OAI22_X1   g07590(.A1(new_n757_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n752_), .ZN(new_n7847_));
  NAND2_X1   g07591(.A1(new_n1182_), .A2(\b[45] ), .ZN(new_n7848_));
  AOI21_X1   g07592(.A1(new_n7847_), .A2(new_n7848_), .B(new_n760_), .ZN(new_n7849_));
  NAND2_X1   g07593(.A1(new_n5004_), .A2(new_n7849_), .ZN(new_n7850_));
  XOR2_X1    g07594(.A1(new_n7850_), .A2(\a[14] ), .Z(new_n7851_));
  INV_X1     g07595(.I(new_n7851_), .ZN(new_n7852_));
  NAND2_X1   g07596(.A1(new_n7846_), .A2(new_n7852_), .ZN(new_n7853_));
  NOR2_X1    g07597(.A1(new_n7846_), .A2(new_n7852_), .ZN(new_n7854_));
  INV_X1     g07598(.I(new_n7854_), .ZN(new_n7855_));
  AOI21_X1   g07599(.A1(new_n7855_), .A2(new_n7853_), .B(new_n7581_), .ZN(new_n7856_));
  NOR2_X1    g07600(.A1(new_n7846_), .A2(new_n7851_), .ZN(new_n7857_));
  INV_X1     g07601(.I(new_n7857_), .ZN(new_n7858_));
  NAND2_X1   g07602(.A1(new_n7846_), .A2(new_n7851_), .ZN(new_n7859_));
  AOI21_X1   g07603(.A1(new_n7858_), .A2(new_n7859_), .B(new_n7580_), .ZN(new_n7860_));
  NOR3_X1    g07604(.A1(new_n7856_), .A2(new_n7860_), .A3(new_n7579_), .ZN(new_n7861_));
  INV_X1     g07605(.I(new_n7853_), .ZN(new_n7862_));
  OAI21_X1   g07606(.A1(new_n7862_), .A2(new_n7854_), .B(new_n7580_), .ZN(new_n7863_));
  INV_X1     g07607(.I(new_n7859_), .ZN(new_n7864_));
  OAI21_X1   g07608(.A1(new_n7864_), .A2(new_n7857_), .B(new_n7581_), .ZN(new_n7865_));
  AOI21_X1   g07609(.A1(new_n7863_), .A2(new_n7865_), .B(new_n7524_), .ZN(new_n7866_));
  NOR2_X1    g07610(.A1(new_n7866_), .A2(new_n7861_), .ZN(new_n7867_));
  OAI22_X1   g07611(.A1(new_n582_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n577_), .ZN(new_n7868_));
  NAND2_X1   g07612(.A1(new_n960_), .A2(\b[48] ), .ZN(new_n7869_));
  AOI21_X1   g07613(.A1(new_n7868_), .A2(new_n7869_), .B(new_n585_), .ZN(new_n7870_));
  NAND2_X1   g07614(.A1(new_n5537_), .A2(new_n7870_), .ZN(new_n7871_));
  XOR2_X1    g07615(.A1(new_n7871_), .A2(\a[11] ), .Z(new_n7872_));
  XOR2_X1    g07616(.A1(new_n7867_), .A2(new_n7872_), .Z(new_n7873_));
  NOR2_X1    g07617(.A1(new_n7873_), .A2(new_n7578_), .ZN(new_n7874_));
  NAND3_X1   g07618(.A1(new_n7863_), .A2(new_n7865_), .A3(new_n7524_), .ZN(new_n7875_));
  OAI21_X1   g07619(.A1(new_n7856_), .A2(new_n7860_), .B(new_n7579_), .ZN(new_n7876_));
  INV_X1     g07620(.I(new_n7872_), .ZN(new_n7877_));
  NAND3_X1   g07621(.A1(new_n7876_), .A2(new_n7875_), .A3(new_n7877_), .ZN(new_n7878_));
  OAI21_X1   g07622(.A1(new_n7866_), .A2(new_n7861_), .B(new_n7872_), .ZN(new_n7879_));
  AOI21_X1   g07623(.A1(new_n7879_), .A2(new_n7878_), .B(new_n7577_), .ZN(new_n7880_));
  NOR2_X1    g07624(.A1(new_n7874_), .A2(new_n7880_), .ZN(new_n7881_));
  OAI22_X1   g07625(.A1(new_n437_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n431_), .ZN(new_n7882_));
  NAND2_X1   g07626(.A1(new_n775_), .A2(\b[51] ), .ZN(new_n7883_));
  AOI21_X1   g07627(.A1(new_n7882_), .A2(new_n7883_), .B(new_n440_), .ZN(new_n7884_));
  NAND2_X1   g07628(.A1(new_n6219_), .A2(new_n7884_), .ZN(new_n7885_));
  XOR2_X1    g07629(.A1(new_n7885_), .A2(\a[8] ), .Z(new_n7886_));
  XNOR2_X1   g07630(.A1(new_n7881_), .A2(new_n7886_), .ZN(new_n7887_));
  NOR2_X1    g07631(.A1(new_n7532_), .A2(new_n7537_), .ZN(new_n7888_));
  XNOR2_X1   g07632(.A1(new_n7887_), .A2(new_n7888_), .ZN(new_n7889_));
  INV_X1     g07633(.I(\b[59] ), .ZN(new_n7890_));
  NOR2_X1    g07634(.A1(new_n7553_), .A2(new_n7305_), .ZN(new_n7891_));
  INV_X1     g07635(.I(new_n7553_), .ZN(new_n7892_));
  NOR2_X1    g07636(.A1(new_n7892_), .A2(\b[57] ), .ZN(new_n7893_));
  OAI21_X1   g07637(.A1(new_n7893_), .A2(new_n7891_), .B(new_n7555_), .ZN(new_n7894_));
  XOR2_X1    g07638(.A1(new_n7894_), .A2(new_n7890_), .Z(new_n7895_));
  OAI22_X1   g07639(.A1(new_n405_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n404_), .ZN(new_n7896_));
  NAND2_X1   g07640(.A1(new_n279_), .A2(\b[57] ), .ZN(new_n7897_));
  AOI21_X1   g07641(.A1(new_n7896_), .A2(new_n7897_), .B(new_n264_), .ZN(new_n7898_));
  NAND2_X1   g07642(.A1(new_n7895_), .A2(new_n7898_), .ZN(new_n7899_));
  XOR2_X1    g07643(.A1(new_n7899_), .A2(\a[2] ), .Z(new_n7900_));
  OAI22_X1   g07644(.A1(new_n364_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n320_), .ZN(new_n7901_));
  NAND2_X1   g07645(.A1(new_n594_), .A2(\b[54] ), .ZN(new_n7902_));
  AOI21_X1   g07646(.A1(new_n7901_), .A2(new_n7902_), .B(new_n312_), .ZN(new_n7903_));
  NAND2_X1   g07647(.A1(new_n6994_), .A2(new_n7903_), .ZN(new_n7904_));
  XOR2_X1    g07648(.A1(new_n7904_), .A2(\a[5] ), .Z(new_n7905_));
  NOR2_X1    g07649(.A1(new_n7900_), .A2(new_n7905_), .ZN(new_n7906_));
  INV_X1     g07650(.I(new_n7906_), .ZN(new_n7907_));
  NAND2_X1   g07651(.A1(new_n7900_), .A2(new_n7905_), .ZN(new_n7908_));
  NAND2_X1   g07652(.A1(new_n7907_), .A2(new_n7908_), .ZN(new_n7909_));
  NAND2_X1   g07653(.A1(new_n7889_), .A2(new_n7909_), .ZN(new_n7910_));
  XNOR2_X1   g07654(.A1(new_n7900_), .A2(new_n7905_), .ZN(new_n7911_));
  OAI21_X1   g07655(.A1(new_n7889_), .A2(new_n7911_), .B(new_n7910_), .ZN(new_n7912_));
  INV_X1     g07656(.I(new_n7538_), .ZN(new_n7913_));
  INV_X1     g07657(.I(new_n7543_), .ZN(new_n7914_));
  NAND2_X1   g07658(.A1(new_n7010_), .A2(new_n7303_), .ZN(new_n7915_));
  NAND2_X1   g07659(.A1(new_n7915_), .A2(new_n7302_), .ZN(new_n7916_));
  XOR2_X1    g07660(.A1(new_n7916_), .A2(new_n7914_), .Z(new_n7917_));
  NAND2_X1   g07661(.A1(new_n7917_), .A2(new_n7913_), .ZN(new_n7918_));
  XOR2_X1    g07662(.A1(new_n7918_), .A2(new_n7912_), .Z(new_n7919_));
  NAND2_X1   g07663(.A1(new_n7916_), .A2(new_n7914_), .ZN(new_n7920_));
  XOR2_X1    g07664(.A1(new_n7919_), .A2(new_n7920_), .Z(\f[59] ));
  OAI21_X1   g07665(.A1(new_n7305_), .A2(new_n7890_), .B(new_n7560_), .ZN(new_n7922_));
  NAND2_X1   g07666(.A1(new_n7892_), .A2(new_n7922_), .ZN(new_n7923_));
  OAI21_X1   g07667(.A1(\b[57] ), .A2(\b[59] ), .B(\b[58] ), .ZN(new_n7924_));
  NAND2_X1   g07668(.A1(new_n7923_), .A2(new_n7924_), .ZN(new_n7925_));
  XOR2_X1    g07669(.A1(\b[59] ), .A2(\b[60] ), .Z(new_n7926_));
  NAND2_X1   g07670(.A1(new_n7925_), .A2(new_n7926_), .ZN(new_n7927_));
  XOR2_X1    g07671(.A1(\b[59] ), .A2(\b[60] ), .Z(new_n7928_));
  OAI21_X1   g07672(.A1(new_n7925_), .A2(new_n7928_), .B(new_n7927_), .ZN(new_n7929_));
  INV_X1     g07673(.I(\b[60] ), .ZN(new_n7930_));
  OAI22_X1   g07674(.A1(new_n405_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n404_), .ZN(new_n7931_));
  NAND2_X1   g07675(.A1(new_n279_), .A2(\b[58] ), .ZN(new_n7932_));
  AOI21_X1   g07676(.A1(new_n7931_), .A2(new_n7932_), .B(new_n264_), .ZN(new_n7933_));
  NAND2_X1   g07677(.A1(new_n7929_), .A2(new_n7933_), .ZN(new_n7934_));
  XOR2_X1    g07678(.A1(new_n7934_), .A2(\a[2] ), .Z(new_n7935_));
  OAI22_X1   g07679(.A1(new_n364_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n320_), .ZN(new_n7936_));
  NAND2_X1   g07680(.A1(new_n594_), .A2(\b[55] ), .ZN(new_n7937_));
  AOI21_X1   g07681(.A1(new_n7936_), .A2(new_n7937_), .B(new_n312_), .ZN(new_n7938_));
  NAND2_X1   g07682(.A1(new_n7308_), .A2(new_n7938_), .ZN(new_n7939_));
  XOR2_X1    g07683(.A1(new_n7939_), .A2(\a[5] ), .Z(new_n7940_));
  AOI21_X1   g07684(.A1(new_n7889_), .A2(new_n7908_), .B(new_n7906_), .ZN(new_n7941_));
  AOI21_X1   g07685(.A1(new_n7876_), .A2(new_n7875_), .B(new_n7877_), .ZN(new_n7942_));
  OAI21_X1   g07686(.A1(new_n7578_), .A2(new_n7942_), .B(new_n7878_), .ZN(new_n7943_));
  AOI21_X1   g07687(.A1(new_n7580_), .A2(new_n7844_), .B(new_n7843_), .ZN(new_n7944_));
  INV_X1     g07688(.I(new_n7944_), .ZN(new_n7945_));
  AOI21_X1   g07689(.A1(new_n7718_), .A2(new_n7719_), .B(new_n7715_), .ZN(new_n7946_));
  NOR2_X1    g07690(.A1(new_n7417_), .A2(new_n7696_), .ZN(new_n7947_));
  INV_X1     g07691(.I(new_n7699_), .ZN(new_n7948_));
  XOR2_X1    g07692(.A1(new_n7691_), .A2(new_n7948_), .Z(new_n7949_));
  AOI21_X1   g07693(.A1(new_n7410_), .A2(new_n7416_), .B(new_n7697_), .ZN(new_n7950_));
  AOI21_X1   g07694(.A1(new_n7949_), .A2(new_n7950_), .B(new_n7947_), .ZN(new_n7951_));
  AOI21_X1   g07695(.A1(new_n7602_), .A2(new_n7640_), .B(new_n7622_), .ZN(new_n7952_));
  NAND2_X1   g07696(.A1(\a[59] ), .A2(\a[60] ), .ZN(new_n7953_));
  OR2_X2     g07697(.A1(\a[59] ), .A2(\a[60] ), .Z(new_n7954_));
  NAND2_X1   g07698(.A1(new_n7954_), .A2(new_n7953_), .ZN(new_n7955_));
  NOR2_X1    g07699(.A1(new_n7955_), .A2(new_n258_), .ZN(new_n7956_));
  INV_X1     g07700(.I(new_n7956_), .ZN(new_n7957_));
  NAND2_X1   g07701(.A1(new_n7614_), .A2(new_n7603_), .ZN(new_n7958_));
  OAI22_X1   g07702(.A1(new_n290_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n292_), .ZN(new_n7959_));
  OAI21_X1   g07703(.A1(new_n267_), .A2(new_n7611_), .B(new_n7959_), .ZN(new_n7960_));
  NAND3_X1   g07704(.A1(new_n7960_), .A2(new_n298_), .A3(new_n7604_), .ZN(new_n7961_));
  XOR2_X1    g07705(.A1(new_n7961_), .A2(\a[59] ), .Z(new_n7962_));
  XOR2_X1    g07706(.A1(new_n7958_), .A2(new_n7962_), .Z(new_n7963_));
  XOR2_X1    g07707(.A1(new_n7963_), .A2(new_n7957_), .Z(new_n7964_));
  AOI22_X1   g07708(.A1(new_n6506_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n6509_), .ZN(new_n7965_));
  NOR2_X1    g07709(.A1(new_n6729_), .A2(new_n393_), .ZN(new_n7966_));
  OAI21_X1   g07710(.A1(new_n7965_), .A2(new_n7966_), .B(new_n6512_), .ZN(new_n7967_));
  NOR2_X1    g07711(.A1(new_n524_), .A2(new_n7967_), .ZN(new_n7968_));
  XOR2_X1    g07712(.A1(new_n7968_), .A2(new_n6516_), .Z(new_n7969_));
  INV_X1     g07713(.I(new_n7969_), .ZN(new_n7970_));
  NAND2_X1   g07714(.A1(new_n7964_), .A2(new_n7970_), .ZN(new_n7971_));
  XOR2_X1    g07715(.A1(new_n7963_), .A2(new_n7956_), .Z(new_n7972_));
  NAND2_X1   g07716(.A1(new_n7972_), .A2(new_n7969_), .ZN(new_n7973_));
  AOI21_X1   g07717(.A1(new_n7971_), .A2(new_n7973_), .B(new_n7952_), .ZN(new_n7974_));
  INV_X1     g07718(.I(new_n7974_), .ZN(new_n7975_));
  XOR2_X1    g07719(.A1(new_n7972_), .A2(new_n7969_), .Z(new_n7976_));
  NAND2_X1   g07720(.A1(new_n7976_), .A2(new_n7952_), .ZN(new_n7977_));
  NAND2_X1   g07721(.A1(new_n7977_), .A2(new_n7975_), .ZN(new_n7978_));
  OAI22_X1   g07722(.A1(new_n5786_), .A2(new_n510_), .B1(new_n495_), .B2(new_n5792_), .ZN(new_n7979_));
  NAND2_X1   g07723(.A1(new_n6745_), .A2(\b[7] ), .ZN(new_n7980_));
  AOI21_X1   g07724(.A1(new_n7980_), .A2(new_n7979_), .B(new_n5796_), .ZN(new_n7981_));
  NAND2_X1   g07725(.A1(new_n518_), .A2(new_n7981_), .ZN(new_n7982_));
  XOR2_X1    g07726(.A1(new_n7982_), .A2(\a[53] ), .Z(new_n7983_));
  NAND2_X1   g07727(.A1(new_n7647_), .A2(new_n7650_), .ZN(new_n7984_));
  NOR2_X1    g07728(.A1(new_n7641_), .A2(new_n7644_), .ZN(new_n7985_));
  NAND2_X1   g07729(.A1(new_n7985_), .A2(new_n7645_), .ZN(new_n7986_));
  NAND2_X1   g07730(.A1(new_n7984_), .A2(new_n7986_), .ZN(new_n7987_));
  XOR2_X1    g07731(.A1(new_n7987_), .A2(new_n7983_), .Z(new_n7988_));
  XOR2_X1    g07732(.A1(new_n7988_), .A2(new_n7978_), .Z(new_n7989_));
  OAI22_X1   g07733(.A1(new_n5228_), .A2(new_n717_), .B1(new_n659_), .B2(new_n5225_), .ZN(new_n7990_));
  NAND2_X1   g07734(.A1(new_n5387_), .A2(\b[10] ), .ZN(new_n7991_));
  AOI21_X1   g07735(.A1(new_n7990_), .A2(new_n7991_), .B(new_n5231_), .ZN(new_n7992_));
  NAND2_X1   g07736(.A1(new_n716_), .A2(new_n7992_), .ZN(new_n7993_));
  XOR2_X1    g07737(.A1(new_n7993_), .A2(\a[50] ), .Z(new_n7994_));
  INV_X1     g07738(.I(new_n7994_), .ZN(new_n7995_));
  NAND2_X1   g07739(.A1(new_n7675_), .A2(new_n7665_), .ZN(new_n7996_));
  NAND3_X1   g07740(.A1(new_n7996_), .A2(new_n7382_), .A3(new_n7668_), .ZN(new_n7997_));
  OAI21_X1   g07741(.A1(new_n7661_), .A2(new_n7662_), .B(new_n7659_), .ZN(new_n7998_));
  AOI21_X1   g07742(.A1(new_n7997_), .A2(new_n7998_), .B(new_n7995_), .ZN(new_n7999_));
  NOR2_X1    g07743(.A1(new_n7670_), .A2(new_n7679_), .ZN(new_n8000_));
  OAI21_X1   g07744(.A1(new_n8000_), .A2(new_n7673_), .B(new_n7998_), .ZN(new_n8001_));
  NOR2_X1    g07745(.A1(new_n8001_), .A2(new_n7994_), .ZN(new_n8002_));
  OAI21_X1   g07746(.A1(new_n8002_), .A2(new_n7999_), .B(new_n7989_), .ZN(new_n8003_));
  XNOR2_X1   g07747(.A1(new_n7988_), .A2(new_n7978_), .ZN(new_n8004_));
  NAND2_X1   g07748(.A1(new_n8001_), .A2(new_n7994_), .ZN(new_n8005_));
  NAND3_X1   g07749(.A1(new_n7997_), .A2(new_n7995_), .A3(new_n7998_), .ZN(new_n8006_));
  NAND3_X1   g07750(.A1(new_n8005_), .A2(new_n8006_), .A3(new_n8004_), .ZN(new_n8007_));
  NAND2_X1   g07751(.A1(new_n8003_), .A2(new_n8007_), .ZN(new_n8008_));
  OAI22_X1   g07752(.A1(new_n4711_), .A2(new_n904_), .B1(new_n848_), .B2(new_n4706_), .ZN(new_n8009_));
  NAND2_X1   g07753(.A1(new_n5814_), .A2(\b[13] ), .ZN(new_n8010_));
  AOI21_X1   g07754(.A1(new_n8009_), .A2(new_n8010_), .B(new_n4714_), .ZN(new_n8011_));
  NAND2_X1   g07755(.A1(new_n907_), .A2(new_n8011_), .ZN(new_n8012_));
  XOR2_X1    g07756(.A1(new_n8012_), .A2(\a[47] ), .Z(new_n8013_));
  NOR3_X1    g07757(.A1(new_n7688_), .A2(new_n7689_), .A3(new_n7685_), .ZN(new_n8014_));
  OAI21_X1   g07758(.A1(new_n8014_), .A2(new_n7948_), .B(new_n7690_), .ZN(new_n8015_));
  NAND2_X1   g07759(.A1(new_n8015_), .A2(new_n8013_), .ZN(new_n8016_));
  INV_X1     g07760(.I(new_n8013_), .ZN(new_n8017_));
  NAND3_X1   g07761(.A1(new_n7690_), .A2(new_n7687_), .A3(new_n7699_), .ZN(new_n8018_));
  NAND3_X1   g07762(.A1(new_n8018_), .A2(new_n7690_), .A3(new_n8017_), .ZN(new_n8019_));
  AOI21_X1   g07763(.A1(new_n8016_), .A2(new_n8019_), .B(new_n8008_), .ZN(new_n8020_));
  AND2_X2    g07764(.A1(new_n8003_), .A2(new_n8007_), .Z(new_n8021_));
  AOI21_X1   g07765(.A1(new_n8018_), .A2(new_n7690_), .B(new_n8017_), .ZN(new_n8022_));
  NOR2_X1    g07766(.A1(new_n8015_), .A2(new_n8013_), .ZN(new_n8023_));
  NOR3_X1    g07767(.A1(new_n8023_), .A2(new_n8022_), .A3(new_n8021_), .ZN(new_n8024_));
  OAI22_X1   g07768(.A1(new_n4208_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n4203_), .ZN(new_n8025_));
  NAND2_X1   g07769(.A1(new_n5244_), .A2(\b[16] ), .ZN(new_n8026_));
  AOI21_X1   g07770(.A1(new_n8025_), .A2(new_n8026_), .B(new_n4211_), .ZN(new_n8027_));
  NAND2_X1   g07771(.A1(new_n1123_), .A2(new_n8027_), .ZN(new_n8028_));
  XOR2_X1    g07772(.A1(new_n8028_), .A2(\a[44] ), .Z(new_n8029_));
  NOR3_X1    g07773(.A1(new_n8024_), .A2(new_n8020_), .A3(new_n8029_), .ZN(new_n8030_));
  OAI21_X1   g07774(.A1(new_n8023_), .A2(new_n8022_), .B(new_n8021_), .ZN(new_n8031_));
  NAND3_X1   g07775(.A1(new_n8016_), .A2(new_n8019_), .A3(new_n8008_), .ZN(new_n8032_));
  INV_X1     g07776(.I(new_n8029_), .ZN(new_n8033_));
  AOI21_X1   g07777(.A1(new_n8031_), .A2(new_n8032_), .B(new_n8033_), .ZN(new_n8034_));
  OAI21_X1   g07778(.A1(new_n8030_), .A2(new_n8034_), .B(new_n7951_), .ZN(new_n8035_));
  NOR2_X1    g07779(.A1(new_n7691_), .A2(new_n7699_), .ZN(new_n8036_));
  AOI21_X1   g07780(.A1(new_n7690_), .A2(new_n7687_), .B(new_n7948_), .ZN(new_n8037_));
  OAI21_X1   g07781(.A1(new_n8036_), .A2(new_n8037_), .B(new_n7950_), .ZN(new_n8038_));
  OAI21_X1   g07782(.A1(new_n7417_), .A2(new_n7696_), .B(new_n8038_), .ZN(new_n8039_));
  NAND3_X1   g07783(.A1(new_n8031_), .A2(new_n8032_), .A3(new_n8033_), .ZN(new_n8040_));
  OAI21_X1   g07784(.A1(new_n8024_), .A2(new_n8020_), .B(new_n8029_), .ZN(new_n8041_));
  NAND3_X1   g07785(.A1(new_n8041_), .A2(new_n8040_), .A3(new_n8039_), .ZN(new_n8042_));
  OAI22_X1   g07786(.A1(new_n3736_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n3731_), .ZN(new_n8043_));
  NAND2_X1   g07787(.A1(new_n4730_), .A2(\b[19] ), .ZN(new_n8044_));
  AOI21_X1   g07788(.A1(new_n8043_), .A2(new_n8044_), .B(new_n3739_), .ZN(new_n8045_));
  NAND2_X1   g07789(.A1(new_n1396_), .A2(new_n8045_), .ZN(new_n8046_));
  XOR2_X1    g07790(.A1(new_n8046_), .A2(\a[41] ), .Z(new_n8047_));
  AOI21_X1   g07791(.A1(new_n8035_), .A2(new_n8042_), .B(new_n8047_), .ZN(new_n8048_));
  NAND2_X1   g07792(.A1(new_n8035_), .A2(new_n8042_), .ZN(new_n8049_));
  INV_X1     g07793(.I(new_n8047_), .ZN(new_n8050_));
  NOR2_X1    g07794(.A1(new_n8049_), .A2(new_n8050_), .ZN(new_n8051_));
  OAI21_X1   g07795(.A1(new_n8051_), .A2(new_n8048_), .B(new_n7946_), .ZN(new_n8052_));
  OAI21_X1   g07796(.A1(new_n7709_), .A2(new_n7705_), .B(new_n7716_), .ZN(new_n8053_));
  NAND3_X1   g07797(.A1(new_n8035_), .A2(new_n8042_), .A3(new_n8050_), .ZN(new_n8054_));
  AOI21_X1   g07798(.A1(new_n8041_), .A2(new_n8040_), .B(new_n8039_), .ZN(new_n8055_));
  NOR3_X1    g07799(.A1(new_n8030_), .A2(new_n8034_), .A3(new_n7951_), .ZN(new_n8056_));
  OAI21_X1   g07800(.A1(new_n8056_), .A2(new_n8055_), .B(new_n8047_), .ZN(new_n8057_));
  NAND2_X1   g07801(.A1(new_n8057_), .A2(new_n8054_), .ZN(new_n8058_));
  NAND2_X1   g07802(.A1(new_n8058_), .A2(new_n8053_), .ZN(new_n8059_));
  NAND2_X1   g07803(.A1(new_n8059_), .A2(new_n8052_), .ZN(new_n8060_));
  NOR2_X1    g07804(.A1(new_n7720_), .A2(new_n7715_), .ZN(new_n8061_));
  NOR2_X1    g07805(.A1(new_n7710_), .A2(new_n7716_), .ZN(new_n8062_));
  NOR2_X1    g07806(.A1(new_n8062_), .A2(new_n8061_), .ZN(new_n8063_));
  NOR2_X1    g07807(.A1(new_n8063_), .A2(new_n7727_), .ZN(new_n8064_));
  INV_X1     g07808(.I(new_n8064_), .ZN(new_n8065_));
  NAND2_X1   g07809(.A1(new_n8063_), .A2(new_n7727_), .ZN(new_n8066_));
  OAI21_X1   g07810(.A1(new_n7741_), .A2(new_n7740_), .B(new_n8066_), .ZN(new_n8067_));
  OAI22_X1   g07811(.A1(new_n3298_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n3293_), .ZN(new_n8068_));
  NAND2_X1   g07812(.A1(new_n4227_), .A2(\b[22] ), .ZN(new_n8069_));
  AOI21_X1   g07813(.A1(new_n8068_), .A2(new_n8069_), .B(new_n3301_), .ZN(new_n8070_));
  NAND2_X1   g07814(.A1(new_n1708_), .A2(new_n8070_), .ZN(new_n8071_));
  XOR2_X1    g07815(.A1(new_n8071_), .A2(\a[38] ), .Z(new_n8072_));
  AOI21_X1   g07816(.A1(new_n8067_), .A2(new_n8065_), .B(new_n8072_), .ZN(new_n8073_));
  NOR2_X1    g07817(.A1(new_n7722_), .A2(new_n7744_), .ZN(new_n8074_));
  AOI21_X1   g07818(.A1(new_n7731_), .A2(new_n7730_), .B(new_n8074_), .ZN(new_n8075_));
  INV_X1     g07819(.I(new_n8072_), .ZN(new_n8076_));
  NOR3_X1    g07820(.A1(new_n8075_), .A2(new_n8064_), .A3(new_n8076_), .ZN(new_n8077_));
  OAI21_X1   g07821(.A1(new_n8077_), .A2(new_n8073_), .B(new_n8060_), .ZN(new_n8078_));
  INV_X1     g07822(.I(new_n8060_), .ZN(new_n8079_));
  NOR3_X1    g07823(.A1(new_n8075_), .A2(new_n8064_), .A3(new_n8072_), .ZN(new_n8080_));
  AOI21_X1   g07824(.A1(new_n8067_), .A2(new_n8065_), .B(new_n8076_), .ZN(new_n8081_));
  OAI21_X1   g07825(.A1(new_n8080_), .A2(new_n8081_), .B(new_n8079_), .ZN(new_n8082_));
  NAND2_X1   g07826(.A1(new_n8078_), .A2(new_n8082_), .ZN(new_n8083_));
  OAI22_X1   g07827(.A1(new_n2846_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n2841_), .ZN(new_n8084_));
  NAND2_X1   g07828(.A1(new_n3755_), .A2(\b[25] ), .ZN(new_n8085_));
  AOI21_X1   g07829(.A1(new_n8084_), .A2(new_n8085_), .B(new_n2849_), .ZN(new_n8086_));
  NAND2_X1   g07830(.A1(new_n2042_), .A2(new_n8086_), .ZN(new_n8087_));
  XOR2_X1    g07831(.A1(new_n8087_), .A2(\a[35] ), .Z(new_n8088_));
  NOR3_X1    g07832(.A1(new_n7743_), .A2(new_n7748_), .A3(new_n7763_), .ZN(new_n8089_));
  NOR2_X1    g07833(.A1(new_n7434_), .A2(new_n7430_), .ZN(new_n8090_));
  NOR3_X1    g07834(.A1(new_n7729_), .A2(new_n7157_), .A3(new_n7440_), .ZN(new_n8091_));
  OAI21_X1   g07835(.A1(new_n8090_), .A2(new_n8091_), .B(new_n7730_), .ZN(new_n8092_));
  NAND2_X1   g07836(.A1(new_n7745_), .A2(new_n8092_), .ZN(new_n8093_));
  NAND2_X1   g07837(.A1(new_n7442_), .A2(new_n7443_), .ZN(new_n8094_));
  NAND3_X1   g07838(.A1(new_n7739_), .A2(new_n7135_), .A3(new_n7439_), .ZN(new_n8095_));
  AOI21_X1   g07839(.A1(new_n8094_), .A2(new_n8095_), .B(new_n7740_), .ZN(new_n8096_));
  NAND2_X1   g07840(.A1(new_n7728_), .A2(new_n8096_), .ZN(new_n8097_));
  AOI21_X1   g07841(.A1(new_n8097_), .A2(new_n8093_), .B(new_n7737_), .ZN(new_n8098_));
  OAI21_X1   g07842(.A1(new_n8089_), .A2(new_n8098_), .B(new_n8088_), .ZN(new_n8099_));
  INV_X1     g07843(.I(new_n8088_), .ZN(new_n8100_));
  NAND3_X1   g07844(.A1(new_n7757_), .A2(new_n7760_), .A3(new_n7753_), .ZN(new_n8101_));
  NOR2_X1    g07845(.A1(new_n7728_), .A2(new_n8096_), .ZN(new_n8102_));
  NOR2_X1    g07846(.A1(new_n7745_), .A2(new_n8092_), .ZN(new_n8103_));
  OAI21_X1   g07847(.A1(new_n8102_), .A2(new_n8103_), .B(new_n7736_), .ZN(new_n8104_));
  NAND3_X1   g07848(.A1(new_n8101_), .A2(new_n8100_), .A3(new_n8104_), .ZN(new_n8105_));
  AOI21_X1   g07849(.A1(new_n8099_), .A2(new_n8105_), .B(new_n8083_), .ZN(new_n8106_));
  OAI21_X1   g07850(.A1(new_n8075_), .A2(new_n8064_), .B(new_n8076_), .ZN(new_n8107_));
  NAND3_X1   g07851(.A1(new_n8067_), .A2(new_n8065_), .A3(new_n8072_), .ZN(new_n8108_));
  AOI21_X1   g07852(.A1(new_n8107_), .A2(new_n8108_), .B(new_n8079_), .ZN(new_n8109_));
  NAND3_X1   g07853(.A1(new_n8067_), .A2(new_n8065_), .A3(new_n8076_), .ZN(new_n8110_));
  OAI21_X1   g07854(.A1(new_n8075_), .A2(new_n8064_), .B(new_n8072_), .ZN(new_n8111_));
  AOI21_X1   g07855(.A1(new_n8111_), .A2(new_n8110_), .B(new_n8060_), .ZN(new_n8112_));
  NOR2_X1    g07856(.A1(new_n8109_), .A2(new_n8112_), .ZN(new_n8113_));
  AOI21_X1   g07857(.A1(new_n8101_), .A2(new_n8104_), .B(new_n8100_), .ZN(new_n8114_));
  NOR3_X1    g07858(.A1(new_n8089_), .A2(new_n8098_), .A3(new_n8088_), .ZN(new_n8115_));
  NOR3_X1    g07859(.A1(new_n8115_), .A2(new_n8114_), .A3(new_n8113_), .ZN(new_n8116_));
  NOR2_X1    g07860(.A1(new_n8106_), .A2(new_n8116_), .ZN(new_n8117_));
  OAI22_X1   g07861(.A1(new_n2452_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n2447_), .ZN(new_n8118_));
  NAND2_X1   g07862(.A1(new_n3312_), .A2(\b[28] ), .ZN(new_n8119_));
  AOI21_X1   g07863(.A1(new_n8118_), .A2(new_n8119_), .B(new_n2455_), .ZN(new_n8120_));
  NAND2_X1   g07864(.A1(new_n2404_), .A2(new_n8120_), .ZN(new_n8121_));
  XOR2_X1    g07865(.A1(new_n8121_), .A2(\a[32] ), .Z(new_n8122_));
  INV_X1     g07866(.I(new_n8122_), .ZN(new_n8123_));
  OAI21_X1   g07867(.A1(new_n7764_), .A2(new_n7754_), .B(new_n7596_), .ZN(new_n8124_));
  AOI21_X1   g07868(.A1(new_n7767_), .A2(new_n7766_), .B(new_n7596_), .ZN(new_n8125_));
  NOR3_X1    g07869(.A1(new_n7764_), .A2(new_n7754_), .A3(new_n7597_), .ZN(new_n8126_));
  OAI21_X1   g07870(.A1(new_n8125_), .A2(new_n8126_), .B(new_n7598_), .ZN(new_n8127_));
  AOI21_X1   g07871(.A1(new_n8127_), .A2(new_n8124_), .B(new_n8123_), .ZN(new_n8128_));
  INV_X1     g07872(.I(new_n8124_), .ZN(new_n8129_));
  OAI21_X1   g07873(.A1(new_n7764_), .A2(new_n7754_), .B(new_n7597_), .ZN(new_n8130_));
  NAND3_X1   g07874(.A1(new_n7767_), .A2(new_n7766_), .A3(new_n7596_), .ZN(new_n8131_));
  AOI21_X1   g07875(.A1(new_n8130_), .A2(new_n8131_), .B(new_n7466_), .ZN(new_n8132_));
  NOR3_X1    g07876(.A1(new_n8132_), .A2(new_n8122_), .A3(new_n8129_), .ZN(new_n8133_));
  OAI21_X1   g07877(.A1(new_n8128_), .A2(new_n8133_), .B(new_n8117_), .ZN(new_n8134_));
  OAI21_X1   g07878(.A1(new_n8115_), .A2(new_n8114_), .B(new_n8113_), .ZN(new_n8135_));
  NAND3_X1   g07879(.A1(new_n8099_), .A2(new_n8105_), .A3(new_n8083_), .ZN(new_n8136_));
  NAND2_X1   g07880(.A1(new_n8135_), .A2(new_n8136_), .ZN(new_n8137_));
  OAI21_X1   g07881(.A1(new_n8132_), .A2(new_n8129_), .B(new_n8122_), .ZN(new_n8138_));
  NAND3_X1   g07882(.A1(new_n8127_), .A2(new_n8123_), .A3(new_n8124_), .ZN(new_n8139_));
  NAND3_X1   g07883(.A1(new_n8139_), .A2(new_n8138_), .A3(new_n8137_), .ZN(new_n8140_));
  NAND2_X1   g07884(.A1(new_n8134_), .A2(new_n8140_), .ZN(new_n8141_));
  OAI22_X1   g07885(.A1(new_n2084_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n2079_), .ZN(new_n8142_));
  NAND2_X1   g07886(.A1(new_n2864_), .A2(\b[31] ), .ZN(new_n8143_));
  AOI21_X1   g07887(.A1(new_n8142_), .A2(new_n8143_), .B(new_n2087_), .ZN(new_n8144_));
  NAND2_X1   g07888(.A1(new_n2797_), .A2(new_n8144_), .ZN(new_n8145_));
  XOR2_X1    g07889(.A1(new_n8145_), .A2(\a[29] ), .Z(new_n8146_));
  AOI21_X1   g07890(.A1(new_n7773_), .A2(new_n7777_), .B(new_n7585_), .ZN(new_n8147_));
  NAND3_X1   g07891(.A1(new_n7767_), .A2(new_n7766_), .A3(new_n7597_), .ZN(new_n8148_));
  AOI21_X1   g07892(.A1(new_n8124_), .A2(new_n8148_), .B(new_n7466_), .ZN(new_n8149_));
  INV_X1     g07893(.I(new_n8149_), .ZN(new_n8150_));
  NAND3_X1   g07894(.A1(new_n8124_), .A2(new_n8148_), .A3(new_n7466_), .ZN(new_n8151_));
  AOI21_X1   g07895(.A1(new_n8150_), .A2(new_n8151_), .B(new_n7774_), .ZN(new_n8152_));
  OAI21_X1   g07896(.A1(new_n8147_), .A2(new_n8152_), .B(new_n8146_), .ZN(new_n8153_));
  INV_X1     g07897(.I(new_n8146_), .ZN(new_n8154_));
  OAI21_X1   g07898(.A1(new_n7780_), .A2(new_n7779_), .B(new_n7586_), .ZN(new_n8155_));
  INV_X1     g07899(.I(new_n8151_), .ZN(new_n8156_));
  OAI21_X1   g07900(.A1(new_n8156_), .A2(new_n8149_), .B(new_n7591_), .ZN(new_n8157_));
  NAND3_X1   g07901(.A1(new_n8155_), .A2(new_n8154_), .A3(new_n8157_), .ZN(new_n8158_));
  AOI21_X1   g07902(.A1(new_n8158_), .A2(new_n8153_), .B(new_n8141_), .ZN(new_n8159_));
  AOI21_X1   g07903(.A1(new_n8139_), .A2(new_n8138_), .B(new_n8137_), .ZN(new_n8160_));
  NOR3_X1    g07904(.A1(new_n8128_), .A2(new_n8133_), .A3(new_n8117_), .ZN(new_n8161_));
  NOR2_X1    g07905(.A1(new_n8160_), .A2(new_n8161_), .ZN(new_n8162_));
  AOI21_X1   g07906(.A1(new_n8155_), .A2(new_n8157_), .B(new_n8154_), .ZN(new_n8163_));
  NOR3_X1    g07907(.A1(new_n8147_), .A2(new_n8146_), .A3(new_n8152_), .ZN(new_n8164_));
  NOR3_X1    g07908(.A1(new_n8163_), .A2(new_n8164_), .A3(new_n8162_), .ZN(new_n8165_));
  NOR2_X1    g07909(.A1(new_n8165_), .A2(new_n8159_), .ZN(new_n8166_));
  OAI22_X1   g07910(.A1(new_n1760_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n1755_), .ZN(new_n8167_));
  NAND2_X1   g07911(.A1(new_n2470_), .A2(\b[34] ), .ZN(new_n8168_));
  AOI21_X1   g07912(.A1(new_n8167_), .A2(new_n8168_), .B(new_n1763_), .ZN(new_n8169_));
  NAND2_X1   g07913(.A1(new_n3246_), .A2(new_n8169_), .ZN(new_n8170_));
  XOR2_X1    g07914(.A1(new_n8170_), .A2(\a[26] ), .Z(new_n8171_));
  NAND3_X1   g07915(.A1(new_n7796_), .A2(new_n7795_), .A3(new_n7793_), .ZN(new_n8172_));
  NAND2_X1   g07916(.A1(new_n8172_), .A2(new_n8171_), .ZN(new_n8173_));
  INV_X1     g07917(.I(new_n8173_), .ZN(new_n8174_));
  NOR2_X1    g07918(.A1(new_n8172_), .A2(new_n8171_), .ZN(new_n8175_));
  OAI21_X1   g07919(.A1(new_n8174_), .A2(new_n8175_), .B(new_n8166_), .ZN(new_n8176_));
  OAI21_X1   g07920(.A1(new_n8163_), .A2(new_n8164_), .B(new_n8162_), .ZN(new_n8177_));
  NAND3_X1   g07921(.A1(new_n8158_), .A2(new_n8153_), .A3(new_n8141_), .ZN(new_n8178_));
  NAND2_X1   g07922(.A1(new_n8177_), .A2(new_n8178_), .ZN(new_n8179_));
  INV_X1     g07923(.I(new_n8175_), .ZN(new_n8180_));
  NAND3_X1   g07924(.A1(new_n8180_), .A2(new_n8179_), .A3(new_n8173_), .ZN(new_n8181_));
  NAND2_X1   g07925(.A1(new_n8176_), .A2(new_n8181_), .ZN(new_n8182_));
  OAI22_X1   g07926(.A1(new_n1444_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n1439_), .ZN(new_n8183_));
  NAND2_X1   g07927(.A1(new_n2098_), .A2(\b[37] ), .ZN(new_n8184_));
  AOI21_X1   g07928(.A1(new_n8183_), .A2(new_n8184_), .B(new_n1447_), .ZN(new_n8185_));
  NAND2_X1   g07929(.A1(new_n3700_), .A2(new_n8185_), .ZN(new_n8186_));
  NOR2_X1    g07930(.A1(new_n8186_), .A2(\a[23] ), .ZN(new_n8187_));
  INV_X1     g07931(.I(new_n8187_), .ZN(new_n8188_));
  NAND2_X1   g07932(.A1(new_n8186_), .A2(\a[23] ), .ZN(new_n8189_));
  NAND2_X1   g07933(.A1(new_n8188_), .A2(new_n8189_), .ZN(new_n8190_));
  INV_X1     g07934(.I(new_n8190_), .ZN(new_n8191_));
  NAND2_X1   g07935(.A1(new_n7814_), .A2(new_n7813_), .ZN(new_n8192_));
  OAI21_X1   g07936(.A1(new_n8192_), .A2(new_n7827_), .B(new_n8191_), .ZN(new_n8193_));
  NAND4_X1   g07937(.A1(new_n7811_), .A2(new_n7813_), .A3(new_n7814_), .A4(new_n8190_), .ZN(new_n8194_));
  AOI21_X1   g07938(.A1(new_n8193_), .A2(new_n8194_), .B(new_n8182_), .ZN(new_n8195_));
  AOI21_X1   g07939(.A1(new_n8180_), .A2(new_n8173_), .B(new_n8179_), .ZN(new_n8196_));
  NOR3_X1    g07940(.A1(new_n8174_), .A2(new_n8166_), .A3(new_n8175_), .ZN(new_n8197_));
  NOR2_X1    g07941(.A1(new_n8196_), .A2(new_n8197_), .ZN(new_n8198_));
  INV_X1     g07942(.I(new_n8193_), .ZN(new_n8199_));
  INV_X1     g07943(.I(new_n8194_), .ZN(new_n8200_));
  NOR3_X1    g07944(.A1(new_n8199_), .A2(new_n8198_), .A3(new_n8200_), .ZN(new_n8201_));
  NOR2_X1    g07945(.A1(new_n8201_), .A2(new_n8195_), .ZN(new_n8202_));
  INV_X1     g07946(.I(new_n7831_), .ZN(new_n8203_));
  OAI22_X1   g07947(.A1(new_n1168_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n1163_), .ZN(new_n8204_));
  NAND2_X1   g07948(.A1(new_n1774_), .A2(\b[40] ), .ZN(new_n8205_));
  AOI21_X1   g07949(.A1(new_n8204_), .A2(new_n8205_), .B(new_n1171_), .ZN(new_n8206_));
  NAND2_X1   g07950(.A1(new_n4017_), .A2(new_n8206_), .ZN(new_n8207_));
  XOR2_X1    g07951(.A1(new_n8207_), .A2(\a[20] ), .Z(new_n8208_));
  INV_X1     g07952(.I(new_n8208_), .ZN(new_n8209_));
  AOI21_X1   g07953(.A1(new_n7837_), .A2(new_n8203_), .B(new_n8209_), .ZN(new_n8210_));
  OAI21_X1   g07954(.A1(new_n7820_), .A2(new_n7812_), .B(new_n7830_), .ZN(new_n8211_));
  NAND3_X1   g07955(.A1(new_n7829_), .A2(new_n7828_), .A3(new_n7825_), .ZN(new_n8212_));
  AOI21_X1   g07956(.A1(new_n8212_), .A2(new_n8211_), .B(new_n7584_), .ZN(new_n8213_));
  NOR3_X1    g07957(.A1(new_n8213_), .A2(new_n7831_), .A3(new_n8208_), .ZN(new_n8214_));
  OAI21_X1   g07958(.A1(new_n8214_), .A2(new_n8210_), .B(new_n8202_), .ZN(new_n8215_));
  OAI21_X1   g07959(.A1(new_n8199_), .A2(new_n8200_), .B(new_n8198_), .ZN(new_n8216_));
  NAND3_X1   g07960(.A1(new_n8182_), .A2(new_n8193_), .A3(new_n8194_), .ZN(new_n8217_));
  NAND2_X1   g07961(.A1(new_n8216_), .A2(new_n8217_), .ZN(new_n8218_));
  OAI21_X1   g07962(.A1(new_n8213_), .A2(new_n7831_), .B(new_n8208_), .ZN(new_n8219_));
  NAND3_X1   g07963(.A1(new_n7837_), .A2(new_n8203_), .A3(new_n8209_), .ZN(new_n8220_));
  NAND3_X1   g07964(.A1(new_n8219_), .A2(new_n8220_), .A3(new_n8218_), .ZN(new_n8221_));
  OAI22_X1   g07965(.A1(new_n940_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n935_), .ZN(new_n8222_));
  NAND2_X1   g07966(.A1(new_n1458_), .A2(\b[43] ), .ZN(new_n8223_));
  AOI21_X1   g07967(.A1(new_n8222_), .A2(new_n8223_), .B(new_n943_), .ZN(new_n8224_));
  NAND2_X1   g07968(.A1(new_n4513_), .A2(new_n8224_), .ZN(new_n8225_));
  XOR2_X1    g07969(.A1(new_n8225_), .A2(\a[17] ), .Z(new_n8226_));
  AOI21_X1   g07970(.A1(new_n8215_), .A2(new_n8221_), .B(new_n8226_), .ZN(new_n8227_));
  NAND2_X1   g07971(.A1(new_n8215_), .A2(new_n8221_), .ZN(new_n8228_));
  INV_X1     g07972(.I(new_n8226_), .ZN(new_n8229_));
  NOR2_X1    g07973(.A1(new_n8228_), .A2(new_n8229_), .ZN(new_n8230_));
  OAI21_X1   g07974(.A1(new_n8230_), .A2(new_n8227_), .B(new_n7945_), .ZN(new_n8231_));
  NAND3_X1   g07975(.A1(new_n8215_), .A2(new_n8221_), .A3(new_n8229_), .ZN(new_n8232_));
  AOI21_X1   g07976(.A1(new_n8219_), .A2(new_n8220_), .B(new_n8218_), .ZN(new_n8233_));
  NOR3_X1    g07977(.A1(new_n8214_), .A2(new_n8210_), .A3(new_n8202_), .ZN(new_n8234_));
  OAI21_X1   g07978(.A1(new_n8234_), .A2(new_n8233_), .B(new_n8226_), .ZN(new_n8235_));
  NAND2_X1   g07979(.A1(new_n8235_), .A2(new_n8232_), .ZN(new_n8236_));
  NAND2_X1   g07980(.A1(new_n8236_), .A2(new_n7944_), .ZN(new_n8237_));
  NAND2_X1   g07981(.A1(new_n8237_), .A2(new_n8231_), .ZN(new_n8238_));
  OAI22_X1   g07982(.A1(new_n757_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n752_), .ZN(new_n8239_));
  NAND2_X1   g07983(.A1(new_n1182_), .A2(\b[46] ), .ZN(new_n8240_));
  AOI21_X1   g07984(.A1(new_n8239_), .A2(new_n8240_), .B(new_n760_), .ZN(new_n8241_));
  NAND2_X1   g07985(.A1(new_n5177_), .A2(new_n8241_), .ZN(new_n8242_));
  XOR2_X1    g07986(.A1(new_n8242_), .A2(\a[14] ), .Z(new_n8243_));
  OAI21_X1   g07987(.A1(new_n7845_), .A2(new_n7843_), .B(new_n7581_), .ZN(new_n8244_));
  INV_X1     g07988(.I(new_n7843_), .ZN(new_n8245_));
  NAND3_X1   g07989(.A1(new_n8245_), .A2(new_n7844_), .A3(new_n7580_), .ZN(new_n8246_));
  AOI21_X1   g07990(.A1(new_n8246_), .A2(new_n8244_), .B(new_n7852_), .ZN(new_n8247_));
  XOR2_X1    g07991(.A1(new_n8247_), .A2(new_n8243_), .Z(new_n8248_));
  XOR2_X1    g07992(.A1(new_n8248_), .A2(new_n8238_), .Z(new_n8249_));
  OAI22_X1   g07993(.A1(new_n582_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n577_), .ZN(new_n8250_));
  NAND2_X1   g07994(.A1(new_n960_), .A2(\b[49] ), .ZN(new_n8251_));
  AOI21_X1   g07995(.A1(new_n8250_), .A2(new_n8251_), .B(new_n585_), .ZN(new_n8252_));
  NAND2_X1   g07996(.A1(new_n5741_), .A2(new_n8252_), .ZN(new_n8253_));
  XOR2_X1    g07997(.A1(new_n8253_), .A2(\a[11] ), .Z(new_n8254_));
  XOR2_X1    g07998(.A1(new_n8249_), .A2(new_n8254_), .Z(new_n8255_));
  INV_X1     g07999(.I(new_n8255_), .ZN(new_n8256_));
  INV_X1     g08000(.I(new_n8254_), .ZN(new_n8257_));
  NAND2_X1   g08001(.A1(new_n8249_), .A2(new_n8257_), .ZN(new_n8258_));
  XNOR2_X1   g08002(.A1(new_n8248_), .A2(new_n8238_), .ZN(new_n8259_));
  NAND2_X1   g08003(.A1(new_n8259_), .A2(new_n8254_), .ZN(new_n8260_));
  AOI21_X1   g08004(.A1(new_n8260_), .A2(new_n8258_), .B(new_n7943_), .ZN(new_n8261_));
  AOI21_X1   g08005(.A1(new_n8256_), .A2(new_n7943_), .B(new_n8261_), .ZN(new_n8262_));
  INV_X1     g08006(.I(new_n8262_), .ZN(new_n8263_));
  OAI22_X1   g08007(.A1(new_n437_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n431_), .ZN(new_n8264_));
  NAND2_X1   g08008(.A1(new_n775_), .A2(\b[52] ), .ZN(new_n8265_));
  AOI21_X1   g08009(.A1(new_n8264_), .A2(new_n8265_), .B(new_n440_), .ZN(new_n8266_));
  NAND2_X1   g08010(.A1(new_n6237_), .A2(new_n8266_), .ZN(new_n8267_));
  XOR2_X1    g08011(.A1(new_n8267_), .A2(\a[8] ), .Z(new_n8268_));
  INV_X1     g08012(.I(new_n7881_), .ZN(new_n8269_));
  AOI22_X1   g08013(.A1(new_n8269_), .A2(new_n7886_), .B1(new_n7532_), .B2(new_n7537_), .ZN(new_n8270_));
  NAND2_X1   g08014(.A1(new_n8270_), .A2(new_n7887_), .ZN(new_n8271_));
  XOR2_X1    g08015(.A1(new_n8271_), .A2(new_n8268_), .Z(new_n8272_));
  NOR2_X1    g08016(.A1(new_n8272_), .A2(new_n8263_), .ZN(new_n8273_));
  NAND2_X1   g08017(.A1(new_n8272_), .A2(new_n8263_), .ZN(new_n8274_));
  INV_X1     g08018(.I(new_n8274_), .ZN(new_n8275_));
  NOR2_X1    g08019(.A1(new_n8275_), .A2(new_n8273_), .ZN(new_n8276_));
  XOR2_X1    g08020(.A1(new_n8276_), .A2(new_n7941_), .Z(new_n8277_));
  XOR2_X1    g08021(.A1(new_n8277_), .A2(new_n7940_), .Z(new_n8278_));
  XOR2_X1    g08022(.A1(new_n8278_), .A2(new_n7935_), .Z(new_n8279_));
  AOI21_X1   g08023(.A1(new_n7538_), .A2(new_n7543_), .B(new_n7912_), .ZN(new_n8281_));
  NAND2_X1   g08024(.A1(\f[59] ), .A2(new_n8281_), .ZN(new_n8282_));
  OR2_X2     g08025(.A1(new_n8282_), .A2(new_n8279_), .Z(new_n8283_));
  NAND2_X1   g08026(.A1(new_n8282_), .A2(new_n8279_), .ZN(new_n8284_));
  NAND2_X1   g08027(.A1(new_n8283_), .A2(new_n8284_), .ZN(\f[60] ));
  OAI21_X1   g08028(.A1(new_n8249_), .A2(new_n8257_), .B(new_n7943_), .ZN(new_n8286_));
  NAND2_X1   g08029(.A1(new_n8286_), .A2(new_n8258_), .ZN(new_n8287_));
  INV_X1     g08030(.I(new_n8232_), .ZN(new_n8288_));
  AOI21_X1   g08031(.A1(new_n8228_), .A2(new_n8226_), .B(new_n7944_), .ZN(new_n8289_));
  NOR2_X1    g08032(.A1(new_n8289_), .A2(new_n8288_), .ZN(new_n8290_));
  INV_X1     g08033(.I(new_n7986_), .ZN(new_n8291_));
  INV_X1     g08034(.I(new_n7983_), .ZN(new_n8292_));
  NAND3_X1   g08035(.A1(new_n7977_), .A2(new_n7975_), .A3(new_n8292_), .ZN(new_n8293_));
  INV_X1     g08036(.I(new_n7952_), .ZN(new_n8294_));
  XOR2_X1    g08037(.A1(new_n7964_), .A2(new_n7969_), .Z(new_n8295_));
  NOR2_X1    g08038(.A1(new_n8295_), .A2(new_n8294_), .ZN(new_n8296_));
  OAI21_X1   g08039(.A1(new_n8296_), .A2(new_n7974_), .B(new_n7983_), .ZN(new_n8297_));
  AOI21_X1   g08040(.A1(new_n8297_), .A2(new_n8293_), .B(new_n8291_), .ZN(new_n8298_));
  AOI22_X1   g08041(.A1(new_n8298_), .A2(new_n7984_), .B1(new_n7978_), .B2(new_n7983_), .ZN(new_n8299_));
  NAND2_X1   g08042(.A1(new_n7973_), .A2(new_n8294_), .ZN(new_n8300_));
  INV_X1     g08043(.I(new_n7603_), .ZN(new_n8301_));
  NOR2_X1    g08044(.A1(new_n7623_), .A2(new_n8301_), .ZN(new_n8302_));
  OAI21_X1   g08045(.A1(new_n8302_), .A2(new_n7962_), .B(new_n7957_), .ZN(new_n8303_));
  INV_X1     g08046(.I(new_n8303_), .ZN(new_n8304_));
  OAI22_X1   g08047(.A1(new_n393_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n290_), .ZN(new_n8305_));
  OAI21_X1   g08048(.A1(new_n292_), .A2(new_n7611_), .B(new_n8305_), .ZN(new_n8306_));
  NAND3_X1   g08049(.A1(new_n8306_), .A2(new_n334_), .A3(new_n7604_), .ZN(new_n8307_));
  XOR2_X1    g08050(.A1(new_n8307_), .A2(\a[59] ), .Z(new_n8308_));
  INV_X1     g08051(.I(\a[62] ), .ZN(new_n8309_));
  XOR2_X1    g08052(.A1(\a[59] ), .A2(\a[60] ), .Z(new_n8310_));
  XNOR2_X1   g08053(.A1(\a[61] ), .A2(\a[62] ), .ZN(new_n8311_));
  NAND2_X1   g08054(.A1(new_n8311_), .A2(new_n8310_), .ZN(new_n8312_));
  NOR2_X1    g08055(.A1(new_n8312_), .A2(new_n267_), .ZN(new_n8313_));
  INV_X1     g08056(.I(\a[61] ), .ZN(new_n8314_));
  NOR2_X1    g08057(.A1(new_n7954_), .A2(new_n8314_), .ZN(new_n8315_));
  NOR2_X1    g08058(.A1(new_n7953_), .A2(\a[61] ), .ZN(new_n8316_));
  NOR2_X1    g08059(.A1(new_n8315_), .A2(new_n8316_), .ZN(new_n8317_));
  NOR2_X1    g08060(.A1(new_n8317_), .A2(new_n258_), .ZN(new_n8318_));
  XNOR2_X1   g08061(.A1(\a[61] ), .A2(\a[62] ), .ZN(new_n8319_));
  NOR2_X1    g08062(.A1(new_n7955_), .A2(new_n8319_), .ZN(new_n8320_));
  INV_X1     g08063(.I(new_n8320_), .ZN(new_n8321_));
  NOR4_X1    g08064(.A1(new_n8318_), .A2(new_n8313_), .A3(new_n8321_), .A4(new_n261_), .ZN(new_n8322_));
  XOR2_X1    g08065(.A1(new_n8322_), .A2(new_n8309_), .Z(new_n8323_));
  NOR2_X1    g08066(.A1(new_n7957_), .A2(\a[62] ), .ZN(new_n8324_));
  XOR2_X1    g08067(.A1(new_n8323_), .A2(new_n8324_), .Z(new_n8325_));
  XOR2_X1    g08068(.A1(new_n8325_), .A2(new_n8308_), .Z(new_n8326_));
  NOR2_X1    g08069(.A1(new_n8326_), .A2(new_n8304_), .ZN(new_n8327_));
  XNOR2_X1   g08070(.A1(new_n8323_), .A2(new_n8324_), .ZN(new_n8328_));
  NAND2_X1   g08071(.A1(new_n8328_), .A2(new_n8308_), .ZN(new_n8329_));
  NOR2_X1    g08072(.A1(new_n8328_), .A2(new_n8308_), .ZN(new_n8330_));
  INV_X1     g08073(.I(new_n8330_), .ZN(new_n8331_));
  AOI21_X1   g08074(.A1(new_n8331_), .A2(new_n8329_), .B(new_n8303_), .ZN(new_n8332_));
  NOR2_X1    g08075(.A1(new_n8327_), .A2(new_n8332_), .ZN(new_n8333_));
  OAI22_X1   g08076(.A1(new_n6721_), .A2(new_n403_), .B1(new_n6723_), .B2(new_n450_), .ZN(new_n8334_));
  NAND2_X1   g08077(.A1(new_n7617_), .A2(\b[5] ), .ZN(new_n8335_));
  AOI21_X1   g08078(.A1(new_n8335_), .A2(new_n8334_), .B(new_n6731_), .ZN(new_n8336_));
  NAND2_X1   g08079(.A1(new_n454_), .A2(new_n8336_), .ZN(new_n8337_));
  XOR2_X1    g08080(.A1(new_n8337_), .A2(\a[56] ), .Z(new_n8338_));
  XOR2_X1    g08081(.A1(new_n8333_), .A2(new_n8338_), .Z(new_n8339_));
  AOI21_X1   g08082(.A1(new_n7971_), .A2(new_n8300_), .B(new_n8339_), .ZN(new_n8340_));
  NOR2_X1    g08083(.A1(new_n7964_), .A2(new_n7970_), .ZN(new_n8341_));
  OAI21_X1   g08084(.A1(new_n7952_), .A2(new_n8341_), .B(new_n7971_), .ZN(new_n8342_));
  INV_X1     g08085(.I(new_n8333_), .ZN(new_n8343_));
  NOR2_X1    g08086(.A1(new_n8343_), .A2(new_n8338_), .ZN(new_n8344_));
  INV_X1     g08087(.I(new_n8344_), .ZN(new_n8345_));
  NAND2_X1   g08088(.A1(new_n8343_), .A2(new_n8338_), .ZN(new_n8346_));
  AOI21_X1   g08089(.A1(new_n8345_), .A2(new_n8346_), .B(new_n8342_), .ZN(new_n8347_));
  NOR2_X1    g08090(.A1(new_n8347_), .A2(new_n8340_), .ZN(new_n8348_));
  OAI22_X1   g08091(.A1(new_n5786_), .A2(new_n617_), .B1(new_n510_), .B2(new_n5792_), .ZN(new_n8349_));
  NAND2_X1   g08092(.A1(new_n6745_), .A2(\b[8] ), .ZN(new_n8350_));
  AOI21_X1   g08093(.A1(new_n8350_), .A2(new_n8349_), .B(new_n5796_), .ZN(new_n8351_));
  NAND2_X1   g08094(.A1(new_n616_), .A2(new_n8351_), .ZN(new_n8352_));
  XOR2_X1    g08095(.A1(new_n8352_), .A2(\a[53] ), .Z(new_n8353_));
  XOR2_X1    g08096(.A1(new_n8348_), .A2(new_n8353_), .Z(new_n8354_));
  NOR2_X1    g08097(.A1(new_n8299_), .A2(new_n8354_), .ZN(new_n8355_));
  INV_X1     g08098(.I(new_n7984_), .ZN(new_n8356_));
  NAND2_X1   g08099(.A1(new_n7978_), .A2(new_n7983_), .ZN(new_n8357_));
  NOR3_X1    g08100(.A1(new_n8296_), .A2(new_n7974_), .A3(new_n7983_), .ZN(new_n8358_));
  AOI21_X1   g08101(.A1(new_n7977_), .A2(new_n7975_), .B(new_n8292_), .ZN(new_n8359_));
  OAI21_X1   g08102(.A1(new_n8358_), .A2(new_n8359_), .B(new_n7986_), .ZN(new_n8360_));
  OAI21_X1   g08103(.A1(new_n8360_), .A2(new_n8356_), .B(new_n8357_), .ZN(new_n8361_));
  INV_X1     g08104(.I(new_n8353_), .ZN(new_n8362_));
  NAND2_X1   g08105(.A1(new_n8348_), .A2(new_n8362_), .ZN(new_n8363_));
  INV_X1     g08106(.I(new_n8363_), .ZN(new_n8364_));
  NOR2_X1    g08107(.A1(new_n8348_), .A2(new_n8362_), .ZN(new_n8365_));
  NOR2_X1    g08108(.A1(new_n8364_), .A2(new_n8365_), .ZN(new_n8366_));
  NOR2_X1    g08109(.A1(new_n8366_), .A2(new_n8361_), .ZN(new_n8367_));
  NOR2_X1    g08110(.A1(new_n8367_), .A2(new_n8355_), .ZN(new_n8368_));
  OAI22_X1   g08111(.A1(new_n5228_), .A2(new_n795_), .B1(new_n717_), .B2(new_n5225_), .ZN(new_n8369_));
  NAND2_X1   g08112(.A1(new_n5387_), .A2(\b[11] ), .ZN(new_n8370_));
  AOI21_X1   g08113(.A1(new_n8369_), .A2(new_n8370_), .B(new_n5231_), .ZN(new_n8371_));
  NAND2_X1   g08114(.A1(new_n799_), .A2(new_n8371_), .ZN(new_n8372_));
  XOR2_X1    g08115(.A1(new_n8372_), .A2(\a[50] ), .Z(new_n8373_));
  INV_X1     g08116(.I(new_n8373_), .ZN(new_n8374_));
  XOR2_X1    g08117(.A1(new_n8368_), .A2(new_n8374_), .Z(new_n8375_));
  OAI22_X1   g08118(.A1(new_n4711_), .A2(new_n992_), .B1(new_n904_), .B2(new_n4706_), .ZN(new_n8376_));
  NAND2_X1   g08119(.A1(new_n5814_), .A2(\b[14] ), .ZN(new_n8377_));
  AOI21_X1   g08120(.A1(new_n8376_), .A2(new_n8377_), .B(new_n4714_), .ZN(new_n8378_));
  NAND2_X1   g08121(.A1(new_n991_), .A2(new_n8378_), .ZN(new_n8379_));
  XOR2_X1    g08122(.A1(new_n8379_), .A2(\a[47] ), .Z(new_n8380_));
  INV_X1     g08123(.I(new_n8380_), .ZN(new_n8381_));
  NAND2_X1   g08124(.A1(new_n8375_), .A2(new_n8381_), .ZN(new_n8382_));
  XOR2_X1    g08125(.A1(new_n8368_), .A2(new_n8373_), .Z(new_n8383_));
  NAND2_X1   g08126(.A1(new_n8383_), .A2(new_n8380_), .ZN(new_n8384_));
  NAND2_X1   g08127(.A1(new_n8382_), .A2(new_n8384_), .ZN(new_n8385_));
  INV_X1     g08128(.I(new_n8385_), .ZN(new_n8386_));
  OAI22_X1   g08129(.A1(new_n4208_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n4203_), .ZN(new_n8387_));
  NAND2_X1   g08130(.A1(new_n5244_), .A2(\b[17] ), .ZN(new_n8388_));
  AOI21_X1   g08131(.A1(new_n8387_), .A2(new_n8388_), .B(new_n4211_), .ZN(new_n8389_));
  NAND2_X1   g08132(.A1(new_n1225_), .A2(new_n8389_), .ZN(new_n8390_));
  XOR2_X1    g08133(.A1(new_n8390_), .A2(\a[44] ), .Z(new_n8391_));
  INV_X1     g08134(.I(new_n8391_), .ZN(new_n8392_));
  NAND3_X1   g08135(.A1(new_n8041_), .A2(new_n8040_), .A3(new_n7951_), .ZN(new_n8393_));
  AOI21_X1   g08136(.A1(new_n8393_), .A2(new_n8041_), .B(new_n8392_), .ZN(new_n8394_));
  OAI21_X1   g08137(.A1(new_n8039_), .A2(new_n8030_), .B(new_n8041_), .ZN(new_n8395_));
  NOR2_X1    g08138(.A1(new_n8395_), .A2(new_n8391_), .ZN(new_n8396_));
  OAI21_X1   g08139(.A1(new_n8396_), .A2(new_n8394_), .B(new_n8386_), .ZN(new_n8397_));
  NAND2_X1   g08140(.A1(new_n8395_), .A2(new_n8391_), .ZN(new_n8398_));
  NAND3_X1   g08141(.A1(new_n8393_), .A2(new_n8041_), .A3(new_n8392_), .ZN(new_n8399_));
  NAND3_X1   g08142(.A1(new_n8398_), .A2(new_n8399_), .A3(new_n8385_), .ZN(new_n8400_));
  OAI22_X1   g08143(.A1(new_n3736_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n3731_), .ZN(new_n8401_));
  NAND2_X1   g08144(.A1(new_n4730_), .A2(\b[20] ), .ZN(new_n8402_));
  AOI21_X1   g08145(.A1(new_n8401_), .A2(new_n8402_), .B(new_n3739_), .ZN(new_n8403_));
  NAND2_X1   g08146(.A1(new_n1517_), .A2(new_n8403_), .ZN(new_n8404_));
  XOR2_X1    g08147(.A1(new_n8404_), .A2(\a[41] ), .Z(new_n8405_));
  AOI21_X1   g08148(.A1(new_n8397_), .A2(new_n8400_), .B(new_n8405_), .ZN(new_n8406_));
  AOI21_X1   g08149(.A1(new_n8398_), .A2(new_n8399_), .B(new_n8385_), .ZN(new_n8407_));
  NOR3_X1    g08150(.A1(new_n8396_), .A2(new_n8394_), .A3(new_n8386_), .ZN(new_n8408_));
  INV_X1     g08151(.I(new_n8405_), .ZN(new_n8409_));
  NOR3_X1    g08152(.A1(new_n8408_), .A2(new_n8407_), .A3(new_n8409_), .ZN(new_n8410_));
  NOR2_X1    g08153(.A1(new_n8410_), .A2(new_n8406_), .ZN(new_n8411_));
  OAI21_X1   g08154(.A1(new_n8408_), .A2(new_n8407_), .B(new_n8409_), .ZN(new_n8412_));
  NAND3_X1   g08155(.A1(new_n8397_), .A2(new_n8400_), .A3(new_n8405_), .ZN(new_n8413_));
  INV_X1     g08156(.I(new_n8054_), .ZN(new_n8414_));
  AOI21_X1   g08157(.A1(new_n8049_), .A2(new_n8047_), .B(new_n8053_), .ZN(new_n8415_));
  OAI22_X1   g08158(.A1(new_n3298_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n3293_), .ZN(new_n8416_));
  NAND2_X1   g08159(.A1(new_n4227_), .A2(\b[23] ), .ZN(new_n8417_));
  AOI21_X1   g08160(.A1(new_n8416_), .A2(new_n8417_), .B(new_n3301_), .ZN(new_n8418_));
  NAND2_X1   g08161(.A1(new_n1828_), .A2(new_n8418_), .ZN(new_n8419_));
  XOR2_X1    g08162(.A1(new_n8419_), .A2(\a[38] ), .Z(new_n8420_));
  INV_X1     g08163(.I(new_n8420_), .ZN(new_n8421_));
  OAI21_X1   g08164(.A1(new_n8415_), .A2(new_n8414_), .B(new_n8421_), .ZN(new_n8422_));
  NAND2_X1   g08165(.A1(new_n8057_), .A2(new_n7946_), .ZN(new_n8423_));
  NAND3_X1   g08166(.A1(new_n8423_), .A2(new_n8054_), .A3(new_n8420_), .ZN(new_n8424_));
  AOI22_X1   g08167(.A1(new_n8412_), .A2(new_n8413_), .B1(new_n8424_), .B2(new_n8422_), .ZN(new_n8425_));
  NAND3_X1   g08168(.A1(new_n8423_), .A2(new_n8054_), .A3(new_n8421_), .ZN(new_n8426_));
  OAI21_X1   g08169(.A1(new_n8415_), .A2(new_n8414_), .B(new_n8420_), .ZN(new_n8427_));
  NAND2_X1   g08170(.A1(new_n8426_), .A2(new_n8427_), .ZN(new_n8428_));
  AOI21_X1   g08171(.A1(new_n8411_), .A2(new_n8428_), .B(new_n8425_), .ZN(new_n8429_));
  AOI21_X1   g08172(.A1(new_n8092_), .A2(new_n8066_), .B(new_n8064_), .ZN(new_n8430_));
  AOI21_X1   g08173(.A1(new_n8430_), .A2(new_n8072_), .B(new_n8060_), .ZN(new_n8431_));
  OAI22_X1   g08174(.A1(new_n2846_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n2841_), .ZN(new_n8432_));
  NAND2_X1   g08175(.A1(new_n3755_), .A2(\b[26] ), .ZN(new_n8433_));
  AOI21_X1   g08176(.A1(new_n8432_), .A2(new_n8433_), .B(new_n2849_), .ZN(new_n8434_));
  NAND2_X1   g08177(.A1(new_n2174_), .A2(new_n8434_), .ZN(new_n8435_));
  XOR2_X1    g08178(.A1(new_n8435_), .A2(\a[35] ), .Z(new_n8436_));
  INV_X1     g08179(.I(new_n8436_), .ZN(new_n8437_));
  OAI21_X1   g08180(.A1(new_n8431_), .A2(new_n8073_), .B(new_n8437_), .ZN(new_n8438_));
  OAI21_X1   g08181(.A1(new_n8096_), .A2(new_n8074_), .B(new_n8065_), .ZN(new_n8439_));
  OAI21_X1   g08182(.A1(new_n8439_), .A2(new_n8076_), .B(new_n8079_), .ZN(new_n8440_));
  NAND3_X1   g08183(.A1(new_n8440_), .A2(new_n8107_), .A3(new_n8436_), .ZN(new_n8441_));
  AOI21_X1   g08184(.A1(new_n8441_), .A2(new_n8438_), .B(new_n8429_), .ZN(new_n8442_));
  NAND2_X1   g08185(.A1(new_n8412_), .A2(new_n8413_), .ZN(new_n8443_));
  NAND2_X1   g08186(.A1(new_n8424_), .A2(new_n8422_), .ZN(new_n8444_));
  NAND2_X1   g08187(.A1(new_n8443_), .A2(new_n8444_), .ZN(new_n8445_));
  NAND2_X1   g08188(.A1(new_n8411_), .A2(new_n8428_), .ZN(new_n8446_));
  NAND2_X1   g08189(.A1(new_n8446_), .A2(new_n8445_), .ZN(new_n8447_));
  NAND3_X1   g08190(.A1(new_n8440_), .A2(new_n8107_), .A3(new_n8437_), .ZN(new_n8448_));
  OAI21_X1   g08191(.A1(new_n8431_), .A2(new_n8073_), .B(new_n8436_), .ZN(new_n8449_));
  AOI21_X1   g08192(.A1(new_n8448_), .A2(new_n8449_), .B(new_n8447_), .ZN(new_n8450_));
  NOR2_X1    g08193(.A1(new_n8442_), .A2(new_n8450_), .ZN(new_n8451_));
  OAI22_X1   g08194(.A1(new_n2452_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n2447_), .ZN(new_n8452_));
  NAND2_X1   g08195(.A1(new_n3312_), .A2(\b[29] ), .ZN(new_n8453_));
  AOI21_X1   g08196(.A1(new_n8452_), .A2(new_n8453_), .B(new_n2455_), .ZN(new_n8454_));
  NAND2_X1   g08197(.A1(new_n2546_), .A2(new_n8454_), .ZN(new_n8455_));
  XOR2_X1    g08198(.A1(new_n8455_), .A2(\a[32] ), .Z(new_n8456_));
  INV_X1     g08199(.I(new_n8456_), .ZN(new_n8457_));
  NAND2_X1   g08200(.A1(new_n8451_), .A2(new_n8457_), .ZN(new_n8458_));
  OAI21_X1   g08201(.A1(new_n8442_), .A2(new_n8450_), .B(new_n8456_), .ZN(new_n8459_));
  NAND2_X1   g08202(.A1(new_n8458_), .A2(new_n8459_), .ZN(new_n8460_));
  OAI22_X1   g08203(.A1(new_n2084_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n2079_), .ZN(new_n8461_));
  NAND2_X1   g08204(.A1(new_n2864_), .A2(\b[32] ), .ZN(new_n8462_));
  AOI21_X1   g08205(.A1(new_n8461_), .A2(new_n8462_), .B(new_n2087_), .ZN(new_n8463_));
  NAND2_X1   g08206(.A1(new_n2963_), .A2(new_n8463_), .ZN(new_n8464_));
  XOR2_X1    g08207(.A1(new_n8464_), .A2(\a[29] ), .Z(new_n8465_));
  XOR2_X1    g08208(.A1(new_n8460_), .A2(new_n8465_), .Z(new_n8466_));
  OAI22_X1   g08209(.A1(new_n1760_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n1755_), .ZN(new_n8467_));
  NAND2_X1   g08210(.A1(new_n2470_), .A2(\b[35] ), .ZN(new_n8468_));
  AOI21_X1   g08211(.A1(new_n8467_), .A2(new_n8468_), .B(new_n1763_), .ZN(new_n8469_));
  NAND2_X1   g08212(.A1(new_n3411_), .A2(new_n8469_), .ZN(new_n8470_));
  XOR2_X1    g08213(.A1(new_n8470_), .A2(\a[26] ), .Z(new_n8471_));
  NOR2_X1    g08214(.A1(new_n8466_), .A2(new_n8471_), .ZN(new_n8472_));
  AOI21_X1   g08215(.A1(new_n8458_), .A2(new_n8459_), .B(new_n8465_), .ZN(new_n8473_));
  INV_X1     g08216(.I(new_n8473_), .ZN(new_n8474_));
  NAND3_X1   g08217(.A1(new_n8458_), .A2(new_n8459_), .A3(new_n8465_), .ZN(new_n8475_));
  INV_X1     g08218(.I(new_n8471_), .ZN(new_n8476_));
  AOI21_X1   g08219(.A1(new_n8474_), .A2(new_n8475_), .B(new_n8476_), .ZN(new_n8477_));
  NOR2_X1    g08220(.A1(new_n8472_), .A2(new_n8477_), .ZN(new_n8478_));
  INV_X1     g08221(.I(new_n8478_), .ZN(new_n8479_));
  INV_X1     g08222(.I(new_n8171_), .ZN(new_n8480_));
  NAND3_X1   g08223(.A1(new_n8177_), .A2(new_n8178_), .A3(new_n8480_), .ZN(new_n8481_));
  OAI21_X1   g08224(.A1(new_n8165_), .A2(new_n8159_), .B(new_n8171_), .ZN(new_n8482_));
  AOI22_X1   g08225(.A1(new_n8482_), .A2(new_n8481_), .B1(new_n8480_), .B2(new_n8172_), .ZN(new_n8483_));
  OAI22_X1   g08226(.A1(new_n1444_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n1439_), .ZN(new_n8484_));
  NAND2_X1   g08227(.A1(new_n2098_), .A2(\b[38] ), .ZN(new_n8485_));
  AOI21_X1   g08228(.A1(new_n8484_), .A2(new_n8485_), .B(new_n1447_), .ZN(new_n8486_));
  NAND2_X1   g08229(.A1(new_n3844_), .A2(new_n8486_), .ZN(new_n8487_));
  XOR2_X1    g08230(.A1(new_n8487_), .A2(\a[23] ), .Z(new_n8488_));
  XOR2_X1    g08231(.A1(new_n8483_), .A2(new_n8488_), .Z(new_n8489_));
  NAND2_X1   g08232(.A1(new_n8489_), .A2(new_n8479_), .ZN(new_n8490_));
  XOR2_X1    g08233(.A1(new_n8483_), .A2(new_n8488_), .Z(new_n8491_));
  OAI21_X1   g08234(.A1(new_n8479_), .A2(new_n8491_), .B(new_n8490_), .ZN(new_n8492_));
  OAI22_X1   g08235(.A1(new_n1168_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n1163_), .ZN(new_n8493_));
  NAND2_X1   g08236(.A1(new_n1774_), .A2(\b[41] ), .ZN(new_n8494_));
  AOI21_X1   g08237(.A1(new_n8493_), .A2(new_n8494_), .B(new_n1171_), .ZN(new_n8495_));
  NAND2_X1   g08238(.A1(new_n4320_), .A2(new_n8495_), .ZN(new_n8496_));
  XOR2_X1    g08239(.A1(new_n8496_), .A2(\a[20] ), .Z(new_n8497_));
  INV_X1     g08240(.I(new_n8497_), .ZN(new_n8498_));
  NAND2_X1   g08241(.A1(new_n8492_), .A2(new_n8498_), .ZN(new_n8499_));
  NOR2_X1    g08242(.A1(new_n8491_), .A2(new_n8479_), .ZN(new_n8500_));
  AOI21_X1   g08243(.A1(new_n8479_), .A2(new_n8489_), .B(new_n8500_), .ZN(new_n8501_));
  NAND2_X1   g08244(.A1(new_n8501_), .A2(new_n8497_), .ZN(new_n8502_));
  NAND2_X1   g08245(.A1(new_n8502_), .A2(new_n8499_), .ZN(new_n8503_));
  OAI22_X1   g08246(.A1(new_n940_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n935_), .ZN(new_n8504_));
  NAND2_X1   g08247(.A1(new_n1458_), .A2(\b[44] ), .ZN(new_n8505_));
  AOI21_X1   g08248(.A1(new_n8504_), .A2(new_n8505_), .B(new_n943_), .ZN(new_n8506_));
  NAND2_X1   g08249(.A1(new_n4833_), .A2(new_n8506_), .ZN(new_n8507_));
  XOR2_X1    g08250(.A1(new_n8507_), .A2(\a[17] ), .Z(new_n8508_));
  XOR2_X1    g08251(.A1(new_n8503_), .A2(new_n8508_), .Z(new_n8509_));
  NOR2_X1    g08252(.A1(new_n8509_), .A2(new_n8290_), .ZN(new_n8510_));
  NAND2_X1   g08253(.A1(new_n8235_), .A2(new_n7945_), .ZN(new_n8511_));
  NAND2_X1   g08254(.A1(new_n8511_), .A2(new_n8232_), .ZN(new_n8512_));
  INV_X1     g08255(.I(new_n8508_), .ZN(new_n8513_));
  XOR2_X1    g08256(.A1(new_n8503_), .A2(new_n8513_), .Z(new_n8514_));
  NOR2_X1    g08257(.A1(new_n8514_), .A2(new_n8512_), .ZN(new_n8515_));
  OAI22_X1   g08258(.A1(new_n757_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n752_), .ZN(new_n8516_));
  NAND2_X1   g08259(.A1(new_n1182_), .A2(\b[47] ), .ZN(new_n8517_));
  AOI21_X1   g08260(.A1(new_n8516_), .A2(new_n8517_), .B(new_n760_), .ZN(new_n8518_));
  NAND2_X1   g08261(.A1(new_n5196_), .A2(new_n8518_), .ZN(new_n8519_));
  XOR2_X1    g08262(.A1(new_n8519_), .A2(\a[14] ), .Z(new_n8520_));
  NOR3_X1    g08263(.A1(new_n8510_), .A2(new_n8515_), .A3(new_n8520_), .ZN(new_n8521_));
  NOR2_X1    g08264(.A1(new_n8510_), .A2(new_n8515_), .ZN(new_n8522_));
  INV_X1     g08265(.I(new_n8520_), .ZN(new_n8523_));
  NOR2_X1    g08266(.A1(new_n8522_), .A2(new_n8523_), .ZN(new_n8524_));
  NOR2_X1    g08267(.A1(new_n8524_), .A2(new_n8521_), .ZN(new_n8525_));
  OAI22_X1   g08268(.A1(new_n582_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n577_), .ZN(new_n8526_));
  NAND2_X1   g08269(.A1(new_n960_), .A2(\b[50] ), .ZN(new_n8527_));
  AOI21_X1   g08270(.A1(new_n8526_), .A2(new_n8527_), .B(new_n585_), .ZN(new_n8528_));
  NAND2_X1   g08271(.A1(new_n5954_), .A2(new_n8528_), .ZN(new_n8529_));
  XOR2_X1    g08272(.A1(new_n8529_), .A2(\a[11] ), .Z(new_n8530_));
  INV_X1     g08273(.I(new_n8530_), .ZN(new_n8531_));
  XOR2_X1    g08274(.A1(new_n8525_), .A2(new_n8531_), .Z(new_n8532_));
  NAND2_X1   g08275(.A1(new_n8532_), .A2(new_n8287_), .ZN(new_n8533_));
  XOR2_X1    g08276(.A1(new_n8525_), .A2(new_n8531_), .Z(new_n8534_));
  OAI21_X1   g08277(.A1(new_n8287_), .A2(new_n8534_), .B(new_n8533_), .ZN(new_n8535_));
  OAI22_X1   g08278(.A1(new_n437_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n431_), .ZN(new_n8536_));
  NAND2_X1   g08279(.A1(new_n775_), .A2(\b[53] ), .ZN(new_n8537_));
  AOI21_X1   g08280(.A1(new_n8536_), .A2(new_n8537_), .B(new_n440_), .ZN(new_n8538_));
  NAND2_X1   g08281(.A1(new_n6471_), .A2(new_n8538_), .ZN(new_n8539_));
  XOR2_X1    g08282(.A1(new_n8539_), .A2(\a[8] ), .Z(new_n8540_));
  NOR2_X1    g08283(.A1(new_n8535_), .A2(new_n8540_), .ZN(new_n8541_));
  INV_X1     g08284(.I(new_n8541_), .ZN(new_n8542_));
  NAND2_X1   g08285(.A1(new_n8535_), .A2(new_n8540_), .ZN(new_n8543_));
  NAND2_X1   g08286(.A1(new_n8542_), .A2(new_n8543_), .ZN(new_n8544_));
  XOR2_X1    g08287(.A1(new_n7925_), .A2(\b[59] ), .Z(new_n8545_));
  NAND2_X1   g08288(.A1(new_n8545_), .A2(new_n7926_), .ZN(new_n8546_));
  NOR2_X1    g08289(.A1(new_n8546_), .A2(\b[61] ), .ZN(new_n8547_));
  INV_X1     g08290(.I(\b[61] ), .ZN(new_n8548_));
  AOI21_X1   g08291(.A1(new_n8545_), .A2(new_n7926_), .B(new_n8548_), .ZN(new_n8549_));
  OR2_X2     g08292(.A1(new_n8547_), .A2(new_n8549_), .Z(new_n8550_));
  OAI22_X1   g08293(.A1(new_n405_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n404_), .ZN(new_n8551_));
  NAND2_X1   g08294(.A1(new_n279_), .A2(\b[59] ), .ZN(new_n8552_));
  AOI21_X1   g08295(.A1(new_n8551_), .A2(new_n8552_), .B(new_n264_), .ZN(new_n8553_));
  NAND2_X1   g08296(.A1(new_n8550_), .A2(new_n8553_), .ZN(new_n8554_));
  XOR2_X1    g08297(.A1(new_n8554_), .A2(\a[2] ), .Z(new_n8555_));
  OAI22_X1   g08298(.A1(new_n364_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n320_), .ZN(new_n8556_));
  NAND2_X1   g08299(.A1(new_n594_), .A2(\b[56] ), .ZN(new_n8557_));
  AOI21_X1   g08300(.A1(new_n8556_), .A2(new_n8557_), .B(new_n312_), .ZN(new_n8558_));
  NAND2_X1   g08301(.A1(new_n7559_), .A2(new_n8558_), .ZN(new_n8559_));
  XOR2_X1    g08302(.A1(new_n8559_), .A2(\a[5] ), .Z(new_n8560_));
  XNOR2_X1   g08303(.A1(new_n8555_), .A2(new_n8560_), .ZN(new_n8561_));
  INV_X1     g08304(.I(new_n8561_), .ZN(new_n8562_));
  NOR2_X1    g08305(.A1(new_n8555_), .A2(new_n8560_), .ZN(new_n8563_));
  INV_X1     g08306(.I(new_n8563_), .ZN(new_n8564_));
  NAND2_X1   g08307(.A1(new_n8555_), .A2(new_n8560_), .ZN(new_n8565_));
  AOI21_X1   g08308(.A1(new_n8564_), .A2(new_n8565_), .B(new_n8544_), .ZN(new_n8566_));
  AOI21_X1   g08309(.A1(new_n8544_), .A2(new_n8562_), .B(new_n8566_), .ZN(new_n8567_));
  NOR2_X1    g08310(.A1(new_n7935_), .A2(new_n7940_), .ZN(new_n8568_));
  INV_X1     g08311(.I(new_n8276_), .ZN(new_n8569_));
  AOI21_X1   g08312(.A1(new_n7935_), .A2(new_n7940_), .B(new_n8569_), .ZN(new_n8570_));
  NOR2_X1    g08313(.A1(new_n8570_), .A2(new_n8568_), .ZN(new_n8571_));
  XNOR2_X1   g08314(.A1(new_n7935_), .A2(new_n7940_), .ZN(new_n8572_));
  XOR2_X1    g08315(.A1(new_n8276_), .A2(new_n8572_), .Z(new_n8573_));
  NAND2_X1   g08316(.A1(new_n8573_), .A2(new_n7941_), .ZN(new_n8574_));
  NAND2_X1   g08317(.A1(new_n8283_), .A2(new_n8574_), .ZN(new_n8575_));
  XOR2_X1    g08318(.A1(new_n8575_), .A2(new_n8571_), .Z(new_n8576_));
  XOR2_X1    g08319(.A1(new_n8576_), .A2(new_n8567_), .Z(\f[61] ));
  INV_X1     g08320(.I(new_n8571_), .ZN(new_n8578_));
  XOR2_X1    g08321(.A1(new_n8571_), .A2(new_n8567_), .Z(new_n8579_));
  NAND3_X1   g08322(.A1(new_n8283_), .A2(new_n8574_), .A3(new_n8579_), .ZN(new_n8580_));
  OAI21_X1   g08323(.A1(new_n8567_), .A2(new_n8578_), .B(new_n8580_), .ZN(new_n8581_));
  INV_X1     g08324(.I(new_n8565_), .ZN(new_n8582_));
  OAI21_X1   g08325(.A1(new_n8544_), .A2(new_n8582_), .B(new_n8564_), .ZN(new_n8583_));
  INV_X1     g08326(.I(new_n8521_), .ZN(new_n8584_));
  NOR2_X1    g08327(.A1(new_n8492_), .A2(new_n8497_), .ZN(new_n8585_));
  INV_X1     g08328(.I(new_n8488_), .ZN(new_n8586_));
  NAND2_X1   g08329(.A1(new_n8179_), .A2(new_n8171_), .ZN(new_n8587_));
  INV_X1     g08330(.I(new_n8172_), .ZN(new_n8588_));
  NOR3_X1    g08331(.A1(new_n8165_), .A2(new_n8159_), .A3(new_n8171_), .ZN(new_n8589_));
  AOI21_X1   g08332(.A1(new_n8177_), .A2(new_n8178_), .B(new_n8480_), .ZN(new_n8590_));
  OAI21_X1   g08333(.A1(new_n8589_), .A2(new_n8590_), .B(new_n8588_), .ZN(new_n8591_));
  NAND3_X1   g08334(.A1(new_n8591_), .A2(new_n8479_), .A3(new_n8587_), .ZN(new_n8592_));
  NAND2_X1   g08335(.A1(new_n8483_), .A2(new_n8478_), .ZN(new_n8593_));
  AOI21_X1   g08336(.A1(new_n8592_), .A2(new_n8593_), .B(new_n8586_), .ZN(new_n8594_));
  OAI22_X1   g08337(.A1(new_n2084_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n2079_), .ZN(new_n8595_));
  NAND2_X1   g08338(.A1(new_n2864_), .A2(\b[33] ), .ZN(new_n8596_));
  AOI21_X1   g08339(.A1(new_n8595_), .A2(new_n8596_), .B(new_n2087_), .ZN(new_n8597_));
  NAND2_X1   g08340(.A1(new_n3101_), .A2(new_n8597_), .ZN(new_n8598_));
  XOR2_X1    g08341(.A1(new_n8598_), .A2(\a[29] ), .Z(new_n8599_));
  INV_X1     g08342(.I(new_n8599_), .ZN(new_n8600_));
  OAI22_X1   g08343(.A1(new_n2452_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n2447_), .ZN(new_n8601_));
  NAND2_X1   g08344(.A1(new_n3312_), .A2(\b[30] ), .ZN(new_n8602_));
  AOI21_X1   g08345(.A1(new_n8601_), .A2(new_n8602_), .B(new_n2455_), .ZN(new_n8603_));
  NAND2_X1   g08346(.A1(new_n2659_), .A2(new_n8603_), .ZN(new_n8604_));
  XOR2_X1    g08347(.A1(new_n8604_), .A2(\a[32] ), .Z(new_n8605_));
  NOR2_X1    g08348(.A1(new_n8415_), .A2(new_n8414_), .ZN(new_n8606_));
  NOR2_X1    g08349(.A1(new_n8410_), .A2(new_n8606_), .ZN(new_n8607_));
  NOR2_X1    g08350(.A1(new_n8383_), .A2(new_n8380_), .ZN(new_n8608_));
  NOR3_X1    g08351(.A1(new_n8367_), .A2(new_n8355_), .A3(new_n8373_), .ZN(new_n8609_));
  INV_X1     g08352(.I(new_n8609_), .ZN(new_n8610_));
  INV_X1     g08353(.I(new_n8365_), .ZN(new_n8611_));
  AOI21_X1   g08354(.A1(new_n8361_), .A2(new_n8611_), .B(new_n8364_), .ZN(new_n8612_));
  AOI21_X1   g08355(.A1(new_n8342_), .A2(new_n8346_), .B(new_n8344_), .ZN(new_n8613_));
  INV_X1     g08356(.I(new_n8613_), .ZN(new_n8614_));
  AOI21_X1   g08357(.A1(new_n8303_), .A2(new_n8329_), .B(new_n8330_), .ZN(new_n8615_));
  NOR4_X1    g08358(.A1(new_n8322_), .A2(\a[62] ), .A3(\b[0] ), .A4(new_n8310_), .ZN(new_n8616_));
  OAI22_X1   g08359(.A1(new_n292_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n267_), .ZN(new_n8617_));
  XNOR2_X1   g08360(.A1(\a[59] ), .A2(\a[60] ), .ZN(new_n8618_));
  XNOR2_X1   g08361(.A1(\a[59] ), .A2(\a[61] ), .ZN(new_n8619_));
  NAND2_X1   g08362(.A1(new_n8618_), .A2(new_n8619_), .ZN(new_n8620_));
  XNOR2_X1   g08363(.A1(\a[59] ), .A2(\a[62] ), .ZN(new_n8621_));
  NAND2_X1   g08364(.A1(new_n8620_), .A2(new_n8621_), .ZN(new_n8622_));
  OAI21_X1   g08365(.A1(new_n258_), .A2(new_n8622_), .B(new_n8617_), .ZN(new_n8623_));
  NAND3_X1   g08366(.A1(new_n8623_), .A2(new_n5389_), .A3(new_n8320_), .ZN(new_n8624_));
  XOR2_X1    g08367(.A1(new_n8624_), .A2(new_n8309_), .Z(new_n8625_));
  XOR2_X1    g08368(.A1(new_n8625_), .A2(new_n8616_), .Z(new_n8626_));
  OAI22_X1   g08369(.A1(new_n347_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n393_), .ZN(new_n8627_));
  INV_X1     g08370(.I(new_n7611_), .ZN(new_n8628_));
  NAND2_X1   g08371(.A1(new_n8628_), .A2(\b[3] ), .ZN(new_n8629_));
  AOI21_X1   g08372(.A1(new_n8629_), .A2(new_n8627_), .B(new_n7354_), .ZN(new_n8630_));
  NAND2_X1   g08373(.A1(new_n352_), .A2(new_n8630_), .ZN(new_n8631_));
  XOR2_X1    g08374(.A1(new_n8631_), .A2(\a[59] ), .Z(new_n8632_));
  INV_X1     g08375(.I(new_n8632_), .ZN(new_n8633_));
  NAND2_X1   g08376(.A1(new_n8633_), .A2(new_n8626_), .ZN(new_n8634_));
  XOR2_X1    g08377(.A1(new_n8624_), .A2(\a[62] ), .Z(new_n8635_));
  XOR2_X1    g08378(.A1(new_n8635_), .A2(new_n8616_), .Z(new_n8636_));
  NAND2_X1   g08379(.A1(new_n8636_), .A2(new_n8632_), .ZN(new_n8637_));
  AOI21_X1   g08380(.A1(new_n8634_), .A2(new_n8637_), .B(new_n8615_), .ZN(new_n8638_));
  INV_X1     g08381(.I(new_n8615_), .ZN(new_n8639_));
  XOR2_X1    g08382(.A1(new_n8626_), .A2(new_n8632_), .Z(new_n8640_));
  NOR2_X1    g08383(.A1(new_n8640_), .A2(new_n8639_), .ZN(new_n8641_));
  NOR2_X1    g08384(.A1(new_n8641_), .A2(new_n8638_), .ZN(new_n8642_));
  OAI22_X1   g08385(.A1(new_n6721_), .A2(new_n450_), .B1(new_n6723_), .B2(new_n495_), .ZN(new_n8643_));
  NAND2_X1   g08386(.A1(new_n7617_), .A2(\b[6] ), .ZN(new_n8644_));
  AOI21_X1   g08387(.A1(new_n8644_), .A2(new_n8643_), .B(new_n6731_), .ZN(new_n8645_));
  NAND2_X1   g08388(.A1(new_n494_), .A2(new_n8645_), .ZN(new_n8646_));
  XOR2_X1    g08389(.A1(new_n8646_), .A2(\a[56] ), .Z(new_n8647_));
  XOR2_X1    g08390(.A1(new_n8642_), .A2(new_n8647_), .Z(new_n8648_));
  NAND2_X1   g08391(.A1(new_n8614_), .A2(new_n8648_), .ZN(new_n8649_));
  NOR2_X1    g08392(.A1(new_n8642_), .A2(new_n8647_), .ZN(new_n8650_));
  AND2_X2    g08393(.A1(new_n8642_), .A2(new_n8647_), .Z(new_n8651_));
  OAI21_X1   g08394(.A1(new_n8650_), .A2(new_n8651_), .B(new_n8613_), .ZN(new_n8652_));
  OAI22_X1   g08395(.A1(new_n5786_), .A2(new_n659_), .B1(new_n617_), .B2(new_n5792_), .ZN(new_n8653_));
  NAND2_X1   g08396(.A1(new_n6745_), .A2(\b[9] ), .ZN(new_n8654_));
  AOI21_X1   g08397(.A1(new_n8654_), .A2(new_n8653_), .B(new_n5796_), .ZN(new_n8655_));
  NAND2_X1   g08398(.A1(new_n663_), .A2(new_n8655_), .ZN(new_n8656_));
  XOR2_X1    g08399(.A1(new_n8656_), .A2(\a[53] ), .Z(new_n8657_));
  AOI21_X1   g08400(.A1(new_n8649_), .A2(new_n8652_), .B(new_n8657_), .ZN(new_n8658_));
  NAND3_X1   g08401(.A1(new_n8649_), .A2(new_n8652_), .A3(new_n8657_), .ZN(new_n8659_));
  INV_X1     g08402(.I(new_n8659_), .ZN(new_n8660_));
  NOR2_X1    g08403(.A1(new_n8660_), .A2(new_n8658_), .ZN(new_n8661_));
  NOR2_X1    g08404(.A1(new_n8612_), .A2(new_n8661_), .ZN(new_n8662_));
  OAI21_X1   g08405(.A1(new_n8299_), .A2(new_n8365_), .B(new_n8363_), .ZN(new_n8663_));
  INV_X1     g08406(.I(new_n8658_), .ZN(new_n8664_));
  NAND2_X1   g08407(.A1(new_n8664_), .A2(new_n8659_), .ZN(new_n8665_));
  NOR2_X1    g08408(.A1(new_n8663_), .A2(new_n8665_), .ZN(new_n8666_));
  OAI22_X1   g08409(.A1(new_n5228_), .A2(new_n848_), .B1(new_n795_), .B2(new_n5225_), .ZN(new_n8667_));
  NAND2_X1   g08410(.A1(new_n5387_), .A2(\b[12] ), .ZN(new_n8668_));
  AOI21_X1   g08411(.A1(new_n8667_), .A2(new_n8668_), .B(new_n5231_), .ZN(new_n8669_));
  NAND2_X1   g08412(.A1(new_n847_), .A2(new_n8669_), .ZN(new_n8670_));
  XOR2_X1    g08413(.A1(new_n8670_), .A2(\a[50] ), .Z(new_n8671_));
  NOR3_X1    g08414(.A1(new_n8666_), .A2(new_n8662_), .A3(new_n8671_), .ZN(new_n8672_));
  NAND2_X1   g08415(.A1(new_n8663_), .A2(new_n8665_), .ZN(new_n8673_));
  NAND2_X1   g08416(.A1(new_n8612_), .A2(new_n8661_), .ZN(new_n8674_));
  INV_X1     g08417(.I(new_n8671_), .ZN(new_n8675_));
  AOI21_X1   g08418(.A1(new_n8673_), .A2(new_n8674_), .B(new_n8675_), .ZN(new_n8676_));
  OAI22_X1   g08419(.A1(new_n4711_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n4706_), .ZN(new_n8677_));
  NAND2_X1   g08420(.A1(new_n5814_), .A2(\b[15] ), .ZN(new_n8678_));
  AOI21_X1   g08421(.A1(new_n8677_), .A2(new_n8678_), .B(new_n4714_), .ZN(new_n8679_));
  NAND2_X1   g08422(.A1(new_n1047_), .A2(new_n8679_), .ZN(new_n8680_));
  XOR2_X1    g08423(.A1(new_n8680_), .A2(\a[47] ), .Z(new_n8681_));
  INV_X1     g08424(.I(new_n8681_), .ZN(new_n8682_));
  OAI21_X1   g08425(.A1(new_n8676_), .A2(new_n8672_), .B(new_n8682_), .ZN(new_n8683_));
  NAND3_X1   g08426(.A1(new_n8673_), .A2(new_n8674_), .A3(new_n8675_), .ZN(new_n8684_));
  OAI21_X1   g08427(.A1(new_n8666_), .A2(new_n8662_), .B(new_n8671_), .ZN(new_n8685_));
  NAND3_X1   g08428(.A1(new_n8685_), .A2(new_n8684_), .A3(new_n8681_), .ZN(new_n8686_));
  AOI21_X1   g08429(.A1(new_n8683_), .A2(new_n8686_), .B(new_n8610_), .ZN(new_n8687_));
  NAND3_X1   g08430(.A1(new_n8685_), .A2(new_n8684_), .A3(new_n8682_), .ZN(new_n8688_));
  OAI21_X1   g08431(.A1(new_n8676_), .A2(new_n8672_), .B(new_n8681_), .ZN(new_n8689_));
  AOI21_X1   g08432(.A1(new_n8689_), .A2(new_n8688_), .B(new_n8609_), .ZN(new_n8690_));
  OAI21_X1   g08433(.A1(new_n8687_), .A2(new_n8690_), .B(new_n8608_), .ZN(new_n8691_));
  AOI21_X1   g08434(.A1(new_n8685_), .A2(new_n8684_), .B(new_n8681_), .ZN(new_n8692_));
  NOR3_X1    g08435(.A1(new_n8676_), .A2(new_n8672_), .A3(new_n8682_), .ZN(new_n8693_));
  OAI21_X1   g08436(.A1(new_n8693_), .A2(new_n8692_), .B(new_n8609_), .ZN(new_n8694_));
  NOR3_X1    g08437(.A1(new_n8676_), .A2(new_n8672_), .A3(new_n8681_), .ZN(new_n8695_));
  AOI21_X1   g08438(.A1(new_n8685_), .A2(new_n8684_), .B(new_n8682_), .ZN(new_n8696_));
  OAI21_X1   g08439(.A1(new_n8695_), .A2(new_n8696_), .B(new_n8610_), .ZN(new_n8697_));
  NAND3_X1   g08440(.A1(new_n8694_), .A2(new_n8697_), .A3(new_n8382_), .ZN(new_n8698_));
  OAI22_X1   g08441(.A1(new_n4208_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n4203_), .ZN(new_n8699_));
  NAND2_X1   g08442(.A1(new_n5244_), .A2(\b[18] ), .ZN(new_n8700_));
  AOI21_X1   g08443(.A1(new_n8699_), .A2(new_n8700_), .B(new_n4211_), .ZN(new_n8701_));
  NAND2_X1   g08444(.A1(new_n1304_), .A2(new_n8701_), .ZN(new_n8702_));
  XOR2_X1    g08445(.A1(new_n8702_), .A2(\a[44] ), .Z(new_n8703_));
  AOI21_X1   g08446(.A1(new_n8691_), .A2(new_n8698_), .B(new_n8703_), .ZN(new_n8704_));
  INV_X1     g08447(.I(new_n8704_), .ZN(new_n8705_));
  NAND3_X1   g08448(.A1(new_n8691_), .A2(new_n8698_), .A3(new_n8703_), .ZN(new_n8706_));
  OAI22_X1   g08449(.A1(new_n3736_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n3731_), .ZN(new_n8707_));
  NAND2_X1   g08450(.A1(new_n4730_), .A2(\b[21] ), .ZN(new_n8708_));
  AOI21_X1   g08451(.A1(new_n8707_), .A2(new_n8708_), .B(new_n3739_), .ZN(new_n8709_));
  NAND2_X1   g08452(.A1(new_n1604_), .A2(new_n8709_), .ZN(new_n8710_));
  XOR2_X1    g08453(.A1(new_n8710_), .A2(\a[41] ), .Z(new_n8711_));
  AOI21_X1   g08454(.A1(new_n8705_), .A2(new_n8706_), .B(new_n8711_), .ZN(new_n8712_));
  INV_X1     g08455(.I(new_n8706_), .ZN(new_n8713_));
  INV_X1     g08456(.I(new_n8711_), .ZN(new_n8714_));
  NOR3_X1    g08457(.A1(new_n8713_), .A2(new_n8704_), .A3(new_n8714_), .ZN(new_n8715_));
  NOR2_X1    g08458(.A1(new_n8712_), .A2(new_n8715_), .ZN(new_n8716_));
  INV_X1     g08459(.I(new_n8716_), .ZN(new_n8717_));
  OAI21_X1   g08460(.A1(new_n8607_), .A2(new_n8406_), .B(new_n8717_), .ZN(new_n8718_));
  NAND2_X1   g08461(.A1(new_n8423_), .A2(new_n8054_), .ZN(new_n8719_));
  NAND2_X1   g08462(.A1(new_n8413_), .A2(new_n8719_), .ZN(new_n8720_));
  NAND3_X1   g08463(.A1(new_n8720_), .A2(new_n8412_), .A3(new_n8716_), .ZN(new_n8721_));
  OAI22_X1   g08464(.A1(new_n3298_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n3293_), .ZN(new_n8722_));
  NAND2_X1   g08465(.A1(new_n4227_), .A2(\b[24] ), .ZN(new_n8723_));
  AOI21_X1   g08466(.A1(new_n8722_), .A2(new_n8723_), .B(new_n3301_), .ZN(new_n8724_));
  NAND2_X1   g08467(.A1(new_n1926_), .A2(new_n8724_), .ZN(new_n8725_));
  XOR2_X1    g08468(.A1(new_n8725_), .A2(\a[38] ), .Z(new_n8726_));
  INV_X1     g08469(.I(new_n8726_), .ZN(new_n8727_));
  NAND3_X1   g08470(.A1(new_n8718_), .A2(new_n8721_), .A3(new_n8727_), .ZN(new_n8728_));
  AOI21_X1   g08471(.A1(new_n8720_), .A2(new_n8412_), .B(new_n8716_), .ZN(new_n8729_));
  NOR3_X1    g08472(.A1(new_n8607_), .A2(new_n8406_), .A3(new_n8717_), .ZN(new_n8730_));
  OAI21_X1   g08473(.A1(new_n8730_), .A2(new_n8729_), .B(new_n8726_), .ZN(new_n8731_));
  NAND2_X1   g08474(.A1(new_n8731_), .A2(new_n8728_), .ZN(new_n8732_));
  NAND2_X1   g08475(.A1(new_n8411_), .A2(new_n8719_), .ZN(new_n8733_));
  NAND2_X1   g08476(.A1(new_n8443_), .A2(new_n8606_), .ZN(new_n8734_));
  AOI21_X1   g08477(.A1(new_n8733_), .A2(new_n8734_), .B(new_n8421_), .ZN(new_n8735_));
  NOR3_X1    g08478(.A1(new_n8431_), .A2(new_n8447_), .A3(new_n8073_), .ZN(new_n8736_));
  NOR3_X1    g08479(.A1(new_n8736_), .A2(new_n8732_), .A3(new_n8735_), .ZN(new_n8737_));
  NOR3_X1    g08480(.A1(new_n8730_), .A2(new_n8729_), .A3(new_n8726_), .ZN(new_n8738_));
  AOI21_X1   g08481(.A1(new_n8718_), .A2(new_n8721_), .B(new_n8727_), .ZN(new_n8739_));
  NOR2_X1    g08482(.A1(new_n8738_), .A2(new_n8739_), .ZN(new_n8740_));
  INV_X1     g08483(.I(new_n8735_), .ZN(new_n8741_));
  NAND3_X1   g08484(.A1(new_n8440_), .A2(new_n8107_), .A3(new_n8429_), .ZN(new_n8742_));
  AOI21_X1   g08485(.A1(new_n8741_), .A2(new_n8742_), .B(new_n8740_), .ZN(new_n8743_));
  OAI22_X1   g08486(.A1(new_n2846_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n2841_), .ZN(new_n8744_));
  NAND2_X1   g08487(.A1(new_n3755_), .A2(\b[27] ), .ZN(new_n8745_));
  AOI21_X1   g08488(.A1(new_n8744_), .A2(new_n8745_), .B(new_n2849_), .ZN(new_n8746_));
  NAND2_X1   g08489(.A1(new_n2276_), .A2(new_n8746_), .ZN(new_n8747_));
  XOR2_X1    g08490(.A1(new_n8747_), .A2(\a[35] ), .Z(new_n8748_));
  NOR3_X1    g08491(.A1(new_n8743_), .A2(new_n8737_), .A3(new_n8748_), .ZN(new_n8749_));
  NAND3_X1   g08492(.A1(new_n8740_), .A2(new_n8742_), .A3(new_n8741_), .ZN(new_n8750_));
  OAI21_X1   g08493(.A1(new_n8735_), .A2(new_n8736_), .B(new_n8732_), .ZN(new_n8751_));
  INV_X1     g08494(.I(new_n8748_), .ZN(new_n8752_));
  AOI21_X1   g08495(.A1(new_n8751_), .A2(new_n8750_), .B(new_n8752_), .ZN(new_n8753_));
  AOI21_X1   g08496(.A1(new_n8440_), .A2(new_n8107_), .B(new_n8447_), .ZN(new_n8754_));
  NOR3_X1    g08497(.A1(new_n8431_), .A2(new_n8073_), .A3(new_n8429_), .ZN(new_n8755_));
  OAI21_X1   g08498(.A1(new_n8754_), .A2(new_n8755_), .B(new_n8436_), .ZN(new_n8756_));
  OAI21_X1   g08499(.A1(new_n8442_), .A2(new_n8450_), .B(new_n8756_), .ZN(new_n8757_));
  NOR3_X1    g08500(.A1(new_n8749_), .A2(new_n8757_), .A3(new_n8753_), .ZN(new_n8758_));
  NAND3_X1   g08501(.A1(new_n8751_), .A2(new_n8750_), .A3(new_n8752_), .ZN(new_n8759_));
  OAI21_X1   g08502(.A1(new_n8743_), .A2(new_n8737_), .B(new_n8748_), .ZN(new_n8760_));
  AOI21_X1   g08503(.A1(new_n8440_), .A2(new_n8107_), .B(new_n8436_), .ZN(new_n8761_));
  NOR3_X1    g08504(.A1(new_n8431_), .A2(new_n8073_), .A3(new_n8437_), .ZN(new_n8762_));
  OAI21_X1   g08505(.A1(new_n8761_), .A2(new_n8762_), .B(new_n8447_), .ZN(new_n8763_));
  NOR3_X1    g08506(.A1(new_n8431_), .A2(new_n8073_), .A3(new_n8436_), .ZN(new_n8764_));
  AOI21_X1   g08507(.A1(new_n8440_), .A2(new_n8107_), .B(new_n8437_), .ZN(new_n8765_));
  OAI21_X1   g08508(.A1(new_n8765_), .A2(new_n8764_), .B(new_n8429_), .ZN(new_n8766_));
  OAI21_X1   g08509(.A1(new_n8431_), .A2(new_n8073_), .B(new_n8429_), .ZN(new_n8767_));
  NAND3_X1   g08510(.A1(new_n8440_), .A2(new_n8447_), .A3(new_n8107_), .ZN(new_n8768_));
  NAND2_X1   g08511(.A1(new_n8768_), .A2(new_n8767_), .ZN(new_n8769_));
  AOI22_X1   g08512(.A1(new_n8763_), .A2(new_n8766_), .B1(new_n8436_), .B2(new_n8769_), .ZN(new_n8770_));
  AOI21_X1   g08513(.A1(new_n8759_), .A2(new_n8760_), .B(new_n8770_), .ZN(new_n8771_));
  NOR3_X1    g08514(.A1(new_n8771_), .A2(new_n8758_), .A3(new_n8459_), .ZN(new_n8772_));
  INV_X1     g08515(.I(new_n8459_), .ZN(new_n8773_));
  NAND3_X1   g08516(.A1(new_n8770_), .A2(new_n8760_), .A3(new_n8759_), .ZN(new_n8774_));
  OAI21_X1   g08517(.A1(new_n8749_), .A2(new_n8753_), .B(new_n8757_), .ZN(new_n8775_));
  AOI21_X1   g08518(.A1(new_n8775_), .A2(new_n8774_), .B(new_n8773_), .ZN(new_n8776_));
  OAI21_X1   g08519(.A1(new_n8772_), .A2(new_n8776_), .B(new_n8605_), .ZN(new_n8777_));
  INV_X1     g08520(.I(new_n8605_), .ZN(new_n8778_));
  NAND3_X1   g08521(.A1(new_n8775_), .A2(new_n8774_), .A3(new_n8773_), .ZN(new_n8779_));
  OAI21_X1   g08522(.A1(new_n8771_), .A2(new_n8758_), .B(new_n8459_), .ZN(new_n8780_));
  NAND3_X1   g08523(.A1(new_n8780_), .A2(new_n8779_), .A3(new_n8778_), .ZN(new_n8781_));
  AOI21_X1   g08524(.A1(new_n8777_), .A2(new_n8781_), .B(new_n8600_), .ZN(new_n8782_));
  AOI21_X1   g08525(.A1(new_n8780_), .A2(new_n8779_), .B(new_n8778_), .ZN(new_n8783_));
  NOR3_X1    g08526(.A1(new_n8772_), .A2(new_n8776_), .A3(new_n8605_), .ZN(new_n8784_));
  NOR3_X1    g08527(.A1(new_n8784_), .A2(new_n8783_), .A3(new_n8599_), .ZN(new_n8785_));
  NOR3_X1    g08528(.A1(new_n8785_), .A2(new_n8782_), .A3(new_n8474_), .ZN(new_n8786_));
  OAI21_X1   g08529(.A1(new_n8784_), .A2(new_n8783_), .B(new_n8599_), .ZN(new_n8787_));
  NAND3_X1   g08530(.A1(new_n8777_), .A2(new_n8781_), .A3(new_n8600_), .ZN(new_n8788_));
  AOI21_X1   g08531(.A1(new_n8787_), .A2(new_n8788_), .B(new_n8473_), .ZN(new_n8789_));
  OAI22_X1   g08532(.A1(new_n1760_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n1755_), .ZN(new_n8790_));
  NAND2_X1   g08533(.A1(new_n2470_), .A2(\b[36] ), .ZN(new_n8791_));
  AOI21_X1   g08534(.A1(new_n8790_), .A2(new_n8791_), .B(new_n1763_), .ZN(new_n8792_));
  NAND2_X1   g08535(.A1(new_n3565_), .A2(new_n8792_), .ZN(new_n8793_));
  XOR2_X1    g08536(.A1(new_n8793_), .A2(\a[26] ), .Z(new_n8794_));
  NOR3_X1    g08537(.A1(new_n8786_), .A2(new_n8789_), .A3(new_n8794_), .ZN(new_n8795_));
  NAND3_X1   g08538(.A1(new_n8787_), .A2(new_n8788_), .A3(new_n8473_), .ZN(new_n8796_));
  OAI21_X1   g08539(.A1(new_n8785_), .A2(new_n8782_), .B(new_n8474_), .ZN(new_n8797_));
  INV_X1     g08540(.I(new_n8794_), .ZN(new_n8798_));
  AOI21_X1   g08541(.A1(new_n8797_), .A2(new_n8796_), .B(new_n8798_), .ZN(new_n8799_));
  INV_X1     g08542(.I(new_n8477_), .ZN(new_n8800_));
  OAI21_X1   g08543(.A1(new_n8483_), .A2(new_n8479_), .B(new_n8800_), .ZN(new_n8801_));
  NOR3_X1    g08544(.A1(new_n8801_), .A2(new_n8795_), .A3(new_n8799_), .ZN(new_n8802_));
  NAND3_X1   g08545(.A1(new_n8797_), .A2(new_n8796_), .A3(new_n8798_), .ZN(new_n8803_));
  OAI21_X1   g08546(.A1(new_n8786_), .A2(new_n8789_), .B(new_n8794_), .ZN(new_n8804_));
  NAND3_X1   g08547(.A1(new_n8591_), .A2(new_n8478_), .A3(new_n8587_), .ZN(new_n8805_));
  AOI22_X1   g08548(.A1(new_n8805_), .A2(new_n8800_), .B1(new_n8803_), .B2(new_n8804_), .ZN(new_n8806_));
  OAI22_X1   g08549(.A1(new_n1444_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n1439_), .ZN(new_n8807_));
  NAND2_X1   g08550(.A1(new_n2098_), .A2(\b[39] ), .ZN(new_n8808_));
  AOI21_X1   g08551(.A1(new_n8807_), .A2(new_n8808_), .B(new_n1447_), .ZN(new_n8809_));
  NAND2_X1   g08552(.A1(new_n3996_), .A2(new_n8809_), .ZN(new_n8810_));
  XOR2_X1    g08553(.A1(new_n8810_), .A2(\a[23] ), .Z(new_n8811_));
  NOR3_X1    g08554(.A1(new_n8806_), .A2(new_n8802_), .A3(new_n8811_), .ZN(new_n8812_));
  NAND4_X1   g08555(.A1(new_n8805_), .A2(new_n8800_), .A3(new_n8803_), .A4(new_n8804_), .ZN(new_n8813_));
  NOR2_X1    g08556(.A1(new_n8483_), .A2(new_n8479_), .ZN(new_n8814_));
  OAI22_X1   g08557(.A1(new_n8814_), .A2(new_n8477_), .B1(new_n8795_), .B2(new_n8799_), .ZN(new_n8815_));
  INV_X1     g08558(.I(new_n8811_), .ZN(new_n8816_));
  AOI21_X1   g08559(.A1(new_n8815_), .A2(new_n8813_), .B(new_n8816_), .ZN(new_n8817_));
  OAI21_X1   g08560(.A1(new_n8812_), .A2(new_n8817_), .B(new_n8594_), .ZN(new_n8818_));
  INV_X1     g08561(.I(new_n8594_), .ZN(new_n8819_));
  AOI21_X1   g08562(.A1(new_n8815_), .A2(new_n8813_), .B(new_n8811_), .ZN(new_n8820_));
  NOR3_X1    g08563(.A1(new_n8806_), .A2(new_n8802_), .A3(new_n8816_), .ZN(new_n8821_));
  OAI21_X1   g08564(.A1(new_n8821_), .A2(new_n8820_), .B(new_n8819_), .ZN(new_n8822_));
  OAI22_X1   g08565(.A1(new_n1168_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n1163_), .ZN(new_n8823_));
  NAND2_X1   g08566(.A1(new_n1774_), .A2(\b[42] ), .ZN(new_n8824_));
  AOI21_X1   g08567(.A1(new_n8823_), .A2(new_n8824_), .B(new_n1171_), .ZN(new_n8825_));
  NAND2_X1   g08568(.A1(new_n4500_), .A2(new_n8825_), .ZN(new_n8826_));
  XOR2_X1    g08569(.A1(new_n8826_), .A2(\a[20] ), .Z(new_n8827_));
  AOI21_X1   g08570(.A1(new_n8818_), .A2(new_n8822_), .B(new_n8827_), .ZN(new_n8828_));
  NAND3_X1   g08571(.A1(new_n8815_), .A2(new_n8813_), .A3(new_n8816_), .ZN(new_n8829_));
  OAI21_X1   g08572(.A1(new_n8806_), .A2(new_n8802_), .B(new_n8811_), .ZN(new_n8830_));
  AOI21_X1   g08573(.A1(new_n8830_), .A2(new_n8829_), .B(new_n8819_), .ZN(new_n8831_));
  OAI21_X1   g08574(.A1(new_n8806_), .A2(new_n8802_), .B(new_n8816_), .ZN(new_n8832_));
  NAND3_X1   g08575(.A1(new_n8815_), .A2(new_n8813_), .A3(new_n8811_), .ZN(new_n8833_));
  AOI21_X1   g08576(.A1(new_n8832_), .A2(new_n8833_), .B(new_n8594_), .ZN(new_n8834_));
  INV_X1     g08577(.I(new_n8827_), .ZN(new_n8835_));
  NOR3_X1    g08578(.A1(new_n8831_), .A2(new_n8834_), .A3(new_n8835_), .ZN(new_n8836_));
  OAI22_X1   g08579(.A1(new_n940_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n935_), .ZN(new_n8837_));
  NAND2_X1   g08580(.A1(new_n1458_), .A2(\b[45] ), .ZN(new_n8838_));
  AOI21_X1   g08581(.A1(new_n8837_), .A2(new_n8838_), .B(new_n943_), .ZN(new_n8839_));
  NAND2_X1   g08582(.A1(new_n5004_), .A2(new_n8839_), .ZN(new_n8840_));
  XOR2_X1    g08583(.A1(new_n8840_), .A2(\a[17] ), .Z(new_n8841_));
  NOR3_X1    g08584(.A1(new_n8828_), .A2(new_n8836_), .A3(new_n8841_), .ZN(new_n8842_));
  OAI21_X1   g08585(.A1(new_n8831_), .A2(new_n8834_), .B(new_n8835_), .ZN(new_n8843_));
  NAND3_X1   g08586(.A1(new_n8818_), .A2(new_n8822_), .A3(new_n8827_), .ZN(new_n8844_));
  INV_X1     g08587(.I(new_n8841_), .ZN(new_n8845_));
  AOI21_X1   g08588(.A1(new_n8843_), .A2(new_n8844_), .B(new_n8845_), .ZN(new_n8846_));
  OAI21_X1   g08589(.A1(new_n8846_), .A2(new_n8842_), .B(new_n8585_), .ZN(new_n8847_));
  INV_X1     g08590(.I(new_n8585_), .ZN(new_n8848_));
  AOI21_X1   g08591(.A1(new_n8843_), .A2(new_n8844_), .B(new_n8841_), .ZN(new_n8849_));
  NOR3_X1    g08592(.A1(new_n8828_), .A2(new_n8836_), .A3(new_n8845_), .ZN(new_n8850_));
  OAI21_X1   g08593(.A1(new_n8849_), .A2(new_n8850_), .B(new_n8848_), .ZN(new_n8851_));
  XOR2_X1    g08594(.A1(new_n8492_), .A2(new_n8498_), .Z(new_n8852_));
  AOI21_X1   g08595(.A1(new_n8511_), .A2(new_n8232_), .B(new_n8852_), .ZN(new_n8853_));
  NAND3_X1   g08596(.A1(new_n8847_), .A2(new_n8851_), .A3(new_n8853_), .ZN(new_n8854_));
  NAND3_X1   g08597(.A1(new_n8843_), .A2(new_n8844_), .A3(new_n8845_), .ZN(new_n8855_));
  OAI21_X1   g08598(.A1(new_n8828_), .A2(new_n8836_), .B(new_n8841_), .ZN(new_n8856_));
  AOI21_X1   g08599(.A1(new_n8856_), .A2(new_n8855_), .B(new_n8848_), .ZN(new_n8857_));
  OAI21_X1   g08600(.A1(new_n8828_), .A2(new_n8836_), .B(new_n8845_), .ZN(new_n8858_));
  NAND3_X1   g08601(.A1(new_n8843_), .A2(new_n8844_), .A3(new_n8841_), .ZN(new_n8859_));
  AOI21_X1   g08602(.A1(new_n8858_), .A2(new_n8859_), .B(new_n8585_), .ZN(new_n8860_));
  OAI21_X1   g08603(.A1(new_n8289_), .A2(new_n8288_), .B(new_n8503_), .ZN(new_n8861_));
  OAI21_X1   g08604(.A1(new_n8857_), .A2(new_n8860_), .B(new_n8861_), .ZN(new_n8862_));
  NAND3_X1   g08605(.A1(new_n8511_), .A2(new_n8232_), .A3(new_n8503_), .ZN(new_n8863_));
  OAI21_X1   g08606(.A1(new_n8289_), .A2(new_n8288_), .B(new_n8852_), .ZN(new_n8864_));
  AOI21_X1   g08607(.A1(new_n8864_), .A2(new_n8863_), .B(new_n8508_), .ZN(new_n8865_));
  NAND3_X1   g08608(.A1(new_n8862_), .A2(new_n8854_), .A3(new_n8865_), .ZN(new_n8866_));
  NOR3_X1    g08609(.A1(new_n8857_), .A2(new_n8860_), .A3(new_n8861_), .ZN(new_n8867_));
  AOI21_X1   g08610(.A1(new_n8847_), .A2(new_n8851_), .B(new_n8853_), .ZN(new_n8868_));
  NOR3_X1    g08611(.A1(new_n8289_), .A2(new_n8852_), .A3(new_n8288_), .ZN(new_n8869_));
  AOI21_X1   g08612(.A1(new_n8511_), .A2(new_n8232_), .B(new_n8503_), .ZN(new_n8870_));
  OAI21_X1   g08613(.A1(new_n8870_), .A2(new_n8869_), .B(new_n8513_), .ZN(new_n8871_));
  OAI21_X1   g08614(.A1(new_n8868_), .A2(new_n8867_), .B(new_n8871_), .ZN(new_n8872_));
  OAI22_X1   g08615(.A1(new_n757_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n752_), .ZN(new_n8873_));
  NAND2_X1   g08616(.A1(new_n1182_), .A2(\b[48] ), .ZN(new_n8874_));
  AOI21_X1   g08617(.A1(new_n8873_), .A2(new_n8874_), .B(new_n760_), .ZN(new_n8875_));
  NAND2_X1   g08618(.A1(new_n5537_), .A2(new_n8875_), .ZN(new_n8876_));
  XOR2_X1    g08619(.A1(new_n8876_), .A2(\a[14] ), .Z(new_n8877_));
  INV_X1     g08620(.I(new_n8877_), .ZN(new_n8878_));
  NAND3_X1   g08621(.A1(new_n8872_), .A2(new_n8866_), .A3(new_n8878_), .ZN(new_n8879_));
  NOR3_X1    g08622(.A1(new_n8868_), .A2(new_n8867_), .A3(new_n8871_), .ZN(new_n8880_));
  AOI21_X1   g08623(.A1(new_n8862_), .A2(new_n8854_), .B(new_n8865_), .ZN(new_n8881_));
  OAI21_X1   g08624(.A1(new_n8881_), .A2(new_n8880_), .B(new_n8877_), .ZN(new_n8882_));
  OAI22_X1   g08625(.A1(new_n582_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n577_), .ZN(new_n8883_));
  NAND2_X1   g08626(.A1(new_n960_), .A2(\b[51] ), .ZN(new_n8884_));
  AOI21_X1   g08627(.A1(new_n8883_), .A2(new_n8884_), .B(new_n585_), .ZN(new_n8885_));
  NAND2_X1   g08628(.A1(new_n6219_), .A2(new_n8885_), .ZN(new_n8886_));
  XOR2_X1    g08629(.A1(new_n8886_), .A2(\a[11] ), .Z(new_n8887_));
  INV_X1     g08630(.I(new_n8887_), .ZN(new_n8888_));
  NAND3_X1   g08631(.A1(new_n8882_), .A2(new_n8879_), .A3(new_n8888_), .ZN(new_n8889_));
  NOR3_X1    g08632(.A1(new_n8881_), .A2(new_n8880_), .A3(new_n8877_), .ZN(new_n8890_));
  AOI21_X1   g08633(.A1(new_n8872_), .A2(new_n8866_), .B(new_n8878_), .ZN(new_n8891_));
  OAI21_X1   g08634(.A1(new_n8890_), .A2(new_n8891_), .B(new_n8887_), .ZN(new_n8892_));
  AOI21_X1   g08635(.A1(new_n8892_), .A2(new_n8889_), .B(new_n8584_), .ZN(new_n8893_));
  OAI21_X1   g08636(.A1(new_n8890_), .A2(new_n8891_), .B(new_n8888_), .ZN(new_n8894_));
  NAND3_X1   g08637(.A1(new_n8882_), .A2(new_n8879_), .A3(new_n8887_), .ZN(new_n8895_));
  AOI21_X1   g08638(.A1(new_n8894_), .A2(new_n8895_), .B(new_n8521_), .ZN(new_n8896_));
  NOR2_X1    g08639(.A1(new_n8893_), .A2(new_n8896_), .ZN(new_n8897_));
  NOR2_X1    g08640(.A1(new_n8259_), .A2(new_n8254_), .ZN(new_n8898_));
  NAND2_X1   g08641(.A1(new_n7879_), .A2(new_n7577_), .ZN(new_n8899_));
  AOI22_X1   g08642(.A1(new_n8259_), .A2(new_n8254_), .B1(new_n8899_), .B2(new_n7878_), .ZN(new_n8900_));
  NOR3_X1    g08643(.A1(new_n8900_), .A2(new_n8898_), .A3(new_n8530_), .ZN(new_n8901_));
  AOI21_X1   g08644(.A1(new_n8286_), .A2(new_n8258_), .B(new_n8531_), .ZN(new_n8902_));
  OAI21_X1   g08645(.A1(new_n8902_), .A2(new_n8901_), .B(new_n8525_), .ZN(new_n8903_));
  XOR2_X1    g08646(.A1(new_n8897_), .A2(new_n8903_), .Z(new_n8904_));
  AOI21_X1   g08647(.A1(new_n8286_), .A2(new_n8258_), .B(new_n8530_), .ZN(new_n8905_));
  XOR2_X1    g08648(.A1(new_n8904_), .A2(new_n8905_), .Z(new_n8906_));
  OAI22_X1   g08649(.A1(new_n364_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n320_), .ZN(new_n8907_));
  NAND2_X1   g08650(.A1(new_n594_), .A2(\b[57] ), .ZN(new_n8908_));
  AOI21_X1   g08651(.A1(new_n8907_), .A2(new_n8908_), .B(new_n312_), .ZN(new_n8909_));
  NAND2_X1   g08652(.A1(new_n7895_), .A2(new_n8909_), .ZN(new_n8910_));
  XOR2_X1    g08653(.A1(new_n8910_), .A2(\a[5] ), .Z(new_n8911_));
  OAI22_X1   g08654(.A1(new_n437_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n431_), .ZN(new_n8912_));
  NAND2_X1   g08655(.A1(new_n775_), .A2(\b[54] ), .ZN(new_n8913_));
  AOI21_X1   g08656(.A1(new_n8912_), .A2(new_n8913_), .B(new_n440_), .ZN(new_n8914_));
  NAND2_X1   g08657(.A1(new_n6994_), .A2(new_n8914_), .ZN(new_n8915_));
  XOR2_X1    g08658(.A1(new_n8915_), .A2(\a[8] ), .Z(new_n8916_));
  XNOR2_X1   g08659(.A1(new_n8911_), .A2(new_n8916_), .ZN(new_n8917_));
  INV_X1     g08660(.I(new_n8917_), .ZN(new_n8918_));
  NOR2_X1    g08661(.A1(new_n8911_), .A2(new_n8916_), .ZN(new_n8919_));
  NAND2_X1   g08662(.A1(new_n8911_), .A2(new_n8916_), .ZN(new_n8920_));
  INV_X1     g08663(.I(new_n8920_), .ZN(new_n8921_));
  NOR2_X1    g08664(.A1(new_n8921_), .A2(new_n8919_), .ZN(new_n8922_));
  NOR2_X1    g08665(.A1(new_n8906_), .A2(new_n8922_), .ZN(new_n8923_));
  AOI21_X1   g08666(.A1(new_n8906_), .A2(new_n8918_), .B(new_n8923_), .ZN(new_n8924_));
  OAI21_X1   g08667(.A1(new_n7890_), .A2(new_n8548_), .B(new_n7930_), .ZN(new_n8925_));
  NAND3_X1   g08668(.A1(new_n7923_), .A2(new_n7924_), .A3(new_n8925_), .ZN(new_n8926_));
  OAI21_X1   g08669(.A1(\b[59] ), .A2(\b[61] ), .B(\b[60] ), .ZN(new_n8927_));
  XNOR2_X1   g08670(.A1(\b[61] ), .A2(\b[62] ), .ZN(new_n8928_));
  AOI21_X1   g08671(.A1(new_n8926_), .A2(new_n8927_), .B(new_n8928_), .ZN(new_n8929_));
  NAND2_X1   g08672(.A1(new_n8926_), .A2(new_n8927_), .ZN(new_n8930_));
  NAND2_X1   g08673(.A1(\b[61] ), .A2(\b[62] ), .ZN(new_n8931_));
  INV_X1     g08674(.I(\b[62] ), .ZN(new_n8932_));
  NAND2_X1   g08675(.A1(new_n8548_), .A2(new_n8932_), .ZN(new_n8933_));
  AOI21_X1   g08676(.A1(new_n8931_), .A2(new_n8933_), .B(new_n8930_), .ZN(new_n8934_));
  OR2_X2     g08677(.A1(new_n8934_), .A2(new_n8929_), .Z(new_n8935_));
  OAI22_X1   g08678(.A1(new_n405_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n404_), .ZN(new_n8936_));
  NAND2_X1   g08679(.A1(new_n279_), .A2(\b[60] ), .ZN(new_n8937_));
  AOI21_X1   g08680(.A1(new_n8936_), .A2(new_n8937_), .B(new_n264_), .ZN(new_n8938_));
  NAND2_X1   g08681(.A1(new_n8935_), .A2(new_n8938_), .ZN(new_n8939_));
  XOR2_X1    g08682(.A1(new_n8939_), .A2(\a[2] ), .Z(new_n8940_));
  XOR2_X1    g08683(.A1(new_n8924_), .A2(new_n8940_), .Z(new_n8941_));
  NAND2_X1   g08684(.A1(new_n8941_), .A2(new_n8541_), .ZN(new_n8942_));
  NOR2_X1    g08685(.A1(new_n8924_), .A2(new_n8940_), .ZN(new_n8943_));
  NAND2_X1   g08686(.A1(new_n8924_), .A2(new_n8940_), .ZN(new_n8944_));
  INV_X1     g08687(.I(new_n8944_), .ZN(new_n8945_));
  OAI21_X1   g08688(.A1(new_n8945_), .A2(new_n8943_), .B(new_n8542_), .ZN(new_n8946_));
  NAND2_X1   g08689(.A1(new_n8942_), .A2(new_n8946_), .ZN(new_n8947_));
  XNOR2_X1   g08690(.A1(new_n8947_), .A2(new_n8583_), .ZN(new_n8948_));
  INV_X1     g08691(.I(new_n8947_), .ZN(new_n8949_));
  OR2_X2     g08692(.A1(new_n8949_), .A2(new_n8583_), .Z(new_n8950_));
  NAND2_X1   g08693(.A1(new_n8949_), .A2(new_n8583_), .ZN(new_n8951_));
  NAND2_X1   g08694(.A1(new_n8950_), .A2(new_n8951_), .ZN(new_n8952_));
  MUX2_X1    g08695(.I0(new_n8952_), .I1(new_n8948_), .S(new_n8581_), .Z(\f[62] ));
  NAND2_X1   g08696(.A1(new_n8930_), .A2(new_n8931_), .ZN(new_n8954_));
  NAND2_X1   g08697(.A1(new_n8954_), .A2(new_n8933_), .ZN(new_n8955_));
  INV_X1     g08698(.I(\b[63] ), .ZN(new_n8956_));
  NOR2_X1    g08699(.A1(new_n8956_), .A2(\b[62] ), .ZN(new_n8957_));
  NOR2_X1    g08700(.A1(new_n8932_), .A2(\b[63] ), .ZN(new_n8958_));
  OR2_X2     g08701(.A1(new_n8957_), .A2(new_n8958_), .Z(new_n8959_));
  XOR2_X1    g08702(.A1(\b[62] ), .A2(\b[63] ), .Z(new_n8960_));
  NOR2_X1    g08703(.A1(new_n8955_), .A2(new_n8960_), .ZN(new_n8961_));
  AOI21_X1   g08704(.A1(new_n8955_), .A2(new_n8959_), .B(new_n8961_), .ZN(new_n8962_));
  INV_X1     g08705(.I(new_n8962_), .ZN(new_n8963_));
  NOR2_X1    g08706(.A1(new_n405_), .A2(new_n8956_), .ZN(new_n8964_));
  NOR2_X1    g08707(.A1(new_n280_), .A2(new_n8548_), .ZN(new_n8965_));
  NOR2_X1    g08708(.A1(new_n404_), .A2(new_n8932_), .ZN(new_n8966_));
  NOR4_X1    g08709(.A1(new_n8964_), .A2(new_n264_), .A3(new_n8965_), .A4(new_n8966_), .ZN(new_n8967_));
  NAND2_X1   g08710(.A1(new_n8963_), .A2(new_n8967_), .ZN(new_n8968_));
  XOR2_X1    g08711(.A1(new_n8968_), .A2(\a[2] ), .Z(new_n8969_));
  OAI22_X1   g08712(.A1(new_n364_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n320_), .ZN(new_n8970_));
  NAND2_X1   g08713(.A1(new_n594_), .A2(\b[58] ), .ZN(new_n8971_));
  AOI21_X1   g08714(.A1(new_n8970_), .A2(new_n8971_), .B(new_n312_), .ZN(new_n8972_));
  NAND2_X1   g08715(.A1(new_n7929_), .A2(new_n8972_), .ZN(new_n8973_));
  XOR2_X1    g08716(.A1(new_n8973_), .A2(new_n308_), .Z(new_n8974_));
  AOI21_X1   g08717(.A1(new_n8585_), .A2(new_n8844_), .B(new_n8828_), .ZN(new_n8975_));
  INV_X1     g08718(.I(new_n8650_), .ZN(new_n8976_));
  OAI21_X1   g08719(.A1(new_n8613_), .A2(new_n8651_), .B(new_n8976_), .ZN(new_n8977_));
  INV_X1     g08720(.I(new_n8977_), .ZN(new_n8978_));
  NAND2_X1   g08721(.A1(new_n8639_), .A2(new_n8637_), .ZN(new_n8979_));
  NAND2_X1   g08722(.A1(new_n8635_), .A2(new_n8616_), .ZN(new_n8980_));
  OAI22_X1   g08723(.A1(new_n290_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n292_), .ZN(new_n8981_));
  OAI21_X1   g08724(.A1(new_n267_), .A2(new_n8622_), .B(new_n8981_), .ZN(new_n8982_));
  NAND3_X1   g08725(.A1(new_n8982_), .A2(new_n298_), .A3(new_n8320_), .ZN(new_n8983_));
  XOR2_X1    g08726(.A1(new_n8983_), .A2(new_n8309_), .Z(new_n8984_));
  XNOR2_X1   g08727(.A1(\a[62] ), .A2(\a[63] ), .ZN(new_n8985_));
  NOR2_X1    g08728(.A1(new_n8985_), .A2(new_n258_), .ZN(new_n8986_));
  XOR2_X1    g08729(.A1(new_n8984_), .A2(new_n8986_), .Z(new_n8987_));
  NOR2_X1    g08730(.A1(new_n8987_), .A2(new_n8980_), .ZN(new_n8988_));
  XOR2_X1    g08731(.A1(new_n8983_), .A2(\a[62] ), .Z(new_n8989_));
  NAND2_X1   g08732(.A1(new_n8989_), .A2(new_n8986_), .ZN(new_n8990_));
  OAI21_X1   g08733(.A1(new_n258_), .A2(new_n8985_), .B(new_n8984_), .ZN(new_n8991_));
  AOI22_X1   g08734(.A1(new_n8990_), .A2(new_n8991_), .B1(new_n8616_), .B2(new_n8635_), .ZN(new_n8992_));
  NOR2_X1    g08735(.A1(new_n8988_), .A2(new_n8992_), .ZN(new_n8993_));
  NOR2_X1    g08736(.A1(new_n7351_), .A2(new_n347_), .ZN(new_n8994_));
  NOR2_X1    g08737(.A1(new_n7346_), .A2(new_n403_), .ZN(new_n8995_));
  OAI22_X1   g08738(.A1(new_n8994_), .A2(new_n8995_), .B1(new_n7611_), .B2(new_n393_), .ZN(new_n8996_));
  AND3_X2    g08739(.A1(new_n402_), .A2(new_n7604_), .A3(new_n8996_), .Z(new_n8997_));
  XOR2_X1    g08740(.A1(new_n8997_), .A2(\a[59] ), .Z(new_n8998_));
  NAND2_X1   g08741(.A1(new_n8993_), .A2(new_n8998_), .ZN(new_n8999_));
  INV_X1     g08742(.I(new_n8993_), .ZN(new_n9000_));
  INV_X1     g08743(.I(new_n8998_), .ZN(new_n9001_));
  NAND2_X1   g08744(.A1(new_n9000_), .A2(new_n9001_), .ZN(new_n9002_));
  AOI22_X1   g08745(.A1(new_n9002_), .A2(new_n8999_), .B1(new_n8634_), .B2(new_n8979_), .ZN(new_n9003_));
  NAND2_X1   g08746(.A1(new_n8979_), .A2(new_n8634_), .ZN(new_n9004_));
  NAND2_X1   g08747(.A1(new_n9000_), .A2(new_n8998_), .ZN(new_n9005_));
  NAND2_X1   g08748(.A1(new_n8993_), .A2(new_n9001_), .ZN(new_n9006_));
  AOI21_X1   g08749(.A1(new_n9005_), .A2(new_n9006_), .B(new_n9004_), .ZN(new_n9007_));
  NOR2_X1    g08750(.A1(new_n9003_), .A2(new_n9007_), .ZN(new_n9008_));
  INV_X1     g08751(.I(new_n9008_), .ZN(new_n9009_));
  OAI22_X1   g08752(.A1(new_n6721_), .A2(new_n495_), .B1(new_n6723_), .B2(new_n510_), .ZN(new_n9010_));
  NAND2_X1   g08753(.A1(new_n7617_), .A2(\b[7] ), .ZN(new_n9011_));
  AOI21_X1   g08754(.A1(new_n9011_), .A2(new_n9010_), .B(new_n6731_), .ZN(new_n9012_));
  NAND2_X1   g08755(.A1(new_n518_), .A2(new_n9012_), .ZN(new_n9013_));
  XOR2_X1    g08756(.A1(new_n9013_), .A2(\a[56] ), .Z(new_n9014_));
  NOR2_X1    g08757(.A1(new_n9009_), .A2(new_n9014_), .ZN(new_n9015_));
  INV_X1     g08758(.I(new_n9015_), .ZN(new_n9016_));
  NAND2_X1   g08759(.A1(new_n9009_), .A2(new_n9014_), .ZN(new_n9017_));
  AOI21_X1   g08760(.A1(new_n9016_), .A2(new_n9017_), .B(new_n8978_), .ZN(new_n9018_));
  XOR2_X1    g08761(.A1(new_n9008_), .A2(new_n9014_), .Z(new_n9019_));
  NOR2_X1    g08762(.A1(new_n9019_), .A2(new_n8977_), .ZN(new_n9020_));
  NOR2_X1    g08763(.A1(new_n9018_), .A2(new_n9020_), .ZN(new_n9021_));
  INV_X1     g08764(.I(new_n9021_), .ZN(new_n9022_));
  OAI22_X1   g08765(.A1(new_n5786_), .A2(new_n717_), .B1(new_n659_), .B2(new_n5792_), .ZN(new_n9023_));
  NAND2_X1   g08766(.A1(new_n6745_), .A2(\b[10] ), .ZN(new_n9024_));
  AOI21_X1   g08767(.A1(new_n9024_), .A2(new_n9023_), .B(new_n5796_), .ZN(new_n9025_));
  NAND2_X1   g08768(.A1(new_n716_), .A2(new_n9025_), .ZN(new_n9026_));
  XOR2_X1    g08769(.A1(new_n9026_), .A2(\a[53] ), .Z(new_n9027_));
  NAND2_X1   g08770(.A1(new_n8649_), .A2(new_n8652_), .ZN(new_n9028_));
  NAND2_X1   g08771(.A1(new_n9028_), .A2(new_n8657_), .ZN(new_n9029_));
  OAI21_X1   g08772(.A1(new_n8663_), .A2(new_n8661_), .B(new_n9029_), .ZN(new_n9030_));
  NAND2_X1   g08773(.A1(new_n9030_), .A2(new_n9027_), .ZN(new_n9031_));
  INV_X1     g08774(.I(new_n9027_), .ZN(new_n9032_));
  NAND2_X1   g08775(.A1(new_n8612_), .A2(new_n8665_), .ZN(new_n9033_));
  NAND3_X1   g08776(.A1(new_n9033_), .A2(new_n9032_), .A3(new_n9029_), .ZN(new_n9034_));
  AOI21_X1   g08777(.A1(new_n9031_), .A2(new_n9034_), .B(new_n9022_), .ZN(new_n9035_));
  AOI21_X1   g08778(.A1(new_n9033_), .A2(new_n9029_), .B(new_n9032_), .ZN(new_n9036_));
  NOR2_X1    g08779(.A1(new_n9030_), .A2(new_n9027_), .ZN(new_n9037_));
  NOR3_X1    g08780(.A1(new_n9037_), .A2(new_n9036_), .A3(new_n9021_), .ZN(new_n9038_));
  NOR2_X1    g08781(.A1(new_n9038_), .A2(new_n9035_), .ZN(new_n9039_));
  OAI22_X1   g08782(.A1(new_n5228_), .A2(new_n904_), .B1(new_n848_), .B2(new_n5225_), .ZN(new_n9040_));
  NAND2_X1   g08783(.A1(new_n5387_), .A2(\b[13] ), .ZN(new_n9041_));
  AOI21_X1   g08784(.A1(new_n9040_), .A2(new_n9041_), .B(new_n5231_), .ZN(new_n9042_));
  NAND2_X1   g08785(.A1(new_n907_), .A2(new_n9042_), .ZN(new_n9043_));
  XOR2_X1    g08786(.A1(new_n9043_), .A2(\a[50] ), .Z(new_n9044_));
  INV_X1     g08787(.I(new_n9044_), .ZN(new_n9045_));
  NAND3_X1   g08788(.A1(new_n8685_), .A2(new_n8684_), .A3(new_n8610_), .ZN(new_n9046_));
  AOI21_X1   g08789(.A1(new_n9046_), .A2(new_n8685_), .B(new_n9045_), .ZN(new_n9047_));
  OAI21_X1   g08790(.A1(new_n8609_), .A2(new_n8672_), .B(new_n8685_), .ZN(new_n9048_));
  NOR2_X1    g08791(.A1(new_n9048_), .A2(new_n9044_), .ZN(new_n9049_));
  OAI21_X1   g08792(.A1(new_n9047_), .A2(new_n9049_), .B(new_n9039_), .ZN(new_n9050_));
  OAI21_X1   g08793(.A1(new_n9037_), .A2(new_n9036_), .B(new_n9021_), .ZN(new_n9051_));
  NAND3_X1   g08794(.A1(new_n9031_), .A2(new_n9034_), .A3(new_n9022_), .ZN(new_n9052_));
  NAND2_X1   g08795(.A1(new_n9051_), .A2(new_n9052_), .ZN(new_n9053_));
  NAND2_X1   g08796(.A1(new_n9048_), .A2(new_n9044_), .ZN(new_n9054_));
  NAND3_X1   g08797(.A1(new_n9046_), .A2(new_n8685_), .A3(new_n9045_), .ZN(new_n9055_));
  NAND3_X1   g08798(.A1(new_n9055_), .A2(new_n9054_), .A3(new_n9053_), .ZN(new_n9056_));
  NAND2_X1   g08799(.A1(new_n9050_), .A2(new_n9056_), .ZN(new_n9057_));
  NOR3_X1    g08800(.A1(new_n8687_), .A2(new_n8690_), .A3(new_n8608_), .ZN(new_n9058_));
  OAI22_X1   g08801(.A1(new_n4711_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n4706_), .ZN(new_n9059_));
  NAND2_X1   g08802(.A1(new_n5814_), .A2(\b[16] ), .ZN(new_n9060_));
  AOI21_X1   g08803(.A1(new_n9059_), .A2(new_n9060_), .B(new_n4714_), .ZN(new_n9061_));
  NAND2_X1   g08804(.A1(new_n1123_), .A2(new_n9061_), .ZN(new_n9062_));
  XOR2_X1    g08805(.A1(new_n9062_), .A2(\a[47] ), .Z(new_n9063_));
  OAI21_X1   g08806(.A1(new_n8676_), .A2(new_n8672_), .B(new_n8610_), .ZN(new_n9064_));
  NAND3_X1   g08807(.A1(new_n8685_), .A2(new_n8684_), .A3(new_n8609_), .ZN(new_n9065_));
  AOI21_X1   g08808(.A1(new_n9064_), .A2(new_n9065_), .B(new_n8682_), .ZN(new_n9066_));
  OAI21_X1   g08809(.A1(new_n9058_), .A2(new_n9066_), .B(new_n9063_), .ZN(new_n9067_));
  INV_X1     g08810(.I(new_n9063_), .ZN(new_n9068_));
  INV_X1     g08811(.I(new_n9066_), .ZN(new_n9069_));
  NAND3_X1   g08812(.A1(new_n8698_), .A2(new_n9068_), .A3(new_n9069_), .ZN(new_n9070_));
  AOI21_X1   g08813(.A1(new_n9067_), .A2(new_n9070_), .B(new_n9057_), .ZN(new_n9071_));
  AOI21_X1   g08814(.A1(new_n9055_), .A2(new_n9054_), .B(new_n9053_), .ZN(new_n9072_));
  NOR3_X1    g08815(.A1(new_n9047_), .A2(new_n9049_), .A3(new_n9039_), .ZN(new_n9073_));
  NOR2_X1    g08816(.A1(new_n9073_), .A2(new_n9072_), .ZN(new_n9074_));
  AOI21_X1   g08817(.A1(new_n8698_), .A2(new_n9069_), .B(new_n9068_), .ZN(new_n9075_));
  NOR3_X1    g08818(.A1(new_n9058_), .A2(new_n9063_), .A3(new_n9066_), .ZN(new_n9076_));
  NOR3_X1    g08819(.A1(new_n9075_), .A2(new_n9076_), .A3(new_n9074_), .ZN(new_n9077_));
  OAI22_X1   g08820(.A1(new_n4208_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n4203_), .ZN(new_n9078_));
  NAND2_X1   g08821(.A1(new_n5244_), .A2(\b[19] ), .ZN(new_n9079_));
  AOI21_X1   g08822(.A1(new_n9078_), .A2(new_n9079_), .B(new_n4211_), .ZN(new_n9080_));
  NAND2_X1   g08823(.A1(new_n1396_), .A2(new_n9080_), .ZN(new_n9081_));
  XOR2_X1    g08824(.A1(new_n9081_), .A2(\a[44] ), .Z(new_n9082_));
  INV_X1     g08825(.I(new_n9082_), .ZN(new_n9083_));
  OAI21_X1   g08826(.A1(new_n9071_), .A2(new_n9077_), .B(new_n9083_), .ZN(new_n9084_));
  OAI21_X1   g08827(.A1(new_n9075_), .A2(new_n9076_), .B(new_n9074_), .ZN(new_n9085_));
  NAND3_X1   g08828(.A1(new_n9067_), .A2(new_n9070_), .A3(new_n9057_), .ZN(new_n9086_));
  NAND3_X1   g08829(.A1(new_n9085_), .A2(new_n9086_), .A3(new_n9082_), .ZN(new_n9087_));
  AOI21_X1   g08830(.A1(new_n9084_), .A2(new_n9087_), .B(new_n8705_), .ZN(new_n9088_));
  NAND3_X1   g08831(.A1(new_n9085_), .A2(new_n9086_), .A3(new_n9083_), .ZN(new_n9089_));
  OAI21_X1   g08832(.A1(new_n9077_), .A2(new_n9071_), .B(new_n9082_), .ZN(new_n9090_));
  AOI21_X1   g08833(.A1(new_n9090_), .A2(new_n9089_), .B(new_n8704_), .ZN(new_n9091_));
  NOR2_X1    g08834(.A1(new_n9088_), .A2(new_n9091_), .ZN(new_n9092_));
  INV_X1     g08835(.I(new_n9092_), .ZN(new_n9093_));
  OAI22_X1   g08836(.A1(new_n3736_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n3731_), .ZN(new_n9094_));
  NAND2_X1   g08837(.A1(new_n4730_), .A2(\b[22] ), .ZN(new_n9095_));
  AOI21_X1   g08838(.A1(new_n9094_), .A2(new_n9095_), .B(new_n3739_), .ZN(new_n9096_));
  NAND2_X1   g08839(.A1(new_n1708_), .A2(new_n9096_), .ZN(new_n9097_));
  XOR2_X1    g08840(.A1(new_n9097_), .A2(\a[41] ), .Z(new_n9098_));
  AOI21_X1   g08841(.A1(new_n8705_), .A2(new_n8706_), .B(new_n8714_), .ZN(new_n9099_));
  NOR3_X1    g08842(.A1(new_n8607_), .A2(new_n8406_), .A3(new_n8716_), .ZN(new_n9100_));
  OAI21_X1   g08843(.A1(new_n9100_), .A2(new_n9099_), .B(new_n9098_), .ZN(new_n9101_));
  INV_X1     g08844(.I(new_n9098_), .ZN(new_n9102_));
  INV_X1     g08845(.I(new_n9099_), .ZN(new_n9103_));
  NAND3_X1   g08846(.A1(new_n8720_), .A2(new_n8412_), .A3(new_n8717_), .ZN(new_n9104_));
  NAND3_X1   g08847(.A1(new_n9104_), .A2(new_n9102_), .A3(new_n9103_), .ZN(new_n9105_));
  AOI21_X1   g08848(.A1(new_n9101_), .A2(new_n9105_), .B(new_n9093_), .ZN(new_n9106_));
  AOI21_X1   g08849(.A1(new_n9104_), .A2(new_n9103_), .B(new_n9102_), .ZN(new_n9107_));
  NOR3_X1    g08850(.A1(new_n9100_), .A2(new_n9098_), .A3(new_n9099_), .ZN(new_n9108_));
  NOR3_X1    g08851(.A1(new_n9108_), .A2(new_n9107_), .A3(new_n9092_), .ZN(new_n9109_));
  NOR2_X1    g08852(.A1(new_n9109_), .A2(new_n9106_), .ZN(new_n9110_));
  INV_X1     g08853(.I(new_n9110_), .ZN(new_n9111_));
  NOR2_X1    g08854(.A1(new_n8736_), .A2(new_n8735_), .ZN(new_n9112_));
  OAI22_X1   g08855(.A1(new_n3298_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n3293_), .ZN(new_n9113_));
  NAND2_X1   g08856(.A1(new_n4227_), .A2(\b[25] ), .ZN(new_n9114_));
  AOI21_X1   g08857(.A1(new_n9113_), .A2(new_n9114_), .B(new_n3301_), .ZN(new_n9115_));
  NAND2_X1   g08858(.A1(new_n2042_), .A2(new_n9115_), .ZN(new_n9116_));
  XOR2_X1    g08859(.A1(new_n9116_), .A2(\a[38] ), .Z(new_n9117_));
  NOR2_X1    g08860(.A1(new_n8738_), .A2(new_n8739_), .ZN(new_n9118_));
  INV_X1     g08861(.I(new_n9118_), .ZN(new_n9119_));
  OAI21_X1   g08862(.A1(new_n9112_), .A2(new_n9119_), .B(new_n9117_), .ZN(new_n9120_));
  NAND2_X1   g08863(.A1(new_n8742_), .A2(new_n8741_), .ZN(new_n9121_));
  INV_X1     g08864(.I(new_n9117_), .ZN(new_n9122_));
  NAND3_X1   g08865(.A1(new_n9121_), .A2(new_n9118_), .A3(new_n9122_), .ZN(new_n9123_));
  AOI21_X1   g08866(.A1(new_n9120_), .A2(new_n9123_), .B(new_n9111_), .ZN(new_n9124_));
  AOI21_X1   g08867(.A1(new_n9121_), .A2(new_n9118_), .B(new_n9122_), .ZN(new_n9125_));
  NOR3_X1    g08868(.A1(new_n9112_), .A2(new_n9119_), .A3(new_n9117_), .ZN(new_n9126_));
  NOR3_X1    g08869(.A1(new_n9126_), .A2(new_n9125_), .A3(new_n9110_), .ZN(new_n9127_));
  NOR2_X1    g08870(.A1(new_n9127_), .A2(new_n9124_), .ZN(new_n9128_));
  OAI22_X1   g08871(.A1(new_n2846_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n2841_), .ZN(new_n9129_));
  NAND2_X1   g08872(.A1(new_n3755_), .A2(\b[28] ), .ZN(new_n9130_));
  AOI21_X1   g08873(.A1(new_n9129_), .A2(new_n9130_), .B(new_n2849_), .ZN(new_n9131_));
  NAND2_X1   g08874(.A1(new_n2404_), .A2(new_n9131_), .ZN(new_n9132_));
  XOR2_X1    g08875(.A1(new_n9132_), .A2(\a[35] ), .Z(new_n9133_));
  INV_X1     g08876(.I(new_n9133_), .ZN(new_n9134_));
  NOR3_X1    g08877(.A1(new_n8770_), .A2(new_n8749_), .A3(new_n8753_), .ZN(new_n9135_));
  NOR2_X1    g08878(.A1(new_n9135_), .A2(new_n9134_), .ZN(new_n9136_));
  NAND4_X1   g08879(.A1(new_n8757_), .A2(new_n8760_), .A3(new_n8759_), .A4(new_n9134_), .ZN(new_n9137_));
  INV_X1     g08880(.I(new_n9137_), .ZN(new_n9138_));
  OAI21_X1   g08881(.A1(new_n9136_), .A2(new_n9138_), .B(new_n9128_), .ZN(new_n9139_));
  OAI21_X1   g08882(.A1(new_n9126_), .A2(new_n9125_), .B(new_n9110_), .ZN(new_n9140_));
  NAND3_X1   g08883(.A1(new_n9120_), .A2(new_n9123_), .A3(new_n9111_), .ZN(new_n9141_));
  NAND2_X1   g08884(.A1(new_n9140_), .A2(new_n9141_), .ZN(new_n9142_));
  NAND3_X1   g08885(.A1(new_n8757_), .A2(new_n8760_), .A3(new_n8759_), .ZN(new_n9143_));
  NAND2_X1   g08886(.A1(new_n9143_), .A2(new_n9133_), .ZN(new_n9144_));
  NAND3_X1   g08887(.A1(new_n9144_), .A2(new_n9142_), .A3(new_n9137_), .ZN(new_n9145_));
  OAI22_X1   g08888(.A1(new_n2452_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n2447_), .ZN(new_n9146_));
  NAND2_X1   g08889(.A1(new_n3312_), .A2(\b[31] ), .ZN(new_n9147_));
  AOI21_X1   g08890(.A1(new_n9146_), .A2(new_n9147_), .B(new_n2455_), .ZN(new_n9148_));
  NAND2_X1   g08891(.A1(new_n2797_), .A2(new_n9148_), .ZN(new_n9149_));
  XOR2_X1    g08892(.A1(new_n9149_), .A2(\a[32] ), .Z(new_n9150_));
  INV_X1     g08893(.I(new_n9150_), .ZN(new_n9151_));
  NAND3_X1   g08894(.A1(new_n9139_), .A2(new_n9145_), .A3(new_n9151_), .ZN(new_n9152_));
  AOI21_X1   g08895(.A1(new_n9144_), .A2(new_n9137_), .B(new_n9142_), .ZN(new_n9153_));
  NOR3_X1    g08896(.A1(new_n9136_), .A2(new_n9138_), .A3(new_n9128_), .ZN(new_n9154_));
  OAI21_X1   g08897(.A1(new_n9154_), .A2(new_n9153_), .B(new_n9150_), .ZN(new_n9155_));
  NAND2_X1   g08898(.A1(new_n9155_), .A2(new_n9152_), .ZN(new_n9156_));
  INV_X1     g08899(.I(new_n9156_), .ZN(new_n9157_));
  OAI22_X1   g08900(.A1(new_n2084_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n2079_), .ZN(new_n9158_));
  NAND2_X1   g08901(.A1(new_n2864_), .A2(\b[34] ), .ZN(new_n9159_));
  AOI21_X1   g08902(.A1(new_n9158_), .A2(new_n9159_), .B(new_n2087_), .ZN(new_n9160_));
  NAND2_X1   g08903(.A1(new_n3246_), .A2(new_n9160_), .ZN(new_n9161_));
  XOR2_X1    g08904(.A1(new_n9161_), .A2(\a[29] ), .Z(new_n9162_));
  AOI21_X1   g08905(.A1(new_n8775_), .A2(new_n8774_), .B(new_n8778_), .ZN(new_n9163_));
  INV_X1     g08906(.I(new_n9163_), .ZN(new_n9164_));
  AOI21_X1   g08907(.A1(new_n8775_), .A2(new_n8774_), .B(new_n8605_), .ZN(new_n9165_));
  NOR3_X1    g08908(.A1(new_n8771_), .A2(new_n8758_), .A3(new_n8778_), .ZN(new_n9166_));
  OAI21_X1   g08909(.A1(new_n9166_), .A2(new_n9165_), .B(new_n8459_), .ZN(new_n9167_));
  NAND2_X1   g08910(.A1(new_n9167_), .A2(new_n9164_), .ZN(new_n9168_));
  NAND2_X1   g08911(.A1(new_n9168_), .A2(new_n9162_), .ZN(new_n9169_));
  INV_X1     g08912(.I(new_n9162_), .ZN(new_n9170_));
  OAI21_X1   g08913(.A1(new_n8771_), .A2(new_n8758_), .B(new_n8778_), .ZN(new_n9171_));
  NAND3_X1   g08914(.A1(new_n8775_), .A2(new_n8774_), .A3(new_n8605_), .ZN(new_n9172_));
  NAND2_X1   g08915(.A1(new_n9171_), .A2(new_n9172_), .ZN(new_n9173_));
  AOI21_X1   g08916(.A1(new_n9173_), .A2(new_n8459_), .B(new_n9163_), .ZN(new_n9174_));
  NAND2_X1   g08917(.A1(new_n9174_), .A2(new_n9170_), .ZN(new_n9175_));
  NAND2_X1   g08918(.A1(new_n9169_), .A2(new_n9175_), .ZN(new_n9176_));
  NAND2_X1   g08919(.A1(new_n9176_), .A2(new_n9157_), .ZN(new_n9177_));
  NAND3_X1   g08920(.A1(new_n9169_), .A2(new_n9175_), .A3(new_n9156_), .ZN(new_n9178_));
  NAND2_X1   g08921(.A1(new_n8775_), .A2(new_n8774_), .ZN(new_n9179_));
  NOR2_X1    g08922(.A1(new_n8773_), .A2(new_n8605_), .ZN(new_n9180_));
  NOR2_X1    g08923(.A1(new_n8459_), .A2(new_n8778_), .ZN(new_n9181_));
  NOR2_X1    g08924(.A1(new_n9180_), .A2(new_n9181_), .ZN(new_n9182_));
  NOR2_X1    g08925(.A1(new_n9182_), .A2(new_n9179_), .ZN(new_n9183_));
  NAND2_X1   g08926(.A1(new_n9182_), .A2(new_n9179_), .ZN(new_n9184_));
  INV_X1     g08927(.I(new_n9184_), .ZN(new_n9185_));
  OAI21_X1   g08928(.A1(new_n9185_), .A2(new_n9183_), .B(new_n8599_), .ZN(new_n9186_));
  NAND4_X1   g08929(.A1(new_n9186_), .A2(new_n8787_), .A3(new_n8788_), .A4(new_n8474_), .ZN(new_n9187_));
  NAND3_X1   g08930(.A1(new_n9177_), .A2(new_n9178_), .A3(new_n9187_), .ZN(new_n9188_));
  AOI21_X1   g08931(.A1(new_n9169_), .A2(new_n9175_), .B(new_n9156_), .ZN(new_n9189_));
  INV_X1     g08932(.I(new_n9178_), .ZN(new_n9190_));
  INV_X1     g08933(.I(new_n9183_), .ZN(new_n9191_));
  AOI21_X1   g08934(.A1(new_n9191_), .A2(new_n9184_), .B(new_n8600_), .ZN(new_n9192_));
  NOR4_X1    g08935(.A1(new_n9192_), .A2(new_n8782_), .A3(new_n8785_), .A4(new_n8473_), .ZN(new_n9193_));
  OAI21_X1   g08936(.A1(new_n9190_), .A2(new_n9189_), .B(new_n9193_), .ZN(new_n9194_));
  NAND2_X1   g08937(.A1(new_n9194_), .A2(new_n9188_), .ZN(new_n9195_));
  OAI22_X1   g08938(.A1(new_n1760_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n1755_), .ZN(new_n9196_));
  NAND2_X1   g08939(.A1(new_n2470_), .A2(\b[37] ), .ZN(new_n9197_));
  AOI21_X1   g08940(.A1(new_n9196_), .A2(new_n9197_), .B(new_n1763_), .ZN(new_n9198_));
  NAND2_X1   g08941(.A1(new_n3700_), .A2(new_n9198_), .ZN(new_n9199_));
  XOR2_X1    g08942(.A1(new_n9199_), .A2(\a[26] ), .Z(new_n9200_));
  INV_X1     g08943(.I(new_n9200_), .ZN(new_n9201_));
  NOR2_X1    g08944(.A1(new_n8795_), .A2(new_n8799_), .ZN(new_n9202_));
  AOI21_X1   g08945(.A1(new_n9202_), .A2(new_n8801_), .B(new_n9201_), .ZN(new_n9203_));
  INV_X1     g08946(.I(new_n9203_), .ZN(new_n9204_));
  NAND3_X1   g08947(.A1(new_n9202_), .A2(new_n8801_), .A3(new_n9201_), .ZN(new_n9205_));
  AOI21_X1   g08948(.A1(new_n9204_), .A2(new_n9205_), .B(new_n9195_), .ZN(new_n9206_));
  AND2_X2    g08949(.A1(new_n9194_), .A2(new_n9188_), .Z(new_n9207_));
  INV_X1     g08950(.I(new_n9205_), .ZN(new_n9208_));
  NOR3_X1    g08951(.A1(new_n9208_), .A2(new_n9207_), .A3(new_n9203_), .ZN(new_n9209_));
  NOR2_X1    g08952(.A1(new_n9209_), .A2(new_n9206_), .ZN(new_n9210_));
  OAI22_X1   g08953(.A1(new_n1444_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n1439_), .ZN(new_n9211_));
  NAND2_X1   g08954(.A1(new_n2098_), .A2(\b[40] ), .ZN(new_n9212_));
  AOI21_X1   g08955(.A1(new_n9211_), .A2(new_n9212_), .B(new_n1447_), .ZN(new_n9213_));
  NAND2_X1   g08956(.A1(new_n4017_), .A2(new_n9213_), .ZN(new_n9214_));
  XOR2_X1    g08957(.A1(new_n9214_), .A2(\a[23] ), .Z(new_n9215_));
  INV_X1     g08958(.I(new_n9215_), .ZN(new_n9216_));
  AOI21_X1   g08959(.A1(new_n8822_), .A2(new_n8830_), .B(new_n9216_), .ZN(new_n9217_));
  NOR3_X1    g08960(.A1(new_n8834_), .A2(new_n8817_), .A3(new_n9215_), .ZN(new_n9218_));
  OAI21_X1   g08961(.A1(new_n9217_), .A2(new_n9218_), .B(new_n9210_), .ZN(new_n9219_));
  OAI21_X1   g08962(.A1(new_n9203_), .A2(new_n9208_), .B(new_n9207_), .ZN(new_n9220_));
  NAND3_X1   g08963(.A1(new_n9204_), .A2(new_n9195_), .A3(new_n9205_), .ZN(new_n9221_));
  NAND2_X1   g08964(.A1(new_n9220_), .A2(new_n9221_), .ZN(new_n9222_));
  OAI21_X1   g08965(.A1(new_n8834_), .A2(new_n8817_), .B(new_n9215_), .ZN(new_n9223_));
  NAND3_X1   g08966(.A1(new_n8822_), .A2(new_n8830_), .A3(new_n9216_), .ZN(new_n9224_));
  NAND3_X1   g08967(.A1(new_n9224_), .A2(new_n9223_), .A3(new_n9222_), .ZN(new_n9225_));
  NAND2_X1   g08968(.A1(new_n9219_), .A2(new_n9225_), .ZN(new_n9226_));
  OAI22_X1   g08969(.A1(new_n1168_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n1163_), .ZN(new_n9227_));
  NAND2_X1   g08970(.A1(new_n1774_), .A2(\b[43] ), .ZN(new_n9228_));
  AOI21_X1   g08971(.A1(new_n9227_), .A2(new_n9228_), .B(new_n1171_), .ZN(new_n9229_));
  NAND2_X1   g08972(.A1(new_n4513_), .A2(new_n9229_), .ZN(new_n9230_));
  XOR2_X1    g08973(.A1(new_n9230_), .A2(\a[20] ), .Z(new_n9231_));
  INV_X1     g08974(.I(new_n9231_), .ZN(new_n9232_));
  NAND2_X1   g08975(.A1(new_n9226_), .A2(new_n9232_), .ZN(new_n9233_));
  NAND3_X1   g08976(.A1(new_n9219_), .A2(new_n9225_), .A3(new_n9231_), .ZN(new_n9234_));
  AOI21_X1   g08977(.A1(new_n9233_), .A2(new_n9234_), .B(new_n8975_), .ZN(new_n9235_));
  INV_X1     g08978(.I(new_n8975_), .ZN(new_n9236_));
  NAND3_X1   g08979(.A1(new_n9219_), .A2(new_n9225_), .A3(new_n9232_), .ZN(new_n9237_));
  AOI21_X1   g08980(.A1(new_n9224_), .A2(new_n9223_), .B(new_n9222_), .ZN(new_n9238_));
  NOR3_X1    g08981(.A1(new_n9217_), .A2(new_n9218_), .A3(new_n9210_), .ZN(new_n9239_));
  OAI21_X1   g08982(.A1(new_n9238_), .A2(new_n9239_), .B(new_n9231_), .ZN(new_n9240_));
  AOI21_X1   g08983(.A1(new_n9240_), .A2(new_n9237_), .B(new_n9236_), .ZN(new_n9241_));
  NOR2_X1    g08984(.A1(new_n9235_), .A2(new_n9241_), .ZN(new_n9242_));
  INV_X1     g08985(.I(new_n9242_), .ZN(new_n9243_));
  OAI22_X1   g08986(.A1(new_n940_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n935_), .ZN(new_n9244_));
  NAND2_X1   g08987(.A1(new_n1458_), .A2(\b[46] ), .ZN(new_n9245_));
  AOI21_X1   g08988(.A1(new_n9244_), .A2(new_n9245_), .B(new_n943_), .ZN(new_n9246_));
  NAND2_X1   g08989(.A1(new_n5177_), .A2(new_n9246_), .ZN(new_n9247_));
  XOR2_X1    g08990(.A1(new_n9247_), .A2(\a[17] ), .Z(new_n9248_));
  NOR2_X1    g08991(.A1(new_n8857_), .A2(new_n8860_), .ZN(new_n9249_));
  AOI21_X1   g08992(.A1(new_n8290_), .A2(new_n8852_), .B(new_n8508_), .ZN(new_n9250_));
  AOI21_X1   g08993(.A1(new_n9249_), .A2(new_n9250_), .B(new_n8861_), .ZN(new_n9251_));
  OAI21_X1   g08994(.A1(new_n8828_), .A2(new_n8836_), .B(new_n8848_), .ZN(new_n9252_));
  NAND3_X1   g08995(.A1(new_n8843_), .A2(new_n8844_), .A3(new_n8585_), .ZN(new_n9253_));
  AOI21_X1   g08996(.A1(new_n9252_), .A2(new_n9253_), .B(new_n8845_), .ZN(new_n9254_));
  OAI21_X1   g08997(.A1(new_n9251_), .A2(new_n9254_), .B(new_n9248_), .ZN(new_n9255_));
  INV_X1     g08998(.I(new_n9248_), .ZN(new_n9256_));
  NAND2_X1   g08999(.A1(new_n8847_), .A2(new_n8851_), .ZN(new_n9257_));
  OAI21_X1   g09000(.A1(new_n8512_), .A2(new_n8503_), .B(new_n8513_), .ZN(new_n9258_));
  OAI21_X1   g09001(.A1(new_n9257_), .A2(new_n9258_), .B(new_n8853_), .ZN(new_n9259_));
  INV_X1     g09002(.I(new_n9254_), .ZN(new_n9260_));
  NAND3_X1   g09003(.A1(new_n9259_), .A2(new_n9256_), .A3(new_n9260_), .ZN(new_n9261_));
  AOI21_X1   g09004(.A1(new_n9255_), .A2(new_n9261_), .B(new_n9243_), .ZN(new_n9262_));
  AOI21_X1   g09005(.A1(new_n9259_), .A2(new_n9260_), .B(new_n9256_), .ZN(new_n9263_));
  NOR3_X1    g09006(.A1(new_n9251_), .A2(new_n9248_), .A3(new_n9254_), .ZN(new_n9264_));
  NOR3_X1    g09007(.A1(new_n9264_), .A2(new_n9263_), .A3(new_n9242_), .ZN(new_n9265_));
  NOR2_X1    g09008(.A1(new_n9262_), .A2(new_n9265_), .ZN(new_n9266_));
  OAI22_X1   g09009(.A1(new_n757_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n752_), .ZN(new_n9267_));
  NAND2_X1   g09010(.A1(new_n1182_), .A2(\b[49] ), .ZN(new_n9268_));
  AOI21_X1   g09011(.A1(new_n9267_), .A2(new_n9268_), .B(new_n760_), .ZN(new_n9269_));
  NAND2_X1   g09012(.A1(new_n5741_), .A2(new_n9269_), .ZN(new_n9270_));
  XOR2_X1    g09013(.A1(new_n9270_), .A2(\a[14] ), .Z(new_n9271_));
  INV_X1     g09014(.I(new_n9271_), .ZN(new_n9272_));
  NAND3_X1   g09015(.A1(new_n8882_), .A2(new_n8879_), .A3(new_n8584_), .ZN(new_n9273_));
  AOI21_X1   g09016(.A1(new_n9273_), .A2(new_n8882_), .B(new_n9272_), .ZN(new_n9274_));
  OAI21_X1   g09017(.A1(new_n8521_), .A2(new_n8890_), .B(new_n8882_), .ZN(new_n9275_));
  NOR2_X1    g09018(.A1(new_n9275_), .A2(new_n9271_), .ZN(new_n9276_));
  OAI21_X1   g09019(.A1(new_n9276_), .A2(new_n9274_), .B(new_n9266_), .ZN(new_n9277_));
  OAI21_X1   g09020(.A1(new_n9264_), .A2(new_n9263_), .B(new_n9242_), .ZN(new_n9278_));
  NAND3_X1   g09021(.A1(new_n9243_), .A2(new_n9255_), .A3(new_n9261_), .ZN(new_n9279_));
  NAND2_X1   g09022(.A1(new_n9279_), .A2(new_n9278_), .ZN(new_n9280_));
  NAND2_X1   g09023(.A1(new_n9275_), .A2(new_n9271_), .ZN(new_n9281_));
  NAND3_X1   g09024(.A1(new_n9273_), .A2(new_n8882_), .A3(new_n9272_), .ZN(new_n9282_));
  NAND3_X1   g09025(.A1(new_n9281_), .A2(new_n9282_), .A3(new_n9280_), .ZN(new_n9283_));
  OAI22_X1   g09026(.A1(new_n582_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n577_), .ZN(new_n9284_));
  NAND2_X1   g09027(.A1(new_n960_), .A2(\b[52] ), .ZN(new_n9285_));
  AOI21_X1   g09028(.A1(new_n9284_), .A2(new_n9285_), .B(new_n585_), .ZN(new_n9286_));
  NAND2_X1   g09029(.A1(new_n6237_), .A2(new_n9286_), .ZN(new_n9287_));
  XOR2_X1    g09030(.A1(new_n9287_), .A2(\a[11] ), .Z(new_n9288_));
  INV_X1     g09031(.I(new_n9288_), .ZN(new_n9289_));
  NAND3_X1   g09032(.A1(new_n9277_), .A2(new_n9283_), .A3(new_n9289_), .ZN(new_n9290_));
  AOI21_X1   g09033(.A1(new_n9281_), .A2(new_n9282_), .B(new_n9280_), .ZN(new_n9291_));
  NOR3_X1    g09034(.A1(new_n9276_), .A2(new_n9274_), .A3(new_n9266_), .ZN(new_n9292_));
  OAI21_X1   g09035(.A1(new_n9292_), .A2(new_n9291_), .B(new_n9288_), .ZN(new_n9293_));
  NAND2_X1   g09036(.A1(new_n9293_), .A2(new_n9290_), .ZN(new_n9294_));
  OAI21_X1   g09037(.A1(new_n8900_), .A2(new_n8898_), .B(new_n8531_), .ZN(new_n9295_));
  NOR3_X1    g09038(.A1(new_n8893_), .A2(new_n8896_), .A3(new_n9295_), .ZN(new_n9296_));
  AOI21_X1   g09039(.A1(new_n8882_), .A2(new_n8879_), .B(new_n8521_), .ZN(new_n9297_));
  NOR3_X1    g09040(.A1(new_n8890_), .A2(new_n8891_), .A3(new_n8584_), .ZN(new_n9298_));
  OAI21_X1   g09041(.A1(new_n9298_), .A2(new_n9297_), .B(new_n8887_), .ZN(new_n9299_));
  OAI21_X1   g09042(.A1(new_n9296_), .A2(new_n8903_), .B(new_n9299_), .ZN(new_n9300_));
  OAI22_X1   g09043(.A1(new_n437_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n431_), .ZN(new_n9301_));
  NAND2_X1   g09044(.A1(new_n775_), .A2(\b[55] ), .ZN(new_n9302_));
  AOI21_X1   g09045(.A1(new_n9301_), .A2(new_n9302_), .B(new_n440_), .ZN(new_n9303_));
  NAND2_X1   g09046(.A1(new_n7308_), .A2(new_n9303_), .ZN(new_n9304_));
  XOR2_X1    g09047(.A1(new_n9304_), .A2(\a[8] ), .Z(new_n9305_));
  INV_X1     g09048(.I(new_n9305_), .ZN(new_n9306_));
  XOR2_X1    g09049(.A1(new_n9300_), .A2(new_n9306_), .Z(new_n9307_));
  NAND2_X1   g09050(.A1(new_n9307_), .A2(new_n9294_), .ZN(new_n9308_));
  XOR2_X1    g09051(.A1(new_n9300_), .A2(new_n9306_), .Z(new_n9309_));
  OAI21_X1   g09052(.A1(new_n9294_), .A2(new_n9309_), .B(new_n9308_), .ZN(new_n9310_));
  NOR2_X1    g09053(.A1(new_n8906_), .A2(new_n8921_), .ZN(new_n9311_));
  NOR2_X1    g09054(.A1(new_n9311_), .A2(new_n8919_), .ZN(new_n9312_));
  XOR2_X1    g09055(.A1(new_n9312_), .A2(new_n9310_), .Z(new_n9313_));
  XNOR2_X1   g09056(.A1(new_n9313_), .A2(new_n8974_), .ZN(new_n9314_));
  XOR2_X1    g09057(.A1(new_n9314_), .A2(new_n8969_), .Z(new_n9315_));
  AOI21_X1   g09058(.A1(new_n8541_), .A2(new_n8944_), .B(new_n8943_), .ZN(new_n9316_));
  XOR2_X1    g09059(.A1(new_n9315_), .A2(new_n9316_), .Z(new_n9317_));
  OAI21_X1   g09060(.A1(new_n8581_), .A2(new_n8949_), .B(new_n8583_), .ZN(new_n9318_));
  XOR2_X1    g09061(.A1(new_n9318_), .A2(new_n9317_), .Z(\f[63] ));
  INV_X1     g09062(.I(new_n8958_), .ZN(new_n9320_));
  NAND2_X1   g09063(.A1(new_n8955_), .A2(new_n8957_), .ZN(new_n9321_));
  OAI21_X1   g09064(.A1(new_n8955_), .A2(new_n9320_), .B(new_n9321_), .ZN(new_n9322_));
  INV_X1     g09065(.I(new_n9322_), .ZN(new_n9323_));
  NOR2_X1    g09066(.A1(new_n280_), .A2(new_n8932_), .ZN(new_n9324_));
  NOR2_X1    g09067(.A1(new_n404_), .A2(new_n8956_), .ZN(new_n9325_));
  NOR4_X1    g09068(.A1(new_n9323_), .A2(new_n264_), .A3(new_n9324_), .A4(new_n9325_), .ZN(new_n9326_));
  XOR2_X1    g09069(.A1(new_n9326_), .A2(new_n271_), .Z(new_n9327_));
  INV_X1     g09070(.I(new_n9327_), .ZN(new_n9328_));
  OAI22_X1   g09071(.A1(new_n364_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n320_), .ZN(new_n9329_));
  NAND2_X1   g09072(.A1(new_n594_), .A2(\b[59] ), .ZN(new_n9330_));
  AOI21_X1   g09073(.A1(new_n9329_), .A2(new_n9330_), .B(new_n312_), .ZN(new_n9331_));
  NAND3_X1   g09074(.A1(new_n8550_), .A2(new_n308_), .A3(new_n9331_), .ZN(new_n9332_));
  NAND2_X1   g09075(.A1(new_n8550_), .A2(new_n9331_), .ZN(new_n9333_));
  NAND2_X1   g09076(.A1(new_n9333_), .A2(\a[5] ), .ZN(new_n9334_));
  NAND2_X1   g09077(.A1(new_n9334_), .A2(new_n9332_), .ZN(new_n9335_));
  AOI21_X1   g09078(.A1(new_n9277_), .A2(new_n9283_), .B(new_n9289_), .ZN(new_n9336_));
  OAI21_X1   g09079(.A1(new_n9300_), .A2(new_n9336_), .B(new_n9290_), .ZN(new_n9337_));
  INV_X1     g09080(.I(new_n9237_), .ZN(new_n9338_));
  AOI21_X1   g09081(.A1(new_n9226_), .A2(new_n9231_), .B(new_n8975_), .ZN(new_n9339_));
  OAI22_X1   g09082(.A1(new_n1168_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n1163_), .ZN(new_n9340_));
  NAND2_X1   g09083(.A1(new_n1774_), .A2(\b[44] ), .ZN(new_n9341_));
  AOI21_X1   g09084(.A1(new_n9340_), .A2(new_n9341_), .B(new_n1171_), .ZN(new_n9342_));
  NAND2_X1   g09085(.A1(new_n4833_), .A2(new_n9342_), .ZN(new_n9343_));
  XOR2_X1    g09086(.A1(new_n9343_), .A2(\a[20] ), .Z(new_n9344_));
  OAI22_X1   g09087(.A1(new_n1444_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n1439_), .ZN(new_n9345_));
  NAND2_X1   g09088(.A1(new_n2098_), .A2(\b[41] ), .ZN(new_n9346_));
  AOI21_X1   g09089(.A1(new_n9345_), .A2(new_n9346_), .B(new_n1447_), .ZN(new_n9347_));
  NAND2_X1   g09090(.A1(new_n4320_), .A2(new_n9347_), .ZN(new_n9348_));
  XOR2_X1    g09091(.A1(new_n9348_), .A2(\a[23] ), .Z(new_n9349_));
  INV_X1     g09092(.I(new_n9349_), .ZN(new_n9350_));
  AOI21_X1   g09093(.A1(new_n9085_), .A2(new_n9086_), .B(new_n9083_), .ZN(new_n9351_));
  OAI21_X1   g09094(.A1(new_n8705_), .A2(new_n9351_), .B(new_n9089_), .ZN(new_n9352_));
  AOI21_X1   g09095(.A1(new_n8977_), .A2(new_n9017_), .B(new_n9015_), .ZN(new_n9353_));
  INV_X1     g09096(.I(new_n9353_), .ZN(new_n9354_));
  NAND2_X1   g09097(.A1(new_n9004_), .A2(new_n9006_), .ZN(new_n9355_));
  NAND2_X1   g09098(.A1(new_n8980_), .A2(new_n8990_), .ZN(new_n9356_));
  OAI22_X1   g09099(.A1(new_n393_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n290_), .ZN(new_n9357_));
  OAI21_X1   g09100(.A1(new_n292_), .A2(new_n8622_), .B(new_n9357_), .ZN(new_n9358_));
  NAND3_X1   g09101(.A1(new_n9358_), .A2(new_n334_), .A3(new_n8320_), .ZN(new_n9359_));
  XOR2_X1    g09102(.A1(new_n9359_), .A2(\a[62] ), .Z(new_n9360_));
  NOR2_X1    g09103(.A1(new_n8985_), .A2(new_n267_), .ZN(new_n9361_));
  INV_X1     g09104(.I(\a[63] ), .ZN(new_n9362_));
  NOR2_X1    g09105(.A1(new_n8309_), .A2(new_n9362_), .ZN(new_n9363_));
  INV_X1     g09106(.I(new_n9363_), .ZN(new_n9364_));
  NOR2_X1    g09107(.A1(new_n9364_), .A2(new_n258_), .ZN(new_n9365_));
  XNOR2_X1   g09108(.A1(new_n9361_), .A2(new_n9365_), .ZN(new_n9366_));
  XNOR2_X1   g09109(.A1(new_n9360_), .A2(new_n9366_), .ZN(new_n9367_));
  AOI21_X1   g09110(.A1(new_n8991_), .A2(new_n9356_), .B(new_n9367_), .ZN(new_n9368_));
  NAND2_X1   g09111(.A1(new_n9356_), .A2(new_n8991_), .ZN(new_n9369_));
  NOR2_X1    g09112(.A1(new_n9360_), .A2(new_n9366_), .ZN(new_n9370_));
  INV_X1     g09113(.I(new_n9370_), .ZN(new_n9371_));
  NAND2_X1   g09114(.A1(new_n9360_), .A2(new_n9366_), .ZN(new_n9372_));
  AOI21_X1   g09115(.A1(new_n9371_), .A2(new_n9372_), .B(new_n9369_), .ZN(new_n9373_));
  NOR2_X1    g09116(.A1(new_n9373_), .A2(new_n9368_), .ZN(new_n9374_));
  OAI22_X1   g09117(.A1(new_n450_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n403_), .ZN(new_n9375_));
  NAND2_X1   g09118(.A1(new_n8628_), .A2(\b[5] ), .ZN(new_n9376_));
  AOI21_X1   g09119(.A1(new_n9376_), .A2(new_n9375_), .B(new_n7354_), .ZN(new_n9377_));
  NAND2_X1   g09120(.A1(new_n454_), .A2(new_n9377_), .ZN(new_n9378_));
  XOR2_X1    g09121(.A1(new_n9378_), .A2(\a[59] ), .Z(new_n9379_));
  XOR2_X1    g09122(.A1(new_n9374_), .A2(new_n9379_), .Z(new_n9380_));
  AOI21_X1   g09123(.A1(new_n9005_), .A2(new_n9355_), .B(new_n9380_), .ZN(new_n9381_));
  NAND2_X1   g09124(.A1(new_n9355_), .A2(new_n9005_), .ZN(new_n9382_));
  INV_X1     g09125(.I(new_n9379_), .ZN(new_n9383_));
  NAND2_X1   g09126(.A1(new_n9374_), .A2(new_n9383_), .ZN(new_n9384_));
  OAI21_X1   g09127(.A1(new_n9373_), .A2(new_n9368_), .B(new_n9379_), .ZN(new_n9385_));
  AOI21_X1   g09128(.A1(new_n9384_), .A2(new_n9385_), .B(new_n9382_), .ZN(new_n9386_));
  NOR2_X1    g09129(.A1(new_n9386_), .A2(new_n9381_), .ZN(new_n9387_));
  OAI22_X1   g09130(.A1(new_n6721_), .A2(new_n510_), .B1(new_n6723_), .B2(new_n617_), .ZN(new_n9388_));
  NAND2_X1   g09131(.A1(new_n7617_), .A2(\b[8] ), .ZN(new_n9389_));
  AOI21_X1   g09132(.A1(new_n9389_), .A2(new_n9388_), .B(new_n6731_), .ZN(new_n9390_));
  NAND2_X1   g09133(.A1(new_n616_), .A2(new_n9390_), .ZN(new_n9391_));
  XOR2_X1    g09134(.A1(new_n9391_), .A2(\a[56] ), .Z(new_n9392_));
  INV_X1     g09135(.I(new_n9392_), .ZN(new_n9393_));
  XOR2_X1    g09136(.A1(new_n9387_), .A2(new_n9393_), .Z(new_n9394_));
  NAND2_X1   g09137(.A1(new_n9394_), .A2(new_n9354_), .ZN(new_n9395_));
  NAND2_X1   g09138(.A1(new_n9387_), .A2(new_n9393_), .ZN(new_n9396_));
  INV_X1     g09139(.I(new_n9396_), .ZN(new_n9397_));
  NOR2_X1    g09140(.A1(new_n9387_), .A2(new_n9393_), .ZN(new_n9398_));
  OAI21_X1   g09141(.A1(new_n9397_), .A2(new_n9398_), .B(new_n9353_), .ZN(new_n9399_));
  NAND2_X1   g09142(.A1(new_n9395_), .A2(new_n9399_), .ZN(new_n9400_));
  OAI22_X1   g09143(.A1(new_n5786_), .A2(new_n795_), .B1(new_n717_), .B2(new_n5792_), .ZN(new_n9401_));
  NAND2_X1   g09144(.A1(new_n6745_), .A2(\b[11] ), .ZN(new_n9402_));
  AOI21_X1   g09145(.A1(new_n9402_), .A2(new_n9401_), .B(new_n5796_), .ZN(new_n9403_));
  NAND2_X1   g09146(.A1(new_n799_), .A2(new_n9403_), .ZN(new_n9404_));
  XOR2_X1    g09147(.A1(new_n9404_), .A2(\a[53] ), .Z(new_n9405_));
  INV_X1     g09148(.I(new_n9405_), .ZN(new_n9406_));
  XOR2_X1    g09149(.A1(new_n9400_), .A2(new_n9406_), .Z(new_n9407_));
  OAI22_X1   g09150(.A1(new_n5228_), .A2(new_n992_), .B1(new_n904_), .B2(new_n5225_), .ZN(new_n9408_));
  NAND2_X1   g09151(.A1(new_n5387_), .A2(\b[14] ), .ZN(new_n9409_));
  AOI21_X1   g09152(.A1(new_n9408_), .A2(new_n9409_), .B(new_n5231_), .ZN(new_n9410_));
  NAND2_X1   g09153(.A1(new_n991_), .A2(new_n9410_), .ZN(new_n9411_));
  XOR2_X1    g09154(.A1(new_n9411_), .A2(\a[50] ), .Z(new_n9412_));
  XOR2_X1    g09155(.A1(new_n9021_), .A2(new_n9032_), .Z(new_n9413_));
  AOI21_X1   g09156(.A1(new_n9032_), .A2(new_n9030_), .B(new_n9413_), .ZN(new_n9414_));
  XOR2_X1    g09157(.A1(new_n9414_), .A2(new_n9412_), .Z(new_n9415_));
  XOR2_X1    g09158(.A1(new_n9415_), .A2(new_n9407_), .Z(new_n9416_));
  OAI22_X1   g09159(.A1(new_n4711_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n4706_), .ZN(new_n9417_));
  NAND2_X1   g09160(.A1(new_n5814_), .A2(\b[17] ), .ZN(new_n9418_));
  AOI21_X1   g09161(.A1(new_n9417_), .A2(new_n9418_), .B(new_n4714_), .ZN(new_n9419_));
  NAND2_X1   g09162(.A1(new_n1225_), .A2(new_n9419_), .ZN(new_n9420_));
  XOR2_X1    g09163(.A1(new_n9420_), .A2(\a[47] ), .Z(new_n9421_));
  XOR2_X1    g09164(.A1(new_n9416_), .A2(new_n9421_), .Z(new_n9422_));
  OAI22_X1   g09165(.A1(new_n4208_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n4203_), .ZN(new_n9423_));
  NAND2_X1   g09166(.A1(new_n5244_), .A2(\b[20] ), .ZN(new_n9424_));
  AOI21_X1   g09167(.A1(new_n9423_), .A2(new_n9424_), .B(new_n4211_), .ZN(new_n9425_));
  NAND2_X1   g09168(.A1(new_n1517_), .A2(new_n9425_), .ZN(new_n9426_));
  XOR2_X1    g09169(.A1(new_n9426_), .A2(\a[44] ), .Z(new_n9427_));
  INV_X1     g09170(.I(new_n9427_), .ZN(new_n9428_));
  NAND2_X1   g09171(.A1(new_n9422_), .A2(new_n9428_), .ZN(new_n9429_));
  INV_X1     g09172(.I(new_n9421_), .ZN(new_n9430_));
  XOR2_X1    g09173(.A1(new_n9416_), .A2(new_n9430_), .Z(new_n9431_));
  NAND2_X1   g09174(.A1(new_n9431_), .A2(new_n9427_), .ZN(new_n9432_));
  NAND2_X1   g09175(.A1(new_n9429_), .A2(new_n9432_), .ZN(new_n9433_));
  OAI22_X1   g09176(.A1(new_n3736_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n3731_), .ZN(new_n9434_));
  NAND2_X1   g09177(.A1(new_n4730_), .A2(\b[23] ), .ZN(new_n9435_));
  AOI21_X1   g09178(.A1(new_n9434_), .A2(new_n9435_), .B(new_n3739_), .ZN(new_n9436_));
  NAND2_X1   g09179(.A1(new_n1828_), .A2(new_n9436_), .ZN(new_n9437_));
  XOR2_X1    g09180(.A1(new_n9437_), .A2(\a[41] ), .Z(new_n9438_));
  XOR2_X1    g09181(.A1(new_n9433_), .A2(new_n9438_), .Z(new_n9439_));
  NAND2_X1   g09182(.A1(new_n9439_), .A2(new_n9352_), .ZN(new_n9440_));
  NOR3_X1    g09183(.A1(new_n9077_), .A2(new_n9071_), .A3(new_n9082_), .ZN(new_n9441_));
  AOI21_X1   g09184(.A1(new_n8704_), .A2(new_n9090_), .B(new_n9441_), .ZN(new_n9442_));
  INV_X1     g09185(.I(new_n9438_), .ZN(new_n9443_));
  XOR2_X1    g09186(.A1(new_n9433_), .A2(new_n9443_), .Z(new_n9444_));
  NAND2_X1   g09187(.A1(new_n9444_), .A2(new_n9442_), .ZN(new_n9445_));
  NAND2_X1   g09188(.A1(new_n9440_), .A2(new_n9445_), .ZN(new_n9446_));
  OAI22_X1   g09189(.A1(new_n3298_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n3293_), .ZN(new_n9447_));
  NAND2_X1   g09190(.A1(new_n4227_), .A2(\b[26] ), .ZN(new_n9448_));
  AOI21_X1   g09191(.A1(new_n9447_), .A2(new_n9448_), .B(new_n3301_), .ZN(new_n9449_));
  NAND2_X1   g09192(.A1(new_n2174_), .A2(new_n9449_), .ZN(new_n9450_));
  XOR2_X1    g09193(.A1(new_n9450_), .A2(\a[38] ), .Z(new_n9451_));
  NOR2_X1    g09194(.A1(new_n9446_), .A2(new_n9451_), .ZN(new_n9452_));
  XOR2_X1    g09195(.A1(new_n9433_), .A2(new_n9443_), .Z(new_n9453_));
  NOR2_X1    g09196(.A1(new_n9453_), .A2(new_n9442_), .ZN(new_n9454_));
  AOI21_X1   g09197(.A1(new_n9442_), .A2(new_n9444_), .B(new_n9454_), .ZN(new_n9455_));
  INV_X1     g09198(.I(new_n9451_), .ZN(new_n9456_));
  NOR2_X1    g09199(.A1(new_n9455_), .A2(new_n9456_), .ZN(new_n9457_));
  NOR2_X1    g09200(.A1(new_n9457_), .A2(new_n9452_), .ZN(new_n9458_));
  OAI22_X1   g09201(.A1(new_n2846_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n2841_), .ZN(new_n9459_));
  NAND2_X1   g09202(.A1(new_n3755_), .A2(\b[29] ), .ZN(new_n9460_));
  AOI21_X1   g09203(.A1(new_n9459_), .A2(new_n9460_), .B(new_n2849_), .ZN(new_n9461_));
  NAND2_X1   g09204(.A1(new_n2546_), .A2(new_n9461_), .ZN(new_n9462_));
  XOR2_X1    g09205(.A1(new_n9462_), .A2(\a[35] ), .Z(new_n9463_));
  NOR2_X1    g09206(.A1(new_n9458_), .A2(new_n9463_), .ZN(new_n9464_));
  NAND2_X1   g09207(.A1(new_n9455_), .A2(new_n9456_), .ZN(new_n9465_));
  NAND2_X1   g09208(.A1(new_n9446_), .A2(new_n9451_), .ZN(new_n9466_));
  NAND2_X1   g09209(.A1(new_n9465_), .A2(new_n9466_), .ZN(new_n9467_));
  INV_X1     g09210(.I(new_n9463_), .ZN(new_n9468_));
  NOR2_X1    g09211(.A1(new_n9467_), .A2(new_n9468_), .ZN(new_n9469_));
  OAI22_X1   g09212(.A1(new_n2452_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n2447_), .ZN(new_n9470_));
  NAND2_X1   g09213(.A1(new_n3312_), .A2(\b[32] ), .ZN(new_n9471_));
  AOI21_X1   g09214(.A1(new_n9470_), .A2(new_n9471_), .B(new_n2455_), .ZN(new_n9472_));
  NAND2_X1   g09215(.A1(new_n2963_), .A2(new_n9472_), .ZN(new_n9473_));
  XOR2_X1    g09216(.A1(new_n9473_), .A2(new_n2442_), .Z(new_n9474_));
  OAI21_X1   g09217(.A1(new_n9464_), .A2(new_n9469_), .B(new_n9474_), .ZN(new_n9475_));
  INV_X1     g09218(.I(new_n9475_), .ZN(new_n9476_));
  NAND2_X1   g09219(.A1(new_n9467_), .A2(new_n9468_), .ZN(new_n9477_));
  NAND2_X1   g09220(.A1(new_n9458_), .A2(new_n9463_), .ZN(new_n9478_));
  NAND2_X1   g09221(.A1(new_n9478_), .A2(new_n9477_), .ZN(new_n9479_));
  NOR2_X1    g09222(.A1(new_n9479_), .A2(new_n9474_), .ZN(new_n9480_));
  OAI22_X1   g09223(.A1(new_n2084_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n2079_), .ZN(new_n9481_));
  NAND2_X1   g09224(.A1(new_n2864_), .A2(\b[35] ), .ZN(new_n9482_));
  AOI21_X1   g09225(.A1(new_n9481_), .A2(new_n9482_), .B(new_n2087_), .ZN(new_n9483_));
  NAND2_X1   g09226(.A1(new_n3411_), .A2(new_n9483_), .ZN(new_n9484_));
  XOR2_X1    g09227(.A1(new_n9484_), .A2(\a[29] ), .Z(new_n9485_));
  OAI21_X1   g09228(.A1(new_n9476_), .A2(new_n9480_), .B(new_n9485_), .ZN(new_n9486_));
  OR3_X2     g09229(.A1(new_n9476_), .A2(new_n9480_), .A3(new_n9485_), .Z(new_n9487_));
  NAND2_X1   g09230(.A1(new_n9487_), .A2(new_n9486_), .ZN(new_n9488_));
  INV_X1     g09231(.I(new_n9488_), .ZN(new_n9489_));
  OAI22_X1   g09232(.A1(new_n1760_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n1755_), .ZN(new_n9490_));
  NAND2_X1   g09233(.A1(new_n2470_), .A2(\b[38] ), .ZN(new_n9491_));
  AOI21_X1   g09234(.A1(new_n9490_), .A2(new_n9491_), .B(new_n1763_), .ZN(new_n9492_));
  NAND2_X1   g09235(.A1(new_n3844_), .A2(new_n9492_), .ZN(new_n9493_));
  XOR2_X1    g09236(.A1(new_n9493_), .A2(\a[26] ), .Z(new_n9494_));
  INV_X1     g09237(.I(new_n9494_), .ZN(new_n9495_));
  NOR3_X1    g09238(.A1(new_n9154_), .A2(new_n9153_), .A3(new_n9150_), .ZN(new_n9496_));
  AOI21_X1   g09239(.A1(new_n9139_), .A2(new_n9145_), .B(new_n9151_), .ZN(new_n9497_));
  NOR3_X1    g09240(.A1(new_n9174_), .A2(new_n9496_), .A3(new_n9497_), .ZN(new_n9498_));
  AOI21_X1   g09241(.A1(new_n9152_), .A2(new_n9155_), .B(new_n9168_), .ZN(new_n9499_));
  OAI21_X1   g09242(.A1(new_n9499_), .A2(new_n9498_), .B(new_n9162_), .ZN(new_n9500_));
  NOR3_X1    g09243(.A1(new_n9499_), .A2(new_n9498_), .A3(new_n9162_), .ZN(new_n9501_));
  NAND3_X1   g09244(.A1(new_n9168_), .A2(new_n9155_), .A3(new_n9152_), .ZN(new_n9502_));
  OAI21_X1   g09245(.A1(new_n9496_), .A2(new_n9497_), .B(new_n9174_), .ZN(new_n9503_));
  AOI21_X1   g09246(.A1(new_n9503_), .A2(new_n9502_), .B(new_n9170_), .ZN(new_n9504_));
  OAI21_X1   g09247(.A1(new_n9501_), .A2(new_n9504_), .B(new_n9193_), .ZN(new_n9505_));
  AOI21_X1   g09248(.A1(new_n9505_), .A2(new_n9500_), .B(new_n9495_), .ZN(new_n9506_));
  NAND3_X1   g09249(.A1(new_n9503_), .A2(new_n9502_), .A3(new_n9170_), .ZN(new_n9507_));
  OAI21_X1   g09250(.A1(new_n9499_), .A2(new_n9498_), .B(new_n9162_), .ZN(new_n9508_));
  AOI22_X1   g09251(.A1(new_n9508_), .A2(new_n9507_), .B1(new_n9170_), .B2(new_n9187_), .ZN(new_n9509_));
  NOR2_X1    g09252(.A1(new_n9509_), .A2(new_n9494_), .ZN(new_n9510_));
  OAI21_X1   g09253(.A1(new_n9506_), .A2(new_n9510_), .B(new_n9489_), .ZN(new_n9511_));
  NAND2_X1   g09254(.A1(new_n9509_), .A2(new_n9494_), .ZN(new_n9512_));
  NAND3_X1   g09255(.A1(new_n9505_), .A2(new_n9495_), .A3(new_n9500_), .ZN(new_n9513_));
  NAND3_X1   g09256(.A1(new_n9512_), .A2(new_n9513_), .A3(new_n9488_), .ZN(new_n9514_));
  AOI21_X1   g09257(.A1(new_n9511_), .A2(new_n9514_), .B(new_n9350_), .ZN(new_n9515_));
  AOI21_X1   g09258(.A1(new_n9512_), .A2(new_n9513_), .B(new_n9488_), .ZN(new_n9516_));
  NOR3_X1    g09259(.A1(new_n9506_), .A2(new_n9510_), .A3(new_n9489_), .ZN(new_n9517_));
  NOR3_X1    g09260(.A1(new_n9516_), .A2(new_n9517_), .A3(new_n9349_), .ZN(new_n9518_));
  OAI21_X1   g09261(.A1(new_n9518_), .A2(new_n9515_), .B(new_n9344_), .ZN(new_n9519_));
  INV_X1     g09262(.I(new_n9344_), .ZN(new_n9520_));
  OAI21_X1   g09263(.A1(new_n9517_), .A2(new_n9516_), .B(new_n9349_), .ZN(new_n9521_));
  NAND3_X1   g09264(.A1(new_n9511_), .A2(new_n9514_), .A3(new_n9350_), .ZN(new_n9522_));
  NAND3_X1   g09265(.A1(new_n9521_), .A2(new_n9522_), .A3(new_n9520_), .ZN(new_n9523_));
  NAND2_X1   g09266(.A1(new_n9519_), .A2(new_n9523_), .ZN(new_n9524_));
  OAI22_X1   g09267(.A1(new_n940_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n935_), .ZN(new_n9525_));
  NAND2_X1   g09268(.A1(new_n1458_), .A2(\b[47] ), .ZN(new_n9526_));
  AOI21_X1   g09269(.A1(new_n9525_), .A2(new_n9526_), .B(new_n943_), .ZN(new_n9527_));
  NAND2_X1   g09270(.A1(new_n5196_), .A2(new_n9527_), .ZN(new_n9528_));
  XOR2_X1    g09271(.A1(new_n9528_), .A2(\a[17] ), .Z(new_n9529_));
  INV_X1     g09272(.I(new_n9529_), .ZN(new_n9530_));
  NAND2_X1   g09273(.A1(new_n9524_), .A2(new_n9530_), .ZN(new_n9531_));
  AOI21_X1   g09274(.A1(new_n9521_), .A2(new_n9522_), .B(new_n9520_), .ZN(new_n9532_));
  NOR3_X1    g09275(.A1(new_n9518_), .A2(new_n9515_), .A3(new_n9344_), .ZN(new_n9533_));
  NOR2_X1    g09276(.A1(new_n9533_), .A2(new_n9532_), .ZN(new_n9534_));
  NAND2_X1   g09277(.A1(new_n9534_), .A2(new_n9529_), .ZN(new_n9535_));
  NAND2_X1   g09278(.A1(new_n9535_), .A2(new_n9531_), .ZN(new_n9536_));
  OAI21_X1   g09279(.A1(new_n9338_), .A2(new_n9339_), .B(new_n9536_), .ZN(new_n9537_));
  NAND2_X1   g09280(.A1(new_n9240_), .A2(new_n9236_), .ZN(new_n9538_));
  NAND2_X1   g09281(.A1(new_n9534_), .A2(new_n9530_), .ZN(new_n9539_));
  AOI21_X1   g09282(.A1(new_n9519_), .A2(new_n9523_), .B(new_n9530_), .ZN(new_n9540_));
  INV_X1     g09283(.I(new_n9540_), .ZN(new_n9541_));
  NAND2_X1   g09284(.A1(new_n9539_), .A2(new_n9541_), .ZN(new_n9542_));
  NAND3_X1   g09285(.A1(new_n9542_), .A2(new_n9538_), .A3(new_n9237_), .ZN(new_n9543_));
  NAND2_X1   g09286(.A1(new_n9537_), .A2(new_n9543_), .ZN(new_n9544_));
  OAI22_X1   g09287(.A1(new_n757_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n752_), .ZN(new_n9545_));
  NAND2_X1   g09288(.A1(new_n1182_), .A2(\b[50] ), .ZN(new_n9546_));
  AOI21_X1   g09289(.A1(new_n9545_), .A2(new_n9546_), .B(new_n760_), .ZN(new_n9547_));
  NAND2_X1   g09290(.A1(new_n5954_), .A2(new_n9547_), .ZN(new_n9548_));
  XOR2_X1    g09291(.A1(new_n9548_), .A2(\a[14] ), .Z(new_n9549_));
  NOR2_X1    g09292(.A1(new_n9544_), .A2(new_n9549_), .ZN(new_n9550_));
  AOI22_X1   g09293(.A1(new_n9538_), .A2(new_n9237_), .B1(new_n9531_), .B2(new_n9535_), .ZN(new_n9551_));
  NOR2_X1    g09294(.A1(new_n9524_), .A2(new_n9529_), .ZN(new_n9552_));
  NOR2_X1    g09295(.A1(new_n9552_), .A2(new_n9540_), .ZN(new_n9553_));
  NOR3_X1    g09296(.A1(new_n9339_), .A2(new_n9553_), .A3(new_n9338_), .ZN(new_n9554_));
  NOR2_X1    g09297(.A1(new_n9551_), .A2(new_n9554_), .ZN(new_n9555_));
  INV_X1     g09298(.I(new_n9549_), .ZN(new_n9556_));
  NOR2_X1    g09299(.A1(new_n9555_), .A2(new_n9556_), .ZN(new_n9557_));
  NOR2_X1    g09300(.A1(new_n9550_), .A2(new_n9557_), .ZN(new_n9558_));
  OAI22_X1   g09301(.A1(new_n582_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n577_), .ZN(new_n9559_));
  NAND2_X1   g09302(.A1(new_n960_), .A2(\b[53] ), .ZN(new_n9560_));
  AOI21_X1   g09303(.A1(new_n9559_), .A2(new_n9560_), .B(new_n585_), .ZN(new_n9561_));
  NAND2_X1   g09304(.A1(new_n6471_), .A2(new_n9561_), .ZN(new_n9562_));
  XOR2_X1    g09305(.A1(new_n9562_), .A2(\a[11] ), .Z(new_n9563_));
  NOR2_X1    g09306(.A1(new_n9558_), .A2(new_n9563_), .ZN(new_n9564_));
  INV_X1     g09307(.I(new_n9558_), .ZN(new_n9565_));
  INV_X1     g09308(.I(new_n9563_), .ZN(new_n9566_));
  NOR2_X1    g09309(.A1(new_n9565_), .A2(new_n9566_), .ZN(new_n9567_));
  NOR2_X1    g09310(.A1(new_n9567_), .A2(new_n9564_), .ZN(new_n9568_));
  OAI22_X1   g09311(.A1(new_n437_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n431_), .ZN(new_n9569_));
  NAND2_X1   g09312(.A1(new_n775_), .A2(\b[56] ), .ZN(new_n9570_));
  AOI21_X1   g09313(.A1(new_n9569_), .A2(new_n9570_), .B(new_n440_), .ZN(new_n9571_));
  NAND2_X1   g09314(.A1(new_n7559_), .A2(new_n9571_), .ZN(new_n9572_));
  XOR2_X1    g09315(.A1(new_n9572_), .A2(\a[8] ), .Z(new_n9573_));
  XOR2_X1    g09316(.A1(new_n9568_), .A2(new_n9573_), .Z(new_n9574_));
  XOR2_X1    g09317(.A1(new_n9568_), .A2(new_n9573_), .Z(new_n9575_));
  NOR2_X1    g09318(.A1(new_n9575_), .A2(new_n9337_), .ZN(new_n9576_));
  AOI21_X1   g09319(.A1(new_n9337_), .A2(new_n9574_), .B(new_n9576_), .ZN(new_n9577_));
  NAND2_X1   g09320(.A1(new_n9306_), .A2(new_n8974_), .ZN(new_n9578_));
  XOR2_X1    g09321(.A1(new_n9294_), .A2(new_n9300_), .Z(new_n9579_));
  OR3_X2     g09322(.A1(new_n9579_), .A2(new_n8974_), .A3(new_n9306_), .Z(new_n9580_));
  NAND2_X1   g09323(.A1(new_n9580_), .A2(new_n9578_), .ZN(new_n9581_));
  XOR2_X1    g09324(.A1(new_n9581_), .A2(new_n9577_), .Z(new_n9582_));
  XOR2_X1    g09325(.A1(new_n9582_), .A2(new_n9335_), .Z(new_n9583_));
  XOR2_X1    g09326(.A1(new_n9583_), .A2(new_n9328_), .Z(new_n9584_));
  XOR2_X1    g09327(.A1(new_n9310_), .A2(new_n8974_), .Z(new_n9585_));
  NAND3_X1   g09328(.A1(new_n9585_), .A2(new_n8969_), .A3(new_n9312_), .ZN(new_n9586_));
  OAI21_X1   g09329(.A1(new_n8969_), .A2(new_n9312_), .B(new_n9586_), .ZN(new_n9587_));
  NOR2_X1    g09330(.A1(new_n8581_), .A2(new_n8950_), .ZN(new_n9588_));
  NAND2_X1   g09331(.A1(new_n9315_), .A2(new_n9316_), .ZN(new_n9589_));
  NAND3_X1   g09332(.A1(new_n9317_), .A2(new_n8950_), .A3(new_n9589_), .ZN(new_n9590_));
  NOR2_X1    g09333(.A1(new_n9588_), .A2(new_n9590_), .ZN(new_n9591_));
  XOR2_X1    g09334(.A1(new_n9591_), .A2(new_n9587_), .Z(new_n9592_));
  XOR2_X1    g09335(.A1(new_n9592_), .A2(new_n9584_), .Z(\f[64] ));
  NAND2_X1   g09336(.A1(new_n8955_), .A2(new_n8932_), .ZN(new_n9594_));
  NAND2_X1   g09337(.A1(new_n9594_), .A2(\b[63] ), .ZN(new_n9595_));
  NOR2_X1    g09338(.A1(new_n9595_), .A2(new_n264_), .ZN(new_n9596_));
  NAND4_X1   g09339(.A1(new_n9596_), .A2(\a[2] ), .A3(\b[63] ), .A4(new_n279_), .ZN(new_n9597_));
  INV_X1     g09340(.I(new_n9597_), .ZN(new_n9598_));
  OAI22_X1   g09341(.A1(new_n364_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n320_), .ZN(new_n9599_));
  NAND2_X1   g09342(.A1(new_n594_), .A2(\b[60] ), .ZN(new_n9600_));
  AOI21_X1   g09343(.A1(new_n9599_), .A2(new_n9600_), .B(new_n312_), .ZN(new_n9601_));
  NAND2_X1   g09344(.A1(new_n8935_), .A2(new_n9601_), .ZN(new_n9602_));
  XOR2_X1    g09345(.A1(new_n9602_), .A2(\a[5] ), .Z(new_n9603_));
  NOR2_X1    g09346(.A1(new_n9565_), .A2(new_n9563_), .ZN(new_n9604_));
  INV_X1     g09347(.I(new_n9604_), .ZN(new_n9605_));
  NOR2_X1    g09348(.A1(new_n9558_), .A2(new_n9566_), .ZN(new_n9606_));
  INV_X1     g09349(.I(new_n9606_), .ZN(new_n9607_));
  NAND2_X1   g09350(.A1(new_n9337_), .A2(new_n9607_), .ZN(new_n9608_));
  NOR3_X1    g09351(.A1(new_n9339_), .A2(new_n9338_), .A3(new_n9534_), .ZN(new_n9609_));
  AOI21_X1   g09352(.A1(new_n9538_), .A2(new_n9237_), .B(new_n9524_), .ZN(new_n9610_));
  OAI21_X1   g09353(.A1(new_n9610_), .A2(new_n9609_), .B(new_n9529_), .ZN(new_n9611_));
  NAND2_X1   g09354(.A1(new_n9611_), .A2(new_n9544_), .ZN(new_n9612_));
  OAI22_X1   g09355(.A1(new_n1444_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n1439_), .ZN(new_n9613_));
  NAND2_X1   g09356(.A1(new_n2098_), .A2(\b[42] ), .ZN(new_n9614_));
  AOI21_X1   g09357(.A1(new_n9613_), .A2(new_n9614_), .B(new_n1447_), .ZN(new_n9615_));
  NAND2_X1   g09358(.A1(new_n4500_), .A2(new_n9615_), .ZN(new_n9616_));
  XOR2_X1    g09359(.A1(new_n9616_), .A2(\a[23] ), .Z(new_n9617_));
  OAI22_X1   g09360(.A1(new_n1760_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n1755_), .ZN(new_n9618_));
  NAND2_X1   g09361(.A1(new_n2470_), .A2(\b[39] ), .ZN(new_n9619_));
  AOI21_X1   g09362(.A1(new_n9618_), .A2(new_n9619_), .B(new_n1763_), .ZN(new_n9620_));
  NAND2_X1   g09363(.A1(new_n3996_), .A2(new_n9620_), .ZN(new_n9621_));
  XOR2_X1    g09364(.A1(new_n9621_), .A2(\a[26] ), .Z(new_n9622_));
  INV_X1     g09365(.I(new_n9622_), .ZN(new_n9623_));
  AOI21_X1   g09366(.A1(new_n9505_), .A2(new_n9500_), .B(new_n9488_), .ZN(new_n9624_));
  NOR2_X1    g09367(.A1(new_n9509_), .A2(new_n9489_), .ZN(new_n9625_));
  OAI21_X1   g09368(.A1(new_n9624_), .A2(new_n9625_), .B(new_n9494_), .ZN(new_n9626_));
  NOR2_X1    g09369(.A1(new_n9467_), .A2(new_n9463_), .ZN(new_n9627_));
  INV_X1     g09370(.I(new_n9627_), .ZN(new_n9628_));
  XOR2_X1    g09371(.A1(new_n9433_), .A2(new_n9442_), .Z(new_n9629_));
  NOR2_X1    g09372(.A1(new_n9629_), .A2(new_n9443_), .ZN(new_n9630_));
  XOR2_X1    g09373(.A1(new_n9407_), .A2(new_n9414_), .Z(new_n9631_));
  NOR2_X1    g09374(.A1(new_n9631_), .A2(new_n9412_), .ZN(new_n9632_));
  INV_X1     g09375(.I(new_n9632_), .ZN(new_n9633_));
  NOR2_X1    g09376(.A1(new_n9400_), .A2(new_n9405_), .ZN(new_n9634_));
  NAND2_X1   g09377(.A1(new_n9400_), .A2(new_n9405_), .ZN(new_n9635_));
  AOI21_X1   g09378(.A1(new_n9414_), .A2(new_n9635_), .B(new_n9634_), .ZN(new_n9636_));
  INV_X1     g09379(.I(new_n9636_), .ZN(new_n9637_));
  OAI21_X1   g09380(.A1(new_n9353_), .A2(new_n9398_), .B(new_n9396_), .ZN(new_n9638_));
  INV_X1     g09381(.I(new_n9638_), .ZN(new_n9639_));
  NAND2_X1   g09382(.A1(new_n9382_), .A2(new_n9385_), .ZN(new_n9640_));
  NAND2_X1   g09383(.A1(new_n9640_), .A2(new_n9384_), .ZN(new_n9641_));
  AOI21_X1   g09384(.A1(new_n9369_), .A2(new_n9372_), .B(new_n9370_), .ZN(new_n9642_));
  OAI22_X1   g09385(.A1(new_n347_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n393_), .ZN(new_n9643_));
  INV_X1     g09386(.I(new_n8622_), .ZN(new_n9644_));
  NAND2_X1   g09387(.A1(new_n9644_), .A2(\b[3] ), .ZN(new_n9645_));
  AOI21_X1   g09388(.A1(new_n9645_), .A2(new_n9643_), .B(new_n8321_), .ZN(new_n9646_));
  NAND2_X1   g09389(.A1(new_n352_), .A2(new_n9646_), .ZN(new_n9647_));
  XOR2_X1    g09390(.A1(new_n9647_), .A2(\a[62] ), .Z(new_n9648_));
  INV_X1     g09391(.I(new_n8985_), .ZN(new_n9649_));
  NAND2_X1   g09392(.A1(new_n9649_), .A2(\b[2] ), .ZN(new_n9650_));
  NOR2_X1    g09393(.A1(new_n9364_), .A2(new_n267_), .ZN(new_n9651_));
  XOR2_X1    g09394(.A1(new_n9650_), .A2(new_n9651_), .Z(new_n9652_));
  INV_X1     g09395(.I(new_n9652_), .ZN(new_n9653_));
  XOR2_X1    g09396(.A1(new_n9648_), .A2(new_n9653_), .Z(new_n9654_));
  NOR2_X1    g09397(.A1(new_n9654_), .A2(new_n9642_), .ZN(new_n9655_));
  INV_X1     g09398(.I(new_n9642_), .ZN(new_n9656_));
  NOR2_X1    g09399(.A1(new_n9648_), .A2(new_n9652_), .ZN(new_n9657_));
  INV_X1     g09400(.I(new_n9648_), .ZN(new_n9658_));
  NOR2_X1    g09401(.A1(new_n9658_), .A2(new_n9653_), .ZN(new_n9659_));
  NOR2_X1    g09402(.A1(new_n9659_), .A2(new_n9657_), .ZN(new_n9660_));
  NOR2_X1    g09403(.A1(new_n9656_), .A2(new_n9660_), .ZN(new_n9661_));
  NOR2_X1    g09404(.A1(new_n9661_), .A2(new_n9655_), .ZN(new_n9662_));
  OAI22_X1   g09405(.A1(new_n495_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n450_), .ZN(new_n9663_));
  NAND2_X1   g09406(.A1(new_n8628_), .A2(\b[6] ), .ZN(new_n9664_));
  AOI21_X1   g09407(.A1(new_n9664_), .A2(new_n9663_), .B(new_n7354_), .ZN(new_n9665_));
  NAND2_X1   g09408(.A1(new_n494_), .A2(new_n9665_), .ZN(new_n9666_));
  XOR2_X1    g09409(.A1(new_n9666_), .A2(\a[59] ), .Z(new_n9667_));
  INV_X1     g09410(.I(new_n9667_), .ZN(new_n9668_));
  NAND2_X1   g09411(.A1(new_n9662_), .A2(new_n9668_), .ZN(new_n9669_));
  OAI21_X1   g09412(.A1(new_n9661_), .A2(new_n9655_), .B(new_n9667_), .ZN(new_n9670_));
  NAND2_X1   g09413(.A1(new_n9669_), .A2(new_n9670_), .ZN(new_n9671_));
  XOR2_X1    g09414(.A1(new_n9662_), .A2(new_n9667_), .Z(new_n9672_));
  NOR2_X1    g09415(.A1(new_n9641_), .A2(new_n9672_), .ZN(new_n9673_));
  AOI21_X1   g09416(.A1(new_n9641_), .A2(new_n9671_), .B(new_n9673_), .ZN(new_n9674_));
  OAI22_X1   g09417(.A1(new_n6721_), .A2(new_n617_), .B1(new_n6723_), .B2(new_n659_), .ZN(new_n9675_));
  NAND2_X1   g09418(.A1(new_n7617_), .A2(\b[9] ), .ZN(new_n9676_));
  AOI21_X1   g09419(.A1(new_n9676_), .A2(new_n9675_), .B(new_n6731_), .ZN(new_n9677_));
  NAND2_X1   g09420(.A1(new_n663_), .A2(new_n9677_), .ZN(new_n9678_));
  XOR2_X1    g09421(.A1(new_n9678_), .A2(\a[56] ), .Z(new_n9679_));
  XNOR2_X1   g09422(.A1(new_n9674_), .A2(new_n9679_), .ZN(new_n9680_));
  NOR2_X1    g09423(.A1(new_n9680_), .A2(new_n9639_), .ZN(new_n9681_));
  OR2_X2     g09424(.A1(new_n9674_), .A2(new_n9679_), .Z(new_n9682_));
  NAND2_X1   g09425(.A1(new_n9674_), .A2(new_n9679_), .ZN(new_n9683_));
  NAND2_X1   g09426(.A1(new_n9682_), .A2(new_n9683_), .ZN(new_n9684_));
  AOI21_X1   g09427(.A1(new_n9639_), .A2(new_n9684_), .B(new_n9681_), .ZN(new_n9685_));
  OAI22_X1   g09428(.A1(new_n5786_), .A2(new_n848_), .B1(new_n795_), .B2(new_n5792_), .ZN(new_n9686_));
  NAND2_X1   g09429(.A1(new_n6745_), .A2(\b[12] ), .ZN(new_n9687_));
  AOI21_X1   g09430(.A1(new_n9687_), .A2(new_n9686_), .B(new_n5796_), .ZN(new_n9688_));
  NAND2_X1   g09431(.A1(new_n847_), .A2(new_n9688_), .ZN(new_n9689_));
  XOR2_X1    g09432(.A1(new_n9689_), .A2(\a[53] ), .Z(new_n9690_));
  INV_X1     g09433(.I(new_n9690_), .ZN(new_n9691_));
  NAND2_X1   g09434(.A1(new_n9685_), .A2(new_n9691_), .ZN(new_n9692_));
  AOI21_X1   g09435(.A1(new_n9682_), .A2(new_n9683_), .B(new_n9638_), .ZN(new_n9693_));
  OAI21_X1   g09436(.A1(new_n9681_), .A2(new_n9693_), .B(new_n9690_), .ZN(new_n9694_));
  NAND2_X1   g09437(.A1(new_n9692_), .A2(new_n9694_), .ZN(new_n9695_));
  NAND2_X1   g09438(.A1(new_n9637_), .A2(new_n9695_), .ZN(new_n9696_));
  XOR2_X1    g09439(.A1(new_n9685_), .A2(new_n9691_), .Z(new_n9697_));
  NAND2_X1   g09440(.A1(new_n9697_), .A2(new_n9636_), .ZN(new_n9698_));
  OAI22_X1   g09441(.A1(new_n5228_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n5225_), .ZN(new_n9699_));
  NAND2_X1   g09442(.A1(new_n5387_), .A2(\b[15] ), .ZN(new_n9700_));
  AOI21_X1   g09443(.A1(new_n9699_), .A2(new_n9700_), .B(new_n5231_), .ZN(new_n9701_));
  NAND2_X1   g09444(.A1(new_n1047_), .A2(new_n9701_), .ZN(new_n9702_));
  XOR2_X1    g09445(.A1(new_n9702_), .A2(\a[50] ), .Z(new_n9703_));
  INV_X1     g09446(.I(new_n9703_), .ZN(new_n9704_));
  NAND3_X1   g09447(.A1(new_n9698_), .A2(new_n9696_), .A3(new_n9704_), .ZN(new_n9705_));
  AOI21_X1   g09448(.A1(new_n9698_), .A2(new_n9696_), .B(new_n9704_), .ZN(new_n9706_));
  INV_X1     g09449(.I(new_n9706_), .ZN(new_n9707_));
  AOI21_X1   g09450(.A1(new_n9707_), .A2(new_n9705_), .B(new_n9633_), .ZN(new_n9708_));
  INV_X1     g09451(.I(new_n9696_), .ZN(new_n9709_));
  XOR2_X1    g09452(.A1(new_n9685_), .A2(new_n9690_), .Z(new_n9710_));
  NOR2_X1    g09453(.A1(new_n9710_), .A2(new_n9637_), .ZN(new_n9711_));
  OAI21_X1   g09454(.A1(new_n9709_), .A2(new_n9711_), .B(new_n9704_), .ZN(new_n9712_));
  NAND3_X1   g09455(.A1(new_n9698_), .A2(new_n9696_), .A3(new_n9703_), .ZN(new_n9713_));
  AOI21_X1   g09456(.A1(new_n9712_), .A2(new_n9713_), .B(new_n9632_), .ZN(new_n9714_));
  OAI22_X1   g09457(.A1(new_n4711_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n4706_), .ZN(new_n9715_));
  NAND2_X1   g09458(.A1(new_n5814_), .A2(\b[18] ), .ZN(new_n9716_));
  AOI21_X1   g09459(.A1(new_n9715_), .A2(new_n9716_), .B(new_n4714_), .ZN(new_n9717_));
  NAND2_X1   g09460(.A1(new_n1304_), .A2(new_n9717_), .ZN(new_n9718_));
  XOR2_X1    g09461(.A1(new_n9718_), .A2(\a[47] ), .Z(new_n9719_));
  NOR3_X1    g09462(.A1(new_n9708_), .A2(new_n9714_), .A3(new_n9719_), .ZN(new_n9720_));
  INV_X1     g09463(.I(new_n9705_), .ZN(new_n9721_));
  OAI21_X1   g09464(.A1(new_n9721_), .A2(new_n9706_), .B(new_n9632_), .ZN(new_n9722_));
  AOI21_X1   g09465(.A1(new_n9698_), .A2(new_n9696_), .B(new_n9703_), .ZN(new_n9723_));
  NOR3_X1    g09466(.A1(new_n9709_), .A2(new_n9711_), .A3(new_n9704_), .ZN(new_n9724_));
  OAI21_X1   g09467(.A1(new_n9724_), .A2(new_n9723_), .B(new_n9633_), .ZN(new_n9725_));
  INV_X1     g09468(.I(new_n9719_), .ZN(new_n9726_));
  AOI21_X1   g09469(.A1(new_n9722_), .A2(new_n9725_), .B(new_n9726_), .ZN(new_n9727_));
  NOR2_X1    g09470(.A1(new_n9720_), .A2(new_n9727_), .ZN(new_n9728_));
  OAI22_X1   g09471(.A1(new_n4208_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n4203_), .ZN(new_n9729_));
  NAND2_X1   g09472(.A1(new_n5244_), .A2(\b[21] ), .ZN(new_n9730_));
  AOI21_X1   g09473(.A1(new_n9729_), .A2(new_n9730_), .B(new_n4211_), .ZN(new_n9731_));
  NAND2_X1   g09474(.A1(new_n1604_), .A2(new_n9731_), .ZN(new_n9732_));
  XOR2_X1    g09475(.A1(new_n9732_), .A2(\a[44] ), .Z(new_n9733_));
  INV_X1     g09476(.I(new_n9733_), .ZN(new_n9734_));
  NAND2_X1   g09477(.A1(new_n9352_), .A2(new_n9428_), .ZN(new_n9735_));
  OAI21_X1   g09478(.A1(new_n9352_), .A2(new_n9428_), .B(new_n9422_), .ZN(new_n9736_));
  NOR2_X1    g09479(.A1(new_n9416_), .A2(new_n9421_), .ZN(new_n9737_));
  NAND3_X1   g09480(.A1(new_n9736_), .A2(new_n9735_), .A3(new_n9737_), .ZN(new_n9738_));
  NOR2_X1    g09481(.A1(new_n9442_), .A2(new_n9427_), .ZN(new_n9739_));
  AOI21_X1   g09482(.A1(new_n9442_), .A2(new_n9427_), .B(new_n9431_), .ZN(new_n9740_));
  INV_X1     g09483(.I(new_n9737_), .ZN(new_n9741_));
  OAI21_X1   g09484(.A1(new_n9740_), .A2(new_n9739_), .B(new_n9741_), .ZN(new_n9742_));
  AOI21_X1   g09485(.A1(new_n9742_), .A2(new_n9738_), .B(new_n9734_), .ZN(new_n9743_));
  NOR3_X1    g09486(.A1(new_n9740_), .A2(new_n9739_), .A3(new_n9741_), .ZN(new_n9744_));
  AOI21_X1   g09487(.A1(new_n9736_), .A2(new_n9735_), .B(new_n9737_), .ZN(new_n9745_));
  NOR3_X1    g09488(.A1(new_n9744_), .A2(new_n9745_), .A3(new_n9733_), .ZN(new_n9746_));
  OAI21_X1   g09489(.A1(new_n9746_), .A2(new_n9743_), .B(new_n9728_), .ZN(new_n9747_));
  NAND3_X1   g09490(.A1(new_n9722_), .A2(new_n9725_), .A3(new_n9726_), .ZN(new_n9748_));
  OAI21_X1   g09491(.A1(new_n9708_), .A2(new_n9714_), .B(new_n9719_), .ZN(new_n9749_));
  NAND2_X1   g09492(.A1(new_n9749_), .A2(new_n9748_), .ZN(new_n9750_));
  OAI21_X1   g09493(.A1(new_n9744_), .A2(new_n9745_), .B(new_n9733_), .ZN(new_n9751_));
  NAND3_X1   g09494(.A1(new_n9742_), .A2(new_n9738_), .A3(new_n9734_), .ZN(new_n9752_));
  NAND3_X1   g09495(.A1(new_n9751_), .A2(new_n9752_), .A3(new_n9750_), .ZN(new_n9753_));
  OAI22_X1   g09496(.A1(new_n3736_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n3731_), .ZN(new_n9754_));
  NAND2_X1   g09497(.A1(new_n4730_), .A2(\b[24] ), .ZN(new_n9755_));
  AOI21_X1   g09498(.A1(new_n9754_), .A2(new_n9755_), .B(new_n3739_), .ZN(new_n9756_));
  NAND2_X1   g09499(.A1(new_n1926_), .A2(new_n9756_), .ZN(new_n9757_));
  XOR2_X1    g09500(.A1(new_n9757_), .A2(\a[41] ), .Z(new_n9758_));
  AOI21_X1   g09501(.A1(new_n9747_), .A2(new_n9753_), .B(new_n9758_), .ZN(new_n9759_));
  AOI21_X1   g09502(.A1(new_n9751_), .A2(new_n9752_), .B(new_n9750_), .ZN(new_n9760_));
  NOR3_X1    g09503(.A1(new_n9746_), .A2(new_n9743_), .A3(new_n9728_), .ZN(new_n9761_));
  INV_X1     g09504(.I(new_n9758_), .ZN(new_n9762_));
  NOR3_X1    g09505(.A1(new_n9761_), .A2(new_n9760_), .A3(new_n9762_), .ZN(new_n9763_));
  OAI21_X1   g09506(.A1(new_n9763_), .A2(new_n9759_), .B(new_n9630_), .ZN(new_n9764_));
  INV_X1     g09507(.I(new_n9630_), .ZN(new_n9765_));
  NOR3_X1    g09508(.A1(new_n9761_), .A2(new_n9760_), .A3(new_n9758_), .ZN(new_n9766_));
  AOI21_X1   g09509(.A1(new_n9747_), .A2(new_n9753_), .B(new_n9762_), .ZN(new_n9767_));
  OAI21_X1   g09510(.A1(new_n9766_), .A2(new_n9767_), .B(new_n9765_), .ZN(new_n9768_));
  OAI22_X1   g09511(.A1(new_n3298_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n3293_), .ZN(new_n9769_));
  NAND2_X1   g09512(.A1(new_n4227_), .A2(\b[27] ), .ZN(new_n9770_));
  AOI21_X1   g09513(.A1(new_n9769_), .A2(new_n9770_), .B(new_n3301_), .ZN(new_n9771_));
  NAND2_X1   g09514(.A1(new_n2276_), .A2(new_n9771_), .ZN(new_n9772_));
  XOR2_X1    g09515(.A1(new_n9772_), .A2(\a[38] ), .Z(new_n9773_));
  AOI21_X1   g09516(.A1(new_n9764_), .A2(new_n9768_), .B(new_n9773_), .ZN(new_n9774_));
  OAI21_X1   g09517(.A1(new_n9761_), .A2(new_n9760_), .B(new_n9762_), .ZN(new_n9775_));
  NAND3_X1   g09518(.A1(new_n9747_), .A2(new_n9753_), .A3(new_n9758_), .ZN(new_n9776_));
  AOI21_X1   g09519(.A1(new_n9775_), .A2(new_n9776_), .B(new_n9765_), .ZN(new_n9777_));
  NAND3_X1   g09520(.A1(new_n9747_), .A2(new_n9753_), .A3(new_n9762_), .ZN(new_n9778_));
  OAI21_X1   g09521(.A1(new_n9761_), .A2(new_n9760_), .B(new_n9758_), .ZN(new_n9779_));
  AOI21_X1   g09522(.A1(new_n9779_), .A2(new_n9778_), .B(new_n9630_), .ZN(new_n9780_));
  INV_X1     g09523(.I(new_n9773_), .ZN(new_n9781_));
  NOR3_X1    g09524(.A1(new_n9777_), .A2(new_n9780_), .A3(new_n9781_), .ZN(new_n9782_));
  OAI21_X1   g09525(.A1(new_n9774_), .A2(new_n9782_), .B(new_n9457_), .ZN(new_n9783_));
  NOR3_X1    g09526(.A1(new_n9777_), .A2(new_n9780_), .A3(new_n9773_), .ZN(new_n9784_));
  AOI21_X1   g09527(.A1(new_n9764_), .A2(new_n9768_), .B(new_n9781_), .ZN(new_n9785_));
  OAI21_X1   g09528(.A1(new_n9785_), .A2(new_n9784_), .B(new_n9466_), .ZN(new_n9786_));
  OAI22_X1   g09529(.A1(new_n2846_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n2841_), .ZN(new_n9787_));
  NAND2_X1   g09530(.A1(new_n3755_), .A2(\b[30] ), .ZN(new_n9788_));
  AOI21_X1   g09531(.A1(new_n9787_), .A2(new_n9788_), .B(new_n2849_), .ZN(new_n9789_));
  NAND2_X1   g09532(.A1(new_n2659_), .A2(new_n9789_), .ZN(new_n9790_));
  XOR2_X1    g09533(.A1(new_n9790_), .A2(\a[35] ), .Z(new_n9791_));
  INV_X1     g09534(.I(new_n9791_), .ZN(new_n9792_));
  NAND3_X1   g09535(.A1(new_n9783_), .A2(new_n9786_), .A3(new_n9792_), .ZN(new_n9793_));
  OAI21_X1   g09536(.A1(new_n9777_), .A2(new_n9780_), .B(new_n9781_), .ZN(new_n9794_));
  NAND3_X1   g09537(.A1(new_n9764_), .A2(new_n9768_), .A3(new_n9773_), .ZN(new_n9795_));
  AOI21_X1   g09538(.A1(new_n9794_), .A2(new_n9795_), .B(new_n9466_), .ZN(new_n9796_));
  NAND3_X1   g09539(.A1(new_n9764_), .A2(new_n9768_), .A3(new_n9781_), .ZN(new_n9797_));
  OAI21_X1   g09540(.A1(new_n9777_), .A2(new_n9780_), .B(new_n9773_), .ZN(new_n9798_));
  AOI21_X1   g09541(.A1(new_n9797_), .A2(new_n9798_), .B(new_n9457_), .ZN(new_n9799_));
  OAI21_X1   g09542(.A1(new_n9796_), .A2(new_n9799_), .B(new_n9791_), .ZN(new_n9800_));
  AOI21_X1   g09543(.A1(new_n9800_), .A2(new_n9793_), .B(new_n9628_), .ZN(new_n9801_));
  OAI21_X1   g09544(.A1(new_n9796_), .A2(new_n9799_), .B(new_n9792_), .ZN(new_n9802_));
  NAND3_X1   g09545(.A1(new_n9783_), .A2(new_n9786_), .A3(new_n9791_), .ZN(new_n9803_));
  AOI21_X1   g09546(.A1(new_n9802_), .A2(new_n9803_), .B(new_n9627_), .ZN(new_n9804_));
  OAI22_X1   g09547(.A1(new_n2452_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n2447_), .ZN(new_n9805_));
  NAND2_X1   g09548(.A1(new_n3312_), .A2(\b[33] ), .ZN(new_n9806_));
  AOI21_X1   g09549(.A1(new_n9805_), .A2(new_n9806_), .B(new_n2455_), .ZN(new_n9807_));
  NAND2_X1   g09550(.A1(new_n3101_), .A2(new_n9807_), .ZN(new_n9808_));
  XOR2_X1    g09551(.A1(new_n9808_), .A2(\a[32] ), .Z(new_n9809_));
  AOI21_X1   g09552(.A1(new_n9479_), .A2(new_n9474_), .B(new_n9809_), .ZN(new_n9810_));
  INV_X1     g09553(.I(new_n9809_), .ZN(new_n9811_));
  NOR2_X1    g09554(.A1(new_n9475_), .A2(new_n9811_), .ZN(new_n9812_));
  OAI22_X1   g09555(.A1(new_n9801_), .A2(new_n9804_), .B1(new_n9810_), .B2(new_n9812_), .ZN(new_n9813_));
  NOR3_X1    g09556(.A1(new_n9796_), .A2(new_n9799_), .A3(new_n9791_), .ZN(new_n9814_));
  AOI21_X1   g09557(.A1(new_n9783_), .A2(new_n9786_), .B(new_n9792_), .ZN(new_n9815_));
  OAI21_X1   g09558(.A1(new_n9814_), .A2(new_n9815_), .B(new_n9627_), .ZN(new_n9816_));
  AOI21_X1   g09559(.A1(new_n9783_), .A2(new_n9786_), .B(new_n9791_), .ZN(new_n9817_));
  NOR3_X1    g09560(.A1(new_n9796_), .A2(new_n9799_), .A3(new_n9792_), .ZN(new_n9818_));
  OAI21_X1   g09561(.A1(new_n9817_), .A2(new_n9818_), .B(new_n9628_), .ZN(new_n9819_));
  NAND3_X1   g09562(.A1(new_n9479_), .A2(new_n9474_), .A3(new_n9811_), .ZN(new_n9820_));
  NAND2_X1   g09563(.A1(new_n9475_), .A2(new_n9809_), .ZN(new_n9821_));
  NAND2_X1   g09564(.A1(new_n9821_), .A2(new_n9820_), .ZN(new_n9822_));
  NAND3_X1   g09565(.A1(new_n9816_), .A2(new_n9819_), .A3(new_n9822_), .ZN(new_n9823_));
  OAI22_X1   g09566(.A1(new_n2084_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n2079_), .ZN(new_n9824_));
  NAND2_X1   g09567(.A1(new_n2864_), .A2(\b[36] ), .ZN(new_n9825_));
  AOI21_X1   g09568(.A1(new_n9824_), .A2(new_n9825_), .B(new_n2087_), .ZN(new_n9826_));
  NAND2_X1   g09569(.A1(new_n3565_), .A2(new_n9826_), .ZN(new_n9827_));
  XOR2_X1    g09570(.A1(new_n9827_), .A2(\a[29] ), .Z(new_n9828_));
  INV_X1     g09571(.I(new_n9828_), .ZN(new_n9829_));
  NAND3_X1   g09572(.A1(new_n9813_), .A2(new_n9823_), .A3(new_n9829_), .ZN(new_n9830_));
  NOR2_X1    g09573(.A1(new_n9812_), .A2(new_n9810_), .ZN(new_n9831_));
  AOI21_X1   g09574(.A1(new_n9816_), .A2(new_n9819_), .B(new_n9831_), .ZN(new_n9832_));
  NOR2_X1    g09575(.A1(new_n9475_), .A2(new_n9809_), .ZN(new_n9833_));
  AOI21_X1   g09576(.A1(new_n9479_), .A2(new_n9474_), .B(new_n9811_), .ZN(new_n9834_));
  NOR2_X1    g09577(.A1(new_n9833_), .A2(new_n9834_), .ZN(new_n9835_));
  NOR3_X1    g09578(.A1(new_n9801_), .A2(new_n9835_), .A3(new_n9804_), .ZN(new_n9836_));
  OAI21_X1   g09579(.A1(new_n9832_), .A2(new_n9836_), .B(new_n9828_), .ZN(new_n9837_));
  NAND2_X1   g09580(.A1(new_n9837_), .A2(new_n9830_), .ZN(new_n9838_));
  INV_X1     g09581(.I(new_n9485_), .ZN(new_n9839_));
  NAND2_X1   g09582(.A1(new_n9509_), .A2(new_n9839_), .ZN(new_n9840_));
  INV_X1     g09583(.I(new_n9486_), .ZN(new_n9841_));
  NAND3_X1   g09584(.A1(new_n9505_), .A2(new_n9841_), .A3(new_n9500_), .ZN(new_n9842_));
  AOI21_X1   g09585(.A1(new_n9840_), .A2(new_n9842_), .B(new_n9838_), .ZN(new_n9843_));
  NOR3_X1    g09586(.A1(new_n9832_), .A2(new_n9836_), .A3(new_n9828_), .ZN(new_n9844_));
  AOI21_X1   g09587(.A1(new_n9813_), .A2(new_n9823_), .B(new_n9829_), .ZN(new_n9845_));
  NOR2_X1    g09588(.A1(new_n9845_), .A2(new_n9844_), .ZN(new_n9846_));
  AOI21_X1   g09589(.A1(new_n9505_), .A2(new_n9500_), .B(new_n9485_), .ZN(new_n9847_));
  NOR2_X1    g09590(.A1(new_n9509_), .A2(new_n9486_), .ZN(new_n9848_));
  NOR3_X1    g09591(.A1(new_n9847_), .A2(new_n9848_), .A3(new_n9846_), .ZN(new_n9849_));
  OAI21_X1   g09592(.A1(new_n9843_), .A2(new_n9849_), .B(new_n9626_), .ZN(new_n9850_));
  NAND2_X1   g09593(.A1(new_n9509_), .A2(new_n9489_), .ZN(new_n9851_));
  NAND3_X1   g09594(.A1(new_n9505_), .A2(new_n9488_), .A3(new_n9500_), .ZN(new_n9852_));
  AOI21_X1   g09595(.A1(new_n9851_), .A2(new_n9852_), .B(new_n9495_), .ZN(new_n9853_));
  OAI21_X1   g09596(.A1(new_n9847_), .A2(new_n9848_), .B(new_n9846_), .ZN(new_n9854_));
  NAND3_X1   g09597(.A1(new_n9840_), .A2(new_n9842_), .A3(new_n9838_), .ZN(new_n9855_));
  NAND3_X1   g09598(.A1(new_n9853_), .A2(new_n9854_), .A3(new_n9855_), .ZN(new_n9856_));
  AOI21_X1   g09599(.A1(new_n9850_), .A2(new_n9856_), .B(new_n9623_), .ZN(new_n9857_));
  AOI21_X1   g09600(.A1(new_n9854_), .A2(new_n9855_), .B(new_n9853_), .ZN(new_n9858_));
  NOR3_X1    g09601(.A1(new_n9626_), .A2(new_n9843_), .A3(new_n9849_), .ZN(new_n9859_));
  NOR3_X1    g09602(.A1(new_n9859_), .A2(new_n9858_), .A3(new_n9622_), .ZN(new_n9860_));
  OAI21_X1   g09603(.A1(new_n9860_), .A2(new_n9857_), .B(new_n9617_), .ZN(new_n9861_));
  INV_X1     g09604(.I(new_n9617_), .ZN(new_n9862_));
  OAI21_X1   g09605(.A1(new_n9859_), .A2(new_n9858_), .B(new_n9622_), .ZN(new_n9863_));
  NAND3_X1   g09606(.A1(new_n9850_), .A2(new_n9856_), .A3(new_n9623_), .ZN(new_n9864_));
  NAND3_X1   g09607(.A1(new_n9863_), .A2(new_n9864_), .A3(new_n9862_), .ZN(new_n9865_));
  AOI21_X1   g09608(.A1(new_n9511_), .A2(new_n9514_), .B(new_n9349_), .ZN(new_n9866_));
  NAND3_X1   g09609(.A1(new_n9861_), .A2(new_n9865_), .A3(new_n9866_), .ZN(new_n9867_));
  AOI21_X1   g09610(.A1(new_n9863_), .A2(new_n9864_), .B(new_n9862_), .ZN(new_n9868_));
  NOR3_X1    g09611(.A1(new_n9860_), .A2(new_n9857_), .A3(new_n9617_), .ZN(new_n9869_));
  INV_X1     g09612(.I(new_n9866_), .ZN(new_n9870_));
  OAI21_X1   g09613(.A1(new_n9869_), .A2(new_n9868_), .B(new_n9870_), .ZN(new_n9871_));
  OAI22_X1   g09614(.A1(new_n1168_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n1163_), .ZN(new_n9872_));
  NAND2_X1   g09615(.A1(new_n1774_), .A2(\b[45] ), .ZN(new_n9873_));
  AOI21_X1   g09616(.A1(new_n9872_), .A2(new_n9873_), .B(new_n1171_), .ZN(new_n9874_));
  NAND2_X1   g09617(.A1(new_n5004_), .A2(new_n9874_), .ZN(new_n9875_));
  XOR2_X1    g09618(.A1(new_n9875_), .A2(\a[20] ), .Z(new_n9876_));
  INV_X1     g09619(.I(new_n9876_), .ZN(new_n9877_));
  NAND3_X1   g09620(.A1(new_n9871_), .A2(new_n9867_), .A3(new_n9877_), .ZN(new_n9878_));
  NOR3_X1    g09621(.A1(new_n9869_), .A2(new_n9868_), .A3(new_n9870_), .ZN(new_n9879_));
  AOI21_X1   g09622(.A1(new_n9861_), .A2(new_n9865_), .B(new_n9866_), .ZN(new_n9880_));
  OAI21_X1   g09623(.A1(new_n9879_), .A2(new_n9880_), .B(new_n9876_), .ZN(new_n9881_));
  NAND3_X1   g09624(.A1(new_n9538_), .A2(new_n9237_), .A3(new_n9534_), .ZN(new_n9882_));
  NOR3_X1    g09625(.A1(new_n9518_), .A2(new_n9515_), .A3(new_n9520_), .ZN(new_n9883_));
  NAND4_X1   g09626(.A1(new_n9882_), .A2(new_n9881_), .A3(new_n9878_), .A4(new_n9883_), .ZN(new_n9884_));
  NOR3_X1    g09627(.A1(new_n9879_), .A2(new_n9880_), .A3(new_n9876_), .ZN(new_n9885_));
  AOI21_X1   g09628(.A1(new_n9871_), .A2(new_n9867_), .B(new_n9877_), .ZN(new_n9886_));
  NOR3_X1    g09629(.A1(new_n9339_), .A2(new_n9338_), .A3(new_n9524_), .ZN(new_n9887_));
  INV_X1     g09630(.I(new_n9883_), .ZN(new_n9888_));
  OAI22_X1   g09631(.A1(new_n9887_), .A2(new_n9888_), .B1(new_n9885_), .B2(new_n9886_), .ZN(new_n9889_));
  OAI22_X1   g09632(.A1(new_n940_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n935_), .ZN(new_n9890_));
  NAND2_X1   g09633(.A1(new_n1458_), .A2(\b[48] ), .ZN(new_n9891_));
  AOI21_X1   g09634(.A1(new_n9890_), .A2(new_n9891_), .B(new_n943_), .ZN(new_n9892_));
  NAND2_X1   g09635(.A1(new_n5537_), .A2(new_n9892_), .ZN(new_n9893_));
  XOR2_X1    g09636(.A1(new_n9893_), .A2(\a[17] ), .Z(new_n9894_));
  INV_X1     g09637(.I(new_n9894_), .ZN(new_n9895_));
  NAND3_X1   g09638(.A1(new_n9889_), .A2(new_n9884_), .A3(new_n9895_), .ZN(new_n9896_));
  NOR4_X1    g09639(.A1(new_n9887_), .A2(new_n9885_), .A3(new_n9886_), .A4(new_n9888_), .ZN(new_n9897_));
  AOI22_X1   g09640(.A1(new_n9882_), .A2(new_n9883_), .B1(new_n9881_), .B2(new_n9878_), .ZN(new_n9898_));
  OAI21_X1   g09641(.A1(new_n9898_), .A2(new_n9897_), .B(new_n9894_), .ZN(new_n9899_));
  AOI21_X1   g09642(.A1(new_n9899_), .A2(new_n9896_), .B(new_n9612_), .ZN(new_n9900_));
  NAND3_X1   g09643(.A1(new_n9538_), .A2(new_n9237_), .A3(new_n9524_), .ZN(new_n9901_));
  OAI21_X1   g09644(.A1(new_n9339_), .A2(new_n9338_), .B(new_n9534_), .ZN(new_n9902_));
  AOI21_X1   g09645(.A1(new_n9901_), .A2(new_n9902_), .B(new_n9530_), .ZN(new_n9903_));
  NOR2_X1    g09646(.A1(new_n9903_), .A2(new_n9555_), .ZN(new_n9904_));
  OAI21_X1   g09647(.A1(new_n9898_), .A2(new_n9897_), .B(new_n9895_), .ZN(new_n9905_));
  NAND3_X1   g09648(.A1(new_n9889_), .A2(new_n9884_), .A3(new_n9894_), .ZN(new_n9906_));
  AOI21_X1   g09649(.A1(new_n9905_), .A2(new_n9906_), .B(new_n9904_), .ZN(new_n9907_));
  OAI22_X1   g09650(.A1(new_n757_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n752_), .ZN(new_n9908_));
  NAND2_X1   g09651(.A1(new_n1182_), .A2(\b[51] ), .ZN(new_n9909_));
  AOI21_X1   g09652(.A1(new_n9908_), .A2(new_n9909_), .B(new_n760_), .ZN(new_n9910_));
  NAND2_X1   g09653(.A1(new_n6219_), .A2(new_n9910_), .ZN(new_n9911_));
  XOR2_X1    g09654(.A1(new_n9911_), .A2(\a[14] ), .Z(new_n9912_));
  NOR3_X1    g09655(.A1(new_n9900_), .A2(new_n9907_), .A3(new_n9912_), .ZN(new_n9913_));
  NOR3_X1    g09656(.A1(new_n9898_), .A2(new_n9897_), .A3(new_n9894_), .ZN(new_n9914_));
  AOI21_X1   g09657(.A1(new_n9889_), .A2(new_n9884_), .B(new_n9895_), .ZN(new_n9915_));
  OAI21_X1   g09658(.A1(new_n9914_), .A2(new_n9915_), .B(new_n9904_), .ZN(new_n9916_));
  AOI21_X1   g09659(.A1(new_n9889_), .A2(new_n9884_), .B(new_n9894_), .ZN(new_n9917_));
  NOR3_X1    g09660(.A1(new_n9898_), .A2(new_n9897_), .A3(new_n9895_), .ZN(new_n9918_));
  OAI21_X1   g09661(.A1(new_n9918_), .A2(new_n9917_), .B(new_n9612_), .ZN(new_n9919_));
  INV_X1     g09662(.I(new_n9912_), .ZN(new_n9920_));
  AOI21_X1   g09663(.A1(new_n9916_), .A2(new_n9919_), .B(new_n9920_), .ZN(new_n9921_));
  NOR2_X1    g09664(.A1(new_n9544_), .A2(new_n9549_), .ZN(new_n9922_));
  INV_X1     g09665(.I(new_n9922_), .ZN(new_n9923_));
  NOR3_X1    g09666(.A1(new_n9921_), .A2(new_n9913_), .A3(new_n9923_), .ZN(new_n9924_));
  NAND3_X1   g09667(.A1(new_n9916_), .A2(new_n9919_), .A3(new_n9920_), .ZN(new_n9925_));
  OAI21_X1   g09668(.A1(new_n9900_), .A2(new_n9907_), .B(new_n9912_), .ZN(new_n9926_));
  AOI21_X1   g09669(.A1(new_n9926_), .A2(new_n9925_), .B(new_n9922_), .ZN(new_n9927_));
  OAI22_X1   g09670(.A1(new_n437_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n431_), .ZN(new_n9928_));
  NAND2_X1   g09671(.A1(new_n775_), .A2(\b[57] ), .ZN(new_n9929_));
  AOI21_X1   g09672(.A1(new_n9928_), .A2(new_n9929_), .B(new_n440_), .ZN(new_n9930_));
  NAND2_X1   g09673(.A1(new_n7895_), .A2(new_n9930_), .ZN(new_n9931_));
  NOR2_X1    g09674(.A1(new_n9931_), .A2(\a[8] ), .ZN(new_n9932_));
  NAND2_X1   g09675(.A1(new_n9931_), .A2(\a[8] ), .ZN(new_n9933_));
  INV_X1     g09676(.I(new_n9933_), .ZN(new_n9934_));
  OAI22_X1   g09677(.A1(new_n582_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n577_), .ZN(new_n9935_));
  NAND2_X1   g09678(.A1(new_n960_), .A2(\b[54] ), .ZN(new_n9936_));
  AOI21_X1   g09679(.A1(new_n9935_), .A2(new_n9936_), .B(new_n585_), .ZN(new_n9937_));
  NAND2_X1   g09680(.A1(new_n6994_), .A2(new_n9937_), .ZN(new_n9938_));
  XOR2_X1    g09681(.A1(new_n9938_), .A2(\a[11] ), .Z(new_n9939_));
  NOR3_X1    g09682(.A1(new_n9934_), .A2(new_n9932_), .A3(new_n9939_), .ZN(new_n9940_));
  INV_X1     g09683(.I(new_n9932_), .ZN(new_n9941_));
  INV_X1     g09684(.I(new_n9939_), .ZN(new_n9942_));
  AOI21_X1   g09685(.A1(new_n9941_), .A2(new_n9933_), .B(new_n9942_), .ZN(new_n9943_));
  OAI22_X1   g09686(.A1(new_n9927_), .A2(new_n9924_), .B1(new_n9940_), .B2(new_n9943_), .ZN(new_n9944_));
  NAND3_X1   g09687(.A1(new_n9926_), .A2(new_n9925_), .A3(new_n9922_), .ZN(new_n9945_));
  OAI21_X1   g09688(.A1(new_n9921_), .A2(new_n9913_), .B(new_n9923_), .ZN(new_n9946_));
  AOI21_X1   g09689(.A1(new_n9941_), .A2(new_n9933_), .B(new_n9939_), .ZN(new_n9947_));
  NOR3_X1    g09690(.A1(new_n9934_), .A2(new_n9932_), .A3(new_n9942_), .ZN(new_n9948_));
  NOR2_X1    g09691(.A1(new_n9947_), .A2(new_n9948_), .ZN(new_n9949_));
  INV_X1     g09692(.I(new_n9949_), .ZN(new_n9950_));
  NAND3_X1   g09693(.A1(new_n9946_), .A2(new_n9945_), .A3(new_n9950_), .ZN(new_n9951_));
  NAND2_X1   g09694(.A1(new_n9944_), .A2(new_n9951_), .ZN(new_n9952_));
  NAND3_X1   g09695(.A1(new_n9608_), .A2(new_n9952_), .A3(new_n9605_), .ZN(new_n9953_));
  INV_X1     g09696(.I(new_n8525_), .ZN(new_n9954_));
  NAND3_X1   g09697(.A1(new_n8286_), .A2(new_n8258_), .A3(new_n8531_), .ZN(new_n9955_));
  OAI21_X1   g09698(.A1(new_n8900_), .A2(new_n8898_), .B(new_n8530_), .ZN(new_n9956_));
  AOI21_X1   g09699(.A1(new_n9955_), .A2(new_n9956_), .B(new_n9954_), .ZN(new_n9957_));
  NOR3_X1    g09700(.A1(new_n8890_), .A2(new_n8891_), .A3(new_n8887_), .ZN(new_n9958_));
  AOI21_X1   g09701(.A1(new_n8882_), .A2(new_n8879_), .B(new_n8888_), .ZN(new_n9959_));
  OAI21_X1   g09702(.A1(new_n9958_), .A2(new_n9959_), .B(new_n8521_), .ZN(new_n9960_));
  AOI21_X1   g09703(.A1(new_n8882_), .A2(new_n8879_), .B(new_n8887_), .ZN(new_n9961_));
  NOR3_X1    g09704(.A1(new_n8890_), .A2(new_n8891_), .A3(new_n8888_), .ZN(new_n9962_));
  OAI21_X1   g09705(.A1(new_n9962_), .A2(new_n9961_), .B(new_n8584_), .ZN(new_n9963_));
  NAND3_X1   g09706(.A1(new_n9960_), .A2(new_n9963_), .A3(new_n8905_), .ZN(new_n9964_));
  NAND2_X1   g09707(.A1(new_n9964_), .A2(new_n9957_), .ZN(new_n9965_));
  NAND3_X1   g09708(.A1(new_n9293_), .A2(new_n9965_), .A3(new_n9299_), .ZN(new_n9966_));
  AOI21_X1   g09709(.A1(new_n9966_), .A2(new_n9290_), .B(new_n9606_), .ZN(new_n9967_));
  NOR2_X1    g09710(.A1(new_n9943_), .A2(new_n9940_), .ZN(new_n9968_));
  AOI21_X1   g09711(.A1(new_n9946_), .A2(new_n9945_), .B(new_n9968_), .ZN(new_n9969_));
  NOR3_X1    g09712(.A1(new_n9927_), .A2(new_n9924_), .A3(new_n9949_), .ZN(new_n9970_));
  NOR2_X1    g09713(.A1(new_n9970_), .A2(new_n9969_), .ZN(new_n9971_));
  OAI21_X1   g09714(.A1(new_n9967_), .A2(new_n9604_), .B(new_n9971_), .ZN(new_n9972_));
  NAND2_X1   g09715(.A1(new_n9972_), .A2(new_n9953_), .ZN(new_n9973_));
  INV_X1     g09716(.I(new_n9335_), .ZN(new_n9974_));
  NOR2_X1    g09717(.A1(new_n9974_), .A2(new_n9573_), .ZN(new_n9975_));
  INV_X1     g09718(.I(new_n9975_), .ZN(new_n9976_));
  NAND2_X1   g09719(.A1(new_n9974_), .A2(new_n9573_), .ZN(new_n9977_));
  NOR2_X1    g09720(.A1(new_n9337_), .A2(new_n9568_), .ZN(new_n9978_));
  INV_X1     g09721(.I(new_n9568_), .ZN(new_n9979_));
  AOI21_X1   g09722(.A1(new_n9966_), .A2(new_n9290_), .B(new_n9979_), .ZN(new_n9980_));
  OAI21_X1   g09723(.A1(new_n9980_), .A2(new_n9978_), .B(new_n9977_), .ZN(new_n9981_));
  NAND2_X1   g09724(.A1(new_n9981_), .A2(new_n9976_), .ZN(new_n9982_));
  XOR2_X1    g09725(.A1(new_n9982_), .A2(new_n9973_), .Z(new_n9983_));
  XOR2_X1    g09726(.A1(new_n9983_), .A2(new_n9603_), .Z(new_n9984_));
  XOR2_X1    g09727(.A1(new_n9984_), .A2(new_n9598_), .Z(new_n9985_));
  AOI21_X1   g09728(.A1(new_n9580_), .A2(new_n9578_), .B(new_n9327_), .ZN(new_n9986_));
  XOR2_X1    g09729(.A1(new_n9577_), .A2(new_n9974_), .Z(new_n9987_));
  NOR2_X1    g09730(.A1(new_n9581_), .A2(new_n9328_), .ZN(new_n9988_));
  AOI21_X1   g09731(.A1(new_n9988_), .A2(new_n9987_), .B(new_n9986_), .ZN(new_n9989_));
  OR2_X2     g09732(.A1(new_n9985_), .A2(new_n9989_), .Z(new_n9990_));
  NAND2_X1   g09733(.A1(new_n9985_), .A2(new_n9989_), .ZN(new_n9991_));
  NAND2_X1   g09734(.A1(new_n9990_), .A2(new_n9991_), .ZN(\f[65] ));
  NOR2_X1    g09735(.A1(new_n9971_), .A2(new_n9603_), .ZN(new_n9993_));
  AOI22_X1   g09736(.A1(new_n9608_), .A2(new_n9605_), .B1(new_n9971_), .B2(new_n9603_), .ZN(new_n9994_));
  AOI22_X1   g09737(.A1(\b[63] ), .A2(new_n315_), .B1(new_n321_), .B2(\b[62] ), .ZN(new_n9995_));
  NOR2_X1    g09738(.A1(new_n362_), .A2(new_n8548_), .ZN(new_n9996_));
  OAI21_X1   g09739(.A1(new_n9995_), .A2(new_n9996_), .B(new_n311_), .ZN(new_n9997_));
  NOR3_X1    g09740(.A1(new_n8962_), .A2(\a[5] ), .A3(new_n9997_), .ZN(new_n9998_));
  OAI21_X1   g09741(.A1(new_n8962_), .A2(new_n9997_), .B(\a[5] ), .ZN(new_n9999_));
  INV_X1     g09742(.I(new_n9999_), .ZN(new_n10000_));
  NOR2_X1    g09743(.A1(new_n10000_), .A2(new_n9998_), .ZN(new_n10001_));
  INV_X1     g09744(.I(new_n10001_), .ZN(new_n10002_));
  OAI21_X1   g09745(.A1(new_n9994_), .A2(new_n9993_), .B(new_n10002_), .ZN(new_n10003_));
  INV_X1     g09746(.I(new_n9603_), .ZN(new_n10004_));
  NAND2_X1   g09747(.A1(new_n9952_), .A2(new_n10004_), .ZN(new_n10005_));
  NAND3_X1   g09748(.A1(new_n9944_), .A2(new_n9603_), .A3(new_n9951_), .ZN(new_n10006_));
  OAI21_X1   g09749(.A1(new_n9604_), .A2(new_n9967_), .B(new_n10006_), .ZN(new_n10007_));
  NAND3_X1   g09750(.A1(new_n10007_), .A2(new_n10005_), .A3(new_n10001_), .ZN(new_n10008_));
  NAND2_X1   g09751(.A1(new_n10003_), .A2(new_n10008_), .ZN(new_n10009_));
  NAND3_X1   g09752(.A1(new_n9972_), .A2(new_n9953_), .A3(new_n10004_), .ZN(new_n10010_));
  NOR3_X1    g09753(.A1(new_n9967_), .A2(new_n9971_), .A3(new_n9604_), .ZN(new_n10011_));
  AOI21_X1   g09754(.A1(new_n9337_), .A2(new_n9607_), .B(new_n9604_), .ZN(new_n10012_));
  NOR2_X1    g09755(.A1(new_n10012_), .A2(new_n9952_), .ZN(new_n10013_));
  OAI21_X1   g09756(.A1(new_n10011_), .A2(new_n10013_), .B(new_n9603_), .ZN(new_n10014_));
  NAND2_X1   g09757(.A1(new_n10014_), .A2(new_n10010_), .ZN(new_n10015_));
  NAND3_X1   g09758(.A1(new_n9966_), .A2(new_n9290_), .A3(new_n9979_), .ZN(new_n10016_));
  NAND2_X1   g09759(.A1(new_n9337_), .A2(new_n9568_), .ZN(new_n10017_));
  NAND2_X1   g09760(.A1(new_n10016_), .A2(new_n10017_), .ZN(new_n10018_));
  AOI21_X1   g09761(.A1(new_n10018_), .A2(new_n9977_), .B(new_n9975_), .ZN(new_n10019_));
  NOR3_X1    g09762(.A1(new_n10011_), .A2(new_n10013_), .A3(new_n9603_), .ZN(new_n10020_));
  AOI21_X1   g09763(.A1(new_n9972_), .A2(new_n9953_), .B(new_n10004_), .ZN(new_n10021_));
  OAI21_X1   g09764(.A1(new_n10021_), .A2(new_n10020_), .B(new_n10019_), .ZN(new_n10022_));
  NAND3_X1   g09765(.A1(new_n10014_), .A2(new_n10010_), .A3(new_n9982_), .ZN(new_n10023_));
  AOI22_X1   g09766(.A1(new_n10022_), .A2(new_n10023_), .B1(new_n10015_), .B2(new_n9598_), .ZN(new_n10024_));
  AOI21_X1   g09767(.A1(new_n9627_), .A2(new_n9800_), .B(new_n9814_), .ZN(new_n10025_));
  AOI21_X1   g09768(.A1(new_n9457_), .A2(new_n9798_), .B(new_n9784_), .ZN(new_n10026_));
  NOR2_X1    g09769(.A1(new_n9767_), .A2(new_n9765_), .ZN(new_n10027_));
  OAI21_X1   g09770(.A1(new_n9740_), .A2(new_n9739_), .B(new_n9734_), .ZN(new_n10028_));
  NAND2_X1   g09771(.A1(new_n9728_), .A2(new_n9737_), .ZN(new_n10029_));
  NAND2_X1   g09772(.A1(new_n9750_), .A2(new_n9741_), .ZN(new_n10030_));
  NAND2_X1   g09773(.A1(new_n10029_), .A2(new_n10030_), .ZN(new_n10031_));
  NAND4_X1   g09774(.A1(new_n10031_), .A2(new_n9733_), .A3(new_n9735_), .A4(new_n9736_), .ZN(new_n10032_));
  NAND2_X1   g09775(.A1(new_n10032_), .A2(new_n10028_), .ZN(new_n10033_));
  AOI21_X1   g09776(.A1(new_n9749_), .A2(new_n9737_), .B(new_n9720_), .ZN(new_n10034_));
  OAI21_X1   g09777(.A1(new_n9633_), .A2(new_n9724_), .B(new_n9712_), .ZN(new_n10035_));
  INV_X1     g09778(.I(new_n9694_), .ZN(new_n10036_));
  OAI21_X1   g09779(.A1(new_n9636_), .A2(new_n10036_), .B(new_n9692_), .ZN(new_n10037_));
  NAND2_X1   g09780(.A1(new_n9683_), .A2(new_n9638_), .ZN(new_n10038_));
  NAND2_X1   g09781(.A1(new_n10038_), .A2(new_n9682_), .ZN(new_n10039_));
  INV_X1     g09782(.I(new_n10039_), .ZN(new_n10040_));
  NAND2_X1   g09783(.A1(new_n9641_), .A2(new_n9670_), .ZN(new_n10041_));
  INV_X1     g09784(.I(new_n9657_), .ZN(new_n10042_));
  OAI21_X1   g09785(.A1(new_n9642_), .A2(new_n9659_), .B(new_n10042_), .ZN(new_n10043_));
  INV_X1     g09786(.I(new_n10043_), .ZN(new_n10044_));
  NOR2_X1    g09787(.A1(new_n8317_), .A2(new_n347_), .ZN(new_n10045_));
  NOR2_X1    g09788(.A1(new_n8312_), .A2(new_n403_), .ZN(new_n10046_));
  OAI22_X1   g09789(.A1(new_n10045_), .A2(new_n10046_), .B1(new_n8622_), .B2(new_n393_), .ZN(new_n10047_));
  NAND3_X1   g09790(.A1(new_n402_), .A2(new_n8320_), .A3(new_n10047_), .ZN(new_n10048_));
  XOR2_X1    g09791(.A1(new_n10048_), .A2(new_n8309_), .Z(new_n10049_));
  NOR3_X1    g09792(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n292_), .ZN(new_n10050_));
  NOR2_X1    g09793(.A1(new_n9364_), .A2(new_n292_), .ZN(new_n10051_));
  NOR3_X1    g09794(.A1(new_n10051_), .A2(new_n290_), .A3(new_n8985_), .ZN(new_n10052_));
  NOR2_X1    g09795(.A1(new_n10052_), .A2(new_n10050_), .ZN(new_n10053_));
  NOR2_X1    g09796(.A1(new_n10053_), .A2(new_n271_), .ZN(new_n10054_));
  INV_X1     g09797(.I(new_n10053_), .ZN(new_n10055_));
  NOR2_X1    g09798(.A1(new_n10055_), .A2(\a[2] ), .ZN(new_n10056_));
  OAI21_X1   g09799(.A1(new_n10054_), .A2(new_n10056_), .B(new_n10049_), .ZN(new_n10057_));
  NOR2_X1    g09800(.A1(new_n10055_), .A2(new_n271_), .ZN(new_n10058_));
  NOR2_X1    g09801(.A1(new_n10053_), .A2(\a[2] ), .ZN(new_n10059_));
  NOR2_X1    g09802(.A1(new_n10058_), .A2(new_n10059_), .ZN(new_n10060_));
  OAI21_X1   g09803(.A1(new_n10049_), .A2(new_n10060_), .B(new_n10057_), .ZN(new_n10061_));
  OAI22_X1   g09804(.A1(new_n510_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n495_), .ZN(new_n10062_));
  NAND2_X1   g09805(.A1(new_n8628_), .A2(\b[7] ), .ZN(new_n10063_));
  AOI21_X1   g09806(.A1(new_n10063_), .A2(new_n10062_), .B(new_n7354_), .ZN(new_n10064_));
  NAND2_X1   g09807(.A1(new_n518_), .A2(new_n10064_), .ZN(new_n10065_));
  XOR2_X1    g09808(.A1(new_n10065_), .A2(new_n7343_), .Z(new_n10066_));
  INV_X1     g09809(.I(new_n10066_), .ZN(new_n10067_));
  NOR2_X1    g09810(.A1(new_n10067_), .A2(new_n10061_), .ZN(new_n10068_));
  INV_X1     g09811(.I(new_n10068_), .ZN(new_n10069_));
  NAND2_X1   g09812(.A1(new_n10067_), .A2(new_n10061_), .ZN(new_n10070_));
  AOI21_X1   g09813(.A1(new_n10069_), .A2(new_n10070_), .B(new_n10044_), .ZN(new_n10071_));
  XOR2_X1    g09814(.A1(new_n10066_), .A2(new_n10061_), .Z(new_n10072_));
  NOR2_X1    g09815(.A1(new_n10072_), .A2(new_n10043_), .ZN(new_n10073_));
  NOR2_X1    g09816(.A1(new_n10071_), .A2(new_n10073_), .ZN(new_n10074_));
  OAI22_X1   g09817(.A1(new_n6721_), .A2(new_n659_), .B1(new_n6723_), .B2(new_n717_), .ZN(new_n10075_));
  NAND2_X1   g09818(.A1(new_n7617_), .A2(\b[10] ), .ZN(new_n10076_));
  AOI21_X1   g09819(.A1(new_n10076_), .A2(new_n10075_), .B(new_n6731_), .ZN(new_n10077_));
  NAND2_X1   g09820(.A1(new_n716_), .A2(new_n10077_), .ZN(new_n10078_));
  XOR2_X1    g09821(.A1(new_n10078_), .A2(new_n6516_), .Z(new_n10079_));
  NAND2_X1   g09822(.A1(new_n10074_), .A2(new_n10079_), .ZN(new_n10080_));
  INV_X1     g09823(.I(new_n10074_), .ZN(new_n10081_));
  INV_X1     g09824(.I(new_n10079_), .ZN(new_n10082_));
  NAND2_X1   g09825(.A1(new_n10081_), .A2(new_n10082_), .ZN(new_n10083_));
  AOI22_X1   g09826(.A1(new_n10083_), .A2(new_n10080_), .B1(new_n9669_), .B2(new_n10041_), .ZN(new_n10084_));
  NAND2_X1   g09827(.A1(new_n10041_), .A2(new_n9669_), .ZN(new_n10085_));
  NAND2_X1   g09828(.A1(new_n10081_), .A2(new_n10079_), .ZN(new_n10086_));
  NAND2_X1   g09829(.A1(new_n10074_), .A2(new_n10082_), .ZN(new_n10087_));
  AOI21_X1   g09830(.A1(new_n10086_), .A2(new_n10087_), .B(new_n10085_), .ZN(new_n10088_));
  NOR2_X1    g09831(.A1(new_n10084_), .A2(new_n10088_), .ZN(new_n10089_));
  INV_X1     g09832(.I(new_n10089_), .ZN(new_n10090_));
  OAI22_X1   g09833(.A1(new_n5786_), .A2(new_n904_), .B1(new_n848_), .B2(new_n5792_), .ZN(new_n10091_));
  NAND2_X1   g09834(.A1(new_n6745_), .A2(\b[13] ), .ZN(new_n10092_));
  AOI21_X1   g09835(.A1(new_n10092_), .A2(new_n10091_), .B(new_n5796_), .ZN(new_n10093_));
  NAND2_X1   g09836(.A1(new_n907_), .A2(new_n10093_), .ZN(new_n10094_));
  XOR2_X1    g09837(.A1(new_n10094_), .A2(\a[53] ), .Z(new_n10095_));
  NOR2_X1    g09838(.A1(new_n10090_), .A2(new_n10095_), .ZN(new_n10096_));
  INV_X1     g09839(.I(new_n10096_), .ZN(new_n10097_));
  NAND2_X1   g09840(.A1(new_n10090_), .A2(new_n10095_), .ZN(new_n10098_));
  AOI21_X1   g09841(.A1(new_n10097_), .A2(new_n10098_), .B(new_n10040_), .ZN(new_n10099_));
  XOR2_X1    g09842(.A1(new_n10089_), .A2(new_n10095_), .Z(new_n10100_));
  NOR2_X1    g09843(.A1(new_n10100_), .A2(new_n10039_), .ZN(new_n10101_));
  OAI22_X1   g09844(.A1(new_n5228_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n5225_), .ZN(new_n10102_));
  NAND2_X1   g09845(.A1(new_n5387_), .A2(\b[16] ), .ZN(new_n10103_));
  AOI21_X1   g09846(.A1(new_n10102_), .A2(new_n10103_), .B(new_n5231_), .ZN(new_n10104_));
  NAND2_X1   g09847(.A1(new_n1123_), .A2(new_n10104_), .ZN(new_n10105_));
  XOR2_X1    g09848(.A1(new_n10105_), .A2(\a[50] ), .Z(new_n10106_));
  INV_X1     g09849(.I(new_n10106_), .ZN(new_n10107_));
  OAI21_X1   g09850(.A1(new_n10099_), .A2(new_n10101_), .B(new_n10107_), .ZN(new_n10108_));
  INV_X1     g09851(.I(new_n10099_), .ZN(new_n10109_));
  INV_X1     g09852(.I(new_n10101_), .ZN(new_n10110_));
  NAND3_X1   g09853(.A1(new_n10109_), .A2(new_n10110_), .A3(new_n10106_), .ZN(new_n10111_));
  NAND2_X1   g09854(.A1(new_n10111_), .A2(new_n10108_), .ZN(new_n10112_));
  NAND2_X1   g09855(.A1(new_n10112_), .A2(new_n10037_), .ZN(new_n10113_));
  NAND3_X1   g09856(.A1(new_n10109_), .A2(new_n10110_), .A3(new_n10107_), .ZN(new_n10114_));
  OAI21_X1   g09857(.A1(new_n10099_), .A2(new_n10101_), .B(new_n10106_), .ZN(new_n10115_));
  AOI21_X1   g09858(.A1(new_n10114_), .A2(new_n10115_), .B(new_n10037_), .ZN(new_n10116_));
  INV_X1     g09859(.I(new_n10116_), .ZN(new_n10117_));
  OAI22_X1   g09860(.A1(new_n4711_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n4706_), .ZN(new_n10118_));
  NAND2_X1   g09861(.A1(new_n5814_), .A2(\b[19] ), .ZN(new_n10119_));
  AOI21_X1   g09862(.A1(new_n10118_), .A2(new_n10119_), .B(new_n4714_), .ZN(new_n10120_));
  NAND2_X1   g09863(.A1(new_n1396_), .A2(new_n10120_), .ZN(new_n10121_));
  XOR2_X1    g09864(.A1(new_n10121_), .A2(\a[47] ), .Z(new_n10122_));
  INV_X1     g09865(.I(new_n10122_), .ZN(new_n10123_));
  NAND3_X1   g09866(.A1(new_n10117_), .A2(new_n10113_), .A3(new_n10123_), .ZN(new_n10124_));
  INV_X1     g09867(.I(new_n10037_), .ZN(new_n10125_));
  AOI21_X1   g09868(.A1(new_n10108_), .A2(new_n10111_), .B(new_n10125_), .ZN(new_n10126_));
  OAI21_X1   g09869(.A1(new_n10126_), .A2(new_n10116_), .B(new_n10122_), .ZN(new_n10127_));
  NAND2_X1   g09870(.A1(new_n10124_), .A2(new_n10127_), .ZN(new_n10128_));
  NAND2_X1   g09871(.A1(new_n10128_), .A2(new_n10035_), .ZN(new_n10129_));
  AOI21_X1   g09872(.A1(new_n9632_), .A2(new_n9713_), .B(new_n9723_), .ZN(new_n10130_));
  OAI21_X1   g09873(.A1(new_n10126_), .A2(new_n10116_), .B(new_n10123_), .ZN(new_n10131_));
  INV_X1     g09874(.I(new_n10131_), .ZN(new_n10132_));
  NOR3_X1    g09875(.A1(new_n10126_), .A2(new_n10116_), .A3(new_n10123_), .ZN(new_n10133_));
  OAI21_X1   g09876(.A1(new_n10132_), .A2(new_n10133_), .B(new_n10130_), .ZN(new_n10134_));
  OAI22_X1   g09877(.A1(new_n4208_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n4203_), .ZN(new_n10135_));
  NAND2_X1   g09878(.A1(new_n5244_), .A2(\b[22] ), .ZN(new_n10136_));
  AOI21_X1   g09879(.A1(new_n10135_), .A2(new_n10136_), .B(new_n4211_), .ZN(new_n10137_));
  NAND2_X1   g09880(.A1(new_n1708_), .A2(new_n10137_), .ZN(new_n10138_));
  XOR2_X1    g09881(.A1(new_n10138_), .A2(\a[44] ), .Z(new_n10139_));
  INV_X1     g09882(.I(new_n10139_), .ZN(new_n10140_));
  NAND3_X1   g09883(.A1(new_n10129_), .A2(new_n10134_), .A3(new_n10140_), .ZN(new_n10141_));
  AOI21_X1   g09884(.A1(new_n10127_), .A2(new_n10124_), .B(new_n10130_), .ZN(new_n10142_));
  INV_X1     g09885(.I(new_n10133_), .ZN(new_n10143_));
  AOI21_X1   g09886(.A1(new_n10143_), .A2(new_n10131_), .B(new_n10035_), .ZN(new_n10144_));
  OAI21_X1   g09887(.A1(new_n10144_), .A2(new_n10142_), .B(new_n10139_), .ZN(new_n10145_));
  AOI21_X1   g09888(.A1(new_n10145_), .A2(new_n10141_), .B(new_n10034_), .ZN(new_n10146_));
  OAI21_X1   g09889(.A1(new_n9727_), .A2(new_n9741_), .B(new_n9748_), .ZN(new_n10147_));
  OAI21_X1   g09890(.A1(new_n10144_), .A2(new_n10142_), .B(new_n10140_), .ZN(new_n10148_));
  NAND3_X1   g09891(.A1(new_n10129_), .A2(new_n10134_), .A3(new_n10139_), .ZN(new_n10149_));
  AOI21_X1   g09892(.A1(new_n10148_), .A2(new_n10149_), .B(new_n10147_), .ZN(new_n10150_));
  OAI22_X1   g09893(.A1(new_n3736_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n3731_), .ZN(new_n10151_));
  NAND2_X1   g09894(.A1(new_n4730_), .A2(\b[25] ), .ZN(new_n10152_));
  AOI21_X1   g09895(.A1(new_n10151_), .A2(new_n10152_), .B(new_n3739_), .ZN(new_n10153_));
  NAND2_X1   g09896(.A1(new_n2042_), .A2(new_n10153_), .ZN(new_n10154_));
  XOR2_X1    g09897(.A1(new_n10154_), .A2(\a[41] ), .Z(new_n10155_));
  INV_X1     g09898(.I(new_n10155_), .ZN(new_n10156_));
  OAI21_X1   g09899(.A1(new_n10146_), .A2(new_n10150_), .B(new_n10156_), .ZN(new_n10157_));
  NOR3_X1    g09900(.A1(new_n10144_), .A2(new_n10142_), .A3(new_n10139_), .ZN(new_n10158_));
  AOI21_X1   g09901(.A1(new_n10129_), .A2(new_n10134_), .B(new_n10140_), .ZN(new_n10159_));
  OAI21_X1   g09902(.A1(new_n10158_), .A2(new_n10159_), .B(new_n10147_), .ZN(new_n10160_));
  AOI21_X1   g09903(.A1(new_n10129_), .A2(new_n10134_), .B(new_n10139_), .ZN(new_n10161_));
  NOR3_X1    g09904(.A1(new_n10144_), .A2(new_n10142_), .A3(new_n10140_), .ZN(new_n10162_));
  OAI21_X1   g09905(.A1(new_n10162_), .A2(new_n10161_), .B(new_n10034_), .ZN(new_n10163_));
  NAND3_X1   g09906(.A1(new_n10163_), .A2(new_n10160_), .A3(new_n10155_), .ZN(new_n10164_));
  NAND2_X1   g09907(.A1(new_n10157_), .A2(new_n10164_), .ZN(new_n10165_));
  NAND2_X1   g09908(.A1(new_n10033_), .A2(new_n10165_), .ZN(new_n10166_));
  NAND3_X1   g09909(.A1(new_n10163_), .A2(new_n10160_), .A3(new_n10156_), .ZN(new_n10167_));
  OAI21_X1   g09910(.A1(new_n10146_), .A2(new_n10150_), .B(new_n10155_), .ZN(new_n10168_));
  NAND2_X1   g09911(.A1(new_n10168_), .A2(new_n10167_), .ZN(new_n10169_));
  NAND3_X1   g09912(.A1(new_n10169_), .A2(new_n10028_), .A3(new_n10032_), .ZN(new_n10170_));
  NAND2_X1   g09913(.A1(new_n10166_), .A2(new_n10170_), .ZN(new_n10171_));
  OAI22_X1   g09914(.A1(new_n3298_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n3293_), .ZN(new_n10172_));
  NAND2_X1   g09915(.A1(new_n4227_), .A2(\b[28] ), .ZN(new_n10173_));
  AOI21_X1   g09916(.A1(new_n10172_), .A2(new_n10173_), .B(new_n3301_), .ZN(new_n10174_));
  NAND2_X1   g09917(.A1(new_n2404_), .A2(new_n10174_), .ZN(new_n10175_));
  XOR2_X1    g09918(.A1(new_n10175_), .A2(\a[38] ), .Z(new_n10176_));
  NOR2_X1    g09919(.A1(new_n10171_), .A2(new_n10176_), .ZN(new_n10177_));
  INV_X1     g09920(.I(new_n10176_), .ZN(new_n10178_));
  AOI21_X1   g09921(.A1(new_n10166_), .A2(new_n10170_), .B(new_n10178_), .ZN(new_n10179_));
  OAI22_X1   g09922(.A1(new_n10177_), .A2(new_n10179_), .B1(new_n9766_), .B2(new_n10027_), .ZN(new_n10180_));
  NOR2_X1    g09923(.A1(new_n10027_), .A2(new_n9766_), .ZN(new_n10181_));
  AOI21_X1   g09924(.A1(new_n10166_), .A2(new_n10170_), .B(new_n10176_), .ZN(new_n10182_));
  NOR2_X1    g09925(.A1(new_n10171_), .A2(new_n10178_), .ZN(new_n10183_));
  OAI21_X1   g09926(.A1(new_n10183_), .A2(new_n10182_), .B(new_n10181_), .ZN(new_n10184_));
  OAI22_X1   g09927(.A1(new_n2846_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n2841_), .ZN(new_n10185_));
  NAND2_X1   g09928(.A1(new_n3755_), .A2(\b[31] ), .ZN(new_n10186_));
  AOI21_X1   g09929(.A1(new_n10185_), .A2(new_n10186_), .B(new_n2849_), .ZN(new_n10187_));
  NAND2_X1   g09930(.A1(new_n2797_), .A2(new_n10187_), .ZN(new_n10188_));
  XOR2_X1    g09931(.A1(new_n10188_), .A2(\a[35] ), .Z(new_n10189_));
  INV_X1     g09932(.I(new_n10189_), .ZN(new_n10190_));
  NAND3_X1   g09933(.A1(new_n10180_), .A2(new_n10184_), .A3(new_n10190_), .ZN(new_n10191_));
  AOI21_X1   g09934(.A1(new_n10180_), .A2(new_n10184_), .B(new_n10190_), .ZN(new_n10192_));
  INV_X1     g09935(.I(new_n10192_), .ZN(new_n10193_));
  AOI21_X1   g09936(.A1(new_n10193_), .A2(new_n10191_), .B(new_n10026_), .ZN(new_n10194_));
  INV_X1     g09937(.I(new_n10026_), .ZN(new_n10195_));
  AOI21_X1   g09938(.A1(new_n10180_), .A2(new_n10184_), .B(new_n10189_), .ZN(new_n10196_));
  INV_X1     g09939(.I(new_n10196_), .ZN(new_n10197_));
  NAND3_X1   g09940(.A1(new_n10180_), .A2(new_n10184_), .A3(new_n10189_), .ZN(new_n10198_));
  AOI21_X1   g09941(.A1(new_n10197_), .A2(new_n10198_), .B(new_n10195_), .ZN(new_n10199_));
  OAI22_X1   g09942(.A1(new_n2452_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n2447_), .ZN(new_n10200_));
  NAND2_X1   g09943(.A1(new_n3312_), .A2(\b[34] ), .ZN(new_n10201_));
  AOI21_X1   g09944(.A1(new_n10200_), .A2(new_n10201_), .B(new_n2455_), .ZN(new_n10202_));
  NAND2_X1   g09945(.A1(new_n3246_), .A2(new_n10202_), .ZN(new_n10203_));
  XOR2_X1    g09946(.A1(new_n10203_), .A2(\a[32] ), .Z(new_n10204_));
  INV_X1     g09947(.I(new_n10204_), .ZN(new_n10205_));
  OAI21_X1   g09948(.A1(new_n10199_), .A2(new_n10194_), .B(new_n10205_), .ZN(new_n10206_));
  INV_X1     g09949(.I(new_n10191_), .ZN(new_n10207_));
  OAI21_X1   g09950(.A1(new_n10207_), .A2(new_n10192_), .B(new_n10195_), .ZN(new_n10208_));
  INV_X1     g09951(.I(new_n10198_), .ZN(new_n10209_));
  OAI21_X1   g09952(.A1(new_n10209_), .A2(new_n10196_), .B(new_n10026_), .ZN(new_n10210_));
  NAND3_X1   g09953(.A1(new_n10210_), .A2(new_n10208_), .A3(new_n10204_), .ZN(new_n10211_));
  AOI21_X1   g09954(.A1(new_n10206_), .A2(new_n10211_), .B(new_n10025_), .ZN(new_n10212_));
  INV_X1     g09955(.I(new_n10025_), .ZN(new_n10213_));
  NAND3_X1   g09956(.A1(new_n10210_), .A2(new_n10208_), .A3(new_n10205_), .ZN(new_n10214_));
  OAI21_X1   g09957(.A1(new_n10199_), .A2(new_n10194_), .B(new_n10204_), .ZN(new_n10215_));
  AOI21_X1   g09958(.A1(new_n10215_), .A2(new_n10214_), .B(new_n10213_), .ZN(new_n10216_));
  NOR2_X1    g09959(.A1(new_n10212_), .A2(new_n10216_), .ZN(new_n10217_));
  OAI22_X1   g09960(.A1(new_n2084_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n2079_), .ZN(new_n10218_));
  NAND2_X1   g09961(.A1(new_n2864_), .A2(\b[37] ), .ZN(new_n10219_));
  AOI21_X1   g09962(.A1(new_n10218_), .A2(new_n10219_), .B(new_n2087_), .ZN(new_n10220_));
  NAND2_X1   g09963(.A1(new_n3700_), .A2(new_n10220_), .ZN(new_n10221_));
  XOR2_X1    g09964(.A1(new_n10221_), .A2(\a[29] ), .Z(new_n10222_));
  INV_X1     g09965(.I(new_n10222_), .ZN(new_n10223_));
  NOR3_X1    g09966(.A1(new_n9801_), .A2(new_n9804_), .A3(new_n9811_), .ZN(new_n10224_));
  INV_X1     g09967(.I(new_n10224_), .ZN(new_n10225_));
  NOR3_X1    g09968(.A1(new_n9801_), .A2(new_n9804_), .A3(new_n9809_), .ZN(new_n10226_));
  AOI21_X1   g09969(.A1(new_n9816_), .A2(new_n9819_), .B(new_n9811_), .ZN(new_n10227_));
  OAI21_X1   g09970(.A1(new_n10227_), .A2(new_n10226_), .B(new_n9475_), .ZN(new_n10228_));
  AOI21_X1   g09971(.A1(new_n10228_), .A2(new_n10225_), .B(new_n10223_), .ZN(new_n10229_));
  NAND3_X1   g09972(.A1(new_n9816_), .A2(new_n9819_), .A3(new_n9811_), .ZN(new_n10230_));
  OAI21_X1   g09973(.A1(new_n9801_), .A2(new_n9804_), .B(new_n9809_), .ZN(new_n10231_));
  AOI21_X1   g09974(.A1(new_n10230_), .A2(new_n10231_), .B(new_n9476_), .ZN(new_n10232_));
  NOR3_X1    g09975(.A1(new_n10232_), .A2(new_n10222_), .A3(new_n10224_), .ZN(new_n10233_));
  OAI21_X1   g09976(.A1(new_n10233_), .A2(new_n10229_), .B(new_n10217_), .ZN(new_n10234_));
  AOI21_X1   g09977(.A1(new_n10210_), .A2(new_n10208_), .B(new_n10204_), .ZN(new_n10235_));
  NOR3_X1    g09978(.A1(new_n10199_), .A2(new_n10194_), .A3(new_n10205_), .ZN(new_n10236_));
  OAI21_X1   g09979(.A1(new_n10236_), .A2(new_n10235_), .B(new_n10213_), .ZN(new_n10237_));
  NOR3_X1    g09980(.A1(new_n10199_), .A2(new_n10194_), .A3(new_n10204_), .ZN(new_n10238_));
  AOI21_X1   g09981(.A1(new_n10210_), .A2(new_n10208_), .B(new_n10205_), .ZN(new_n10239_));
  OAI21_X1   g09982(.A1(new_n10238_), .A2(new_n10239_), .B(new_n10025_), .ZN(new_n10240_));
  NAND2_X1   g09983(.A1(new_n10240_), .A2(new_n10237_), .ZN(new_n10241_));
  OAI21_X1   g09984(.A1(new_n10232_), .A2(new_n10224_), .B(new_n10222_), .ZN(new_n10242_));
  NAND3_X1   g09985(.A1(new_n10228_), .A2(new_n10223_), .A3(new_n10225_), .ZN(new_n10243_));
  NAND3_X1   g09986(.A1(new_n10242_), .A2(new_n10241_), .A3(new_n10243_), .ZN(new_n10244_));
  NAND2_X1   g09987(.A1(new_n10234_), .A2(new_n10244_), .ZN(new_n10245_));
  OAI22_X1   g09988(.A1(new_n1760_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n1755_), .ZN(new_n10246_));
  NAND2_X1   g09989(.A1(new_n2470_), .A2(\b[40] ), .ZN(new_n10247_));
  AOI21_X1   g09990(.A1(new_n10246_), .A2(new_n10247_), .B(new_n1763_), .ZN(new_n10248_));
  NAND2_X1   g09991(.A1(new_n4017_), .A2(new_n10248_), .ZN(new_n10249_));
  XOR2_X1    g09992(.A1(new_n10249_), .A2(\a[26] ), .Z(new_n10250_));
  NOR3_X1    g09993(.A1(new_n9847_), .A2(new_n9848_), .A3(new_n9838_), .ZN(new_n10251_));
  OAI21_X1   g09994(.A1(new_n10251_), .A2(new_n9845_), .B(new_n10250_), .ZN(new_n10252_));
  INV_X1     g09995(.I(new_n10250_), .ZN(new_n10253_));
  NAND3_X1   g09996(.A1(new_n9840_), .A2(new_n9842_), .A3(new_n9846_), .ZN(new_n10254_));
  NAND3_X1   g09997(.A1(new_n10254_), .A2(new_n9837_), .A3(new_n10253_), .ZN(new_n10255_));
  AOI21_X1   g09998(.A1(new_n10252_), .A2(new_n10255_), .B(new_n10245_), .ZN(new_n10256_));
  AOI21_X1   g09999(.A1(new_n10242_), .A2(new_n10243_), .B(new_n10241_), .ZN(new_n10257_));
  NOR3_X1    g10000(.A1(new_n10233_), .A2(new_n10217_), .A3(new_n10229_), .ZN(new_n10258_));
  NOR2_X1    g10001(.A1(new_n10257_), .A2(new_n10258_), .ZN(new_n10259_));
  AOI21_X1   g10002(.A1(new_n10254_), .A2(new_n9837_), .B(new_n10253_), .ZN(new_n10260_));
  NOR3_X1    g10003(.A1(new_n10251_), .A2(new_n9845_), .A3(new_n10250_), .ZN(new_n10261_));
  NOR3_X1    g10004(.A1(new_n10261_), .A2(new_n10260_), .A3(new_n10259_), .ZN(new_n10262_));
  NOR2_X1    g10005(.A1(new_n10262_), .A2(new_n10256_), .ZN(new_n10263_));
  OAI22_X1   g10006(.A1(new_n1444_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n1439_), .ZN(new_n10264_));
  NAND2_X1   g10007(.A1(new_n2098_), .A2(\b[43] ), .ZN(new_n10265_));
  AOI21_X1   g10008(.A1(new_n10264_), .A2(new_n10265_), .B(new_n1447_), .ZN(new_n10266_));
  NAND2_X1   g10009(.A1(new_n4513_), .A2(new_n10266_), .ZN(new_n10267_));
  XOR2_X1    g10010(.A1(new_n10267_), .A2(\a[23] ), .Z(new_n10268_));
  INV_X1     g10011(.I(new_n10268_), .ZN(new_n10269_));
  AOI21_X1   g10012(.A1(new_n9854_), .A2(new_n9855_), .B(new_n9623_), .ZN(new_n10270_));
  INV_X1     g10013(.I(new_n10270_), .ZN(new_n10271_));
  AOI21_X1   g10014(.A1(new_n9854_), .A2(new_n9855_), .B(new_n9622_), .ZN(new_n10272_));
  NOR3_X1    g10015(.A1(new_n9843_), .A2(new_n9849_), .A3(new_n9623_), .ZN(new_n10273_));
  OAI21_X1   g10016(.A1(new_n10273_), .A2(new_n10272_), .B(new_n9626_), .ZN(new_n10274_));
  AOI21_X1   g10017(.A1(new_n10274_), .A2(new_n10271_), .B(new_n10269_), .ZN(new_n10275_));
  OAI21_X1   g10018(.A1(new_n9843_), .A2(new_n9849_), .B(new_n9623_), .ZN(new_n10276_));
  NAND3_X1   g10019(.A1(new_n9854_), .A2(new_n9855_), .A3(new_n9622_), .ZN(new_n10277_));
  AOI21_X1   g10020(.A1(new_n10276_), .A2(new_n10277_), .B(new_n9853_), .ZN(new_n10278_));
  NOR3_X1    g10021(.A1(new_n10278_), .A2(new_n10268_), .A3(new_n10270_), .ZN(new_n10279_));
  OAI21_X1   g10022(.A1(new_n10275_), .A2(new_n10279_), .B(new_n10263_), .ZN(new_n10280_));
  OAI21_X1   g10023(.A1(new_n10261_), .A2(new_n10260_), .B(new_n10259_), .ZN(new_n10281_));
  NAND3_X1   g10024(.A1(new_n10252_), .A2(new_n10255_), .A3(new_n10245_), .ZN(new_n10282_));
  NAND2_X1   g10025(.A1(new_n10281_), .A2(new_n10282_), .ZN(new_n10283_));
  OAI21_X1   g10026(.A1(new_n10278_), .A2(new_n10270_), .B(new_n10268_), .ZN(new_n10284_));
  NAND3_X1   g10027(.A1(new_n10274_), .A2(new_n10269_), .A3(new_n10271_), .ZN(new_n10285_));
  NAND3_X1   g10028(.A1(new_n10285_), .A2(new_n10284_), .A3(new_n10283_), .ZN(new_n10286_));
  NAND2_X1   g10029(.A1(new_n10280_), .A2(new_n10286_), .ZN(new_n10287_));
  OAI22_X1   g10030(.A1(new_n1168_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n1163_), .ZN(new_n10288_));
  NAND2_X1   g10031(.A1(new_n1774_), .A2(\b[46] ), .ZN(new_n10289_));
  AOI21_X1   g10032(.A1(new_n10288_), .A2(new_n10289_), .B(new_n1171_), .ZN(new_n10290_));
  NAND2_X1   g10033(.A1(new_n5177_), .A2(new_n10290_), .ZN(new_n10291_));
  XOR2_X1    g10034(.A1(new_n10291_), .A2(\a[20] ), .Z(new_n10292_));
  NAND3_X1   g10035(.A1(new_n9861_), .A2(new_n9865_), .A3(new_n9870_), .ZN(new_n10293_));
  NAND3_X1   g10036(.A1(new_n9854_), .A2(new_n9855_), .A3(new_n9623_), .ZN(new_n10294_));
  INV_X1     g10037(.I(new_n10294_), .ZN(new_n10295_));
  OAI21_X1   g10038(.A1(new_n10295_), .A2(new_n10270_), .B(new_n9626_), .ZN(new_n10296_));
  NAND3_X1   g10039(.A1(new_n10271_), .A2(new_n10294_), .A3(new_n9853_), .ZN(new_n10297_));
  AOI21_X1   g10040(.A1(new_n10297_), .A2(new_n10296_), .B(new_n9862_), .ZN(new_n10298_));
  OAI21_X1   g10041(.A1(new_n10293_), .A2(new_n10298_), .B(new_n10292_), .ZN(new_n10299_));
  INV_X1     g10042(.I(new_n10292_), .ZN(new_n10300_));
  NOR3_X1    g10043(.A1(new_n9869_), .A2(new_n9868_), .A3(new_n9866_), .ZN(new_n10301_));
  INV_X1     g10044(.I(new_n10298_), .ZN(new_n10302_));
  NAND3_X1   g10045(.A1(new_n10301_), .A2(new_n10302_), .A3(new_n10300_), .ZN(new_n10303_));
  AOI21_X1   g10046(.A1(new_n10303_), .A2(new_n10299_), .B(new_n10287_), .ZN(new_n10304_));
  AOI21_X1   g10047(.A1(new_n10285_), .A2(new_n10284_), .B(new_n10283_), .ZN(new_n10305_));
  NOR3_X1    g10048(.A1(new_n10275_), .A2(new_n10279_), .A3(new_n10263_), .ZN(new_n10306_));
  NOR2_X1    g10049(.A1(new_n10305_), .A2(new_n10306_), .ZN(new_n10307_));
  AOI21_X1   g10050(.A1(new_n10301_), .A2(new_n10302_), .B(new_n10300_), .ZN(new_n10308_));
  NOR3_X1    g10051(.A1(new_n10293_), .A2(new_n10292_), .A3(new_n10298_), .ZN(new_n10309_));
  NOR3_X1    g10052(.A1(new_n10308_), .A2(new_n10309_), .A3(new_n10307_), .ZN(new_n10310_));
  NOR2_X1    g10053(.A1(new_n10310_), .A2(new_n10304_), .ZN(new_n10311_));
  NAND2_X1   g10054(.A1(new_n9882_), .A2(new_n9883_), .ZN(new_n10312_));
  OAI22_X1   g10055(.A1(new_n940_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n935_), .ZN(new_n10313_));
  NAND2_X1   g10056(.A1(new_n1458_), .A2(\b[49] ), .ZN(new_n10314_));
  AOI21_X1   g10057(.A1(new_n10313_), .A2(new_n10314_), .B(new_n943_), .ZN(new_n10315_));
  NAND2_X1   g10058(.A1(new_n5741_), .A2(new_n10315_), .ZN(new_n10316_));
  XOR2_X1    g10059(.A1(new_n10316_), .A2(\a[17] ), .Z(new_n10317_));
  INV_X1     g10060(.I(new_n10317_), .ZN(new_n10318_));
  NOR2_X1    g10061(.A1(new_n9885_), .A2(new_n9886_), .ZN(new_n10319_));
  AOI21_X1   g10062(.A1(new_n10312_), .A2(new_n10319_), .B(new_n10318_), .ZN(new_n10320_));
  NOR2_X1    g10063(.A1(new_n9887_), .A2(new_n9888_), .ZN(new_n10321_));
  NAND2_X1   g10064(.A1(new_n9881_), .A2(new_n9878_), .ZN(new_n10322_));
  NOR3_X1    g10065(.A1(new_n10321_), .A2(new_n10322_), .A3(new_n10317_), .ZN(new_n10323_));
  OAI21_X1   g10066(.A1(new_n10320_), .A2(new_n10323_), .B(new_n10311_), .ZN(new_n10324_));
  OAI21_X1   g10067(.A1(new_n10308_), .A2(new_n10309_), .B(new_n10307_), .ZN(new_n10325_));
  NAND3_X1   g10068(.A1(new_n10303_), .A2(new_n10299_), .A3(new_n10287_), .ZN(new_n10326_));
  NAND2_X1   g10069(.A1(new_n10325_), .A2(new_n10326_), .ZN(new_n10327_));
  OAI21_X1   g10070(.A1(new_n10321_), .A2(new_n10322_), .B(new_n10317_), .ZN(new_n10328_));
  NAND3_X1   g10071(.A1(new_n10312_), .A2(new_n10319_), .A3(new_n10318_), .ZN(new_n10329_));
  NAND3_X1   g10072(.A1(new_n10328_), .A2(new_n10329_), .A3(new_n10327_), .ZN(new_n10330_));
  NAND2_X1   g10073(.A1(new_n10324_), .A2(new_n10330_), .ZN(new_n10331_));
  AOI21_X1   g10074(.A1(new_n9904_), .A2(new_n9906_), .B(new_n9917_), .ZN(new_n10332_));
  OAI22_X1   g10075(.A1(new_n757_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n752_), .ZN(new_n10333_));
  NAND2_X1   g10076(.A1(new_n1182_), .A2(\b[52] ), .ZN(new_n10334_));
  AOI21_X1   g10077(.A1(new_n10333_), .A2(new_n10334_), .B(new_n760_), .ZN(new_n10335_));
  NAND2_X1   g10078(.A1(new_n6237_), .A2(new_n10335_), .ZN(new_n10336_));
  XOR2_X1    g10079(.A1(new_n10336_), .A2(\a[14] ), .Z(new_n10337_));
  NOR2_X1    g10080(.A1(new_n10332_), .A2(new_n10337_), .ZN(new_n10338_));
  OAI21_X1   g10081(.A1(new_n9612_), .A2(new_n9918_), .B(new_n9905_), .ZN(new_n10339_));
  INV_X1     g10082(.I(new_n10337_), .ZN(new_n10340_));
  NOR2_X1    g10083(.A1(new_n10339_), .A2(new_n10340_), .ZN(new_n10341_));
  OAI21_X1   g10084(.A1(new_n10341_), .A2(new_n10338_), .B(new_n10331_), .ZN(new_n10342_));
  AOI21_X1   g10085(.A1(new_n10328_), .A2(new_n10329_), .B(new_n10327_), .ZN(new_n10343_));
  NOR3_X1    g10086(.A1(new_n10320_), .A2(new_n10323_), .A3(new_n10311_), .ZN(new_n10344_));
  NOR2_X1    g10087(.A1(new_n10344_), .A2(new_n10343_), .ZN(new_n10345_));
  NOR2_X1    g10088(.A1(new_n10339_), .A2(new_n10337_), .ZN(new_n10346_));
  NAND2_X1   g10089(.A1(new_n9906_), .A2(new_n9904_), .ZN(new_n10347_));
  AOI21_X1   g10090(.A1(new_n10347_), .A2(new_n9905_), .B(new_n10340_), .ZN(new_n10348_));
  OAI21_X1   g10091(.A1(new_n10346_), .A2(new_n10348_), .B(new_n10345_), .ZN(new_n10349_));
  NAND2_X1   g10092(.A1(new_n10342_), .A2(new_n10349_), .ZN(new_n10350_));
  OAI22_X1   g10093(.A1(new_n582_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n577_), .ZN(new_n10351_));
  NAND2_X1   g10094(.A1(new_n960_), .A2(\b[55] ), .ZN(new_n10352_));
  AOI21_X1   g10095(.A1(new_n10351_), .A2(new_n10352_), .B(new_n585_), .ZN(new_n10353_));
  NAND2_X1   g10096(.A1(new_n7308_), .A2(new_n10353_), .ZN(new_n10354_));
  XOR2_X1    g10097(.A1(new_n10354_), .A2(\a[11] ), .Z(new_n10355_));
  INV_X1     g10098(.I(new_n9557_), .ZN(new_n10356_));
  NAND3_X1   g10099(.A1(new_n9926_), .A2(new_n9925_), .A3(new_n10356_), .ZN(new_n10357_));
  NAND2_X1   g10100(.A1(new_n10357_), .A2(new_n10355_), .ZN(new_n10358_));
  INV_X1     g10101(.I(new_n10355_), .ZN(new_n10359_));
  NAND4_X1   g10102(.A1(new_n9926_), .A2(new_n9925_), .A3(new_n10356_), .A4(new_n10359_), .ZN(new_n10360_));
  AOI21_X1   g10103(.A1(new_n10358_), .A2(new_n10360_), .B(new_n10350_), .ZN(new_n10361_));
  NAND2_X1   g10104(.A1(new_n10339_), .A2(new_n10340_), .ZN(new_n10362_));
  NAND2_X1   g10105(.A1(new_n10332_), .A2(new_n10337_), .ZN(new_n10363_));
  AOI21_X1   g10106(.A1(new_n10362_), .A2(new_n10363_), .B(new_n10345_), .ZN(new_n10364_));
  NAND3_X1   g10107(.A1(new_n10347_), .A2(new_n9905_), .A3(new_n10340_), .ZN(new_n10365_));
  NAND2_X1   g10108(.A1(new_n10339_), .A2(new_n10337_), .ZN(new_n10366_));
  AOI21_X1   g10109(.A1(new_n10366_), .A2(new_n10365_), .B(new_n10331_), .ZN(new_n10367_));
  NOR2_X1    g10110(.A1(new_n10364_), .A2(new_n10367_), .ZN(new_n10368_));
  NOR3_X1    g10111(.A1(new_n9921_), .A2(new_n9913_), .A3(new_n9557_), .ZN(new_n10369_));
  NOR2_X1    g10112(.A1(new_n10369_), .A2(new_n10359_), .ZN(new_n10370_));
  NOR4_X1    g10113(.A1(new_n9921_), .A2(new_n9913_), .A3(new_n9557_), .A4(new_n10355_), .ZN(new_n10371_));
  NOR3_X1    g10114(.A1(new_n10370_), .A2(new_n10368_), .A3(new_n10371_), .ZN(new_n10372_));
  INV_X1     g10115(.I(new_n9947_), .ZN(new_n10373_));
  INV_X1     g10116(.I(new_n9948_), .ZN(new_n10374_));
  NAND3_X1   g10117(.A1(new_n9946_), .A2(new_n9945_), .A3(new_n10374_), .ZN(new_n10375_));
  OAI22_X1   g10118(.A1(new_n437_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n431_), .ZN(new_n10376_));
  NAND2_X1   g10119(.A1(new_n775_), .A2(\b[58] ), .ZN(new_n10377_));
  AOI21_X1   g10120(.A1(new_n10376_), .A2(new_n10377_), .B(new_n440_), .ZN(new_n10378_));
  NAND2_X1   g10121(.A1(new_n7929_), .A2(new_n10378_), .ZN(new_n10379_));
  XOR2_X1    g10122(.A1(new_n10379_), .A2(\a[8] ), .Z(new_n10380_));
  AOI21_X1   g10123(.A1(new_n10375_), .A2(new_n10373_), .B(new_n10380_), .ZN(new_n10381_));
  NOR3_X1    g10124(.A1(new_n9927_), .A2(new_n9924_), .A3(new_n9948_), .ZN(new_n10382_));
  INV_X1     g10125(.I(new_n10380_), .ZN(new_n10383_));
  NOR3_X1    g10126(.A1(new_n10382_), .A2(new_n9947_), .A3(new_n10383_), .ZN(new_n10384_));
  OAI22_X1   g10127(.A1(new_n10384_), .A2(new_n10381_), .B1(new_n10361_), .B2(new_n10372_), .ZN(new_n10385_));
  NOR2_X1    g10128(.A1(new_n10361_), .A2(new_n10372_), .ZN(new_n10386_));
  NAND3_X1   g10129(.A1(new_n10375_), .A2(new_n10373_), .A3(new_n10383_), .ZN(new_n10387_));
  OAI21_X1   g10130(.A1(new_n10382_), .A2(new_n9947_), .B(new_n10380_), .ZN(new_n10388_));
  NAND2_X1   g10131(.A1(new_n10388_), .A2(new_n10387_), .ZN(new_n10389_));
  NAND2_X1   g10132(.A1(new_n10389_), .A2(new_n10386_), .ZN(new_n10390_));
  NAND2_X1   g10133(.A1(new_n10390_), .A2(new_n10385_), .ZN(new_n10391_));
  XOR2_X1    g10134(.A1(new_n10024_), .A2(new_n10391_), .Z(new_n10392_));
  XOR2_X1    g10135(.A1(new_n10024_), .A2(new_n10391_), .Z(new_n10393_));
  NOR2_X1    g10136(.A1(new_n10393_), .A2(new_n10009_), .ZN(new_n10394_));
  AOI21_X1   g10137(.A1(new_n10009_), .A2(new_n10392_), .B(new_n10394_), .ZN(new_n10395_));
  XOR2_X1    g10138(.A1(new_n9990_), .A2(new_n10395_), .Z(\f[66] ));
  NAND2_X1   g10139(.A1(new_n10007_), .A2(new_n10005_), .ZN(new_n10397_));
  OAI21_X1   g10140(.A1(new_n10370_), .A2(new_n10371_), .B(new_n10368_), .ZN(new_n10398_));
  NAND3_X1   g10141(.A1(new_n10358_), .A2(new_n10350_), .A3(new_n10360_), .ZN(new_n10399_));
  OAI21_X1   g10142(.A1(new_n10382_), .A2(new_n9947_), .B(new_n10383_), .ZN(new_n10400_));
  NAND3_X1   g10143(.A1(new_n10375_), .A2(new_n10373_), .A3(new_n10380_), .ZN(new_n10401_));
  AOI22_X1   g10144(.A1(new_n10400_), .A2(new_n10401_), .B1(new_n10398_), .B2(new_n10399_), .ZN(new_n10402_));
  AOI21_X1   g10145(.A1(new_n10386_), .A2(new_n10389_), .B(new_n10402_), .ZN(new_n10403_));
  NOR2_X1    g10146(.A1(new_n10403_), .A2(new_n10001_), .ZN(new_n10404_));
  NAND2_X1   g10147(.A1(new_n10403_), .A2(new_n10001_), .ZN(new_n10405_));
  AOI21_X1   g10148(.A1(new_n10397_), .A2(new_n10405_), .B(new_n10404_), .ZN(new_n10406_));
  NAND3_X1   g10149(.A1(new_n10342_), .A2(new_n10349_), .A3(new_n10359_), .ZN(new_n10407_));
  OAI21_X1   g10150(.A1(new_n10364_), .A2(new_n10367_), .B(new_n10355_), .ZN(new_n10408_));
  AOI22_X1   g10151(.A1(new_n10408_), .A2(new_n10407_), .B1(new_n10359_), .B2(new_n10357_), .ZN(new_n10409_));
  NAND2_X1   g10152(.A1(new_n10259_), .A2(new_n10253_), .ZN(new_n10410_));
  NAND2_X1   g10153(.A1(new_n10245_), .A2(new_n10250_), .ZN(new_n10411_));
  AOI21_X1   g10154(.A1(new_n10410_), .A2(new_n10411_), .B(new_n9845_), .ZN(new_n10412_));
  AOI22_X1   g10155(.A1(new_n10412_), .A2(new_n10254_), .B1(new_n10245_), .B2(new_n10250_), .ZN(new_n10413_));
  NOR2_X1    g10156(.A1(new_n10232_), .A2(new_n10224_), .ZN(new_n10414_));
  NOR3_X1    g10157(.A1(new_n10212_), .A2(new_n10216_), .A3(new_n10222_), .ZN(new_n10415_));
  AOI21_X1   g10158(.A1(new_n10240_), .A2(new_n10237_), .B(new_n10223_), .ZN(new_n10416_));
  OAI22_X1   g10159(.A1(new_n10416_), .A2(new_n10415_), .B1(new_n10222_), .B2(new_n10414_), .ZN(new_n10417_));
  AOI21_X1   g10160(.A1(new_n10213_), .A2(new_n10211_), .B(new_n10235_), .ZN(new_n10418_));
  OAI21_X1   g10161(.A1(new_n10026_), .A2(new_n10192_), .B(new_n10191_), .ZN(new_n10419_));
  INV_X1     g10162(.I(new_n10182_), .ZN(new_n10420_));
  OAI22_X1   g10163(.A1(new_n10171_), .A2(new_n10178_), .B1(new_n10027_), .B2(new_n9766_), .ZN(new_n10421_));
  INV_X1     g10164(.I(new_n10157_), .ZN(new_n10422_));
  NOR2_X1    g10165(.A1(new_n10146_), .A2(new_n10150_), .ZN(new_n10423_));
  AOI22_X1   g10166(.A1(new_n10032_), .A2(new_n10028_), .B1(new_n10423_), .B2(new_n10155_), .ZN(new_n10424_));
  AOI21_X1   g10167(.A1(new_n10147_), .A2(new_n10145_), .B(new_n10158_), .ZN(new_n10425_));
  OAI21_X1   g10168(.A1(new_n10130_), .A2(new_n10133_), .B(new_n10131_), .ZN(new_n10426_));
  INV_X1     g10169(.I(new_n10426_), .ZN(new_n10427_));
  INV_X1     g10170(.I(new_n10108_), .ZN(new_n10428_));
  AOI21_X1   g10171(.A1(new_n10037_), .A2(new_n10111_), .B(new_n10428_), .ZN(new_n10429_));
  AOI21_X1   g10172(.A1(new_n10039_), .A2(new_n10098_), .B(new_n10096_), .ZN(new_n10430_));
  NAND2_X1   g10173(.A1(new_n10085_), .A2(new_n10087_), .ZN(new_n10431_));
  NAND2_X1   g10174(.A1(new_n10431_), .A2(new_n10086_), .ZN(new_n10432_));
  INV_X1     g10175(.I(new_n10432_), .ZN(new_n10433_));
  AOI21_X1   g10176(.A1(new_n10043_), .A2(new_n10070_), .B(new_n10068_), .ZN(new_n10434_));
  OAI22_X1   g10177(.A1(new_n450_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n403_), .ZN(new_n10435_));
  NAND2_X1   g10178(.A1(new_n9644_), .A2(\b[5] ), .ZN(new_n10436_));
  AOI21_X1   g10179(.A1(new_n10436_), .A2(new_n10435_), .B(new_n8321_), .ZN(new_n10437_));
  NAND2_X1   g10180(.A1(new_n454_), .A2(new_n10437_), .ZN(new_n10438_));
  XOR2_X1    g10181(.A1(new_n10438_), .A2(\a[62] ), .Z(new_n10439_));
  NOR3_X1    g10182(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n290_), .ZN(new_n10440_));
  NOR2_X1    g10183(.A1(new_n9364_), .A2(new_n290_), .ZN(new_n10441_));
  NOR3_X1    g10184(.A1(new_n10441_), .A2(new_n393_), .A3(new_n8985_), .ZN(new_n10442_));
  NOR2_X1    g10185(.A1(new_n10442_), .A2(new_n10440_), .ZN(new_n10443_));
  INV_X1     g10186(.I(new_n10443_), .ZN(new_n10444_));
  NOR2_X1    g10187(.A1(new_n10444_), .A2(new_n271_), .ZN(new_n10445_));
  NOR2_X1    g10188(.A1(new_n10443_), .A2(\a[2] ), .ZN(new_n10446_));
  NOR2_X1    g10189(.A1(new_n10445_), .A2(new_n10446_), .ZN(new_n10447_));
  NOR2_X1    g10190(.A1(new_n10439_), .A2(new_n10447_), .ZN(new_n10448_));
  XOR2_X1    g10191(.A1(new_n10443_), .A2(new_n271_), .Z(new_n10449_));
  INV_X1     g10192(.I(new_n10449_), .ZN(new_n10450_));
  AOI21_X1   g10193(.A1(new_n10439_), .A2(new_n10450_), .B(new_n10448_), .ZN(new_n10451_));
  INV_X1     g10194(.I(new_n10058_), .ZN(new_n10452_));
  AOI21_X1   g10195(.A1(new_n10049_), .A2(new_n10452_), .B(new_n10059_), .ZN(new_n10453_));
  OAI22_X1   g10196(.A1(new_n617_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n510_), .ZN(new_n10454_));
  NAND2_X1   g10197(.A1(new_n8628_), .A2(\b[8] ), .ZN(new_n10455_));
  AOI21_X1   g10198(.A1(new_n10455_), .A2(new_n10454_), .B(new_n7354_), .ZN(new_n10456_));
  NAND2_X1   g10199(.A1(new_n616_), .A2(new_n10456_), .ZN(new_n10457_));
  XOR2_X1    g10200(.A1(new_n10457_), .A2(\a[59] ), .Z(new_n10458_));
  NOR2_X1    g10201(.A1(new_n10458_), .A2(new_n10453_), .ZN(new_n10459_));
  INV_X1     g10202(.I(new_n10453_), .ZN(new_n10460_));
  INV_X1     g10203(.I(new_n10458_), .ZN(new_n10461_));
  NOR2_X1    g10204(.A1(new_n10461_), .A2(new_n10460_), .ZN(new_n10462_));
  NOR2_X1    g10205(.A1(new_n10462_), .A2(new_n10459_), .ZN(new_n10463_));
  XOR2_X1    g10206(.A1(new_n10458_), .A2(new_n10453_), .Z(new_n10464_));
  NAND2_X1   g10207(.A1(new_n10464_), .A2(new_n10451_), .ZN(new_n10465_));
  OAI21_X1   g10208(.A1(new_n10451_), .A2(new_n10463_), .B(new_n10465_), .ZN(new_n10466_));
  OAI22_X1   g10209(.A1(new_n6721_), .A2(new_n717_), .B1(new_n6723_), .B2(new_n795_), .ZN(new_n10467_));
  NAND2_X1   g10210(.A1(new_n7617_), .A2(\b[11] ), .ZN(new_n10468_));
  AOI21_X1   g10211(.A1(new_n10468_), .A2(new_n10467_), .B(new_n6731_), .ZN(new_n10469_));
  NAND2_X1   g10212(.A1(new_n799_), .A2(new_n10469_), .ZN(new_n10470_));
  XOR2_X1    g10213(.A1(new_n10470_), .A2(new_n6516_), .Z(new_n10471_));
  XNOR2_X1   g10214(.A1(new_n10471_), .A2(new_n10466_), .ZN(new_n10472_));
  NOR2_X1    g10215(.A1(new_n10472_), .A2(new_n10434_), .ZN(new_n10473_));
  INV_X1     g10216(.I(new_n10473_), .ZN(new_n10474_));
  INV_X1     g10217(.I(new_n10466_), .ZN(new_n10475_));
  INV_X1     g10218(.I(new_n10471_), .ZN(new_n10476_));
  NOR2_X1    g10219(.A1(new_n10476_), .A2(new_n10475_), .ZN(new_n10477_));
  NOR2_X1    g10220(.A1(new_n10471_), .A2(new_n10466_), .ZN(new_n10478_));
  OAI21_X1   g10221(.A1(new_n10477_), .A2(new_n10478_), .B(new_n10434_), .ZN(new_n10479_));
  OAI22_X1   g10222(.A1(new_n5786_), .A2(new_n992_), .B1(new_n904_), .B2(new_n5792_), .ZN(new_n10480_));
  NAND2_X1   g10223(.A1(new_n6745_), .A2(\b[14] ), .ZN(new_n10481_));
  AOI21_X1   g10224(.A1(new_n10481_), .A2(new_n10480_), .B(new_n5796_), .ZN(new_n10482_));
  NAND2_X1   g10225(.A1(new_n991_), .A2(new_n10482_), .ZN(new_n10483_));
  XOR2_X1    g10226(.A1(new_n10483_), .A2(\a[53] ), .Z(new_n10484_));
  INV_X1     g10227(.I(new_n10484_), .ZN(new_n10485_));
  NAND3_X1   g10228(.A1(new_n10474_), .A2(new_n10479_), .A3(new_n10485_), .ZN(new_n10486_));
  AOI21_X1   g10229(.A1(new_n10474_), .A2(new_n10479_), .B(new_n10485_), .ZN(new_n10487_));
  INV_X1     g10230(.I(new_n10487_), .ZN(new_n10488_));
  AOI21_X1   g10231(.A1(new_n10488_), .A2(new_n10486_), .B(new_n10433_), .ZN(new_n10489_));
  INV_X1     g10232(.I(new_n10479_), .ZN(new_n10490_));
  OAI21_X1   g10233(.A1(new_n10490_), .A2(new_n10473_), .B(new_n10485_), .ZN(new_n10491_));
  NOR3_X1    g10234(.A1(new_n10490_), .A2(new_n10473_), .A3(new_n10485_), .ZN(new_n10492_));
  INV_X1     g10235(.I(new_n10492_), .ZN(new_n10493_));
  AOI21_X1   g10236(.A1(new_n10493_), .A2(new_n10491_), .B(new_n10432_), .ZN(new_n10494_));
  OAI22_X1   g10237(.A1(new_n5228_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n5225_), .ZN(new_n10495_));
  NAND2_X1   g10238(.A1(new_n5387_), .A2(\b[17] ), .ZN(new_n10496_));
  AOI21_X1   g10239(.A1(new_n10495_), .A2(new_n10496_), .B(new_n5231_), .ZN(new_n10497_));
  AND3_X2    g10240(.A1(new_n1225_), .A2(new_n5220_), .A3(new_n10497_), .Z(new_n10498_));
  AOI21_X1   g10241(.A1(new_n1225_), .A2(new_n10497_), .B(new_n5220_), .ZN(new_n10499_));
  NOR2_X1    g10242(.A1(new_n10498_), .A2(new_n10499_), .ZN(new_n10500_));
  INV_X1     g10243(.I(new_n10500_), .ZN(new_n10501_));
  OAI21_X1   g10244(.A1(new_n10489_), .A2(new_n10494_), .B(new_n10501_), .ZN(new_n10502_));
  INV_X1     g10245(.I(new_n10486_), .ZN(new_n10503_));
  OAI21_X1   g10246(.A1(new_n10503_), .A2(new_n10487_), .B(new_n10432_), .ZN(new_n10504_));
  INV_X1     g10247(.I(new_n10491_), .ZN(new_n10505_));
  OAI21_X1   g10248(.A1(new_n10505_), .A2(new_n10492_), .B(new_n10433_), .ZN(new_n10506_));
  NAND3_X1   g10249(.A1(new_n10504_), .A2(new_n10506_), .A3(new_n10500_), .ZN(new_n10507_));
  AOI21_X1   g10250(.A1(new_n10502_), .A2(new_n10507_), .B(new_n10430_), .ZN(new_n10508_));
  INV_X1     g10251(.I(new_n10430_), .ZN(new_n10509_));
  NAND3_X1   g10252(.A1(new_n10504_), .A2(new_n10506_), .A3(new_n10501_), .ZN(new_n10510_));
  OAI21_X1   g10253(.A1(new_n10489_), .A2(new_n10494_), .B(new_n10500_), .ZN(new_n10511_));
  AOI21_X1   g10254(.A1(new_n10511_), .A2(new_n10510_), .B(new_n10509_), .ZN(new_n10512_));
  OAI22_X1   g10255(.A1(new_n4711_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n4706_), .ZN(new_n10513_));
  NAND2_X1   g10256(.A1(new_n5814_), .A2(\b[20] ), .ZN(new_n10514_));
  AOI21_X1   g10257(.A1(new_n10513_), .A2(new_n10514_), .B(new_n4714_), .ZN(new_n10515_));
  NAND2_X1   g10258(.A1(new_n1517_), .A2(new_n10515_), .ZN(new_n10516_));
  XOR2_X1    g10259(.A1(new_n10516_), .A2(\a[47] ), .Z(new_n10517_));
  INV_X1     g10260(.I(new_n10517_), .ZN(new_n10518_));
  OAI21_X1   g10261(.A1(new_n10508_), .A2(new_n10512_), .B(new_n10518_), .ZN(new_n10519_));
  AOI21_X1   g10262(.A1(new_n10504_), .A2(new_n10506_), .B(new_n10500_), .ZN(new_n10520_));
  NOR3_X1    g10263(.A1(new_n10489_), .A2(new_n10494_), .A3(new_n10501_), .ZN(new_n10521_));
  OAI21_X1   g10264(.A1(new_n10521_), .A2(new_n10520_), .B(new_n10509_), .ZN(new_n10522_));
  NOR3_X1    g10265(.A1(new_n10489_), .A2(new_n10494_), .A3(new_n10500_), .ZN(new_n10523_));
  AOI21_X1   g10266(.A1(new_n10504_), .A2(new_n10506_), .B(new_n10501_), .ZN(new_n10524_));
  OAI21_X1   g10267(.A1(new_n10523_), .A2(new_n10524_), .B(new_n10430_), .ZN(new_n10525_));
  NAND3_X1   g10268(.A1(new_n10522_), .A2(new_n10525_), .A3(new_n10517_), .ZN(new_n10526_));
  AOI21_X1   g10269(.A1(new_n10519_), .A2(new_n10526_), .B(new_n10429_), .ZN(new_n10527_));
  INV_X1     g10270(.I(new_n10429_), .ZN(new_n10528_));
  NAND3_X1   g10271(.A1(new_n10522_), .A2(new_n10525_), .A3(new_n10518_), .ZN(new_n10529_));
  OAI21_X1   g10272(.A1(new_n10508_), .A2(new_n10512_), .B(new_n10517_), .ZN(new_n10530_));
  AOI21_X1   g10273(.A1(new_n10529_), .A2(new_n10530_), .B(new_n10528_), .ZN(new_n10531_));
  OAI22_X1   g10274(.A1(new_n4208_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n4203_), .ZN(new_n10532_));
  NAND2_X1   g10275(.A1(new_n5244_), .A2(\b[23] ), .ZN(new_n10533_));
  AOI21_X1   g10276(.A1(new_n10532_), .A2(new_n10533_), .B(new_n4211_), .ZN(new_n10534_));
  NAND2_X1   g10277(.A1(new_n1828_), .A2(new_n10534_), .ZN(new_n10535_));
  XOR2_X1    g10278(.A1(new_n10535_), .A2(\a[44] ), .Z(new_n10536_));
  INV_X1     g10279(.I(new_n10536_), .ZN(new_n10537_));
  OAI21_X1   g10280(.A1(new_n10531_), .A2(new_n10527_), .B(new_n10537_), .ZN(new_n10538_));
  NOR3_X1    g10281(.A1(new_n10531_), .A2(new_n10527_), .A3(new_n10537_), .ZN(new_n10539_));
  INV_X1     g10282(.I(new_n10539_), .ZN(new_n10540_));
  AOI21_X1   g10283(.A1(new_n10540_), .A2(new_n10538_), .B(new_n10427_), .ZN(new_n10541_));
  INV_X1     g10284(.I(new_n10527_), .ZN(new_n10542_));
  NAND2_X1   g10285(.A1(new_n10530_), .A2(new_n10529_), .ZN(new_n10543_));
  NAND2_X1   g10286(.A1(new_n10543_), .A2(new_n10429_), .ZN(new_n10544_));
  NAND3_X1   g10287(.A1(new_n10542_), .A2(new_n10544_), .A3(new_n10537_), .ZN(new_n10545_));
  OAI21_X1   g10288(.A1(new_n10531_), .A2(new_n10527_), .B(new_n10536_), .ZN(new_n10546_));
  AOI21_X1   g10289(.A1(new_n10545_), .A2(new_n10546_), .B(new_n10426_), .ZN(new_n10547_));
  OAI22_X1   g10290(.A1(new_n3736_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n3731_), .ZN(new_n10548_));
  NAND2_X1   g10291(.A1(new_n4730_), .A2(\b[26] ), .ZN(new_n10549_));
  AOI21_X1   g10292(.A1(new_n10548_), .A2(new_n10549_), .B(new_n3739_), .ZN(new_n10550_));
  NAND2_X1   g10293(.A1(new_n2174_), .A2(new_n10550_), .ZN(new_n10551_));
  XOR2_X1    g10294(.A1(new_n10551_), .A2(new_n3726_), .Z(new_n10552_));
  OAI21_X1   g10295(.A1(new_n10541_), .A2(new_n10547_), .B(new_n10552_), .ZN(new_n10553_));
  INV_X1     g10296(.I(new_n10538_), .ZN(new_n10554_));
  OAI21_X1   g10297(.A1(new_n10554_), .A2(new_n10539_), .B(new_n10426_), .ZN(new_n10555_));
  INV_X1     g10298(.I(new_n10547_), .ZN(new_n10556_));
  INV_X1     g10299(.I(new_n10552_), .ZN(new_n10557_));
  NAND3_X1   g10300(.A1(new_n10556_), .A2(new_n10555_), .A3(new_n10557_), .ZN(new_n10558_));
  AOI21_X1   g10301(.A1(new_n10558_), .A2(new_n10553_), .B(new_n10425_), .ZN(new_n10559_));
  OAI21_X1   g10302(.A1(new_n10034_), .A2(new_n10159_), .B(new_n10141_), .ZN(new_n10560_));
  NAND3_X1   g10303(.A1(new_n10556_), .A2(new_n10555_), .A3(new_n10552_), .ZN(new_n10561_));
  OAI21_X1   g10304(.A1(new_n10541_), .A2(new_n10547_), .B(new_n10557_), .ZN(new_n10562_));
  AOI21_X1   g10305(.A1(new_n10561_), .A2(new_n10562_), .B(new_n10560_), .ZN(new_n10563_));
  OAI22_X1   g10306(.A1(new_n3298_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n3293_), .ZN(new_n10564_));
  NAND2_X1   g10307(.A1(new_n4227_), .A2(\b[29] ), .ZN(new_n10565_));
  AOI21_X1   g10308(.A1(new_n10564_), .A2(new_n10565_), .B(new_n3301_), .ZN(new_n10566_));
  NAND2_X1   g10309(.A1(new_n2546_), .A2(new_n10566_), .ZN(new_n10567_));
  XOR2_X1    g10310(.A1(new_n10567_), .A2(\a[38] ), .Z(new_n10568_));
  NOR3_X1    g10311(.A1(new_n10563_), .A2(new_n10559_), .A3(new_n10568_), .ZN(new_n10569_));
  AOI21_X1   g10312(.A1(new_n10556_), .A2(new_n10555_), .B(new_n10557_), .ZN(new_n10570_));
  NOR3_X1    g10313(.A1(new_n10541_), .A2(new_n10547_), .A3(new_n10552_), .ZN(new_n10571_));
  OAI21_X1   g10314(.A1(new_n10570_), .A2(new_n10571_), .B(new_n10560_), .ZN(new_n10572_));
  NOR3_X1    g10315(.A1(new_n10541_), .A2(new_n10547_), .A3(new_n10557_), .ZN(new_n10573_));
  AOI21_X1   g10316(.A1(new_n10556_), .A2(new_n10555_), .B(new_n10552_), .ZN(new_n10574_));
  OAI21_X1   g10317(.A1(new_n10574_), .A2(new_n10573_), .B(new_n10425_), .ZN(new_n10575_));
  INV_X1     g10318(.I(new_n10568_), .ZN(new_n10576_));
  AOI21_X1   g10319(.A1(new_n10572_), .A2(new_n10575_), .B(new_n10576_), .ZN(new_n10577_));
  OAI22_X1   g10320(.A1(new_n10422_), .A2(new_n10424_), .B1(new_n10577_), .B2(new_n10569_), .ZN(new_n10578_));
  NOR2_X1    g10321(.A1(new_n10424_), .A2(new_n10422_), .ZN(new_n10579_));
  OAI21_X1   g10322(.A1(new_n10563_), .A2(new_n10559_), .B(new_n10576_), .ZN(new_n10580_));
  NAND3_X1   g10323(.A1(new_n10572_), .A2(new_n10575_), .A3(new_n10568_), .ZN(new_n10581_));
  NAND2_X1   g10324(.A1(new_n10580_), .A2(new_n10581_), .ZN(new_n10582_));
  NAND2_X1   g10325(.A1(new_n10579_), .A2(new_n10582_), .ZN(new_n10583_));
  OAI22_X1   g10326(.A1(new_n2846_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n2841_), .ZN(new_n10584_));
  NAND2_X1   g10327(.A1(new_n3755_), .A2(\b[32] ), .ZN(new_n10585_));
  AOI21_X1   g10328(.A1(new_n10584_), .A2(new_n10585_), .B(new_n2849_), .ZN(new_n10586_));
  NAND2_X1   g10329(.A1(new_n2963_), .A2(new_n10586_), .ZN(new_n10587_));
  XOR2_X1    g10330(.A1(new_n10587_), .A2(\a[35] ), .Z(new_n10588_));
  INV_X1     g10331(.I(new_n10588_), .ZN(new_n10589_));
  NAND3_X1   g10332(.A1(new_n10583_), .A2(new_n10578_), .A3(new_n10589_), .ZN(new_n10590_));
  AOI21_X1   g10333(.A1(new_n10583_), .A2(new_n10578_), .B(new_n10589_), .ZN(new_n10591_));
  INV_X1     g10334(.I(new_n10591_), .ZN(new_n10592_));
  AOI22_X1   g10335(.A1(new_n10592_), .A2(new_n10590_), .B1(new_n10420_), .B2(new_n10421_), .ZN(new_n10593_));
  NAND2_X1   g10336(.A1(new_n10421_), .A2(new_n10420_), .ZN(new_n10594_));
  INV_X1     g10337(.I(new_n10578_), .ZN(new_n10595_));
  AOI21_X1   g10338(.A1(new_n10572_), .A2(new_n10575_), .B(new_n10568_), .ZN(new_n10596_));
  NOR3_X1    g10339(.A1(new_n10563_), .A2(new_n10559_), .A3(new_n10576_), .ZN(new_n10597_));
  NOR2_X1    g10340(.A1(new_n10596_), .A2(new_n10597_), .ZN(new_n10598_));
  NOR3_X1    g10341(.A1(new_n10598_), .A2(new_n10422_), .A3(new_n10424_), .ZN(new_n10599_));
  OAI21_X1   g10342(.A1(new_n10595_), .A2(new_n10599_), .B(new_n10589_), .ZN(new_n10600_));
  NAND3_X1   g10343(.A1(new_n10583_), .A2(new_n10578_), .A3(new_n10588_), .ZN(new_n10601_));
  AOI21_X1   g10344(.A1(new_n10600_), .A2(new_n10601_), .B(new_n10594_), .ZN(new_n10602_));
  OAI22_X1   g10345(.A1(new_n2452_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n2447_), .ZN(new_n10603_));
  NAND2_X1   g10346(.A1(new_n3312_), .A2(\b[35] ), .ZN(new_n10604_));
  AOI21_X1   g10347(.A1(new_n10603_), .A2(new_n10604_), .B(new_n2455_), .ZN(new_n10605_));
  NAND2_X1   g10348(.A1(new_n3411_), .A2(new_n10605_), .ZN(new_n10606_));
  XOR2_X1    g10349(.A1(new_n10606_), .A2(\a[32] ), .Z(new_n10607_));
  NOR3_X1    g10350(.A1(new_n10602_), .A2(new_n10593_), .A3(new_n10607_), .ZN(new_n10608_));
  INV_X1     g10351(.I(new_n10590_), .ZN(new_n10609_));
  OAI21_X1   g10352(.A1(new_n10609_), .A2(new_n10591_), .B(new_n10594_), .ZN(new_n10610_));
  NAND2_X1   g10353(.A1(new_n10600_), .A2(new_n10601_), .ZN(new_n10611_));
  NAND3_X1   g10354(.A1(new_n10611_), .A2(new_n10420_), .A3(new_n10421_), .ZN(new_n10612_));
  INV_X1     g10355(.I(new_n10607_), .ZN(new_n10613_));
  AOI21_X1   g10356(.A1(new_n10612_), .A2(new_n10610_), .B(new_n10613_), .ZN(new_n10614_));
  OAI21_X1   g10357(.A1(new_n10614_), .A2(new_n10608_), .B(new_n10419_), .ZN(new_n10615_));
  OAI21_X1   g10358(.A1(new_n10602_), .A2(new_n10593_), .B(new_n10613_), .ZN(new_n10616_));
  NAND3_X1   g10359(.A1(new_n10612_), .A2(new_n10610_), .A3(new_n10607_), .ZN(new_n10617_));
  AOI21_X1   g10360(.A1(new_n10617_), .A2(new_n10616_), .B(new_n10419_), .ZN(new_n10618_));
  INV_X1     g10361(.I(new_n10618_), .ZN(new_n10619_));
  OAI22_X1   g10362(.A1(new_n2084_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n2079_), .ZN(new_n10620_));
  NAND2_X1   g10363(.A1(new_n2864_), .A2(\b[38] ), .ZN(new_n10621_));
  AOI21_X1   g10364(.A1(new_n10620_), .A2(new_n10621_), .B(new_n2087_), .ZN(new_n10622_));
  NAND2_X1   g10365(.A1(new_n3844_), .A2(new_n10622_), .ZN(new_n10623_));
  XOR2_X1    g10366(.A1(new_n10623_), .A2(\a[29] ), .Z(new_n10624_));
  INV_X1     g10367(.I(new_n10624_), .ZN(new_n10625_));
  NAND3_X1   g10368(.A1(new_n10619_), .A2(new_n10615_), .A3(new_n10625_), .ZN(new_n10626_));
  INV_X1     g10369(.I(new_n10615_), .ZN(new_n10627_));
  OAI21_X1   g10370(.A1(new_n10627_), .A2(new_n10618_), .B(new_n10624_), .ZN(new_n10628_));
  AOI21_X1   g10371(.A1(new_n10628_), .A2(new_n10626_), .B(new_n10418_), .ZN(new_n10629_));
  OAI21_X1   g10372(.A1(new_n10025_), .A2(new_n10236_), .B(new_n10206_), .ZN(new_n10630_));
  OAI21_X1   g10373(.A1(new_n10627_), .A2(new_n10618_), .B(new_n10625_), .ZN(new_n10631_));
  NAND3_X1   g10374(.A1(new_n10619_), .A2(new_n10615_), .A3(new_n10624_), .ZN(new_n10632_));
  AOI21_X1   g10375(.A1(new_n10631_), .A2(new_n10632_), .B(new_n10630_), .ZN(new_n10633_));
  OAI22_X1   g10376(.A1(new_n1760_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n1755_), .ZN(new_n10634_));
  NAND2_X1   g10377(.A1(new_n2470_), .A2(\b[41] ), .ZN(new_n10635_));
  AOI21_X1   g10378(.A1(new_n10634_), .A2(new_n10635_), .B(new_n1763_), .ZN(new_n10636_));
  NAND2_X1   g10379(.A1(new_n4320_), .A2(new_n10636_), .ZN(new_n10637_));
  XOR2_X1    g10380(.A1(new_n10637_), .A2(\a[26] ), .Z(new_n10638_));
  INV_X1     g10381(.I(new_n10638_), .ZN(new_n10639_));
  OAI21_X1   g10382(.A1(new_n10633_), .A2(new_n10629_), .B(new_n10639_), .ZN(new_n10640_));
  NOR3_X1    g10383(.A1(new_n10633_), .A2(new_n10629_), .A3(new_n10639_), .ZN(new_n10641_));
  INV_X1     g10384(.I(new_n10641_), .ZN(new_n10642_));
  AOI21_X1   g10385(.A1(new_n10642_), .A2(new_n10640_), .B(new_n10417_), .ZN(new_n10643_));
  INV_X1     g10386(.I(new_n10417_), .ZN(new_n10644_));
  NOR3_X1    g10387(.A1(new_n10627_), .A2(new_n10618_), .A3(new_n10624_), .ZN(new_n10645_));
  AOI21_X1   g10388(.A1(new_n10619_), .A2(new_n10615_), .B(new_n10625_), .ZN(new_n10646_));
  OAI21_X1   g10389(.A1(new_n10645_), .A2(new_n10646_), .B(new_n10630_), .ZN(new_n10647_));
  INV_X1     g10390(.I(new_n10633_), .ZN(new_n10648_));
  NAND3_X1   g10391(.A1(new_n10648_), .A2(new_n10647_), .A3(new_n10639_), .ZN(new_n10649_));
  OAI21_X1   g10392(.A1(new_n10633_), .A2(new_n10629_), .B(new_n10638_), .ZN(new_n10650_));
  AOI21_X1   g10393(.A1(new_n10649_), .A2(new_n10650_), .B(new_n10644_), .ZN(new_n10651_));
  OAI22_X1   g10394(.A1(new_n1444_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n1439_), .ZN(new_n10652_));
  NAND2_X1   g10395(.A1(new_n2098_), .A2(\b[44] ), .ZN(new_n10653_));
  AOI21_X1   g10396(.A1(new_n10652_), .A2(new_n10653_), .B(new_n1447_), .ZN(new_n10654_));
  NAND2_X1   g10397(.A1(new_n4833_), .A2(new_n10654_), .ZN(new_n10655_));
  XOR2_X1    g10398(.A1(new_n10655_), .A2(\a[23] ), .Z(new_n10656_));
  INV_X1     g10399(.I(new_n10656_), .ZN(new_n10657_));
  OAI21_X1   g10400(.A1(new_n10651_), .A2(new_n10643_), .B(new_n10657_), .ZN(new_n10658_));
  INV_X1     g10401(.I(new_n10643_), .ZN(new_n10659_));
  INV_X1     g10402(.I(new_n10651_), .ZN(new_n10660_));
  NAND3_X1   g10403(.A1(new_n10660_), .A2(new_n10659_), .A3(new_n10656_), .ZN(new_n10661_));
  AOI21_X1   g10404(.A1(new_n10658_), .A2(new_n10661_), .B(new_n10413_), .ZN(new_n10662_));
  NAND2_X1   g10405(.A1(new_n10245_), .A2(new_n10250_), .ZN(new_n10663_));
  NOR2_X1    g10406(.A1(new_n10245_), .A2(new_n10250_), .ZN(new_n10664_));
  NOR2_X1    g10407(.A1(new_n10259_), .A2(new_n10253_), .ZN(new_n10665_));
  OAI21_X1   g10408(.A1(new_n10665_), .A2(new_n10664_), .B(new_n9837_), .ZN(new_n10666_));
  OAI21_X1   g10409(.A1(new_n10666_), .A2(new_n10251_), .B(new_n10663_), .ZN(new_n10667_));
  NOR3_X1    g10410(.A1(new_n10651_), .A2(new_n10643_), .A3(new_n10656_), .ZN(new_n10668_));
  AOI21_X1   g10411(.A1(new_n10660_), .A2(new_n10659_), .B(new_n10657_), .ZN(new_n10669_));
  NOR2_X1    g10412(.A1(new_n10669_), .A2(new_n10668_), .ZN(new_n10670_));
  NOR2_X1    g10413(.A1(new_n10670_), .A2(new_n10667_), .ZN(new_n10671_));
  OAI22_X1   g10414(.A1(new_n1168_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n1163_), .ZN(new_n10672_));
  NAND2_X1   g10415(.A1(new_n1774_), .A2(\b[47] ), .ZN(new_n10673_));
  AOI21_X1   g10416(.A1(new_n10672_), .A2(new_n10673_), .B(new_n1171_), .ZN(new_n10674_));
  NAND2_X1   g10417(.A1(new_n5196_), .A2(new_n10674_), .ZN(new_n10675_));
  XOR2_X1    g10418(.A1(new_n10675_), .A2(\a[20] ), .Z(new_n10676_));
  NOR3_X1    g10419(.A1(new_n10671_), .A2(new_n10662_), .A3(new_n10676_), .ZN(new_n10677_));
  NAND2_X1   g10420(.A1(new_n10661_), .A2(new_n10658_), .ZN(new_n10678_));
  NAND2_X1   g10421(.A1(new_n10678_), .A2(new_n10667_), .ZN(new_n10679_));
  OAI21_X1   g10422(.A1(new_n10668_), .A2(new_n10669_), .B(new_n10413_), .ZN(new_n10680_));
  INV_X1     g10423(.I(new_n10676_), .ZN(new_n10681_));
  AOI21_X1   g10424(.A1(new_n10679_), .A2(new_n10680_), .B(new_n10681_), .ZN(new_n10682_));
  NOR2_X1    g10425(.A1(new_n10677_), .A2(new_n10682_), .ZN(new_n10683_));
  INV_X1     g10426(.I(new_n10683_), .ZN(new_n10684_));
  NOR2_X1    g10427(.A1(new_n10293_), .A2(new_n10298_), .ZN(new_n10685_));
  NAND3_X1   g10428(.A1(new_n10280_), .A2(new_n10286_), .A3(new_n10300_), .ZN(new_n10686_));
  INV_X1     g10429(.I(new_n10686_), .ZN(new_n10687_));
  NOR2_X1    g10430(.A1(new_n10307_), .A2(new_n10300_), .ZN(new_n10688_));
  OAI22_X1   g10431(.A1(new_n10688_), .A2(new_n10687_), .B1(new_n10292_), .B2(new_n10685_), .ZN(new_n10689_));
  OAI22_X1   g10432(.A1(new_n940_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n935_), .ZN(new_n10690_));
  NAND2_X1   g10433(.A1(new_n1458_), .A2(\b[50] ), .ZN(new_n10691_));
  AOI21_X1   g10434(.A1(new_n10690_), .A2(new_n10691_), .B(new_n943_), .ZN(new_n10692_));
  NAND2_X1   g10435(.A1(new_n5954_), .A2(new_n10692_), .ZN(new_n10693_));
  XOR2_X1    g10436(.A1(new_n10693_), .A2(\a[17] ), .Z(new_n10694_));
  NOR2_X1    g10437(.A1(new_n10689_), .A2(new_n10694_), .ZN(new_n10695_));
  NAND2_X1   g10438(.A1(new_n10301_), .A2(new_n10302_), .ZN(new_n10696_));
  NAND2_X1   g10439(.A1(new_n10287_), .A2(new_n10292_), .ZN(new_n10697_));
  AOI22_X1   g10440(.A1(new_n10697_), .A2(new_n10686_), .B1(new_n10300_), .B2(new_n10696_), .ZN(new_n10698_));
  INV_X1     g10441(.I(new_n10694_), .ZN(new_n10699_));
  NOR2_X1    g10442(.A1(new_n10698_), .A2(new_n10699_), .ZN(new_n10700_));
  OAI21_X1   g10443(.A1(new_n10695_), .A2(new_n10700_), .B(new_n10684_), .ZN(new_n10701_));
  NOR2_X1    g10444(.A1(new_n10698_), .A2(new_n10694_), .ZN(new_n10702_));
  NOR2_X1    g10445(.A1(new_n10689_), .A2(new_n10699_), .ZN(new_n10703_));
  OAI21_X1   g10446(.A1(new_n10703_), .A2(new_n10702_), .B(new_n10683_), .ZN(new_n10704_));
  OAI22_X1   g10447(.A1(new_n757_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n752_), .ZN(new_n10705_));
  NAND2_X1   g10448(.A1(new_n1182_), .A2(\b[53] ), .ZN(new_n10706_));
  AOI21_X1   g10449(.A1(new_n10705_), .A2(new_n10706_), .B(new_n760_), .ZN(new_n10707_));
  NAND2_X1   g10450(.A1(new_n6471_), .A2(new_n10707_), .ZN(new_n10708_));
  XOR2_X1    g10451(.A1(new_n10708_), .A2(\a[14] ), .Z(new_n10709_));
  INV_X1     g10452(.I(new_n10709_), .ZN(new_n10710_));
  NAND3_X1   g10453(.A1(new_n10701_), .A2(new_n10704_), .A3(new_n10710_), .ZN(new_n10711_));
  NAND2_X1   g10454(.A1(new_n10698_), .A2(new_n10699_), .ZN(new_n10712_));
  NAND2_X1   g10455(.A1(new_n10689_), .A2(new_n10694_), .ZN(new_n10713_));
  AOI21_X1   g10456(.A1(new_n10713_), .A2(new_n10712_), .B(new_n10683_), .ZN(new_n10714_));
  NAND2_X1   g10457(.A1(new_n10689_), .A2(new_n10699_), .ZN(new_n10715_));
  NAND2_X1   g10458(.A1(new_n10698_), .A2(new_n10694_), .ZN(new_n10716_));
  AOI21_X1   g10459(.A1(new_n10715_), .A2(new_n10716_), .B(new_n10684_), .ZN(new_n10717_));
  OAI21_X1   g10460(.A1(new_n10717_), .A2(new_n10714_), .B(new_n10709_), .ZN(new_n10718_));
  NAND2_X1   g10461(.A1(new_n10718_), .A2(new_n10711_), .ZN(new_n10719_));
  OAI22_X1   g10462(.A1(new_n10339_), .A2(new_n10340_), .B1(new_n10343_), .B2(new_n10344_), .ZN(new_n10720_));
  OAI22_X1   g10463(.A1(new_n582_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n577_), .ZN(new_n10721_));
  NAND2_X1   g10464(.A1(new_n960_), .A2(\b[56] ), .ZN(new_n10722_));
  AOI21_X1   g10465(.A1(new_n10721_), .A2(new_n10722_), .B(new_n585_), .ZN(new_n10723_));
  NAND2_X1   g10466(.A1(new_n7559_), .A2(new_n10723_), .ZN(new_n10724_));
  XOR2_X1    g10467(.A1(new_n10724_), .A2(\a[11] ), .Z(new_n10725_));
  AOI21_X1   g10468(.A1(new_n10720_), .A2(new_n10362_), .B(new_n10725_), .ZN(new_n10726_));
  AOI22_X1   g10469(.A1(new_n10332_), .A2(new_n10337_), .B1(new_n10324_), .B2(new_n10330_), .ZN(new_n10727_));
  INV_X1     g10470(.I(new_n10725_), .ZN(new_n10728_));
  NOR3_X1    g10471(.A1(new_n10727_), .A2(new_n10338_), .A3(new_n10728_), .ZN(new_n10729_));
  OAI21_X1   g10472(.A1(new_n10726_), .A2(new_n10729_), .B(new_n10719_), .ZN(new_n10730_));
  NOR3_X1    g10473(.A1(new_n10717_), .A2(new_n10714_), .A3(new_n10709_), .ZN(new_n10731_));
  AOI21_X1   g10474(.A1(new_n10701_), .A2(new_n10704_), .B(new_n10710_), .ZN(new_n10732_));
  NOR2_X1    g10475(.A1(new_n10732_), .A2(new_n10731_), .ZN(new_n10733_));
  NOR3_X1    g10476(.A1(new_n10727_), .A2(new_n10338_), .A3(new_n10725_), .ZN(new_n10734_));
  AOI21_X1   g10477(.A1(new_n10720_), .A2(new_n10362_), .B(new_n10728_), .ZN(new_n10735_));
  OAI21_X1   g10478(.A1(new_n10735_), .A2(new_n10734_), .B(new_n10733_), .ZN(new_n10736_));
  OAI22_X1   g10479(.A1(new_n437_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n431_), .ZN(new_n10737_));
  NAND2_X1   g10480(.A1(new_n775_), .A2(\b[59] ), .ZN(new_n10738_));
  AOI21_X1   g10481(.A1(new_n10737_), .A2(new_n10738_), .B(new_n440_), .ZN(new_n10739_));
  NAND2_X1   g10482(.A1(new_n8550_), .A2(new_n10739_), .ZN(new_n10740_));
  XOR2_X1    g10483(.A1(new_n10740_), .A2(\a[8] ), .Z(new_n10741_));
  AOI21_X1   g10484(.A1(new_n10730_), .A2(new_n10736_), .B(new_n10741_), .ZN(new_n10742_));
  OAI21_X1   g10485(.A1(new_n10727_), .A2(new_n10338_), .B(new_n10728_), .ZN(new_n10743_));
  NAND3_X1   g10486(.A1(new_n10720_), .A2(new_n10362_), .A3(new_n10725_), .ZN(new_n10744_));
  AOI21_X1   g10487(.A1(new_n10743_), .A2(new_n10744_), .B(new_n10733_), .ZN(new_n10745_));
  NAND3_X1   g10488(.A1(new_n10720_), .A2(new_n10362_), .A3(new_n10728_), .ZN(new_n10746_));
  OAI21_X1   g10489(.A1(new_n10727_), .A2(new_n10338_), .B(new_n10725_), .ZN(new_n10747_));
  AOI21_X1   g10490(.A1(new_n10747_), .A2(new_n10746_), .B(new_n10719_), .ZN(new_n10748_));
  INV_X1     g10491(.I(new_n10741_), .ZN(new_n10749_));
  NOR3_X1    g10492(.A1(new_n10745_), .A2(new_n10748_), .A3(new_n10749_), .ZN(new_n10750_));
  OAI21_X1   g10493(.A1(new_n10742_), .A2(new_n10750_), .B(new_n10409_), .ZN(new_n10751_));
  NOR3_X1    g10494(.A1(new_n10364_), .A2(new_n10367_), .A3(new_n10355_), .ZN(new_n10752_));
  AOI21_X1   g10495(.A1(new_n10342_), .A2(new_n10349_), .B(new_n10359_), .ZN(new_n10753_));
  OAI22_X1   g10496(.A1(new_n10753_), .A2(new_n10752_), .B1(new_n10355_), .B2(new_n10369_), .ZN(new_n10754_));
  NOR3_X1    g10497(.A1(new_n10745_), .A2(new_n10748_), .A3(new_n10741_), .ZN(new_n10755_));
  AOI21_X1   g10498(.A1(new_n10730_), .A2(new_n10736_), .B(new_n10749_), .ZN(new_n10756_));
  OAI21_X1   g10499(.A1(new_n10756_), .A2(new_n10755_), .B(new_n10754_), .ZN(new_n10757_));
  NAND2_X1   g10500(.A1(new_n10751_), .A2(new_n10757_), .ZN(new_n10758_));
  OAI21_X1   g10501(.A1(new_n10361_), .A2(new_n10372_), .B(new_n10401_), .ZN(new_n10759_));
  OAI21_X1   g10502(.A1(new_n8956_), .A2(new_n320_), .B(new_n311_), .ZN(new_n10760_));
  AOI21_X1   g10503(.A1(new_n594_), .A2(\b[62] ), .B(new_n10760_), .ZN(new_n10761_));
  NAND3_X1   g10504(.A1(new_n9322_), .A2(new_n308_), .A3(new_n10761_), .ZN(new_n10762_));
  INV_X1     g10505(.I(new_n10762_), .ZN(new_n10763_));
  AOI21_X1   g10506(.A1(new_n9322_), .A2(new_n10761_), .B(new_n308_), .ZN(new_n10764_));
  NOR2_X1    g10507(.A1(new_n10763_), .A2(new_n10764_), .ZN(new_n10765_));
  INV_X1     g10508(.I(new_n10765_), .ZN(new_n10766_));
  NAND3_X1   g10509(.A1(new_n10759_), .A2(new_n10766_), .A3(new_n10400_), .ZN(new_n10767_));
  INV_X1     g10510(.I(new_n10767_), .ZN(new_n10768_));
  AOI21_X1   g10511(.A1(new_n10759_), .A2(new_n10400_), .B(new_n10766_), .ZN(new_n10769_));
  OAI21_X1   g10512(.A1(new_n10768_), .A2(new_n10769_), .B(new_n10758_), .ZN(new_n10770_));
  OAI21_X1   g10513(.A1(new_n10745_), .A2(new_n10748_), .B(new_n10749_), .ZN(new_n10771_));
  NAND3_X1   g10514(.A1(new_n10730_), .A2(new_n10736_), .A3(new_n10741_), .ZN(new_n10772_));
  AOI21_X1   g10515(.A1(new_n10771_), .A2(new_n10772_), .B(new_n10754_), .ZN(new_n10773_));
  NAND3_X1   g10516(.A1(new_n10730_), .A2(new_n10736_), .A3(new_n10749_), .ZN(new_n10774_));
  OAI21_X1   g10517(.A1(new_n10745_), .A2(new_n10748_), .B(new_n10741_), .ZN(new_n10775_));
  AOI21_X1   g10518(.A1(new_n10775_), .A2(new_n10774_), .B(new_n10409_), .ZN(new_n10776_));
  NOR2_X1    g10519(.A1(new_n10773_), .A2(new_n10776_), .ZN(new_n10777_));
  AOI21_X1   g10520(.A1(new_n10759_), .A2(new_n10400_), .B(new_n10765_), .ZN(new_n10778_));
  OAI21_X1   g10521(.A1(new_n10386_), .A2(new_n10384_), .B(new_n10400_), .ZN(new_n10779_));
  NOR2_X1    g10522(.A1(new_n10779_), .A2(new_n10766_), .ZN(new_n10780_));
  OAI21_X1   g10523(.A1(new_n10780_), .A2(new_n10778_), .B(new_n10777_), .ZN(new_n10781_));
  NAND2_X1   g10524(.A1(new_n10770_), .A2(new_n10781_), .ZN(new_n10782_));
  AOI21_X1   g10525(.A1(new_n10007_), .A2(new_n10005_), .B(new_n10001_), .ZN(new_n10783_));
  NOR3_X1    g10526(.A1(new_n9994_), .A2(new_n9993_), .A3(new_n10002_), .ZN(new_n10784_));
  NOR3_X1    g10527(.A1(new_n10784_), .A2(new_n10403_), .A3(new_n10783_), .ZN(new_n10785_));
  AOI21_X1   g10528(.A1(new_n10003_), .A2(new_n10008_), .B(new_n10391_), .ZN(new_n10786_));
  NOR2_X1    g10529(.A1(new_n10786_), .A2(new_n10785_), .ZN(new_n10787_));
  NOR3_X1    g10530(.A1(new_n10024_), .A2(new_n10787_), .A3(new_n10782_), .ZN(new_n10788_));
  NOR2_X1    g10531(.A1(new_n10021_), .A2(new_n10020_), .ZN(new_n10789_));
  AOI21_X1   g10532(.A1(new_n10014_), .A2(new_n10010_), .B(new_n9982_), .ZN(new_n10790_));
  NOR3_X1    g10533(.A1(new_n10021_), .A2(new_n10020_), .A3(new_n10019_), .ZN(new_n10791_));
  OAI22_X1   g10534(.A1(new_n10791_), .A2(new_n10790_), .B1(new_n10789_), .B2(new_n9597_), .ZN(new_n10792_));
  NOR2_X1    g10535(.A1(new_n10382_), .A2(new_n9947_), .ZN(new_n10793_));
  AOI22_X1   g10536(.A1(new_n10793_), .A2(new_n10380_), .B1(new_n10398_), .B2(new_n10399_), .ZN(new_n10794_));
  OAI21_X1   g10537(.A1(new_n10794_), .A2(new_n10381_), .B(new_n10765_), .ZN(new_n10795_));
  AOI22_X1   g10538(.A1(new_n10795_), .A2(new_n10767_), .B1(new_n10751_), .B2(new_n10757_), .ZN(new_n10796_));
  NAND2_X1   g10539(.A1(new_n10779_), .A2(new_n10766_), .ZN(new_n10797_));
  NAND3_X1   g10540(.A1(new_n10759_), .A2(new_n10765_), .A3(new_n10400_), .ZN(new_n10798_));
  AOI21_X1   g10541(.A1(new_n10797_), .A2(new_n10798_), .B(new_n10758_), .ZN(new_n10799_));
  NOR2_X1    g10542(.A1(new_n10799_), .A2(new_n10796_), .ZN(new_n10800_));
  NAND3_X1   g10543(.A1(new_n10391_), .A2(new_n10003_), .A3(new_n10008_), .ZN(new_n10801_));
  OAI21_X1   g10544(.A1(new_n10783_), .A2(new_n10784_), .B(new_n10403_), .ZN(new_n10802_));
  NAND2_X1   g10545(.A1(new_n10802_), .A2(new_n10801_), .ZN(new_n10803_));
  AOI21_X1   g10546(.A1(new_n10792_), .A2(new_n10803_), .B(new_n10800_), .ZN(new_n10804_));
  OAI21_X1   g10547(.A1(new_n10788_), .A2(new_n10804_), .B(new_n10406_), .ZN(new_n10805_));
  INV_X1     g10548(.I(new_n10406_), .ZN(new_n10806_));
  NAND3_X1   g10549(.A1(new_n10792_), .A2(new_n10803_), .A3(new_n10800_), .ZN(new_n10807_));
  OAI21_X1   g10550(.A1(new_n10024_), .A2(new_n10787_), .B(new_n10782_), .ZN(new_n10808_));
  NAND3_X1   g10551(.A1(new_n10808_), .A2(new_n10807_), .A3(new_n10806_), .ZN(new_n10809_));
  NAND2_X1   g10552(.A1(new_n10805_), .A2(new_n10809_), .ZN(\f[67] ));
  NOR2_X1    g10553(.A1(new_n10024_), .A2(new_n10787_), .ZN(new_n10811_));
  AOI22_X1   g10554(.A1(new_n10808_), .A2(new_n10807_), .B1(new_n10811_), .B2(new_n10806_), .ZN(new_n10812_));
  AOI21_X1   g10555(.A1(new_n10758_), .A2(new_n10798_), .B(new_n10778_), .ZN(new_n10813_));
  INV_X1     g10556(.I(new_n9595_), .ZN(new_n10814_));
  AOI22_X1   g10557(.A1(new_n10814_), .A2(new_n311_), .B1(\b[63] ), .B2(new_n594_), .ZN(new_n10815_));
  AOI21_X1   g10558(.A1(new_n10409_), .A2(new_n10772_), .B(new_n10742_), .ZN(new_n10816_));
  AOI21_X1   g10559(.A1(new_n10701_), .A2(new_n10704_), .B(new_n10709_), .ZN(new_n10817_));
  NAND2_X1   g10560(.A1(new_n10713_), .A2(new_n10684_), .ZN(new_n10818_));
  NAND2_X1   g10561(.A1(new_n10818_), .A2(new_n10712_), .ZN(new_n10819_));
  AOI21_X1   g10562(.A1(new_n10679_), .A2(new_n10680_), .B(new_n10676_), .ZN(new_n10820_));
  INV_X1     g10563(.I(new_n10820_), .ZN(new_n10821_));
  NAND2_X1   g10564(.A1(new_n10667_), .A2(new_n10661_), .ZN(new_n10822_));
  AOI21_X1   g10565(.A1(new_n10648_), .A2(new_n10647_), .B(new_n10638_), .ZN(new_n10823_));
  AOI21_X1   g10566(.A1(new_n10642_), .A2(new_n10644_), .B(new_n10823_), .ZN(new_n10824_));
  AOI21_X1   g10567(.A1(new_n10630_), .A2(new_n10628_), .B(new_n10645_), .ZN(new_n10825_));
  INV_X1     g10568(.I(new_n10616_), .ZN(new_n10826_));
  AOI21_X1   g10569(.A1(new_n10419_), .A2(new_n10617_), .B(new_n10826_), .ZN(new_n10827_));
  AOI21_X1   g10570(.A1(new_n10594_), .A2(new_n10592_), .B(new_n10609_), .ZN(new_n10828_));
  OAI21_X1   g10571(.A1(new_n10579_), .A2(new_n10597_), .B(new_n10580_), .ZN(new_n10829_));
  INV_X1     g10572(.I(new_n10829_), .ZN(new_n10830_));
  AOI21_X1   g10573(.A1(new_n10560_), .A2(new_n10558_), .B(new_n10570_), .ZN(new_n10831_));
  AOI21_X1   g10574(.A1(new_n10426_), .A2(new_n10540_), .B(new_n10554_), .ZN(new_n10832_));
  INV_X1     g10575(.I(new_n10832_), .ZN(new_n10833_));
  OAI22_X1   g10576(.A1(new_n4208_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n4203_), .ZN(new_n10834_));
  OAI21_X1   g10577(.A1(new_n1709_), .A2(new_n4362_), .B(new_n10834_), .ZN(new_n10835_));
  AOI21_X1   g10578(.A1(new_n1926_), .A2(new_n4210_), .B(new_n10835_), .ZN(new_n10836_));
  INV_X1     g10579(.I(new_n10836_), .ZN(new_n10837_));
  AOI21_X1   g10580(.A1(new_n10522_), .A2(new_n10525_), .B(new_n10517_), .ZN(new_n10838_));
  AOI21_X1   g10581(.A1(new_n10528_), .A2(new_n10526_), .B(new_n10838_), .ZN(new_n10839_));
  AOI21_X1   g10582(.A1(new_n10509_), .A2(new_n10507_), .B(new_n10520_), .ZN(new_n10840_));
  AOI21_X1   g10583(.A1(new_n10432_), .A2(new_n10488_), .B(new_n10503_), .ZN(new_n10841_));
  INV_X1     g10584(.I(new_n10434_), .ZN(new_n10842_));
  INV_X1     g10585(.I(new_n10478_), .ZN(new_n10843_));
  AOI21_X1   g10586(.A1(new_n10842_), .A2(new_n10843_), .B(new_n10477_), .ZN(new_n10844_));
  INV_X1     g10587(.I(new_n10844_), .ZN(new_n10845_));
  OAI22_X1   g10588(.A1(new_n6721_), .A2(new_n795_), .B1(new_n6723_), .B2(new_n848_), .ZN(new_n10846_));
  NAND2_X1   g10589(.A1(new_n7617_), .A2(\b[12] ), .ZN(new_n10847_));
  AOI21_X1   g10590(.A1(new_n10847_), .A2(new_n10846_), .B(new_n6731_), .ZN(new_n10848_));
  NAND2_X1   g10591(.A1(new_n847_), .A2(new_n10848_), .ZN(new_n10849_));
  XOR2_X1    g10592(.A1(new_n10849_), .A2(\a[56] ), .Z(new_n10850_));
  INV_X1     g10593(.I(new_n10850_), .ZN(new_n10851_));
  OAI22_X1   g10594(.A1(new_n495_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n450_), .ZN(new_n10852_));
  NAND2_X1   g10595(.A1(new_n9644_), .A2(\b[6] ), .ZN(new_n10853_));
  AOI21_X1   g10596(.A1(new_n10853_), .A2(new_n10852_), .B(new_n8321_), .ZN(new_n10854_));
  NAND2_X1   g10597(.A1(new_n494_), .A2(new_n10854_), .ZN(new_n10855_));
  XOR2_X1    g10598(.A1(new_n10855_), .A2(new_n8309_), .Z(new_n10856_));
  NOR3_X1    g10599(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n393_), .ZN(new_n10857_));
  NOR2_X1    g10600(.A1(new_n9364_), .A2(new_n393_), .ZN(new_n10858_));
  NOR3_X1    g10601(.A1(new_n10858_), .A2(new_n347_), .A3(new_n8985_), .ZN(new_n10859_));
  NOR2_X1    g10602(.A1(new_n10859_), .A2(new_n10857_), .ZN(new_n10860_));
  INV_X1     g10603(.I(new_n10860_), .ZN(new_n10861_));
  NOR2_X1    g10604(.A1(new_n10861_), .A2(new_n271_), .ZN(new_n10862_));
  NOR2_X1    g10605(.A1(new_n10860_), .A2(\a[2] ), .ZN(new_n10863_));
  NOR2_X1    g10606(.A1(new_n10862_), .A2(new_n10863_), .ZN(new_n10864_));
  INV_X1     g10607(.I(new_n10864_), .ZN(new_n10865_));
  XOR2_X1    g10608(.A1(new_n10860_), .A2(new_n271_), .Z(new_n10866_));
  NOR2_X1    g10609(.A1(new_n10856_), .A2(new_n10866_), .ZN(new_n10867_));
  AOI21_X1   g10610(.A1(new_n10856_), .A2(new_n10865_), .B(new_n10867_), .ZN(new_n10868_));
  INV_X1     g10611(.I(new_n10868_), .ZN(new_n10869_));
  INV_X1     g10612(.I(new_n10446_), .ZN(new_n10870_));
  OAI21_X1   g10613(.A1(new_n10439_), .A2(new_n10445_), .B(new_n10870_), .ZN(new_n10871_));
  INV_X1     g10614(.I(new_n10871_), .ZN(new_n10872_));
  OAI22_X1   g10615(.A1(new_n659_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n617_), .ZN(new_n10873_));
  NAND2_X1   g10616(.A1(new_n8628_), .A2(\b[9] ), .ZN(new_n10874_));
  AOI21_X1   g10617(.A1(new_n10874_), .A2(new_n10873_), .B(new_n7354_), .ZN(new_n10875_));
  NAND2_X1   g10618(.A1(new_n663_), .A2(new_n10875_), .ZN(new_n10876_));
  XOR2_X1    g10619(.A1(new_n10876_), .A2(\a[59] ), .Z(new_n10877_));
  XOR2_X1    g10620(.A1(new_n10877_), .A2(new_n10872_), .Z(new_n10878_));
  NAND2_X1   g10621(.A1(new_n10878_), .A2(new_n10869_), .ZN(new_n10879_));
  NOR2_X1    g10622(.A1(new_n10877_), .A2(new_n10872_), .ZN(new_n10880_));
  XOR2_X1    g10623(.A1(new_n10876_), .A2(new_n7343_), .Z(new_n10881_));
  NOR2_X1    g10624(.A1(new_n10881_), .A2(new_n10871_), .ZN(new_n10882_));
  OAI21_X1   g10625(.A1(new_n10880_), .A2(new_n10882_), .B(new_n10868_), .ZN(new_n10883_));
  INV_X1     g10626(.I(new_n10459_), .ZN(new_n10884_));
  OAI21_X1   g10627(.A1(new_n10451_), .A2(new_n10462_), .B(new_n10884_), .ZN(new_n10885_));
  NAND3_X1   g10628(.A1(new_n10879_), .A2(new_n10883_), .A3(new_n10885_), .ZN(new_n10886_));
  INV_X1     g10629(.I(new_n10886_), .ZN(new_n10887_));
  AOI21_X1   g10630(.A1(new_n10879_), .A2(new_n10883_), .B(new_n10885_), .ZN(new_n10888_));
  OAI21_X1   g10631(.A1(new_n10887_), .A2(new_n10888_), .B(new_n10851_), .ZN(new_n10889_));
  INV_X1     g10632(.I(new_n10885_), .ZN(new_n10890_));
  AOI21_X1   g10633(.A1(new_n10879_), .A2(new_n10883_), .B(new_n10890_), .ZN(new_n10891_));
  NAND3_X1   g10634(.A1(new_n10879_), .A2(new_n10883_), .A3(new_n10890_), .ZN(new_n10892_));
  INV_X1     g10635(.I(new_n10892_), .ZN(new_n10893_));
  OAI21_X1   g10636(.A1(new_n10893_), .A2(new_n10891_), .B(new_n10850_), .ZN(new_n10894_));
  OAI22_X1   g10637(.A1(new_n5786_), .A2(new_n1044_), .B1(new_n992_), .B2(new_n5792_), .ZN(new_n10895_));
  NAND2_X1   g10638(.A1(new_n6745_), .A2(\b[15] ), .ZN(new_n10896_));
  AOI21_X1   g10639(.A1(new_n10896_), .A2(new_n10895_), .B(new_n5796_), .ZN(new_n10897_));
  AND3_X2    g10640(.A1(new_n1047_), .A2(new_n5783_), .A3(new_n10897_), .Z(new_n10898_));
  AOI21_X1   g10641(.A1(new_n1047_), .A2(new_n10897_), .B(new_n5783_), .ZN(new_n10899_));
  NOR2_X1    g10642(.A1(new_n10898_), .A2(new_n10899_), .ZN(new_n10900_));
  AOI21_X1   g10643(.A1(new_n10889_), .A2(new_n10894_), .B(new_n10900_), .ZN(new_n10901_));
  INV_X1     g10644(.I(new_n10888_), .ZN(new_n10902_));
  AOI21_X1   g10645(.A1(new_n10902_), .A2(new_n10886_), .B(new_n10850_), .ZN(new_n10903_));
  XOR2_X1    g10646(.A1(new_n10881_), .A2(new_n10872_), .Z(new_n10904_));
  NOR2_X1    g10647(.A1(new_n10904_), .A2(new_n10868_), .ZN(new_n10905_));
  INV_X1     g10648(.I(new_n10883_), .ZN(new_n10906_));
  OAI21_X1   g10649(.A1(new_n10905_), .A2(new_n10906_), .B(new_n10885_), .ZN(new_n10907_));
  AOI21_X1   g10650(.A1(new_n10907_), .A2(new_n10892_), .B(new_n10851_), .ZN(new_n10908_));
  INV_X1     g10651(.I(new_n10900_), .ZN(new_n10909_));
  NOR3_X1    g10652(.A1(new_n10903_), .A2(new_n10908_), .A3(new_n10909_), .ZN(new_n10910_));
  OAI21_X1   g10653(.A1(new_n10901_), .A2(new_n10910_), .B(new_n10845_), .ZN(new_n10911_));
  NOR3_X1    g10654(.A1(new_n10903_), .A2(new_n10908_), .A3(new_n10900_), .ZN(new_n10912_));
  AOI21_X1   g10655(.A1(new_n10889_), .A2(new_n10894_), .B(new_n10909_), .ZN(new_n10913_));
  OAI21_X1   g10656(.A1(new_n10913_), .A2(new_n10912_), .B(new_n10844_), .ZN(new_n10914_));
  OAI22_X1   g10657(.A1(new_n5228_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n5225_), .ZN(new_n10915_));
  NAND2_X1   g10658(.A1(new_n5387_), .A2(\b[18] ), .ZN(new_n10916_));
  AOI21_X1   g10659(.A1(new_n10915_), .A2(new_n10916_), .B(new_n5231_), .ZN(new_n10917_));
  NAND2_X1   g10660(.A1(new_n1304_), .A2(new_n10917_), .ZN(new_n10918_));
  XOR2_X1    g10661(.A1(new_n10918_), .A2(\a[50] ), .Z(new_n10919_));
  INV_X1     g10662(.I(new_n10919_), .ZN(new_n10920_));
  NAND3_X1   g10663(.A1(new_n10911_), .A2(new_n10914_), .A3(new_n10920_), .ZN(new_n10921_));
  OAI21_X1   g10664(.A1(new_n10903_), .A2(new_n10908_), .B(new_n10909_), .ZN(new_n10922_));
  NAND3_X1   g10665(.A1(new_n10889_), .A2(new_n10894_), .A3(new_n10900_), .ZN(new_n10923_));
  AOI21_X1   g10666(.A1(new_n10923_), .A2(new_n10922_), .B(new_n10844_), .ZN(new_n10924_));
  NAND3_X1   g10667(.A1(new_n10889_), .A2(new_n10894_), .A3(new_n10909_), .ZN(new_n10925_));
  OAI21_X1   g10668(.A1(new_n10903_), .A2(new_n10908_), .B(new_n10900_), .ZN(new_n10926_));
  AOI21_X1   g10669(.A1(new_n10925_), .A2(new_n10926_), .B(new_n10845_), .ZN(new_n10927_));
  OAI21_X1   g10670(.A1(new_n10927_), .A2(new_n10924_), .B(new_n10919_), .ZN(new_n10928_));
  AOI21_X1   g10671(.A1(new_n10928_), .A2(new_n10921_), .B(new_n10841_), .ZN(new_n10929_));
  INV_X1     g10672(.I(new_n10841_), .ZN(new_n10930_));
  OAI21_X1   g10673(.A1(new_n10927_), .A2(new_n10924_), .B(new_n10920_), .ZN(new_n10931_));
  NAND3_X1   g10674(.A1(new_n10911_), .A2(new_n10914_), .A3(new_n10919_), .ZN(new_n10932_));
  AOI21_X1   g10675(.A1(new_n10931_), .A2(new_n10932_), .B(new_n10930_), .ZN(new_n10933_));
  OAI22_X1   g10676(.A1(new_n4711_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n4706_), .ZN(new_n10934_));
  NAND2_X1   g10677(.A1(new_n5814_), .A2(\b[21] ), .ZN(new_n10935_));
  AOI21_X1   g10678(.A1(new_n10934_), .A2(new_n10935_), .B(new_n4714_), .ZN(new_n10936_));
  NAND2_X1   g10679(.A1(new_n1604_), .A2(new_n10936_), .ZN(new_n10937_));
  XOR2_X1    g10680(.A1(new_n10937_), .A2(\a[47] ), .Z(new_n10938_));
  NOR3_X1    g10681(.A1(new_n10933_), .A2(new_n10929_), .A3(new_n10938_), .ZN(new_n10939_));
  INV_X1     g10682(.I(new_n10939_), .ZN(new_n10940_));
  OAI21_X1   g10683(.A1(new_n10933_), .A2(new_n10929_), .B(new_n10938_), .ZN(new_n10941_));
  AOI21_X1   g10684(.A1(new_n10940_), .A2(new_n10941_), .B(new_n10840_), .ZN(new_n10942_));
  INV_X1     g10685(.I(new_n10840_), .ZN(new_n10943_));
  XOR2_X1    g10686(.A1(new_n10937_), .A2(new_n4701_), .Z(new_n10944_));
  OAI21_X1   g10687(.A1(new_n10933_), .A2(new_n10929_), .B(new_n10944_), .ZN(new_n10945_));
  NAND2_X1   g10688(.A1(new_n10928_), .A2(new_n10921_), .ZN(new_n10946_));
  NAND2_X1   g10689(.A1(new_n10946_), .A2(new_n10930_), .ZN(new_n10947_));
  AOI21_X1   g10690(.A1(new_n10911_), .A2(new_n10914_), .B(new_n10919_), .ZN(new_n10948_));
  NOR3_X1    g10691(.A1(new_n10927_), .A2(new_n10924_), .A3(new_n10920_), .ZN(new_n10949_));
  OAI21_X1   g10692(.A1(new_n10948_), .A2(new_n10949_), .B(new_n10841_), .ZN(new_n10950_));
  NAND3_X1   g10693(.A1(new_n10947_), .A2(new_n10950_), .A3(new_n10938_), .ZN(new_n10951_));
  AOI21_X1   g10694(.A1(new_n10951_), .A2(new_n10945_), .B(new_n10943_), .ZN(new_n10952_));
  OAI21_X1   g10695(.A1(new_n10942_), .A2(new_n10952_), .B(new_n10839_), .ZN(new_n10953_));
  NOR3_X1    g10696(.A1(new_n10508_), .A2(new_n10512_), .A3(new_n10518_), .ZN(new_n10954_));
  OAI21_X1   g10697(.A1(new_n10429_), .A2(new_n10954_), .B(new_n10519_), .ZN(new_n10955_));
  AOI21_X1   g10698(.A1(new_n10947_), .A2(new_n10950_), .B(new_n10944_), .ZN(new_n10956_));
  OAI21_X1   g10699(.A1(new_n10956_), .A2(new_n10939_), .B(new_n10943_), .ZN(new_n10957_));
  AOI21_X1   g10700(.A1(new_n10947_), .A2(new_n10950_), .B(new_n10938_), .ZN(new_n10958_));
  NOR3_X1    g10701(.A1(new_n10933_), .A2(new_n10929_), .A3(new_n10944_), .ZN(new_n10959_));
  OAI21_X1   g10702(.A1(new_n10958_), .A2(new_n10959_), .B(new_n10840_), .ZN(new_n10960_));
  NAND3_X1   g10703(.A1(new_n10960_), .A2(new_n10957_), .A3(new_n10955_), .ZN(new_n10961_));
  AOI21_X1   g10704(.A1(new_n10953_), .A2(new_n10961_), .B(\a[44] ), .ZN(new_n10962_));
  AOI21_X1   g10705(.A1(new_n10960_), .A2(new_n10957_), .B(new_n10955_), .ZN(new_n10963_));
  NOR3_X1    g10706(.A1(new_n10942_), .A2(new_n10839_), .A3(new_n10952_), .ZN(new_n10964_));
  NOR3_X1    g10707(.A1(new_n10964_), .A2(new_n10963_), .A3(new_n4198_), .ZN(new_n10965_));
  OAI21_X1   g10708(.A1(new_n10965_), .A2(new_n10962_), .B(new_n10837_), .ZN(new_n10966_));
  OAI21_X1   g10709(.A1(new_n10964_), .A2(new_n10963_), .B(new_n4198_), .ZN(new_n10967_));
  NAND3_X1   g10710(.A1(new_n10953_), .A2(new_n10961_), .A3(\a[44] ), .ZN(new_n10968_));
  NAND3_X1   g10711(.A1(new_n10967_), .A2(new_n10968_), .A3(new_n10836_), .ZN(new_n10969_));
  OAI22_X1   g10712(.A1(new_n3736_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n3731_), .ZN(new_n10970_));
  NAND2_X1   g10713(.A1(new_n4730_), .A2(\b[27] ), .ZN(new_n10971_));
  AOI21_X1   g10714(.A1(new_n10970_), .A2(new_n10971_), .B(new_n3739_), .ZN(new_n10972_));
  AND3_X2    g10715(.A1(new_n2276_), .A2(new_n3726_), .A3(new_n10972_), .Z(new_n10973_));
  AOI21_X1   g10716(.A1(new_n2276_), .A2(new_n10972_), .B(new_n3726_), .ZN(new_n10974_));
  NOR2_X1    g10717(.A1(new_n10973_), .A2(new_n10974_), .ZN(new_n10975_));
  AOI21_X1   g10718(.A1(new_n10966_), .A2(new_n10969_), .B(new_n10975_), .ZN(new_n10976_));
  AOI21_X1   g10719(.A1(new_n10967_), .A2(new_n10968_), .B(new_n10836_), .ZN(new_n10977_));
  NOR3_X1    g10720(.A1(new_n10965_), .A2(new_n10962_), .A3(new_n10837_), .ZN(new_n10978_));
  INV_X1     g10721(.I(new_n10975_), .ZN(new_n10979_));
  NOR3_X1    g10722(.A1(new_n10978_), .A2(new_n10977_), .A3(new_n10979_), .ZN(new_n10980_));
  OAI21_X1   g10723(.A1(new_n10980_), .A2(new_n10976_), .B(new_n10833_), .ZN(new_n10981_));
  NOR3_X1    g10724(.A1(new_n10978_), .A2(new_n10977_), .A3(new_n10975_), .ZN(new_n10982_));
  AOI21_X1   g10725(.A1(new_n10966_), .A2(new_n10969_), .B(new_n10979_), .ZN(new_n10983_));
  OAI21_X1   g10726(.A1(new_n10982_), .A2(new_n10983_), .B(new_n10832_), .ZN(new_n10984_));
  OAI22_X1   g10727(.A1(new_n3298_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n3293_), .ZN(new_n10985_));
  NAND2_X1   g10728(.A1(new_n4227_), .A2(\b[30] ), .ZN(new_n10986_));
  AOI21_X1   g10729(.A1(new_n10985_), .A2(new_n10986_), .B(new_n3301_), .ZN(new_n10987_));
  NAND2_X1   g10730(.A1(new_n2659_), .A2(new_n10987_), .ZN(new_n10988_));
  XOR2_X1    g10731(.A1(new_n10988_), .A2(\a[38] ), .Z(new_n10989_));
  INV_X1     g10732(.I(new_n10989_), .ZN(new_n10990_));
  NAND3_X1   g10733(.A1(new_n10981_), .A2(new_n10984_), .A3(new_n10990_), .ZN(new_n10991_));
  OAI21_X1   g10734(.A1(new_n10978_), .A2(new_n10977_), .B(new_n10979_), .ZN(new_n10992_));
  NAND3_X1   g10735(.A1(new_n10966_), .A2(new_n10969_), .A3(new_n10975_), .ZN(new_n10993_));
  AOI21_X1   g10736(.A1(new_n10992_), .A2(new_n10993_), .B(new_n10832_), .ZN(new_n10994_));
  NAND3_X1   g10737(.A1(new_n10966_), .A2(new_n10969_), .A3(new_n10979_), .ZN(new_n10995_));
  OAI21_X1   g10738(.A1(new_n10978_), .A2(new_n10977_), .B(new_n10975_), .ZN(new_n10996_));
  AOI21_X1   g10739(.A1(new_n10996_), .A2(new_n10995_), .B(new_n10833_), .ZN(new_n10997_));
  OAI21_X1   g10740(.A1(new_n10994_), .A2(new_n10997_), .B(new_n10989_), .ZN(new_n10998_));
  AOI21_X1   g10741(.A1(new_n10998_), .A2(new_n10991_), .B(new_n10831_), .ZN(new_n10999_));
  INV_X1     g10742(.I(new_n10831_), .ZN(new_n11000_));
  OAI21_X1   g10743(.A1(new_n10994_), .A2(new_n10997_), .B(new_n10990_), .ZN(new_n11001_));
  NAND3_X1   g10744(.A1(new_n10981_), .A2(new_n10984_), .A3(new_n10989_), .ZN(new_n11002_));
  AOI21_X1   g10745(.A1(new_n11001_), .A2(new_n11002_), .B(new_n11000_), .ZN(new_n11003_));
  OAI22_X1   g10746(.A1(new_n2846_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n2841_), .ZN(new_n11004_));
  NAND2_X1   g10747(.A1(new_n3755_), .A2(\b[33] ), .ZN(new_n11005_));
  AOI21_X1   g10748(.A1(new_n11004_), .A2(new_n11005_), .B(new_n2849_), .ZN(new_n11006_));
  AND3_X2    g10749(.A1(new_n3101_), .A2(new_n2836_), .A3(new_n11006_), .Z(new_n11007_));
  AOI21_X1   g10750(.A1(new_n3101_), .A2(new_n11006_), .B(new_n2836_), .ZN(new_n11008_));
  NOR2_X1    g10751(.A1(new_n11007_), .A2(new_n11008_), .ZN(new_n11009_));
  NOR3_X1    g10752(.A1(new_n10999_), .A2(new_n11003_), .A3(new_n11009_), .ZN(new_n11010_));
  INV_X1     g10753(.I(new_n11010_), .ZN(new_n11011_));
  OAI21_X1   g10754(.A1(new_n10999_), .A2(new_n11003_), .B(new_n11009_), .ZN(new_n11012_));
  AOI21_X1   g10755(.A1(new_n11011_), .A2(new_n11012_), .B(new_n10830_), .ZN(new_n11013_));
  OAI22_X1   g10756(.A1(new_n10999_), .A2(new_n11003_), .B1(new_n11007_), .B2(new_n11008_), .ZN(new_n11014_));
  NOR3_X1    g10757(.A1(new_n10994_), .A2(new_n10997_), .A3(new_n10989_), .ZN(new_n11015_));
  AOI21_X1   g10758(.A1(new_n10981_), .A2(new_n10984_), .B(new_n10990_), .ZN(new_n11016_));
  OAI21_X1   g10759(.A1(new_n11016_), .A2(new_n11015_), .B(new_n11000_), .ZN(new_n11017_));
  AOI21_X1   g10760(.A1(new_n10981_), .A2(new_n10984_), .B(new_n10989_), .ZN(new_n11018_));
  NOR3_X1    g10761(.A1(new_n10994_), .A2(new_n10997_), .A3(new_n10990_), .ZN(new_n11019_));
  OAI21_X1   g10762(.A1(new_n11018_), .A2(new_n11019_), .B(new_n10831_), .ZN(new_n11020_));
  NAND3_X1   g10763(.A1(new_n11017_), .A2(new_n11020_), .A3(new_n11009_), .ZN(new_n11021_));
  AOI21_X1   g10764(.A1(new_n11014_), .A2(new_n11021_), .B(new_n10829_), .ZN(new_n11022_));
  AOI22_X1   g10765(.A1(\b[38] ), .A2(new_n2451_), .B1(new_n3116_), .B2(\b[37] ), .ZN(new_n11023_));
  NOR2_X1    g10766(.A1(new_n2602_), .A2(new_n3247_), .ZN(new_n11024_));
  OAI21_X1   g10767(.A1(new_n11023_), .A2(new_n11024_), .B(new_n2454_), .ZN(new_n11025_));
  NOR3_X1    g10768(.A1(new_n3564_), .A2(\a[32] ), .A3(new_n11025_), .ZN(new_n11026_));
  OAI21_X1   g10769(.A1(new_n3564_), .A2(new_n11025_), .B(\a[32] ), .ZN(new_n11027_));
  INV_X1     g10770(.I(new_n11027_), .ZN(new_n11028_));
  NOR2_X1    g10771(.A1(new_n11028_), .A2(new_n11026_), .ZN(new_n11029_));
  INV_X1     g10772(.I(new_n11029_), .ZN(new_n11030_));
  OAI21_X1   g10773(.A1(new_n11013_), .A2(new_n11022_), .B(new_n11030_), .ZN(new_n11031_));
  INV_X1     g10774(.I(new_n11012_), .ZN(new_n11032_));
  OAI21_X1   g10775(.A1(new_n11032_), .A2(new_n11010_), .B(new_n10829_), .ZN(new_n11033_));
  INV_X1     g10776(.I(new_n11022_), .ZN(new_n11034_));
  NAND3_X1   g10777(.A1(new_n11034_), .A2(new_n11033_), .A3(new_n11029_), .ZN(new_n11035_));
  AOI21_X1   g10778(.A1(new_n11035_), .A2(new_n11031_), .B(new_n10828_), .ZN(new_n11036_));
  INV_X1     g10779(.I(new_n10828_), .ZN(new_n11037_));
  NOR3_X1    g10780(.A1(new_n11013_), .A2(new_n11022_), .A3(new_n11029_), .ZN(new_n11038_));
  INV_X1     g10781(.I(new_n11038_), .ZN(new_n11039_));
  OAI21_X1   g10782(.A1(new_n11013_), .A2(new_n11022_), .B(new_n11029_), .ZN(new_n11040_));
  AOI21_X1   g10783(.A1(new_n11039_), .A2(new_n11040_), .B(new_n11037_), .ZN(new_n11041_));
  OAI22_X1   g10784(.A1(new_n2084_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n2079_), .ZN(new_n11042_));
  NAND2_X1   g10785(.A1(new_n2864_), .A2(\b[39] ), .ZN(new_n11043_));
  AOI21_X1   g10786(.A1(new_n11042_), .A2(new_n11043_), .B(new_n2087_), .ZN(new_n11044_));
  NAND2_X1   g10787(.A1(new_n3996_), .A2(new_n11044_), .ZN(new_n11045_));
  XOR2_X1    g10788(.A1(new_n11045_), .A2(\a[29] ), .Z(new_n11046_));
  INV_X1     g10789(.I(new_n11046_), .ZN(new_n11047_));
  OAI21_X1   g10790(.A1(new_n11041_), .A2(new_n11036_), .B(new_n11047_), .ZN(new_n11048_));
  AOI21_X1   g10791(.A1(new_n11034_), .A2(new_n11033_), .B(new_n11029_), .ZN(new_n11049_));
  NOR3_X1    g10792(.A1(new_n11013_), .A2(new_n11022_), .A3(new_n11030_), .ZN(new_n11050_));
  OAI21_X1   g10793(.A1(new_n11049_), .A2(new_n11050_), .B(new_n11037_), .ZN(new_n11051_));
  AOI21_X1   g10794(.A1(new_n11034_), .A2(new_n11033_), .B(new_n11030_), .ZN(new_n11052_));
  OAI21_X1   g10795(.A1(new_n11052_), .A2(new_n11038_), .B(new_n10828_), .ZN(new_n11053_));
  NAND3_X1   g10796(.A1(new_n11051_), .A2(new_n11053_), .A3(new_n11046_), .ZN(new_n11054_));
  AOI21_X1   g10797(.A1(new_n11048_), .A2(new_n11054_), .B(new_n10827_), .ZN(new_n11055_));
  NAND2_X1   g10798(.A1(new_n10617_), .A2(new_n10419_), .ZN(new_n11056_));
  NAND2_X1   g10799(.A1(new_n11056_), .A2(new_n10616_), .ZN(new_n11057_));
  NAND3_X1   g10800(.A1(new_n11051_), .A2(new_n11053_), .A3(new_n11047_), .ZN(new_n11058_));
  OAI21_X1   g10801(.A1(new_n11041_), .A2(new_n11036_), .B(new_n11046_), .ZN(new_n11059_));
  AOI21_X1   g10802(.A1(new_n11059_), .A2(new_n11058_), .B(new_n11057_), .ZN(new_n11060_));
  AOI22_X1   g10803(.A1(\b[44] ), .A2(new_n1759_), .B1(new_n2289_), .B2(\b[43] ), .ZN(new_n11061_));
  NOR2_X1    g10804(.A1(new_n1857_), .A2(new_n4018_), .ZN(new_n11062_));
  OAI21_X1   g10805(.A1(new_n11061_), .A2(new_n11062_), .B(new_n1762_), .ZN(new_n11063_));
  NOR3_X1    g10806(.A1(new_n4499_), .A2(\a[26] ), .A3(new_n11063_), .ZN(new_n11064_));
  NOR2_X1    g10807(.A1(new_n4499_), .A2(new_n11063_), .ZN(new_n11065_));
  NOR2_X1    g10808(.A1(new_n11065_), .A2(new_n1750_), .ZN(new_n11066_));
  NOR2_X1    g10809(.A1(new_n11066_), .A2(new_n11064_), .ZN(new_n11067_));
  INV_X1     g10810(.I(new_n11067_), .ZN(new_n11068_));
  OAI21_X1   g10811(.A1(new_n11060_), .A2(new_n11055_), .B(new_n11068_), .ZN(new_n11069_));
  AOI21_X1   g10812(.A1(new_n11051_), .A2(new_n11053_), .B(new_n11046_), .ZN(new_n11070_));
  INV_X1     g10813(.I(new_n11054_), .ZN(new_n11071_));
  OAI21_X1   g10814(.A1(new_n11071_), .A2(new_n11070_), .B(new_n11057_), .ZN(new_n11072_));
  NOR3_X1    g10815(.A1(new_n11041_), .A2(new_n11046_), .A3(new_n11036_), .ZN(new_n11073_));
  AOI21_X1   g10816(.A1(new_n11051_), .A2(new_n11053_), .B(new_n11047_), .ZN(new_n11074_));
  OAI21_X1   g10817(.A1(new_n11073_), .A2(new_n11074_), .B(new_n10827_), .ZN(new_n11075_));
  NAND3_X1   g10818(.A1(new_n11072_), .A2(new_n11075_), .A3(new_n11067_), .ZN(new_n11076_));
  AOI21_X1   g10819(.A1(new_n11076_), .A2(new_n11069_), .B(new_n10825_), .ZN(new_n11077_));
  OAI21_X1   g10820(.A1(new_n10418_), .A2(new_n10646_), .B(new_n10626_), .ZN(new_n11078_));
  NAND3_X1   g10821(.A1(new_n11072_), .A2(new_n11075_), .A3(new_n11068_), .ZN(new_n11079_));
  OAI21_X1   g10822(.A1(new_n11060_), .A2(new_n11055_), .B(new_n11067_), .ZN(new_n11080_));
  AOI21_X1   g10823(.A1(new_n11079_), .A2(new_n11080_), .B(new_n11078_), .ZN(new_n11081_));
  OAI22_X1   g10824(.A1(new_n1444_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n1439_), .ZN(new_n11082_));
  NAND2_X1   g10825(.A1(new_n2098_), .A2(\b[45] ), .ZN(new_n11083_));
  AOI21_X1   g10826(.A1(new_n11082_), .A2(new_n11083_), .B(new_n1447_), .ZN(new_n11084_));
  NAND2_X1   g10827(.A1(new_n5004_), .A2(new_n11084_), .ZN(new_n11085_));
  XOR2_X1    g10828(.A1(new_n11085_), .A2(\a[23] ), .Z(new_n11086_));
  INV_X1     g10829(.I(new_n11086_), .ZN(new_n11087_));
  OAI21_X1   g10830(.A1(new_n11077_), .A2(new_n11081_), .B(new_n11087_), .ZN(new_n11088_));
  AOI21_X1   g10831(.A1(new_n11072_), .A2(new_n11075_), .B(new_n11067_), .ZN(new_n11089_));
  NOR3_X1    g10832(.A1(new_n11060_), .A2(new_n11055_), .A3(new_n11068_), .ZN(new_n11090_));
  OAI21_X1   g10833(.A1(new_n11089_), .A2(new_n11090_), .B(new_n11078_), .ZN(new_n11091_));
  NOR3_X1    g10834(.A1(new_n11060_), .A2(new_n11055_), .A3(new_n11067_), .ZN(new_n11092_));
  AOI21_X1   g10835(.A1(new_n11072_), .A2(new_n11075_), .B(new_n11068_), .ZN(new_n11093_));
  OAI21_X1   g10836(.A1(new_n11093_), .A2(new_n11092_), .B(new_n10825_), .ZN(new_n11094_));
  NAND3_X1   g10837(.A1(new_n11094_), .A2(new_n11091_), .A3(new_n11086_), .ZN(new_n11095_));
  AOI21_X1   g10838(.A1(new_n11088_), .A2(new_n11095_), .B(new_n10824_), .ZN(new_n11096_));
  OAI21_X1   g10839(.A1(new_n10417_), .A2(new_n10641_), .B(new_n10640_), .ZN(new_n11097_));
  NAND3_X1   g10840(.A1(new_n11094_), .A2(new_n11091_), .A3(new_n11087_), .ZN(new_n11098_));
  OAI21_X1   g10841(.A1(new_n11077_), .A2(new_n11081_), .B(new_n11086_), .ZN(new_n11099_));
  AOI21_X1   g10842(.A1(new_n11099_), .A2(new_n11098_), .B(new_n11097_), .ZN(new_n11100_));
  OAI22_X1   g10843(.A1(new_n1168_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n1163_), .ZN(new_n11101_));
  NAND2_X1   g10844(.A1(new_n1774_), .A2(\b[48] ), .ZN(new_n11102_));
  AOI21_X1   g10845(.A1(new_n11101_), .A2(new_n11102_), .B(new_n1171_), .ZN(new_n11103_));
  NAND2_X1   g10846(.A1(new_n5537_), .A2(new_n11103_), .ZN(new_n11104_));
  XOR2_X1    g10847(.A1(new_n11104_), .A2(\a[20] ), .Z(new_n11105_));
  INV_X1     g10848(.I(new_n11105_), .ZN(new_n11106_));
  OAI21_X1   g10849(.A1(new_n11096_), .A2(new_n11100_), .B(new_n11106_), .ZN(new_n11107_));
  INV_X1     g10850(.I(new_n11088_), .ZN(new_n11108_));
  NOR3_X1    g10851(.A1(new_n11077_), .A2(new_n11081_), .A3(new_n11087_), .ZN(new_n11109_));
  OAI21_X1   g10852(.A1(new_n11108_), .A2(new_n11109_), .B(new_n11097_), .ZN(new_n11110_));
  INV_X1     g10853(.I(new_n11100_), .ZN(new_n11111_));
  NAND3_X1   g10854(.A1(new_n11111_), .A2(new_n11110_), .A3(new_n11105_), .ZN(new_n11112_));
  AOI22_X1   g10855(.A1(new_n10822_), .A2(new_n10658_), .B1(new_n11112_), .B2(new_n11107_), .ZN(new_n11113_));
  NAND2_X1   g10856(.A1(new_n10822_), .A2(new_n10658_), .ZN(new_n11114_));
  NOR3_X1    g10857(.A1(new_n11096_), .A2(new_n11105_), .A3(new_n11100_), .ZN(new_n11115_));
  AOI21_X1   g10858(.A1(new_n11111_), .A2(new_n11110_), .B(new_n11106_), .ZN(new_n11116_));
  NOR2_X1    g10859(.A1(new_n11116_), .A2(new_n11115_), .ZN(new_n11117_));
  NOR2_X1    g10860(.A1(new_n11114_), .A2(new_n11117_), .ZN(new_n11118_));
  OAI22_X1   g10861(.A1(new_n940_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n935_), .ZN(new_n11119_));
  NAND2_X1   g10862(.A1(new_n1458_), .A2(\b[51] ), .ZN(new_n11120_));
  AOI21_X1   g10863(.A1(new_n11119_), .A2(new_n11120_), .B(new_n943_), .ZN(new_n11121_));
  NAND2_X1   g10864(.A1(new_n6219_), .A2(new_n11121_), .ZN(new_n11122_));
  XOR2_X1    g10865(.A1(new_n11122_), .A2(\a[17] ), .Z(new_n11123_));
  INV_X1     g10866(.I(new_n11123_), .ZN(new_n11124_));
  OAI21_X1   g10867(.A1(new_n11118_), .A2(new_n11113_), .B(new_n11124_), .ZN(new_n11125_));
  NAND2_X1   g10868(.A1(new_n11112_), .A2(new_n11107_), .ZN(new_n11126_));
  NAND2_X1   g10869(.A1(new_n11114_), .A2(new_n11126_), .ZN(new_n11127_));
  NAND3_X1   g10870(.A1(new_n11111_), .A2(new_n11110_), .A3(new_n11106_), .ZN(new_n11128_));
  OAI21_X1   g10871(.A1(new_n11096_), .A2(new_n11100_), .B(new_n11105_), .ZN(new_n11129_));
  NAND2_X1   g10872(.A1(new_n11128_), .A2(new_n11129_), .ZN(new_n11130_));
  NAND3_X1   g10873(.A1(new_n11130_), .A2(new_n10822_), .A3(new_n10658_), .ZN(new_n11131_));
  NAND3_X1   g10874(.A1(new_n11127_), .A2(new_n11131_), .A3(new_n11123_), .ZN(new_n11132_));
  AOI21_X1   g10875(.A1(new_n11125_), .A2(new_n11132_), .B(new_n10821_), .ZN(new_n11133_));
  NAND3_X1   g10876(.A1(new_n11127_), .A2(new_n11131_), .A3(new_n11124_), .ZN(new_n11134_));
  OAI21_X1   g10877(.A1(new_n11118_), .A2(new_n11113_), .B(new_n11123_), .ZN(new_n11135_));
  AOI21_X1   g10878(.A1(new_n11135_), .A2(new_n11134_), .B(new_n10820_), .ZN(new_n11136_));
  OAI22_X1   g10879(.A1(new_n757_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n752_), .ZN(new_n11137_));
  NAND2_X1   g10880(.A1(new_n1182_), .A2(\b[54] ), .ZN(new_n11138_));
  AOI21_X1   g10881(.A1(new_n11137_), .A2(new_n11138_), .B(new_n760_), .ZN(new_n11139_));
  NAND2_X1   g10882(.A1(new_n6994_), .A2(new_n11139_), .ZN(new_n11140_));
  XOR2_X1    g10883(.A1(new_n11140_), .A2(\a[14] ), .Z(new_n11141_));
  INV_X1     g10884(.I(new_n11141_), .ZN(new_n11142_));
  OAI21_X1   g10885(.A1(new_n11133_), .A2(new_n11136_), .B(new_n11142_), .ZN(new_n11143_));
  INV_X1     g10886(.I(new_n11143_), .ZN(new_n11144_));
  NOR3_X1    g10887(.A1(new_n11133_), .A2(new_n11136_), .A3(new_n11142_), .ZN(new_n11145_));
  OAI21_X1   g10888(.A1(new_n11144_), .A2(new_n11145_), .B(new_n10819_), .ZN(new_n11146_));
  AOI21_X1   g10889(.A1(new_n11127_), .A2(new_n11131_), .B(new_n11123_), .ZN(new_n11147_));
  NOR3_X1    g10890(.A1(new_n11118_), .A2(new_n11124_), .A3(new_n11113_), .ZN(new_n11148_));
  OAI21_X1   g10891(.A1(new_n11147_), .A2(new_n11148_), .B(new_n10820_), .ZN(new_n11149_));
  NOR3_X1    g10892(.A1(new_n11118_), .A2(new_n11123_), .A3(new_n11113_), .ZN(new_n11150_));
  AOI21_X1   g10893(.A1(new_n11127_), .A2(new_n11131_), .B(new_n11124_), .ZN(new_n11151_));
  OAI21_X1   g10894(.A1(new_n11151_), .A2(new_n11150_), .B(new_n10821_), .ZN(new_n11152_));
  NAND3_X1   g10895(.A1(new_n11149_), .A2(new_n11152_), .A3(new_n11142_), .ZN(new_n11153_));
  OAI21_X1   g10896(.A1(new_n11133_), .A2(new_n11136_), .B(new_n11141_), .ZN(new_n11154_));
  NAND2_X1   g10897(.A1(new_n11154_), .A2(new_n11153_), .ZN(new_n11155_));
  NAND3_X1   g10898(.A1(new_n11155_), .A2(new_n10712_), .A3(new_n10818_), .ZN(new_n11156_));
  OAI22_X1   g10899(.A1(new_n582_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n577_), .ZN(new_n11157_));
  NAND2_X1   g10900(.A1(new_n960_), .A2(\b[57] ), .ZN(new_n11158_));
  AOI21_X1   g10901(.A1(new_n11157_), .A2(new_n11158_), .B(new_n585_), .ZN(new_n11159_));
  NAND2_X1   g10902(.A1(new_n7895_), .A2(new_n11159_), .ZN(new_n11160_));
  XOR2_X1    g10903(.A1(new_n11160_), .A2(\a[11] ), .Z(new_n11161_));
  AOI21_X1   g10904(.A1(new_n11156_), .A2(new_n11146_), .B(new_n11161_), .ZN(new_n11162_));
  NAND3_X1   g10905(.A1(new_n11149_), .A2(new_n11152_), .A3(new_n11141_), .ZN(new_n11163_));
  AOI22_X1   g10906(.A1(new_n11143_), .A2(new_n11163_), .B1(new_n10712_), .B2(new_n10818_), .ZN(new_n11164_));
  AOI21_X1   g10907(.A1(new_n11153_), .A2(new_n11154_), .B(new_n10819_), .ZN(new_n11165_));
  INV_X1     g10908(.I(new_n11161_), .ZN(new_n11166_));
  NOR3_X1    g10909(.A1(new_n11165_), .A2(new_n11164_), .A3(new_n11166_), .ZN(new_n11167_));
  OAI21_X1   g10910(.A1(new_n11162_), .A2(new_n11167_), .B(new_n10817_), .ZN(new_n11168_));
  INV_X1     g10911(.I(new_n10817_), .ZN(new_n11169_));
  NOR3_X1    g10912(.A1(new_n11165_), .A2(new_n11164_), .A3(new_n11161_), .ZN(new_n11170_));
  AOI21_X1   g10913(.A1(new_n11156_), .A2(new_n11146_), .B(new_n11166_), .ZN(new_n11171_));
  OAI21_X1   g10914(.A1(new_n11171_), .A2(new_n11170_), .B(new_n11169_), .ZN(new_n11172_));
  NAND2_X1   g10915(.A1(new_n11172_), .A2(new_n11168_), .ZN(new_n11173_));
  OAI21_X1   g10916(.A1(new_n10733_), .A2(new_n10729_), .B(new_n10743_), .ZN(new_n11174_));
  OAI22_X1   g10917(.A1(new_n437_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n431_), .ZN(new_n11175_));
  NAND2_X1   g10918(.A1(new_n775_), .A2(\b[60] ), .ZN(new_n11176_));
  AOI21_X1   g10919(.A1(new_n11175_), .A2(new_n11176_), .B(new_n440_), .ZN(new_n11177_));
  NAND2_X1   g10920(.A1(new_n8935_), .A2(new_n11177_), .ZN(new_n11178_));
  XOR2_X1    g10921(.A1(new_n11178_), .A2(\a[8] ), .Z(new_n11179_));
  NOR2_X1    g10922(.A1(new_n11174_), .A2(new_n11179_), .ZN(new_n11180_));
  AOI21_X1   g10923(.A1(new_n10719_), .A2(new_n10744_), .B(new_n10726_), .ZN(new_n11181_));
  INV_X1     g10924(.I(new_n11179_), .ZN(new_n11182_));
  NOR2_X1    g10925(.A1(new_n11181_), .A2(new_n11182_), .ZN(new_n11183_));
  OAI21_X1   g10926(.A1(new_n11180_), .A2(new_n11183_), .B(new_n11173_), .ZN(new_n11184_));
  NAND2_X1   g10927(.A1(new_n11174_), .A2(new_n11182_), .ZN(new_n11185_));
  NAND2_X1   g10928(.A1(new_n11181_), .A2(new_n11179_), .ZN(new_n11186_));
  NAND2_X1   g10929(.A1(new_n11186_), .A2(new_n11185_), .ZN(new_n11187_));
  NAND3_X1   g10930(.A1(new_n11187_), .A2(new_n11168_), .A3(new_n11172_), .ZN(new_n11188_));
  NAND2_X1   g10931(.A1(new_n11184_), .A2(new_n11188_), .ZN(new_n11189_));
  NAND2_X1   g10932(.A1(new_n11189_), .A2(new_n10816_), .ZN(new_n11190_));
  NOR2_X1    g10933(.A1(new_n11189_), .A2(new_n10816_), .ZN(new_n11191_));
  INV_X1     g10934(.I(new_n11191_), .ZN(new_n11192_));
  AOI21_X1   g10935(.A1(new_n11192_), .A2(new_n11190_), .B(\a[5] ), .ZN(new_n11193_));
  INV_X1     g10936(.I(new_n11190_), .ZN(new_n11194_));
  NOR3_X1    g10937(.A1(new_n11194_), .A2(new_n308_), .A3(new_n11191_), .ZN(new_n11195_));
  OAI21_X1   g10938(.A1(new_n11193_), .A2(new_n11195_), .B(new_n10815_), .ZN(new_n11196_));
  INV_X1     g10939(.I(new_n10815_), .ZN(new_n11197_));
  OAI21_X1   g10940(.A1(new_n11194_), .A2(new_n11191_), .B(new_n308_), .ZN(new_n11198_));
  NAND3_X1   g10941(.A1(new_n11192_), .A2(new_n11190_), .A3(\a[5] ), .ZN(new_n11199_));
  NAND3_X1   g10942(.A1(new_n11198_), .A2(new_n11199_), .A3(new_n11197_), .ZN(new_n11200_));
  NAND2_X1   g10943(.A1(new_n11196_), .A2(new_n11200_), .ZN(new_n11201_));
  XOR2_X1    g10944(.A1(new_n11201_), .A2(new_n10813_), .Z(new_n11202_));
  NAND2_X1   g10945(.A1(new_n11202_), .A2(new_n10812_), .ZN(new_n11203_));
  XOR2_X1    g10946(.A1(new_n11201_), .A2(new_n10813_), .Z(new_n11204_));
  OAI21_X1   g10947(.A1(new_n10812_), .A2(new_n11204_), .B(new_n11203_), .ZN(\f[68] ));
  INV_X1     g10948(.I(new_n11189_), .ZN(new_n11206_));
  XOR2_X1    g10949(.A1(new_n10815_), .A2(\a[5] ), .Z(new_n11207_));
  XOR2_X1    g10950(.A1(new_n10816_), .A2(new_n11207_), .Z(new_n11208_));
  OAI21_X1   g10951(.A1(new_n11206_), .A2(new_n11207_), .B(new_n11208_), .ZN(new_n11209_));
  NAND2_X1   g10952(.A1(new_n11173_), .A2(new_n11186_), .ZN(new_n11210_));
  NAND2_X1   g10953(.A1(new_n11210_), .A2(new_n11185_), .ZN(new_n11211_));
  NOR2_X1    g10954(.A1(new_n11167_), .A2(new_n11169_), .ZN(new_n11212_));
  NOR2_X1    g10955(.A1(new_n11212_), .A2(new_n11162_), .ZN(new_n11213_));
  INV_X1     g10956(.I(new_n11213_), .ZN(new_n11214_));
  AOI21_X1   g10957(.A1(new_n10820_), .A2(new_n11132_), .B(new_n11147_), .ZN(new_n11215_));
  NAND2_X1   g10958(.A1(new_n11114_), .A2(new_n11112_), .ZN(new_n11216_));
  AOI21_X1   g10959(.A1(new_n11097_), .A2(new_n11095_), .B(new_n11108_), .ZN(new_n11217_));
  AOI21_X1   g10960(.A1(new_n11078_), .A2(new_n11076_), .B(new_n11089_), .ZN(new_n11218_));
  AOI21_X1   g10961(.A1(new_n11057_), .A2(new_n11054_), .B(new_n11070_), .ZN(new_n11219_));
  INV_X1     g10962(.I(new_n11219_), .ZN(new_n11220_));
  AOI21_X1   g10963(.A1(new_n11037_), .A2(new_n11035_), .B(new_n11049_), .ZN(new_n11221_));
  INV_X1     g10964(.I(new_n11221_), .ZN(new_n11222_));
  AOI21_X1   g10965(.A1(new_n10833_), .A2(new_n10993_), .B(new_n10976_), .ZN(new_n11223_));
  OAI21_X1   g10966(.A1(new_n10942_), .A2(new_n10952_), .B(new_n10955_), .ZN(new_n11224_));
  NAND2_X1   g10967(.A1(new_n10957_), .A2(new_n10960_), .ZN(new_n11225_));
  XOR2_X1    g10968(.A1(new_n10836_), .A2(new_n4198_), .Z(new_n11226_));
  INV_X1     g10969(.I(new_n11226_), .ZN(new_n11227_));
  OAI21_X1   g10970(.A1(new_n11225_), .A2(new_n10955_), .B(new_n11227_), .ZN(new_n11228_));
  NAND2_X1   g10971(.A1(new_n11228_), .A2(new_n11224_), .ZN(new_n11229_));
  AOI21_X1   g10972(.A1(new_n10941_), .A2(new_n10943_), .B(new_n10939_), .ZN(new_n11230_));
  OAI21_X1   g10973(.A1(new_n10841_), .A2(new_n10949_), .B(new_n10931_), .ZN(new_n11231_));
  AOI21_X1   g10974(.A1(new_n10845_), .A2(new_n10923_), .B(new_n10901_), .ZN(new_n11232_));
  OAI21_X1   g10975(.A1(new_n10850_), .A2(new_n10888_), .B(new_n10886_), .ZN(new_n11233_));
  INV_X1     g10976(.I(new_n11233_), .ZN(new_n11234_));
  NOR2_X1    g10977(.A1(new_n10882_), .A2(new_n10868_), .ZN(new_n11235_));
  NOR2_X1    g10978(.A1(new_n11235_), .A2(new_n10880_), .ZN(new_n11236_));
  OAI22_X1   g10979(.A1(new_n717_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n659_), .ZN(new_n11237_));
  NAND2_X1   g10980(.A1(new_n8628_), .A2(\b[10] ), .ZN(new_n11238_));
  AOI21_X1   g10981(.A1(new_n11238_), .A2(new_n11237_), .B(new_n7354_), .ZN(new_n11239_));
  NAND2_X1   g10982(.A1(new_n716_), .A2(new_n11239_), .ZN(new_n11240_));
  XOR2_X1    g10983(.A1(new_n11240_), .A2(\a[59] ), .Z(new_n11241_));
  INV_X1     g10984(.I(new_n10862_), .ZN(new_n11242_));
  AOI21_X1   g10985(.A1(new_n10856_), .A2(new_n11242_), .B(new_n10863_), .ZN(new_n11243_));
  INV_X1     g10986(.I(new_n11243_), .ZN(new_n11244_));
  OAI22_X1   g10987(.A1(new_n510_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n495_), .ZN(new_n11245_));
  NAND2_X1   g10988(.A1(new_n9644_), .A2(\b[7] ), .ZN(new_n11246_));
  AOI21_X1   g10989(.A1(new_n11246_), .A2(new_n11245_), .B(new_n8321_), .ZN(new_n11247_));
  NAND2_X1   g10990(.A1(new_n518_), .A2(new_n11247_), .ZN(new_n11248_));
  XOR2_X1    g10991(.A1(new_n11248_), .A2(new_n8309_), .Z(new_n11249_));
  NOR2_X1    g10992(.A1(new_n8985_), .A2(new_n403_), .ZN(new_n11250_));
  NOR2_X1    g10993(.A1(new_n9364_), .A2(new_n347_), .ZN(new_n11251_));
  XNOR2_X1   g10994(.A1(new_n11250_), .A2(new_n11251_), .ZN(new_n11252_));
  NOR2_X1    g10995(.A1(new_n11252_), .A2(new_n359_), .ZN(new_n11253_));
  NOR2_X1    g10996(.A1(new_n271_), .A2(new_n308_), .ZN(new_n11254_));
  NOR2_X1    g10997(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n11255_));
  NOR2_X1    g10998(.A1(new_n11254_), .A2(new_n11255_), .ZN(new_n11256_));
  INV_X1     g10999(.I(new_n11256_), .ZN(new_n11257_));
  AOI21_X1   g11000(.A1(new_n11252_), .A2(new_n11257_), .B(new_n11253_), .ZN(new_n11258_));
  XOR2_X1    g11001(.A1(new_n11249_), .A2(new_n11258_), .Z(new_n11259_));
  NAND2_X1   g11002(.A1(new_n11259_), .A2(new_n11244_), .ZN(new_n11260_));
  NOR2_X1    g11003(.A1(new_n11249_), .A2(new_n11258_), .ZN(new_n11261_));
  AND2_X2    g11004(.A1(new_n11249_), .A2(new_n11258_), .Z(new_n11262_));
  OAI21_X1   g11005(.A1(new_n11262_), .A2(new_n11261_), .B(new_n11243_), .ZN(new_n11263_));
  NAND2_X1   g11006(.A1(new_n11260_), .A2(new_n11263_), .ZN(new_n11264_));
  NAND2_X1   g11007(.A1(new_n11264_), .A2(new_n11241_), .ZN(new_n11265_));
  NOR2_X1    g11008(.A1(new_n11264_), .A2(new_n11241_), .ZN(new_n11266_));
  INV_X1     g11009(.I(new_n11266_), .ZN(new_n11267_));
  AOI21_X1   g11010(.A1(new_n11267_), .A2(new_n11265_), .B(new_n11236_), .ZN(new_n11268_));
  INV_X1     g11011(.I(new_n10880_), .ZN(new_n11269_));
  OAI21_X1   g11012(.A1(new_n10868_), .A2(new_n10882_), .B(new_n11269_), .ZN(new_n11270_));
  XNOR2_X1   g11013(.A1(new_n11264_), .A2(new_n11241_), .ZN(new_n11271_));
  NOR2_X1    g11014(.A1(new_n11271_), .A2(new_n11270_), .ZN(new_n11272_));
  NOR2_X1    g11015(.A1(new_n11272_), .A2(new_n11268_), .ZN(new_n11273_));
  OAI22_X1   g11016(.A1(new_n6721_), .A2(new_n848_), .B1(new_n6723_), .B2(new_n904_), .ZN(new_n11274_));
  NAND2_X1   g11017(.A1(new_n7617_), .A2(\b[13] ), .ZN(new_n11275_));
  AOI21_X1   g11018(.A1(new_n11275_), .A2(new_n11274_), .B(new_n6731_), .ZN(new_n11276_));
  NAND2_X1   g11019(.A1(new_n907_), .A2(new_n11276_), .ZN(new_n11277_));
  XOR2_X1    g11020(.A1(new_n11277_), .A2(\a[56] ), .Z(new_n11278_));
  INV_X1     g11021(.I(new_n11278_), .ZN(new_n11279_));
  NAND2_X1   g11022(.A1(new_n11273_), .A2(new_n11279_), .ZN(new_n11280_));
  INV_X1     g11023(.I(new_n11265_), .ZN(new_n11281_));
  OAI21_X1   g11024(.A1(new_n11281_), .A2(new_n11266_), .B(new_n11270_), .ZN(new_n11282_));
  OAI21_X1   g11025(.A1(new_n11270_), .A2(new_n11271_), .B(new_n11282_), .ZN(new_n11283_));
  NAND2_X1   g11026(.A1(new_n11283_), .A2(new_n11278_), .ZN(new_n11284_));
  AOI21_X1   g11027(.A1(new_n11284_), .A2(new_n11280_), .B(new_n11234_), .ZN(new_n11285_));
  NAND2_X1   g11028(.A1(new_n11283_), .A2(new_n11279_), .ZN(new_n11286_));
  NAND2_X1   g11029(.A1(new_n11273_), .A2(new_n11278_), .ZN(new_n11287_));
  AOI21_X1   g11030(.A1(new_n11286_), .A2(new_n11287_), .B(new_n11233_), .ZN(new_n11288_));
  OAI22_X1   g11031(.A1(new_n5786_), .A2(new_n1124_), .B1(new_n1044_), .B2(new_n5792_), .ZN(new_n11289_));
  NAND2_X1   g11032(.A1(new_n6745_), .A2(\b[16] ), .ZN(new_n11290_));
  AOI21_X1   g11033(.A1(new_n11290_), .A2(new_n11289_), .B(new_n5796_), .ZN(new_n11291_));
  NAND2_X1   g11034(.A1(new_n1123_), .A2(new_n11291_), .ZN(new_n11292_));
  XOR2_X1    g11035(.A1(new_n11292_), .A2(\a[53] ), .Z(new_n11293_));
  INV_X1     g11036(.I(new_n11293_), .ZN(new_n11294_));
  OAI21_X1   g11037(.A1(new_n11285_), .A2(new_n11288_), .B(new_n11294_), .ZN(new_n11295_));
  NOR2_X1    g11038(.A1(new_n11283_), .A2(new_n11278_), .ZN(new_n11296_));
  NOR2_X1    g11039(.A1(new_n11273_), .A2(new_n11279_), .ZN(new_n11297_));
  OAI21_X1   g11040(.A1(new_n11296_), .A2(new_n11297_), .B(new_n11233_), .ZN(new_n11298_));
  NOR2_X1    g11041(.A1(new_n11273_), .A2(new_n11278_), .ZN(new_n11299_));
  NOR2_X1    g11042(.A1(new_n11283_), .A2(new_n11279_), .ZN(new_n11300_));
  OAI21_X1   g11043(.A1(new_n11300_), .A2(new_n11299_), .B(new_n11234_), .ZN(new_n11301_));
  NAND3_X1   g11044(.A1(new_n11298_), .A2(new_n11301_), .A3(new_n11293_), .ZN(new_n11302_));
  AOI21_X1   g11045(.A1(new_n11295_), .A2(new_n11302_), .B(new_n11232_), .ZN(new_n11303_));
  OAI21_X1   g11046(.A1(new_n10844_), .A2(new_n10910_), .B(new_n10922_), .ZN(new_n11304_));
  NAND3_X1   g11047(.A1(new_n11298_), .A2(new_n11301_), .A3(new_n11294_), .ZN(new_n11305_));
  OAI21_X1   g11048(.A1(new_n11285_), .A2(new_n11288_), .B(new_n11293_), .ZN(new_n11306_));
  AOI21_X1   g11049(.A1(new_n11306_), .A2(new_n11305_), .B(new_n11304_), .ZN(new_n11307_));
  OAI22_X1   g11050(.A1(new_n5228_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n5225_), .ZN(new_n11308_));
  NAND2_X1   g11051(.A1(new_n5387_), .A2(\b[19] ), .ZN(new_n11309_));
  AOI21_X1   g11052(.A1(new_n11308_), .A2(new_n11309_), .B(new_n5231_), .ZN(new_n11310_));
  AND3_X2    g11053(.A1(new_n1396_), .A2(new_n5220_), .A3(new_n11310_), .Z(new_n11311_));
  AOI21_X1   g11054(.A1(new_n1396_), .A2(new_n11310_), .B(new_n5220_), .ZN(new_n11312_));
  NOR2_X1    g11055(.A1(new_n11311_), .A2(new_n11312_), .ZN(new_n11313_));
  NOR3_X1    g11056(.A1(new_n11303_), .A2(new_n11307_), .A3(new_n11313_), .ZN(new_n11314_));
  AOI21_X1   g11057(.A1(new_n11298_), .A2(new_n11301_), .B(new_n11293_), .ZN(new_n11315_));
  NOR3_X1    g11058(.A1(new_n11285_), .A2(new_n11288_), .A3(new_n11294_), .ZN(new_n11316_));
  OAI21_X1   g11059(.A1(new_n11315_), .A2(new_n11316_), .B(new_n11304_), .ZN(new_n11317_));
  NOR3_X1    g11060(.A1(new_n11285_), .A2(new_n11288_), .A3(new_n11293_), .ZN(new_n11318_));
  AOI21_X1   g11061(.A1(new_n11298_), .A2(new_n11301_), .B(new_n11294_), .ZN(new_n11319_));
  OAI21_X1   g11062(.A1(new_n11319_), .A2(new_n11318_), .B(new_n11232_), .ZN(new_n11320_));
  INV_X1     g11063(.I(new_n11313_), .ZN(new_n11321_));
  AOI21_X1   g11064(.A1(new_n11317_), .A2(new_n11320_), .B(new_n11321_), .ZN(new_n11322_));
  OAI21_X1   g11065(.A1(new_n11322_), .A2(new_n11314_), .B(new_n11231_), .ZN(new_n11323_));
  AOI21_X1   g11066(.A1(new_n10930_), .A2(new_n10932_), .B(new_n10948_), .ZN(new_n11324_));
  AOI21_X1   g11067(.A1(new_n11317_), .A2(new_n11320_), .B(new_n11313_), .ZN(new_n11325_));
  NOR3_X1    g11068(.A1(new_n11303_), .A2(new_n11307_), .A3(new_n11321_), .ZN(new_n11326_));
  OAI21_X1   g11069(.A1(new_n11325_), .A2(new_n11326_), .B(new_n11324_), .ZN(new_n11327_));
  OAI22_X1   g11070(.A1(new_n4711_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n4706_), .ZN(new_n11328_));
  NAND2_X1   g11071(.A1(new_n5814_), .A2(\b[22] ), .ZN(new_n11329_));
  AOI21_X1   g11072(.A1(new_n11328_), .A2(new_n11329_), .B(new_n4714_), .ZN(new_n11330_));
  NAND2_X1   g11073(.A1(new_n1708_), .A2(new_n11330_), .ZN(new_n11331_));
  XOR2_X1    g11074(.A1(new_n11331_), .A2(\a[47] ), .Z(new_n11332_));
  INV_X1     g11075(.I(new_n11332_), .ZN(new_n11333_));
  NAND3_X1   g11076(.A1(new_n11323_), .A2(new_n11327_), .A3(new_n11333_), .ZN(new_n11334_));
  NAND3_X1   g11077(.A1(new_n11317_), .A2(new_n11320_), .A3(new_n11321_), .ZN(new_n11335_));
  OAI21_X1   g11078(.A1(new_n11303_), .A2(new_n11307_), .B(new_n11313_), .ZN(new_n11336_));
  AOI21_X1   g11079(.A1(new_n11336_), .A2(new_n11335_), .B(new_n11324_), .ZN(new_n11337_));
  OAI21_X1   g11080(.A1(new_n11303_), .A2(new_n11307_), .B(new_n11321_), .ZN(new_n11338_));
  NAND3_X1   g11081(.A1(new_n11317_), .A2(new_n11320_), .A3(new_n11313_), .ZN(new_n11339_));
  AOI21_X1   g11082(.A1(new_n11338_), .A2(new_n11339_), .B(new_n11231_), .ZN(new_n11340_));
  OAI21_X1   g11083(.A1(new_n11340_), .A2(new_n11337_), .B(new_n11332_), .ZN(new_n11341_));
  AOI21_X1   g11084(.A1(new_n11341_), .A2(new_n11334_), .B(new_n11230_), .ZN(new_n11342_));
  AOI21_X1   g11085(.A1(new_n11323_), .A2(new_n11327_), .B(new_n11332_), .ZN(new_n11343_));
  NOR3_X1    g11086(.A1(new_n11340_), .A2(new_n11337_), .A3(new_n11333_), .ZN(new_n11344_));
  OAI21_X1   g11087(.A1(new_n11343_), .A2(new_n11344_), .B(new_n11230_), .ZN(new_n11345_));
  INV_X1     g11088(.I(new_n11345_), .ZN(new_n11346_));
  OAI22_X1   g11089(.A1(new_n4208_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n4203_), .ZN(new_n11347_));
  NAND2_X1   g11090(.A1(new_n5244_), .A2(\b[25] ), .ZN(new_n11348_));
  AOI21_X1   g11091(.A1(new_n11347_), .A2(new_n11348_), .B(new_n4211_), .ZN(new_n11349_));
  NAND2_X1   g11092(.A1(new_n2042_), .A2(new_n11349_), .ZN(new_n11350_));
  XOR2_X1    g11093(.A1(new_n11350_), .A2(\a[44] ), .Z(new_n11351_));
  INV_X1     g11094(.I(new_n11351_), .ZN(new_n11352_));
  OAI21_X1   g11095(.A1(new_n11346_), .A2(new_n11342_), .B(new_n11352_), .ZN(new_n11353_));
  INV_X1     g11096(.I(new_n11342_), .ZN(new_n11354_));
  NAND3_X1   g11097(.A1(new_n11354_), .A2(new_n11345_), .A3(new_n11351_), .ZN(new_n11355_));
  NAND2_X1   g11098(.A1(new_n11353_), .A2(new_n11355_), .ZN(new_n11356_));
  NAND2_X1   g11099(.A1(new_n11356_), .A2(new_n11229_), .ZN(new_n11357_));
  INV_X1     g11100(.I(new_n11229_), .ZN(new_n11358_));
  NAND3_X1   g11101(.A1(new_n11354_), .A2(new_n11345_), .A3(new_n11352_), .ZN(new_n11359_));
  INV_X1     g11102(.I(new_n11359_), .ZN(new_n11360_));
  AOI21_X1   g11103(.A1(new_n11354_), .A2(new_n11345_), .B(new_n11352_), .ZN(new_n11361_));
  OAI21_X1   g11104(.A1(new_n11361_), .A2(new_n11360_), .B(new_n11358_), .ZN(new_n11362_));
  OAI22_X1   g11105(.A1(new_n3736_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n3731_), .ZN(new_n11363_));
  NAND2_X1   g11106(.A1(new_n4730_), .A2(\b[28] ), .ZN(new_n11364_));
  AOI21_X1   g11107(.A1(new_n11363_), .A2(new_n11364_), .B(new_n3739_), .ZN(new_n11365_));
  NAND2_X1   g11108(.A1(new_n2404_), .A2(new_n11365_), .ZN(new_n11366_));
  XOR2_X1    g11109(.A1(new_n11366_), .A2(\a[41] ), .Z(new_n11367_));
  INV_X1     g11110(.I(new_n11367_), .ZN(new_n11368_));
  NAND3_X1   g11111(.A1(new_n11362_), .A2(new_n11357_), .A3(new_n11368_), .ZN(new_n11369_));
  AOI21_X1   g11112(.A1(new_n11353_), .A2(new_n11355_), .B(new_n11358_), .ZN(new_n11370_));
  INV_X1     g11113(.I(new_n11361_), .ZN(new_n11371_));
  AOI21_X1   g11114(.A1(new_n11371_), .A2(new_n11359_), .B(new_n11229_), .ZN(new_n11372_));
  OAI21_X1   g11115(.A1(new_n11370_), .A2(new_n11372_), .B(new_n11367_), .ZN(new_n11373_));
  AOI21_X1   g11116(.A1(new_n11369_), .A2(new_n11373_), .B(new_n11223_), .ZN(new_n11374_));
  OAI21_X1   g11117(.A1(new_n10832_), .A2(new_n10980_), .B(new_n10992_), .ZN(new_n11375_));
  OAI21_X1   g11118(.A1(new_n11370_), .A2(new_n11372_), .B(new_n11368_), .ZN(new_n11376_));
  NAND3_X1   g11119(.A1(new_n11362_), .A2(new_n11357_), .A3(new_n11367_), .ZN(new_n11377_));
  AOI21_X1   g11120(.A1(new_n11376_), .A2(new_n11377_), .B(new_n11375_), .ZN(new_n11378_));
  OAI22_X1   g11121(.A1(new_n3298_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n3293_), .ZN(new_n11379_));
  NAND2_X1   g11122(.A1(new_n4227_), .A2(\b[31] ), .ZN(new_n11380_));
  AOI21_X1   g11123(.A1(new_n11379_), .A2(new_n11380_), .B(new_n3301_), .ZN(new_n11381_));
  NAND2_X1   g11124(.A1(new_n2797_), .A2(new_n11381_), .ZN(new_n11382_));
  XOR2_X1    g11125(.A1(new_n11382_), .A2(\a[38] ), .Z(new_n11383_));
  INV_X1     g11126(.I(new_n11383_), .ZN(new_n11384_));
  OAI21_X1   g11127(.A1(new_n11378_), .A2(new_n11374_), .B(new_n11384_), .ZN(new_n11385_));
  INV_X1     g11128(.I(new_n11385_), .ZN(new_n11386_));
  NOR3_X1    g11129(.A1(new_n11378_), .A2(new_n11374_), .A3(new_n11384_), .ZN(new_n11387_));
  NOR2_X1    g11130(.A1(new_n11386_), .A2(new_n11387_), .ZN(new_n11388_));
  OAI22_X1   g11131(.A1(new_n2846_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n2841_), .ZN(new_n11389_));
  NAND2_X1   g11132(.A1(new_n3755_), .A2(\b[34] ), .ZN(new_n11390_));
  AOI21_X1   g11133(.A1(new_n11389_), .A2(new_n11390_), .B(new_n2849_), .ZN(new_n11391_));
  NAND2_X1   g11134(.A1(new_n3246_), .A2(new_n11391_), .ZN(new_n11392_));
  XOR2_X1    g11135(.A1(new_n11392_), .A2(\a[35] ), .Z(new_n11393_));
  INV_X1     g11136(.I(new_n11393_), .ZN(new_n11394_));
  NAND2_X1   g11137(.A1(new_n11012_), .A2(new_n10829_), .ZN(new_n11395_));
  AOI21_X1   g11138(.A1(new_n11000_), .A2(new_n11002_), .B(new_n11018_), .ZN(new_n11396_));
  INV_X1     g11139(.I(new_n11396_), .ZN(new_n11397_));
  NAND3_X1   g11140(.A1(new_n11395_), .A2(new_n11011_), .A3(new_n11397_), .ZN(new_n11398_));
  AOI21_X1   g11141(.A1(new_n11395_), .A2(new_n11011_), .B(new_n11397_), .ZN(new_n11399_));
  INV_X1     g11142(.I(new_n11399_), .ZN(new_n11400_));
  AOI21_X1   g11143(.A1(new_n11400_), .A2(new_n11398_), .B(new_n11394_), .ZN(new_n11401_));
  INV_X1     g11144(.I(new_n11398_), .ZN(new_n11402_));
  NOR3_X1    g11145(.A1(new_n11402_), .A2(new_n11393_), .A3(new_n11399_), .ZN(new_n11403_));
  OAI21_X1   g11146(.A1(new_n11401_), .A2(new_n11403_), .B(new_n11388_), .ZN(new_n11404_));
  INV_X1     g11147(.I(new_n11387_), .ZN(new_n11405_));
  NAND2_X1   g11148(.A1(new_n11405_), .A2(new_n11385_), .ZN(new_n11406_));
  OAI21_X1   g11149(.A1(new_n11402_), .A2(new_n11399_), .B(new_n11393_), .ZN(new_n11407_));
  NAND3_X1   g11150(.A1(new_n11400_), .A2(new_n11394_), .A3(new_n11398_), .ZN(new_n11408_));
  NAND3_X1   g11151(.A1(new_n11408_), .A2(new_n11407_), .A3(new_n11406_), .ZN(new_n11409_));
  OAI22_X1   g11152(.A1(new_n2452_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n2447_), .ZN(new_n11410_));
  NAND2_X1   g11153(.A1(new_n3312_), .A2(\b[37] ), .ZN(new_n11411_));
  AOI21_X1   g11154(.A1(new_n11410_), .A2(new_n11411_), .B(new_n2455_), .ZN(new_n11412_));
  NAND2_X1   g11155(.A1(new_n3700_), .A2(new_n11412_), .ZN(new_n11413_));
  XOR2_X1    g11156(.A1(new_n11413_), .A2(\a[32] ), .Z(new_n11414_));
  AOI21_X1   g11157(.A1(new_n11404_), .A2(new_n11409_), .B(new_n11414_), .ZN(new_n11415_));
  AOI21_X1   g11158(.A1(new_n11408_), .A2(new_n11407_), .B(new_n11406_), .ZN(new_n11416_));
  NOR3_X1    g11159(.A1(new_n11401_), .A2(new_n11403_), .A3(new_n11388_), .ZN(new_n11417_));
  INV_X1     g11160(.I(new_n11414_), .ZN(new_n11418_));
  NOR3_X1    g11161(.A1(new_n11416_), .A2(new_n11417_), .A3(new_n11418_), .ZN(new_n11419_));
  OAI21_X1   g11162(.A1(new_n11419_), .A2(new_n11415_), .B(new_n11222_), .ZN(new_n11420_));
  NOR3_X1    g11163(.A1(new_n11416_), .A2(new_n11417_), .A3(new_n11414_), .ZN(new_n11421_));
  AOI21_X1   g11164(.A1(new_n11404_), .A2(new_n11409_), .B(new_n11418_), .ZN(new_n11422_));
  OAI21_X1   g11165(.A1(new_n11421_), .A2(new_n11422_), .B(new_n11221_), .ZN(new_n11423_));
  OAI22_X1   g11166(.A1(new_n2084_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n2079_), .ZN(new_n11424_));
  NAND2_X1   g11167(.A1(new_n2864_), .A2(\b[40] ), .ZN(new_n11425_));
  AOI21_X1   g11168(.A1(new_n11424_), .A2(new_n11425_), .B(new_n2087_), .ZN(new_n11426_));
  NAND2_X1   g11169(.A1(new_n4017_), .A2(new_n11426_), .ZN(new_n11427_));
  XOR2_X1    g11170(.A1(new_n11427_), .A2(\a[29] ), .Z(new_n11428_));
  AOI21_X1   g11171(.A1(new_n11420_), .A2(new_n11423_), .B(new_n11428_), .ZN(new_n11429_));
  OAI21_X1   g11172(.A1(new_n11416_), .A2(new_n11417_), .B(new_n11418_), .ZN(new_n11430_));
  NAND3_X1   g11173(.A1(new_n11404_), .A2(new_n11409_), .A3(new_n11414_), .ZN(new_n11431_));
  AOI21_X1   g11174(.A1(new_n11430_), .A2(new_n11431_), .B(new_n11221_), .ZN(new_n11432_));
  NAND3_X1   g11175(.A1(new_n11404_), .A2(new_n11409_), .A3(new_n11418_), .ZN(new_n11433_));
  OAI21_X1   g11176(.A1(new_n11416_), .A2(new_n11417_), .B(new_n11414_), .ZN(new_n11434_));
  AOI21_X1   g11177(.A1(new_n11434_), .A2(new_n11433_), .B(new_n11222_), .ZN(new_n11435_));
  INV_X1     g11178(.I(new_n11428_), .ZN(new_n11436_));
  NOR3_X1    g11179(.A1(new_n11432_), .A2(new_n11435_), .A3(new_n11436_), .ZN(new_n11437_));
  OAI21_X1   g11180(.A1(new_n11429_), .A2(new_n11437_), .B(new_n11220_), .ZN(new_n11438_));
  NOR3_X1    g11181(.A1(new_n11432_), .A2(new_n11435_), .A3(new_n11428_), .ZN(new_n11439_));
  AOI21_X1   g11182(.A1(new_n11420_), .A2(new_n11423_), .B(new_n11436_), .ZN(new_n11440_));
  OAI21_X1   g11183(.A1(new_n11440_), .A2(new_n11439_), .B(new_n11219_), .ZN(new_n11441_));
  OAI22_X1   g11184(.A1(new_n1760_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n1755_), .ZN(new_n11442_));
  NAND2_X1   g11185(.A1(new_n2470_), .A2(\b[43] ), .ZN(new_n11443_));
  AOI21_X1   g11186(.A1(new_n11442_), .A2(new_n11443_), .B(new_n1763_), .ZN(new_n11444_));
  NAND3_X1   g11187(.A1(new_n4513_), .A2(new_n1750_), .A3(new_n11444_), .ZN(new_n11445_));
  INV_X1     g11188(.I(new_n11445_), .ZN(new_n11446_));
  AOI21_X1   g11189(.A1(new_n4513_), .A2(new_n11444_), .B(new_n1750_), .ZN(new_n11447_));
  NOR2_X1    g11190(.A1(new_n11446_), .A2(new_n11447_), .ZN(new_n11448_));
  INV_X1     g11191(.I(new_n11448_), .ZN(new_n11449_));
  NAND3_X1   g11192(.A1(new_n11438_), .A2(new_n11441_), .A3(new_n11449_), .ZN(new_n11450_));
  OAI21_X1   g11193(.A1(new_n11432_), .A2(new_n11435_), .B(new_n11436_), .ZN(new_n11451_));
  NAND3_X1   g11194(.A1(new_n11420_), .A2(new_n11423_), .A3(new_n11428_), .ZN(new_n11452_));
  AOI21_X1   g11195(.A1(new_n11451_), .A2(new_n11452_), .B(new_n11219_), .ZN(new_n11453_));
  NAND3_X1   g11196(.A1(new_n11420_), .A2(new_n11423_), .A3(new_n11436_), .ZN(new_n11454_));
  OAI21_X1   g11197(.A1(new_n11432_), .A2(new_n11435_), .B(new_n11428_), .ZN(new_n11455_));
  AOI21_X1   g11198(.A1(new_n11455_), .A2(new_n11454_), .B(new_n11220_), .ZN(new_n11456_));
  OAI21_X1   g11199(.A1(new_n11453_), .A2(new_n11456_), .B(new_n11448_), .ZN(new_n11457_));
  AOI21_X1   g11200(.A1(new_n11457_), .A2(new_n11450_), .B(new_n11218_), .ZN(new_n11458_));
  INV_X1     g11201(.I(new_n11218_), .ZN(new_n11459_));
  OAI21_X1   g11202(.A1(new_n11453_), .A2(new_n11456_), .B(new_n11449_), .ZN(new_n11460_));
  NAND3_X1   g11203(.A1(new_n11438_), .A2(new_n11441_), .A3(new_n11448_), .ZN(new_n11461_));
  AOI21_X1   g11204(.A1(new_n11460_), .A2(new_n11461_), .B(new_n11459_), .ZN(new_n11462_));
  OAI22_X1   g11205(.A1(new_n1444_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n1439_), .ZN(new_n11463_));
  NAND2_X1   g11206(.A1(new_n2098_), .A2(\b[46] ), .ZN(new_n11464_));
  AOI21_X1   g11207(.A1(new_n11463_), .A2(new_n11464_), .B(new_n1447_), .ZN(new_n11465_));
  NAND2_X1   g11208(.A1(new_n5177_), .A2(new_n11465_), .ZN(new_n11466_));
  XOR2_X1    g11209(.A1(new_n11466_), .A2(\a[23] ), .Z(new_n11467_));
  INV_X1     g11210(.I(new_n11467_), .ZN(new_n11468_));
  OAI21_X1   g11211(.A1(new_n11458_), .A2(new_n11462_), .B(new_n11468_), .ZN(new_n11469_));
  NOR3_X1    g11212(.A1(new_n11453_), .A2(new_n11456_), .A3(new_n11448_), .ZN(new_n11470_));
  AOI21_X1   g11213(.A1(new_n11438_), .A2(new_n11441_), .B(new_n11449_), .ZN(new_n11471_));
  OAI21_X1   g11214(.A1(new_n11471_), .A2(new_n11470_), .B(new_n11459_), .ZN(new_n11472_));
  AOI21_X1   g11215(.A1(new_n11438_), .A2(new_n11441_), .B(new_n11448_), .ZN(new_n11473_));
  NOR3_X1    g11216(.A1(new_n11453_), .A2(new_n11456_), .A3(new_n11449_), .ZN(new_n11474_));
  OAI21_X1   g11217(.A1(new_n11473_), .A2(new_n11474_), .B(new_n11218_), .ZN(new_n11475_));
  NAND3_X1   g11218(.A1(new_n11472_), .A2(new_n11475_), .A3(new_n11467_), .ZN(new_n11476_));
  AOI21_X1   g11219(.A1(new_n11469_), .A2(new_n11476_), .B(new_n11217_), .ZN(new_n11477_));
  INV_X1     g11220(.I(new_n11217_), .ZN(new_n11478_));
  NAND3_X1   g11221(.A1(new_n11472_), .A2(new_n11475_), .A3(new_n11468_), .ZN(new_n11479_));
  OAI21_X1   g11222(.A1(new_n11458_), .A2(new_n11462_), .B(new_n11467_), .ZN(new_n11480_));
  AOI21_X1   g11223(.A1(new_n11480_), .A2(new_n11479_), .B(new_n11478_), .ZN(new_n11481_));
  OAI22_X1   g11224(.A1(new_n1168_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n1163_), .ZN(new_n11482_));
  NAND2_X1   g11225(.A1(new_n1774_), .A2(\b[49] ), .ZN(new_n11483_));
  AOI21_X1   g11226(.A1(new_n11482_), .A2(new_n11483_), .B(new_n1171_), .ZN(new_n11484_));
  NAND2_X1   g11227(.A1(new_n5741_), .A2(new_n11484_), .ZN(new_n11485_));
  XOR2_X1    g11228(.A1(new_n11485_), .A2(\a[20] ), .Z(new_n11486_));
  INV_X1     g11229(.I(new_n11486_), .ZN(new_n11487_));
  OAI21_X1   g11230(.A1(new_n11477_), .A2(new_n11481_), .B(new_n11487_), .ZN(new_n11488_));
  AOI21_X1   g11231(.A1(new_n11472_), .A2(new_n11475_), .B(new_n11467_), .ZN(new_n11489_));
  NOR3_X1    g11232(.A1(new_n11458_), .A2(new_n11462_), .A3(new_n11468_), .ZN(new_n11490_));
  OAI21_X1   g11233(.A1(new_n11489_), .A2(new_n11490_), .B(new_n11478_), .ZN(new_n11491_));
  INV_X1     g11234(.I(new_n11481_), .ZN(new_n11492_));
  NAND3_X1   g11235(.A1(new_n11492_), .A2(new_n11491_), .A3(new_n11486_), .ZN(new_n11493_));
  AOI22_X1   g11236(.A1(new_n11493_), .A2(new_n11488_), .B1(new_n11107_), .B2(new_n11216_), .ZN(new_n11494_));
  NAND2_X1   g11237(.A1(new_n11216_), .A2(new_n11107_), .ZN(new_n11495_));
  NAND3_X1   g11238(.A1(new_n11492_), .A2(new_n11491_), .A3(new_n11487_), .ZN(new_n11496_));
  OAI21_X1   g11239(.A1(new_n11477_), .A2(new_n11481_), .B(new_n11486_), .ZN(new_n11497_));
  AOI21_X1   g11240(.A1(new_n11496_), .A2(new_n11497_), .B(new_n11495_), .ZN(new_n11498_));
  OAI22_X1   g11241(.A1(new_n940_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n935_), .ZN(new_n11499_));
  NAND2_X1   g11242(.A1(new_n1458_), .A2(\b[52] ), .ZN(new_n11500_));
  AOI21_X1   g11243(.A1(new_n11499_), .A2(new_n11500_), .B(new_n943_), .ZN(new_n11501_));
  NAND2_X1   g11244(.A1(new_n6237_), .A2(new_n11501_), .ZN(new_n11502_));
  XOR2_X1    g11245(.A1(new_n11502_), .A2(\a[17] ), .Z(new_n11503_));
  INV_X1     g11246(.I(new_n11503_), .ZN(new_n11504_));
  OAI21_X1   g11247(.A1(new_n11494_), .A2(new_n11498_), .B(new_n11504_), .ZN(new_n11505_));
  NAND2_X1   g11248(.A1(new_n11493_), .A2(new_n11488_), .ZN(new_n11506_));
  NAND2_X1   g11249(.A1(new_n11506_), .A2(new_n11495_), .ZN(new_n11507_));
  NAND2_X1   g11250(.A1(new_n11496_), .A2(new_n11497_), .ZN(new_n11508_));
  NAND3_X1   g11251(.A1(new_n11508_), .A2(new_n11107_), .A3(new_n11216_), .ZN(new_n11509_));
  NAND3_X1   g11252(.A1(new_n11509_), .A2(new_n11507_), .A3(new_n11503_), .ZN(new_n11510_));
  AOI21_X1   g11253(.A1(new_n11510_), .A2(new_n11505_), .B(new_n11215_), .ZN(new_n11511_));
  INV_X1     g11254(.I(new_n11215_), .ZN(new_n11512_));
  NAND3_X1   g11255(.A1(new_n11509_), .A2(new_n11507_), .A3(new_n11504_), .ZN(new_n11513_));
  OAI21_X1   g11256(.A1(new_n11494_), .A2(new_n11498_), .B(new_n11503_), .ZN(new_n11514_));
  AOI21_X1   g11257(.A1(new_n11513_), .A2(new_n11514_), .B(new_n11512_), .ZN(new_n11515_));
  OR2_X2     g11258(.A1(new_n11511_), .A2(new_n11515_), .Z(new_n11516_));
  AOI21_X1   g11259(.A1(new_n10819_), .A2(new_n11163_), .B(new_n11144_), .ZN(new_n11517_));
  OAI22_X1   g11260(.A1(new_n757_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n752_), .ZN(new_n11518_));
  NAND2_X1   g11261(.A1(new_n1182_), .A2(\b[55] ), .ZN(new_n11519_));
  AOI21_X1   g11262(.A1(new_n11518_), .A2(new_n11519_), .B(new_n760_), .ZN(new_n11520_));
  NAND2_X1   g11263(.A1(new_n7308_), .A2(new_n11520_), .ZN(new_n11521_));
  XOR2_X1    g11264(.A1(new_n11521_), .A2(\a[14] ), .Z(new_n11522_));
  NOR2_X1    g11265(.A1(new_n11517_), .A2(new_n11522_), .ZN(new_n11523_));
  NAND2_X1   g11266(.A1(new_n10819_), .A2(new_n11163_), .ZN(new_n11524_));
  NAND2_X1   g11267(.A1(new_n11524_), .A2(new_n11143_), .ZN(new_n11525_));
  INV_X1     g11268(.I(new_n11522_), .ZN(new_n11526_));
  NOR2_X1    g11269(.A1(new_n11525_), .A2(new_n11526_), .ZN(new_n11527_));
  OAI21_X1   g11270(.A1(new_n11523_), .A2(new_n11527_), .B(new_n11516_), .ZN(new_n11528_));
  NOR2_X1    g11271(.A1(new_n11511_), .A2(new_n11515_), .ZN(new_n11529_));
  NOR2_X1    g11272(.A1(new_n11525_), .A2(new_n11522_), .ZN(new_n11530_));
  NOR2_X1    g11273(.A1(new_n11517_), .A2(new_n11526_), .ZN(new_n11531_));
  OAI21_X1   g11274(.A1(new_n11531_), .A2(new_n11530_), .B(new_n11529_), .ZN(new_n11532_));
  OAI22_X1   g11275(.A1(new_n582_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n577_), .ZN(new_n11533_));
  NAND2_X1   g11276(.A1(new_n960_), .A2(\b[58] ), .ZN(new_n11534_));
  AOI21_X1   g11277(.A1(new_n11533_), .A2(new_n11534_), .B(new_n585_), .ZN(new_n11535_));
  NAND2_X1   g11278(.A1(new_n7929_), .A2(new_n11535_), .ZN(new_n11536_));
  XOR2_X1    g11279(.A1(new_n11536_), .A2(\a[11] ), .Z(new_n11537_));
  AOI21_X1   g11280(.A1(new_n11528_), .A2(new_n11532_), .B(new_n11537_), .ZN(new_n11538_));
  NAND2_X1   g11281(.A1(new_n11525_), .A2(new_n11526_), .ZN(new_n11539_));
  NAND2_X1   g11282(.A1(new_n11517_), .A2(new_n11522_), .ZN(new_n11540_));
  AOI21_X1   g11283(.A1(new_n11540_), .A2(new_n11539_), .B(new_n11529_), .ZN(new_n11541_));
  NAND2_X1   g11284(.A1(new_n11517_), .A2(new_n11526_), .ZN(new_n11542_));
  NAND2_X1   g11285(.A1(new_n11525_), .A2(new_n11522_), .ZN(new_n11543_));
  AOI21_X1   g11286(.A1(new_n11542_), .A2(new_n11543_), .B(new_n11516_), .ZN(new_n11544_));
  INV_X1     g11287(.I(new_n11537_), .ZN(new_n11545_));
  NOR3_X1    g11288(.A1(new_n11544_), .A2(new_n11541_), .A3(new_n11545_), .ZN(new_n11546_));
  OAI21_X1   g11289(.A1(new_n11546_), .A2(new_n11538_), .B(new_n11214_), .ZN(new_n11547_));
  NOR3_X1    g11290(.A1(new_n11544_), .A2(new_n11541_), .A3(new_n11537_), .ZN(new_n11548_));
  AOI21_X1   g11291(.A1(new_n11528_), .A2(new_n11532_), .B(new_n11545_), .ZN(new_n11549_));
  OAI21_X1   g11292(.A1(new_n11548_), .A2(new_n11549_), .B(new_n11213_), .ZN(new_n11550_));
  AOI22_X1   g11293(.A1(new_n436_), .A2(\b[63] ), .B1(new_n686_), .B2(\b[62] ), .ZN(new_n11551_));
  NOR2_X1    g11294(.A1(new_n474_), .A2(new_n8548_), .ZN(new_n11552_));
  OAI21_X1   g11295(.A1(new_n11551_), .A2(new_n11552_), .B(new_n439_), .ZN(new_n11553_));
  NOR2_X1    g11296(.A1(new_n8962_), .A2(new_n11553_), .ZN(new_n11554_));
  XOR2_X1    g11297(.A1(new_n11554_), .A2(new_n429_), .Z(new_n11555_));
  AOI21_X1   g11298(.A1(new_n11547_), .A2(new_n11550_), .B(new_n11555_), .ZN(new_n11556_));
  OAI21_X1   g11299(.A1(new_n11544_), .A2(new_n11541_), .B(new_n11545_), .ZN(new_n11557_));
  NAND3_X1   g11300(.A1(new_n11528_), .A2(new_n11532_), .A3(new_n11537_), .ZN(new_n11558_));
  AOI21_X1   g11301(.A1(new_n11557_), .A2(new_n11558_), .B(new_n11213_), .ZN(new_n11559_));
  NAND3_X1   g11302(.A1(new_n11528_), .A2(new_n11532_), .A3(new_n11545_), .ZN(new_n11560_));
  OAI21_X1   g11303(.A1(new_n11544_), .A2(new_n11541_), .B(new_n11537_), .ZN(new_n11561_));
  AOI21_X1   g11304(.A1(new_n11561_), .A2(new_n11560_), .B(new_n11214_), .ZN(new_n11562_));
  INV_X1     g11305(.I(new_n11555_), .ZN(new_n11563_));
  NOR3_X1    g11306(.A1(new_n11559_), .A2(new_n11562_), .A3(new_n11563_), .ZN(new_n11564_));
  OAI21_X1   g11307(.A1(new_n11556_), .A2(new_n11564_), .B(new_n11211_), .ZN(new_n11565_));
  INV_X1     g11308(.I(new_n11211_), .ZN(new_n11566_));
  NOR3_X1    g11309(.A1(new_n11562_), .A2(new_n11559_), .A3(new_n11555_), .ZN(new_n11567_));
  AOI21_X1   g11310(.A1(new_n11547_), .A2(new_n11550_), .B(new_n11563_), .ZN(new_n11568_));
  OAI21_X1   g11311(.A1(new_n11568_), .A2(new_n11567_), .B(new_n11566_), .ZN(new_n11569_));
  NAND2_X1   g11312(.A1(new_n11565_), .A2(new_n11569_), .ZN(new_n11570_));
  XNOR2_X1   g11313(.A1(new_n11570_), .A2(new_n11209_), .ZN(new_n11571_));
  AOI21_X1   g11314(.A1(new_n11198_), .A2(new_n11199_), .B(new_n11197_), .ZN(new_n11572_));
  NOR3_X1    g11315(.A1(new_n11193_), .A2(new_n11195_), .A3(new_n10815_), .ZN(new_n11573_));
  NOR2_X1    g11316(.A1(new_n11572_), .A2(new_n11573_), .ZN(new_n11574_));
  AOI21_X1   g11317(.A1(new_n10808_), .A2(new_n10807_), .B(new_n10806_), .ZN(new_n11575_));
  OAI21_X1   g11318(.A1(new_n10024_), .A2(new_n10787_), .B(new_n10782_), .ZN(new_n11576_));
  INV_X1     g11319(.I(new_n11576_), .ZN(new_n11577_));
  NOR3_X1    g11320(.A1(new_n11575_), .A2(new_n11577_), .A3(new_n10813_), .ZN(new_n11578_));
  INV_X1     g11321(.I(new_n10813_), .ZN(new_n11579_));
  AOI21_X1   g11322(.A1(new_n10805_), .A2(new_n11576_), .B(new_n11579_), .ZN(new_n11580_));
  OAI21_X1   g11323(.A1(new_n11580_), .A2(new_n11578_), .B(new_n11574_), .ZN(new_n11581_));
  XOR2_X1    g11324(.A1(new_n11581_), .A2(new_n11571_), .Z(new_n11582_));
  NAND2_X1   g11325(.A1(new_n10812_), .A2(new_n11579_), .ZN(new_n11583_));
  XOR2_X1    g11326(.A1(new_n11582_), .A2(new_n11583_), .Z(\f[69] ));
  AOI21_X1   g11327(.A1(new_n11214_), .A2(new_n11558_), .B(new_n11538_), .ZN(new_n11585_));
  AOI21_X1   g11328(.A1(new_n11516_), .A2(new_n11540_), .B(new_n11523_), .ZN(new_n11586_));
  NAND2_X1   g11329(.A1(new_n11510_), .A2(new_n11512_), .ZN(new_n11587_));
  NAND2_X1   g11330(.A1(new_n11587_), .A2(new_n11505_), .ZN(new_n11588_));
  NAND2_X1   g11331(.A1(new_n11493_), .A2(new_n11495_), .ZN(new_n11589_));
  OAI21_X1   g11332(.A1(new_n11217_), .A2(new_n11490_), .B(new_n11469_), .ZN(new_n11590_));
  OAI21_X1   g11333(.A1(new_n11218_), .A2(new_n11471_), .B(new_n11450_), .ZN(new_n11591_));
  OAI21_X1   g11334(.A1(new_n11219_), .A2(new_n11440_), .B(new_n11454_), .ZN(new_n11592_));
  OAI21_X1   g11335(.A1(new_n11221_), .A2(new_n11422_), .B(new_n11433_), .ZN(new_n11593_));
  AOI21_X1   g11336(.A1(new_n11395_), .A2(new_n11011_), .B(new_n11393_), .ZN(new_n11594_));
  NAND2_X1   g11337(.A1(new_n11395_), .A2(new_n11011_), .ZN(new_n11595_));
  NOR2_X1    g11338(.A1(new_n11406_), .A2(new_n11396_), .ZN(new_n11596_));
  NOR2_X1    g11339(.A1(new_n11388_), .A2(new_n11397_), .ZN(new_n11597_));
  OAI21_X1   g11340(.A1(new_n11597_), .A2(new_n11596_), .B(new_n11393_), .ZN(new_n11598_));
  NOR2_X1    g11341(.A1(new_n11598_), .A2(new_n11595_), .ZN(new_n11599_));
  NOR2_X1    g11342(.A1(new_n11599_), .A2(new_n11594_), .ZN(new_n11600_));
  INV_X1     g11343(.I(new_n11600_), .ZN(new_n11601_));
  AOI21_X1   g11344(.A1(new_n11405_), .A2(new_n11397_), .B(new_n11386_), .ZN(new_n11602_));
  INV_X1     g11345(.I(new_n11602_), .ZN(new_n11603_));
  OAI22_X1   g11346(.A1(new_n3298_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n3293_), .ZN(new_n11604_));
  OAI21_X1   g11347(.A1(new_n2660_), .A2(new_n3447_), .B(new_n11604_), .ZN(new_n11605_));
  AOI21_X1   g11348(.A1(new_n2963_), .A2(new_n3300_), .B(new_n11605_), .ZN(new_n11606_));
  INV_X1     g11349(.I(new_n11606_), .ZN(new_n11607_));
  NOR3_X1    g11350(.A1(new_n11370_), .A2(new_n11372_), .A3(new_n11367_), .ZN(new_n11608_));
  AOI21_X1   g11351(.A1(new_n11375_), .A2(new_n11373_), .B(new_n11608_), .ZN(new_n11609_));
  AOI21_X1   g11352(.A1(new_n11229_), .A2(new_n11371_), .B(new_n11360_), .ZN(new_n11610_));
  OAI22_X1   g11353(.A1(new_n4208_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n4203_), .ZN(new_n11611_));
  OAI21_X1   g11354(.A1(new_n1927_), .A2(new_n4362_), .B(new_n11611_), .ZN(new_n11612_));
  AOI21_X1   g11355(.A1(new_n2174_), .A2(new_n4210_), .B(new_n11612_), .ZN(new_n11613_));
  INV_X1     g11356(.I(new_n11613_), .ZN(new_n11614_));
  INV_X1     g11357(.I(new_n11230_), .ZN(new_n11615_));
  NAND3_X1   g11358(.A1(new_n11323_), .A2(new_n11327_), .A3(new_n11332_), .ZN(new_n11616_));
  AOI21_X1   g11359(.A1(new_n11615_), .A2(new_n11616_), .B(new_n11343_), .ZN(new_n11617_));
  AOI21_X1   g11360(.A1(new_n11231_), .A2(new_n11336_), .B(new_n11314_), .ZN(new_n11618_));
  AOI21_X1   g11361(.A1(new_n11304_), .A2(new_n11306_), .B(new_n11318_), .ZN(new_n11619_));
  OAI22_X1   g11362(.A1(new_n5228_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n5225_), .ZN(new_n11620_));
  NAND2_X1   g11363(.A1(new_n5387_), .A2(\b[20] ), .ZN(new_n11621_));
  AOI21_X1   g11364(.A1(new_n11620_), .A2(new_n11621_), .B(new_n5231_), .ZN(new_n11622_));
  NAND2_X1   g11365(.A1(new_n1517_), .A2(new_n11622_), .ZN(new_n11623_));
  XOR2_X1    g11366(.A1(new_n11623_), .A2(\a[50] ), .Z(new_n11624_));
  INV_X1     g11367(.I(new_n11624_), .ZN(new_n11625_));
  OAI22_X1   g11368(.A1(new_n6721_), .A2(new_n904_), .B1(new_n6723_), .B2(new_n992_), .ZN(new_n11626_));
  NAND2_X1   g11369(.A1(new_n7617_), .A2(\b[14] ), .ZN(new_n11627_));
  AOI21_X1   g11370(.A1(new_n11627_), .A2(new_n11626_), .B(new_n6731_), .ZN(new_n11628_));
  NAND2_X1   g11371(.A1(new_n991_), .A2(new_n11628_), .ZN(new_n11629_));
  XOR2_X1    g11372(.A1(new_n11629_), .A2(\a[56] ), .Z(new_n11630_));
  NOR2_X1    g11373(.A1(new_n11261_), .A2(new_n11243_), .ZN(new_n11631_));
  NOR2_X1    g11374(.A1(new_n11631_), .A2(new_n11262_), .ZN(new_n11632_));
  OAI22_X1   g11375(.A1(new_n617_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n510_), .ZN(new_n11633_));
  NAND2_X1   g11376(.A1(new_n9644_), .A2(\b[8] ), .ZN(new_n11634_));
  AOI21_X1   g11377(.A1(new_n11634_), .A2(new_n11633_), .B(new_n8321_), .ZN(new_n11635_));
  NAND2_X1   g11378(.A1(new_n616_), .A2(new_n11635_), .ZN(new_n11636_));
  XOR2_X1    g11379(.A1(new_n11636_), .A2(new_n8309_), .Z(new_n11637_));
  NOR2_X1    g11380(.A1(new_n11252_), .A2(new_n11255_), .ZN(new_n11638_));
  NOR2_X1    g11381(.A1(new_n11638_), .A2(new_n11254_), .ZN(new_n11639_));
  NOR3_X1    g11382(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n403_), .ZN(new_n11640_));
  NOR2_X1    g11383(.A1(new_n9364_), .A2(new_n403_), .ZN(new_n11641_));
  NOR3_X1    g11384(.A1(new_n11641_), .A2(new_n450_), .A3(new_n8985_), .ZN(new_n11642_));
  NOR2_X1    g11385(.A1(new_n11642_), .A2(new_n11640_), .ZN(new_n11643_));
  XOR2_X1    g11386(.A1(new_n11639_), .A2(new_n11643_), .Z(new_n11644_));
  INV_X1     g11387(.I(new_n11644_), .ZN(new_n11645_));
  INV_X1     g11388(.I(new_n11643_), .ZN(new_n11646_));
  XOR2_X1    g11389(.A1(new_n11639_), .A2(new_n11646_), .Z(new_n11647_));
  NOR2_X1    g11390(.A1(new_n11637_), .A2(new_n11647_), .ZN(new_n11648_));
  AOI21_X1   g11391(.A1(new_n11637_), .A2(new_n11645_), .B(new_n11648_), .ZN(new_n11649_));
  OAI22_X1   g11392(.A1(new_n795_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n717_), .ZN(new_n11650_));
  NAND2_X1   g11393(.A1(new_n8628_), .A2(\b[11] ), .ZN(new_n11651_));
  AOI21_X1   g11394(.A1(new_n11651_), .A2(new_n11650_), .B(new_n7354_), .ZN(new_n11652_));
  NAND2_X1   g11395(.A1(new_n799_), .A2(new_n11652_), .ZN(new_n11653_));
  XOR2_X1    g11396(.A1(new_n11653_), .A2(new_n7343_), .Z(new_n11654_));
  NAND2_X1   g11397(.A1(new_n11654_), .A2(new_n11649_), .ZN(new_n11655_));
  INV_X1     g11398(.I(new_n11649_), .ZN(new_n11656_));
  XOR2_X1    g11399(.A1(new_n11653_), .A2(\a[59] ), .Z(new_n11657_));
  NAND2_X1   g11400(.A1(new_n11657_), .A2(new_n11656_), .ZN(new_n11658_));
  AOI21_X1   g11401(.A1(new_n11655_), .A2(new_n11658_), .B(new_n11632_), .ZN(new_n11659_));
  INV_X1     g11402(.I(new_n11632_), .ZN(new_n11660_));
  NAND2_X1   g11403(.A1(new_n11654_), .A2(new_n11656_), .ZN(new_n11661_));
  NAND2_X1   g11404(.A1(new_n11657_), .A2(new_n11649_), .ZN(new_n11662_));
  AOI21_X1   g11405(.A1(new_n11661_), .A2(new_n11662_), .B(new_n11660_), .ZN(new_n11663_));
  NOR2_X1    g11406(.A1(new_n11659_), .A2(new_n11663_), .ZN(new_n11664_));
  AOI21_X1   g11407(.A1(new_n11270_), .A2(new_n11265_), .B(new_n11266_), .ZN(new_n11665_));
  NOR2_X1    g11408(.A1(new_n11664_), .A2(new_n11665_), .ZN(new_n11666_));
  INV_X1     g11409(.I(new_n11666_), .ZN(new_n11667_));
  NAND2_X1   g11410(.A1(new_n11664_), .A2(new_n11665_), .ZN(new_n11668_));
  AOI21_X1   g11411(.A1(new_n11667_), .A2(new_n11668_), .B(new_n11630_), .ZN(new_n11669_));
  INV_X1     g11412(.I(new_n11630_), .ZN(new_n11670_));
  INV_X1     g11413(.I(new_n11665_), .ZN(new_n11671_));
  NAND2_X1   g11414(.A1(new_n11664_), .A2(new_n11671_), .ZN(new_n11672_));
  OAI21_X1   g11415(.A1(new_n11659_), .A2(new_n11663_), .B(new_n11665_), .ZN(new_n11673_));
  AOI21_X1   g11416(.A1(new_n11672_), .A2(new_n11673_), .B(new_n11670_), .ZN(new_n11674_));
  NOR2_X1    g11417(.A1(new_n11669_), .A2(new_n11674_), .ZN(new_n11675_));
  AOI21_X1   g11418(.A1(new_n11233_), .A2(new_n11287_), .B(new_n11299_), .ZN(new_n11676_));
  OAI22_X1   g11419(.A1(new_n5786_), .A2(new_n1222_), .B1(new_n1124_), .B2(new_n5792_), .ZN(new_n11677_));
  NAND2_X1   g11420(.A1(new_n6745_), .A2(\b[17] ), .ZN(new_n11678_));
  AOI21_X1   g11421(.A1(new_n11678_), .A2(new_n11677_), .B(new_n5796_), .ZN(new_n11679_));
  AND3_X2    g11422(.A1(new_n1225_), .A2(new_n5783_), .A3(new_n11679_), .Z(new_n11680_));
  AOI21_X1   g11423(.A1(new_n1225_), .A2(new_n11679_), .B(new_n5783_), .ZN(new_n11681_));
  NOR2_X1    g11424(.A1(new_n11680_), .A2(new_n11681_), .ZN(new_n11682_));
  NOR2_X1    g11425(.A1(new_n11676_), .A2(new_n11682_), .ZN(new_n11683_));
  INV_X1     g11426(.I(new_n11683_), .ZN(new_n11684_));
  NAND2_X1   g11427(.A1(new_n11676_), .A2(new_n11682_), .ZN(new_n11685_));
  AOI21_X1   g11428(.A1(new_n11684_), .A2(new_n11685_), .B(new_n11675_), .ZN(new_n11686_));
  INV_X1     g11429(.I(new_n11675_), .ZN(new_n11687_));
  INV_X1     g11430(.I(new_n11682_), .ZN(new_n11688_));
  NAND2_X1   g11431(.A1(new_n11676_), .A2(new_n11688_), .ZN(new_n11689_));
  NOR2_X1    g11432(.A1(new_n11676_), .A2(new_n11688_), .ZN(new_n11690_));
  INV_X1     g11433(.I(new_n11690_), .ZN(new_n11691_));
  AOI21_X1   g11434(.A1(new_n11689_), .A2(new_n11691_), .B(new_n11687_), .ZN(new_n11692_));
  OAI21_X1   g11435(.A1(new_n11692_), .A2(new_n11686_), .B(new_n11625_), .ZN(new_n11693_));
  INV_X1     g11436(.I(new_n11685_), .ZN(new_n11694_));
  OAI21_X1   g11437(.A1(new_n11683_), .A2(new_n11694_), .B(new_n11687_), .ZN(new_n11695_));
  INV_X1     g11438(.I(new_n11689_), .ZN(new_n11696_));
  OAI21_X1   g11439(.A1(new_n11696_), .A2(new_n11690_), .B(new_n11675_), .ZN(new_n11697_));
  NAND3_X1   g11440(.A1(new_n11695_), .A2(new_n11697_), .A3(new_n11624_), .ZN(new_n11698_));
  AOI21_X1   g11441(.A1(new_n11693_), .A2(new_n11698_), .B(new_n11619_), .ZN(new_n11699_));
  INV_X1     g11442(.I(new_n11619_), .ZN(new_n11700_));
  OAI21_X1   g11443(.A1(new_n11692_), .A2(new_n11686_), .B(new_n11624_), .ZN(new_n11701_));
  NAND3_X1   g11444(.A1(new_n11695_), .A2(new_n11697_), .A3(new_n11625_), .ZN(new_n11702_));
  AOI21_X1   g11445(.A1(new_n11701_), .A2(new_n11702_), .B(new_n11700_), .ZN(new_n11703_));
  OAI22_X1   g11446(.A1(new_n4711_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n4706_), .ZN(new_n11704_));
  NAND2_X1   g11447(.A1(new_n5814_), .A2(\b[23] ), .ZN(new_n11705_));
  AOI21_X1   g11448(.A1(new_n11704_), .A2(new_n11705_), .B(new_n4714_), .ZN(new_n11706_));
  NAND3_X1   g11449(.A1(new_n1828_), .A2(new_n4701_), .A3(new_n11706_), .ZN(new_n11707_));
  INV_X1     g11450(.I(new_n11707_), .ZN(new_n11708_));
  AOI21_X1   g11451(.A1(new_n1828_), .A2(new_n11706_), .B(new_n4701_), .ZN(new_n11709_));
  NOR2_X1    g11452(.A1(new_n11708_), .A2(new_n11709_), .ZN(new_n11710_));
  INV_X1     g11453(.I(new_n11710_), .ZN(new_n11711_));
  OAI21_X1   g11454(.A1(new_n11699_), .A2(new_n11703_), .B(new_n11711_), .ZN(new_n11712_));
  AOI21_X1   g11455(.A1(new_n11695_), .A2(new_n11697_), .B(new_n11624_), .ZN(new_n11713_));
  NOR3_X1    g11456(.A1(new_n11692_), .A2(new_n11686_), .A3(new_n11625_), .ZN(new_n11714_));
  OAI21_X1   g11457(.A1(new_n11714_), .A2(new_n11713_), .B(new_n11700_), .ZN(new_n11715_));
  AOI21_X1   g11458(.A1(new_n11695_), .A2(new_n11697_), .B(new_n11625_), .ZN(new_n11716_));
  NOR3_X1    g11459(.A1(new_n11692_), .A2(new_n11686_), .A3(new_n11624_), .ZN(new_n11717_));
  OAI21_X1   g11460(.A1(new_n11717_), .A2(new_n11716_), .B(new_n11619_), .ZN(new_n11718_));
  NAND3_X1   g11461(.A1(new_n11715_), .A2(new_n11718_), .A3(new_n11710_), .ZN(new_n11719_));
  AOI21_X1   g11462(.A1(new_n11712_), .A2(new_n11719_), .B(new_n11618_), .ZN(new_n11720_));
  INV_X1     g11463(.I(new_n11618_), .ZN(new_n11721_));
  NAND3_X1   g11464(.A1(new_n11715_), .A2(new_n11718_), .A3(new_n11711_), .ZN(new_n11722_));
  OAI21_X1   g11465(.A1(new_n11699_), .A2(new_n11703_), .B(new_n11710_), .ZN(new_n11723_));
  AOI21_X1   g11466(.A1(new_n11723_), .A2(new_n11722_), .B(new_n11721_), .ZN(new_n11724_));
  OAI21_X1   g11467(.A1(new_n11720_), .A2(new_n11724_), .B(new_n11617_), .ZN(new_n11725_));
  OAI21_X1   g11468(.A1(new_n11340_), .A2(new_n11337_), .B(new_n11333_), .ZN(new_n11726_));
  OAI21_X1   g11469(.A1(new_n11230_), .A2(new_n11344_), .B(new_n11726_), .ZN(new_n11727_));
  AOI21_X1   g11470(.A1(new_n11715_), .A2(new_n11718_), .B(new_n11710_), .ZN(new_n11728_));
  NOR3_X1    g11471(.A1(new_n11699_), .A2(new_n11703_), .A3(new_n11711_), .ZN(new_n11729_));
  OAI21_X1   g11472(.A1(new_n11728_), .A2(new_n11729_), .B(new_n11721_), .ZN(new_n11730_));
  NOR3_X1    g11473(.A1(new_n11699_), .A2(new_n11703_), .A3(new_n11710_), .ZN(new_n11731_));
  AOI21_X1   g11474(.A1(new_n11715_), .A2(new_n11718_), .B(new_n11711_), .ZN(new_n11732_));
  OAI21_X1   g11475(.A1(new_n11732_), .A2(new_n11731_), .B(new_n11618_), .ZN(new_n11733_));
  NAND3_X1   g11476(.A1(new_n11730_), .A2(new_n11733_), .A3(new_n11727_), .ZN(new_n11734_));
  AOI21_X1   g11477(.A1(new_n11725_), .A2(new_n11734_), .B(\a[44] ), .ZN(new_n11735_));
  AOI21_X1   g11478(.A1(new_n11730_), .A2(new_n11733_), .B(new_n11727_), .ZN(new_n11736_));
  NOR3_X1    g11479(.A1(new_n11720_), .A2(new_n11724_), .A3(new_n11617_), .ZN(new_n11737_));
  NOR3_X1    g11480(.A1(new_n11736_), .A2(new_n11737_), .A3(new_n4198_), .ZN(new_n11738_));
  OAI21_X1   g11481(.A1(new_n11738_), .A2(new_n11735_), .B(new_n11614_), .ZN(new_n11739_));
  OAI21_X1   g11482(.A1(new_n11736_), .A2(new_n11737_), .B(new_n4198_), .ZN(new_n11740_));
  NAND3_X1   g11483(.A1(new_n11725_), .A2(new_n11734_), .A3(\a[44] ), .ZN(new_n11741_));
  NAND3_X1   g11484(.A1(new_n11740_), .A2(new_n11741_), .A3(new_n11613_), .ZN(new_n11742_));
  OAI22_X1   g11485(.A1(new_n3736_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n3731_), .ZN(new_n11743_));
  NAND2_X1   g11486(.A1(new_n4730_), .A2(\b[29] ), .ZN(new_n11744_));
  AOI21_X1   g11487(.A1(new_n11743_), .A2(new_n11744_), .B(new_n3739_), .ZN(new_n11745_));
  NAND2_X1   g11488(.A1(new_n2546_), .A2(new_n11745_), .ZN(new_n11746_));
  XOR2_X1    g11489(.A1(new_n11746_), .A2(\a[41] ), .Z(new_n11747_));
  INV_X1     g11490(.I(new_n11747_), .ZN(new_n11748_));
  NAND3_X1   g11491(.A1(new_n11739_), .A2(new_n11742_), .A3(new_n11748_), .ZN(new_n11749_));
  AOI21_X1   g11492(.A1(new_n11740_), .A2(new_n11741_), .B(new_n11613_), .ZN(new_n11750_));
  NOR3_X1    g11493(.A1(new_n11738_), .A2(new_n11735_), .A3(new_n11614_), .ZN(new_n11751_));
  OAI21_X1   g11494(.A1(new_n11751_), .A2(new_n11750_), .B(new_n11747_), .ZN(new_n11752_));
  AOI21_X1   g11495(.A1(new_n11752_), .A2(new_n11749_), .B(new_n11610_), .ZN(new_n11753_));
  INV_X1     g11496(.I(new_n11610_), .ZN(new_n11754_));
  OAI21_X1   g11497(.A1(new_n11751_), .A2(new_n11750_), .B(new_n11748_), .ZN(new_n11755_));
  NAND3_X1   g11498(.A1(new_n11739_), .A2(new_n11742_), .A3(new_n11747_), .ZN(new_n11756_));
  AOI21_X1   g11499(.A1(new_n11755_), .A2(new_n11756_), .B(new_n11754_), .ZN(new_n11757_));
  OAI21_X1   g11500(.A1(new_n11753_), .A2(new_n11757_), .B(new_n11609_), .ZN(new_n11758_));
  AOI21_X1   g11501(.A1(new_n11362_), .A2(new_n11357_), .B(new_n11368_), .ZN(new_n11759_));
  OAI21_X1   g11502(.A1(new_n11223_), .A2(new_n11759_), .B(new_n11369_), .ZN(new_n11760_));
  NOR3_X1    g11503(.A1(new_n11751_), .A2(new_n11750_), .A3(new_n11747_), .ZN(new_n11761_));
  AOI21_X1   g11504(.A1(new_n11739_), .A2(new_n11742_), .B(new_n11748_), .ZN(new_n11762_));
  OAI21_X1   g11505(.A1(new_n11761_), .A2(new_n11762_), .B(new_n11754_), .ZN(new_n11763_));
  AOI21_X1   g11506(.A1(new_n11739_), .A2(new_n11742_), .B(new_n11747_), .ZN(new_n11764_));
  NOR3_X1    g11507(.A1(new_n11751_), .A2(new_n11750_), .A3(new_n11748_), .ZN(new_n11765_));
  OAI21_X1   g11508(.A1(new_n11765_), .A2(new_n11764_), .B(new_n11610_), .ZN(new_n11766_));
  NAND3_X1   g11509(.A1(new_n11763_), .A2(new_n11766_), .A3(new_n11760_), .ZN(new_n11767_));
  AOI21_X1   g11510(.A1(new_n11758_), .A2(new_n11767_), .B(\a[38] ), .ZN(new_n11768_));
  AOI21_X1   g11511(.A1(new_n11763_), .A2(new_n11766_), .B(new_n11760_), .ZN(new_n11769_));
  NOR3_X1    g11512(.A1(new_n11753_), .A2(new_n11757_), .A3(new_n11609_), .ZN(new_n11770_));
  NOR3_X1    g11513(.A1(new_n11769_), .A2(new_n11770_), .A3(new_n3288_), .ZN(new_n11771_));
  OAI21_X1   g11514(.A1(new_n11768_), .A2(new_n11771_), .B(new_n11607_), .ZN(new_n11772_));
  OAI21_X1   g11515(.A1(new_n11769_), .A2(new_n11770_), .B(new_n3288_), .ZN(new_n11773_));
  NAND3_X1   g11516(.A1(new_n11758_), .A2(new_n11767_), .A3(\a[38] ), .ZN(new_n11774_));
  NAND3_X1   g11517(.A1(new_n11773_), .A2(new_n11774_), .A3(new_n11606_), .ZN(new_n11775_));
  OAI22_X1   g11518(.A1(new_n2846_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n2841_), .ZN(new_n11776_));
  NAND2_X1   g11519(.A1(new_n3755_), .A2(\b[35] ), .ZN(new_n11777_));
  AOI21_X1   g11520(.A1(new_n11776_), .A2(new_n11777_), .B(new_n2849_), .ZN(new_n11778_));
  NAND2_X1   g11521(.A1(new_n3411_), .A2(new_n11778_), .ZN(new_n11779_));
  XOR2_X1    g11522(.A1(new_n11779_), .A2(\a[35] ), .Z(new_n11780_));
  INV_X1     g11523(.I(new_n11780_), .ZN(new_n11781_));
  NAND3_X1   g11524(.A1(new_n11772_), .A2(new_n11775_), .A3(new_n11781_), .ZN(new_n11782_));
  INV_X1     g11525(.I(new_n11782_), .ZN(new_n11783_));
  AOI21_X1   g11526(.A1(new_n11772_), .A2(new_n11775_), .B(new_n11781_), .ZN(new_n11784_));
  OAI21_X1   g11527(.A1(new_n11783_), .A2(new_n11784_), .B(new_n11603_), .ZN(new_n11785_));
  AOI21_X1   g11528(.A1(new_n11772_), .A2(new_n11775_), .B(new_n11780_), .ZN(new_n11786_));
  AOI21_X1   g11529(.A1(new_n11773_), .A2(new_n11774_), .B(new_n11606_), .ZN(new_n11787_));
  NOR3_X1    g11530(.A1(new_n11768_), .A2(new_n11771_), .A3(new_n11607_), .ZN(new_n11788_));
  NOR3_X1    g11531(.A1(new_n11788_), .A2(new_n11787_), .A3(new_n11781_), .ZN(new_n11789_));
  OAI21_X1   g11532(.A1(new_n11789_), .A2(new_n11786_), .B(new_n11602_), .ZN(new_n11790_));
  OAI22_X1   g11533(.A1(new_n2452_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n2447_), .ZN(new_n11791_));
  NAND2_X1   g11534(.A1(new_n3312_), .A2(\b[38] ), .ZN(new_n11792_));
  AOI21_X1   g11535(.A1(new_n11791_), .A2(new_n11792_), .B(new_n2455_), .ZN(new_n11793_));
  NAND2_X1   g11536(.A1(new_n3844_), .A2(new_n11793_), .ZN(new_n11794_));
  XOR2_X1    g11537(.A1(new_n11794_), .A2(\a[32] ), .Z(new_n11795_));
  AOI21_X1   g11538(.A1(new_n11785_), .A2(new_n11790_), .B(new_n11795_), .ZN(new_n11796_));
  OAI21_X1   g11539(.A1(new_n11788_), .A2(new_n11787_), .B(new_n11780_), .ZN(new_n11797_));
  AOI21_X1   g11540(.A1(new_n11797_), .A2(new_n11782_), .B(new_n11602_), .ZN(new_n11798_));
  OAI21_X1   g11541(.A1(new_n11788_), .A2(new_n11787_), .B(new_n11781_), .ZN(new_n11799_));
  NAND3_X1   g11542(.A1(new_n11772_), .A2(new_n11775_), .A3(new_n11780_), .ZN(new_n11800_));
  AOI21_X1   g11543(.A1(new_n11799_), .A2(new_n11800_), .B(new_n11603_), .ZN(new_n11801_));
  INV_X1     g11544(.I(new_n11795_), .ZN(new_n11802_));
  NOR3_X1    g11545(.A1(new_n11798_), .A2(new_n11801_), .A3(new_n11802_), .ZN(new_n11803_));
  OAI21_X1   g11546(.A1(new_n11796_), .A2(new_n11803_), .B(new_n11601_), .ZN(new_n11804_));
  NOR3_X1    g11547(.A1(new_n11798_), .A2(new_n11801_), .A3(new_n11795_), .ZN(new_n11805_));
  AOI21_X1   g11548(.A1(new_n11785_), .A2(new_n11790_), .B(new_n11802_), .ZN(new_n11806_));
  OAI21_X1   g11549(.A1(new_n11806_), .A2(new_n11805_), .B(new_n11600_), .ZN(new_n11807_));
  OAI22_X1   g11550(.A1(new_n2084_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n2079_), .ZN(new_n11808_));
  NAND2_X1   g11551(.A1(new_n2864_), .A2(\b[41] ), .ZN(new_n11809_));
  AOI21_X1   g11552(.A1(new_n11808_), .A2(new_n11809_), .B(new_n2087_), .ZN(new_n11810_));
  NAND2_X1   g11553(.A1(new_n4320_), .A2(new_n11810_), .ZN(new_n11811_));
  XOR2_X1    g11554(.A1(new_n11811_), .A2(\a[29] ), .Z(new_n11812_));
  AOI21_X1   g11555(.A1(new_n11804_), .A2(new_n11807_), .B(new_n11812_), .ZN(new_n11813_));
  OAI21_X1   g11556(.A1(new_n11798_), .A2(new_n11801_), .B(new_n11802_), .ZN(new_n11814_));
  NAND3_X1   g11557(.A1(new_n11785_), .A2(new_n11790_), .A3(new_n11795_), .ZN(new_n11815_));
  AOI21_X1   g11558(.A1(new_n11815_), .A2(new_n11814_), .B(new_n11600_), .ZN(new_n11816_));
  NAND3_X1   g11559(.A1(new_n11785_), .A2(new_n11790_), .A3(new_n11802_), .ZN(new_n11817_));
  OAI21_X1   g11560(.A1(new_n11798_), .A2(new_n11801_), .B(new_n11795_), .ZN(new_n11818_));
  AOI21_X1   g11561(.A1(new_n11817_), .A2(new_n11818_), .B(new_n11601_), .ZN(new_n11819_));
  INV_X1     g11562(.I(new_n11812_), .ZN(new_n11820_));
  NOR3_X1    g11563(.A1(new_n11819_), .A2(new_n11816_), .A3(new_n11820_), .ZN(new_n11821_));
  OAI21_X1   g11564(.A1(new_n11813_), .A2(new_n11821_), .B(new_n11593_), .ZN(new_n11822_));
  AOI21_X1   g11565(.A1(new_n11222_), .A2(new_n11434_), .B(new_n11421_), .ZN(new_n11823_));
  NOR3_X1    g11566(.A1(new_n11819_), .A2(new_n11816_), .A3(new_n11812_), .ZN(new_n11824_));
  AOI21_X1   g11567(.A1(new_n11807_), .A2(new_n11804_), .B(new_n11820_), .ZN(new_n11825_));
  OAI21_X1   g11568(.A1(new_n11825_), .A2(new_n11824_), .B(new_n11823_), .ZN(new_n11826_));
  OAI22_X1   g11569(.A1(new_n1760_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n1755_), .ZN(new_n11827_));
  NAND2_X1   g11570(.A1(new_n2470_), .A2(\b[44] ), .ZN(new_n11828_));
  AOI21_X1   g11571(.A1(new_n11827_), .A2(new_n11828_), .B(new_n1763_), .ZN(new_n11829_));
  NAND2_X1   g11572(.A1(new_n4833_), .A2(new_n11829_), .ZN(new_n11830_));
  XOR2_X1    g11573(.A1(new_n11830_), .A2(\a[26] ), .Z(new_n11831_));
  AOI21_X1   g11574(.A1(new_n11826_), .A2(new_n11822_), .B(new_n11831_), .ZN(new_n11832_));
  OAI21_X1   g11575(.A1(new_n11819_), .A2(new_n11816_), .B(new_n11820_), .ZN(new_n11833_));
  NAND3_X1   g11576(.A1(new_n11804_), .A2(new_n11807_), .A3(new_n11812_), .ZN(new_n11834_));
  AOI21_X1   g11577(.A1(new_n11833_), .A2(new_n11834_), .B(new_n11823_), .ZN(new_n11835_));
  NAND3_X1   g11578(.A1(new_n11807_), .A2(new_n11804_), .A3(new_n11820_), .ZN(new_n11836_));
  OAI21_X1   g11579(.A1(new_n11819_), .A2(new_n11816_), .B(new_n11812_), .ZN(new_n11837_));
  AOI21_X1   g11580(.A1(new_n11837_), .A2(new_n11836_), .B(new_n11593_), .ZN(new_n11838_));
  INV_X1     g11581(.I(new_n11831_), .ZN(new_n11839_));
  NOR3_X1    g11582(.A1(new_n11835_), .A2(new_n11838_), .A3(new_n11839_), .ZN(new_n11840_));
  OAI21_X1   g11583(.A1(new_n11832_), .A2(new_n11840_), .B(new_n11592_), .ZN(new_n11841_));
  AOI21_X1   g11584(.A1(new_n11220_), .A2(new_n11455_), .B(new_n11439_), .ZN(new_n11842_));
  NOR3_X1    g11585(.A1(new_n11835_), .A2(new_n11838_), .A3(new_n11831_), .ZN(new_n11843_));
  AOI21_X1   g11586(.A1(new_n11826_), .A2(new_n11822_), .B(new_n11839_), .ZN(new_n11844_));
  OAI21_X1   g11587(.A1(new_n11844_), .A2(new_n11843_), .B(new_n11842_), .ZN(new_n11845_));
  OAI22_X1   g11588(.A1(new_n1444_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n1439_), .ZN(new_n11846_));
  NAND2_X1   g11589(.A1(new_n2098_), .A2(\b[47] ), .ZN(new_n11847_));
  AOI21_X1   g11590(.A1(new_n11846_), .A2(new_n11847_), .B(new_n1447_), .ZN(new_n11848_));
  NAND2_X1   g11591(.A1(new_n5196_), .A2(new_n11848_), .ZN(new_n11849_));
  XOR2_X1    g11592(.A1(new_n11849_), .A2(\a[23] ), .Z(new_n11850_));
  AOI21_X1   g11593(.A1(new_n11841_), .A2(new_n11845_), .B(new_n11850_), .ZN(new_n11851_));
  OAI21_X1   g11594(.A1(new_n11835_), .A2(new_n11838_), .B(new_n11839_), .ZN(new_n11852_));
  NAND3_X1   g11595(.A1(new_n11826_), .A2(new_n11822_), .A3(new_n11831_), .ZN(new_n11853_));
  AOI21_X1   g11596(.A1(new_n11852_), .A2(new_n11853_), .B(new_n11842_), .ZN(new_n11854_));
  NAND3_X1   g11597(.A1(new_n11826_), .A2(new_n11822_), .A3(new_n11839_), .ZN(new_n11855_));
  OAI21_X1   g11598(.A1(new_n11835_), .A2(new_n11838_), .B(new_n11831_), .ZN(new_n11856_));
  AOI21_X1   g11599(.A1(new_n11856_), .A2(new_n11855_), .B(new_n11592_), .ZN(new_n11857_));
  INV_X1     g11600(.I(new_n11850_), .ZN(new_n11858_));
  NOR3_X1    g11601(.A1(new_n11854_), .A2(new_n11857_), .A3(new_n11858_), .ZN(new_n11859_));
  OAI21_X1   g11602(.A1(new_n11851_), .A2(new_n11859_), .B(new_n11591_), .ZN(new_n11860_));
  AOI21_X1   g11603(.A1(new_n11459_), .A2(new_n11457_), .B(new_n11470_), .ZN(new_n11861_));
  NOR3_X1    g11604(.A1(new_n11854_), .A2(new_n11857_), .A3(new_n11850_), .ZN(new_n11862_));
  AOI21_X1   g11605(.A1(new_n11841_), .A2(new_n11845_), .B(new_n11858_), .ZN(new_n11863_));
  OAI21_X1   g11606(.A1(new_n11863_), .A2(new_n11862_), .B(new_n11861_), .ZN(new_n11864_));
  OAI22_X1   g11607(.A1(new_n1168_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n1163_), .ZN(new_n11865_));
  NAND2_X1   g11608(.A1(new_n1774_), .A2(\b[50] ), .ZN(new_n11866_));
  AOI21_X1   g11609(.A1(new_n11865_), .A2(new_n11866_), .B(new_n1171_), .ZN(new_n11867_));
  NAND2_X1   g11610(.A1(new_n5954_), .A2(new_n11867_), .ZN(new_n11868_));
  XOR2_X1    g11611(.A1(new_n11868_), .A2(\a[20] ), .Z(new_n11869_));
  AOI21_X1   g11612(.A1(new_n11860_), .A2(new_n11864_), .B(new_n11869_), .ZN(new_n11870_));
  OAI21_X1   g11613(.A1(new_n11854_), .A2(new_n11857_), .B(new_n11858_), .ZN(new_n11871_));
  NAND3_X1   g11614(.A1(new_n11841_), .A2(new_n11845_), .A3(new_n11850_), .ZN(new_n11872_));
  AOI21_X1   g11615(.A1(new_n11871_), .A2(new_n11872_), .B(new_n11861_), .ZN(new_n11873_));
  NAND3_X1   g11616(.A1(new_n11841_), .A2(new_n11845_), .A3(new_n11858_), .ZN(new_n11874_));
  OAI21_X1   g11617(.A1(new_n11854_), .A2(new_n11857_), .B(new_n11850_), .ZN(new_n11875_));
  AOI21_X1   g11618(.A1(new_n11875_), .A2(new_n11874_), .B(new_n11591_), .ZN(new_n11876_));
  INV_X1     g11619(.I(new_n11869_), .ZN(new_n11877_));
  NOR3_X1    g11620(.A1(new_n11873_), .A2(new_n11876_), .A3(new_n11877_), .ZN(new_n11878_));
  OAI21_X1   g11621(.A1(new_n11870_), .A2(new_n11878_), .B(new_n11590_), .ZN(new_n11879_));
  AOI21_X1   g11622(.A1(new_n11478_), .A2(new_n11476_), .B(new_n11489_), .ZN(new_n11880_));
  NOR3_X1    g11623(.A1(new_n11873_), .A2(new_n11876_), .A3(new_n11869_), .ZN(new_n11881_));
  AOI21_X1   g11624(.A1(new_n11860_), .A2(new_n11864_), .B(new_n11877_), .ZN(new_n11882_));
  OAI21_X1   g11625(.A1(new_n11882_), .A2(new_n11881_), .B(new_n11880_), .ZN(new_n11883_));
  OAI22_X1   g11626(.A1(new_n940_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n935_), .ZN(new_n11884_));
  NAND2_X1   g11627(.A1(new_n1458_), .A2(\b[53] ), .ZN(new_n11885_));
  AOI21_X1   g11628(.A1(new_n11884_), .A2(new_n11885_), .B(new_n943_), .ZN(new_n11886_));
  NAND2_X1   g11629(.A1(new_n6471_), .A2(new_n11886_), .ZN(new_n11887_));
  XOR2_X1    g11630(.A1(new_n11887_), .A2(\a[17] ), .Z(new_n11888_));
  INV_X1     g11631(.I(new_n11888_), .ZN(new_n11889_));
  NAND3_X1   g11632(.A1(new_n11879_), .A2(new_n11883_), .A3(new_n11889_), .ZN(new_n11890_));
  OAI21_X1   g11633(.A1(new_n11873_), .A2(new_n11876_), .B(new_n11877_), .ZN(new_n11891_));
  NAND3_X1   g11634(.A1(new_n11860_), .A2(new_n11864_), .A3(new_n11869_), .ZN(new_n11892_));
  AOI21_X1   g11635(.A1(new_n11891_), .A2(new_n11892_), .B(new_n11880_), .ZN(new_n11893_));
  NAND3_X1   g11636(.A1(new_n11860_), .A2(new_n11864_), .A3(new_n11877_), .ZN(new_n11894_));
  OAI21_X1   g11637(.A1(new_n11873_), .A2(new_n11876_), .B(new_n11869_), .ZN(new_n11895_));
  AOI21_X1   g11638(.A1(new_n11895_), .A2(new_n11894_), .B(new_n11590_), .ZN(new_n11896_));
  OAI21_X1   g11639(.A1(new_n11893_), .A2(new_n11896_), .B(new_n11888_), .ZN(new_n11897_));
  AOI22_X1   g11640(.A1(new_n11897_), .A2(new_n11890_), .B1(new_n11589_), .B2(new_n11488_), .ZN(new_n11898_));
  NAND2_X1   g11641(.A1(new_n11589_), .A2(new_n11488_), .ZN(new_n11899_));
  OAI21_X1   g11642(.A1(new_n11893_), .A2(new_n11896_), .B(new_n11889_), .ZN(new_n11900_));
  NAND3_X1   g11643(.A1(new_n11879_), .A2(new_n11883_), .A3(new_n11888_), .ZN(new_n11901_));
  AOI21_X1   g11644(.A1(new_n11900_), .A2(new_n11901_), .B(new_n11899_), .ZN(new_n11902_));
  NOR2_X1    g11645(.A1(new_n11902_), .A2(new_n11898_), .ZN(new_n11903_));
  OAI22_X1   g11646(.A1(new_n757_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n752_), .ZN(new_n11904_));
  NAND2_X1   g11647(.A1(new_n1182_), .A2(\b[56] ), .ZN(new_n11905_));
  AOI21_X1   g11648(.A1(new_n11904_), .A2(new_n11905_), .B(new_n760_), .ZN(new_n11906_));
  NAND2_X1   g11649(.A1(new_n7559_), .A2(new_n11906_), .ZN(new_n11907_));
  XOR2_X1    g11650(.A1(new_n11907_), .A2(\a[14] ), .Z(new_n11908_));
  INV_X1     g11651(.I(new_n11908_), .ZN(new_n11909_));
  NAND2_X1   g11652(.A1(new_n11903_), .A2(new_n11909_), .ZN(new_n11910_));
  NAND2_X1   g11653(.A1(new_n11897_), .A2(new_n11890_), .ZN(new_n11911_));
  NAND2_X1   g11654(.A1(new_n11900_), .A2(new_n11901_), .ZN(new_n11912_));
  MUX2_X1    g11655(.I0(new_n11912_), .I1(new_n11911_), .S(new_n11899_), .Z(new_n11913_));
  NAND2_X1   g11656(.A1(new_n11913_), .A2(new_n11908_), .ZN(new_n11914_));
  NAND2_X1   g11657(.A1(new_n11914_), .A2(new_n11910_), .ZN(new_n11915_));
  NAND2_X1   g11658(.A1(new_n11915_), .A2(new_n11588_), .ZN(new_n11916_));
  AND2_X2    g11659(.A1(new_n11587_), .A2(new_n11505_), .Z(new_n11917_));
  NOR2_X1    g11660(.A1(new_n11903_), .A2(new_n11908_), .ZN(new_n11918_));
  NAND2_X1   g11661(.A1(new_n11903_), .A2(new_n11908_), .ZN(new_n11919_));
  INV_X1     g11662(.I(new_n11919_), .ZN(new_n11920_));
  OAI21_X1   g11663(.A1(new_n11920_), .A2(new_n11918_), .B(new_n11917_), .ZN(new_n11921_));
  OAI22_X1   g11664(.A1(new_n582_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n577_), .ZN(new_n11922_));
  NAND2_X1   g11665(.A1(new_n960_), .A2(\b[59] ), .ZN(new_n11923_));
  AOI21_X1   g11666(.A1(new_n11922_), .A2(new_n11923_), .B(new_n585_), .ZN(new_n11924_));
  NAND2_X1   g11667(.A1(new_n8550_), .A2(new_n11924_), .ZN(new_n11925_));
  NOR2_X1    g11668(.A1(new_n11925_), .A2(\a[11] ), .ZN(new_n11926_));
  NAND2_X1   g11669(.A1(new_n11925_), .A2(\a[11] ), .ZN(new_n11927_));
  INV_X1     g11670(.I(new_n11927_), .ZN(new_n11928_));
  NOR2_X1    g11671(.A1(new_n11928_), .A2(new_n11926_), .ZN(new_n11929_));
  INV_X1     g11672(.I(new_n11929_), .ZN(new_n11930_));
  NAND3_X1   g11673(.A1(new_n11916_), .A2(new_n11921_), .A3(new_n11930_), .ZN(new_n11931_));
  AOI21_X1   g11674(.A1(new_n11914_), .A2(new_n11910_), .B(new_n11917_), .ZN(new_n11932_));
  NAND2_X1   g11675(.A1(new_n11913_), .A2(new_n11909_), .ZN(new_n11933_));
  AOI21_X1   g11676(.A1(new_n11933_), .A2(new_n11919_), .B(new_n11588_), .ZN(new_n11934_));
  OAI21_X1   g11677(.A1(new_n11932_), .A2(new_n11934_), .B(new_n11929_), .ZN(new_n11935_));
  AOI21_X1   g11678(.A1(new_n11931_), .A2(new_n11935_), .B(new_n11586_), .ZN(new_n11936_));
  INV_X1     g11679(.I(new_n11936_), .ZN(new_n11937_));
  AOI21_X1   g11680(.A1(new_n11916_), .A2(new_n11921_), .B(new_n11929_), .ZN(new_n11938_));
  NOR3_X1    g11681(.A1(new_n11932_), .A2(new_n11930_), .A3(new_n11934_), .ZN(new_n11939_));
  OAI21_X1   g11682(.A1(new_n11938_), .A2(new_n11939_), .B(new_n11586_), .ZN(new_n11940_));
  NOR2_X1    g11683(.A1(new_n474_), .A2(new_n8932_), .ZN(new_n11941_));
  NOR2_X1    g11684(.A1(new_n431_), .A2(new_n8956_), .ZN(new_n11942_));
  NOR4_X1    g11685(.A1(new_n9323_), .A2(new_n440_), .A3(new_n11941_), .A4(new_n11942_), .ZN(new_n11943_));
  XOR2_X1    g11686(.A1(new_n11943_), .A2(new_n429_), .Z(new_n11944_));
  INV_X1     g11687(.I(new_n11944_), .ZN(new_n11945_));
  NAND3_X1   g11688(.A1(new_n11937_), .A2(new_n11940_), .A3(new_n11945_), .ZN(new_n11946_));
  INV_X1     g11689(.I(new_n11940_), .ZN(new_n11947_));
  OAI21_X1   g11690(.A1(new_n11947_), .A2(new_n11936_), .B(new_n11944_), .ZN(new_n11948_));
  AOI21_X1   g11691(.A1(new_n11948_), .A2(new_n11946_), .B(new_n11585_), .ZN(new_n11949_));
  INV_X1     g11692(.I(new_n11585_), .ZN(new_n11950_));
  OAI21_X1   g11693(.A1(new_n11947_), .A2(new_n11936_), .B(new_n11945_), .ZN(new_n11951_));
  NAND3_X1   g11694(.A1(new_n11937_), .A2(new_n11940_), .A3(new_n11944_), .ZN(new_n11952_));
  AOI21_X1   g11695(.A1(new_n11951_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n11953_));
  NOR2_X1    g11696(.A1(new_n11953_), .A2(new_n11949_), .ZN(new_n11954_));
  INV_X1     g11697(.I(new_n11556_), .ZN(new_n11955_));
  OR2_X2     g11698(.A1(new_n11564_), .A2(new_n11566_), .Z(new_n11956_));
  NAND2_X1   g11699(.A1(new_n11956_), .A2(new_n11955_), .ZN(new_n11957_));
  XNOR2_X1   g11700(.A1(new_n11954_), .A2(new_n11957_), .ZN(new_n11958_));
  NAND3_X1   g11701(.A1(new_n10805_), .A2(new_n11576_), .A3(new_n11579_), .ZN(new_n11959_));
  NAND2_X1   g11702(.A1(new_n10812_), .A2(new_n10813_), .ZN(new_n11960_));
  AOI21_X1   g11703(.A1(new_n11960_), .A2(new_n11959_), .B(new_n11201_), .ZN(new_n11961_));
  XOR2_X1    g11704(.A1(new_n11570_), .A2(new_n11209_), .Z(new_n11962_));
  NAND3_X1   g11705(.A1(new_n11962_), .A2(new_n10812_), .A3(new_n11579_), .ZN(new_n11963_));
  AND2_X2    g11706(.A1(new_n11565_), .A2(new_n11569_), .Z(new_n11964_));
  NAND2_X1   g11707(.A1(new_n11964_), .A2(new_n11209_), .ZN(new_n11965_));
  INV_X1     g11708(.I(new_n11965_), .ZN(new_n11966_));
  AOI21_X1   g11709(.A1(new_n11961_), .A2(new_n11963_), .B(new_n11966_), .ZN(new_n11967_));
  NAND2_X1   g11710(.A1(new_n11961_), .A2(new_n11963_), .ZN(new_n11968_));
  NAND3_X1   g11711(.A1(new_n11968_), .A2(new_n11958_), .A3(new_n11965_), .ZN(new_n11969_));
  OAI21_X1   g11712(.A1(new_n11967_), .A2(new_n11958_), .B(new_n11969_), .ZN(\f[70] ));
  NOR2_X1    g11713(.A1(new_n11954_), .A2(new_n11957_), .ZN(new_n11971_));
  NAND2_X1   g11714(.A1(new_n11954_), .A2(new_n11957_), .ZN(new_n11972_));
  INV_X1     g11715(.I(new_n11972_), .ZN(new_n11973_));
  NOR2_X1    g11716(.A1(new_n11954_), .A2(new_n11957_), .ZN(new_n11974_));
  OAI21_X1   g11717(.A1(new_n11973_), .A2(new_n11974_), .B(new_n11965_), .ZN(new_n11975_));
  AOI21_X1   g11718(.A1(new_n11961_), .A2(new_n11963_), .B(new_n11975_), .ZN(new_n11976_));
  NOR2_X1    g11719(.A1(new_n11976_), .A2(new_n11971_), .ZN(new_n11977_));
  NAND2_X1   g11720(.A1(new_n11948_), .A2(new_n11950_), .ZN(new_n11978_));
  NAND2_X1   g11721(.A1(new_n11978_), .A2(new_n11946_), .ZN(new_n11979_));
  INV_X1     g11722(.I(new_n11979_), .ZN(new_n11980_));
  AOI22_X1   g11723(.A1(new_n10814_), .A2(new_n439_), .B1(\b[63] ), .B2(new_n775_), .ZN(new_n11981_));
  INV_X1     g11724(.I(new_n11981_), .ZN(new_n11982_));
  NOR2_X1    g11725(.A1(new_n11939_), .A2(new_n11586_), .ZN(new_n11983_));
  NOR2_X1    g11726(.A1(new_n11983_), .A2(new_n11938_), .ZN(new_n11984_));
  NAND2_X1   g11727(.A1(new_n11899_), .A2(new_n11901_), .ZN(new_n11985_));
  NAND2_X1   g11728(.A1(new_n11985_), .A2(new_n11900_), .ZN(new_n11986_));
  AOI21_X1   g11729(.A1(new_n11590_), .A2(new_n11892_), .B(new_n11870_), .ZN(new_n11987_));
  AOI21_X1   g11730(.A1(new_n11591_), .A2(new_n11872_), .B(new_n11851_), .ZN(new_n11988_));
  AOI21_X1   g11731(.A1(new_n11592_), .A2(new_n11853_), .B(new_n11832_), .ZN(new_n11989_));
  INV_X1     g11732(.I(new_n11989_), .ZN(new_n11990_));
  AOI21_X1   g11733(.A1(new_n11593_), .A2(new_n11834_), .B(new_n11813_), .ZN(new_n11991_));
  NOR2_X1    g11734(.A1(new_n11803_), .A2(new_n11600_), .ZN(new_n11992_));
  NOR2_X1    g11735(.A1(new_n11992_), .A2(new_n11796_), .ZN(new_n11993_));
  AOI21_X1   g11736(.A1(new_n11603_), .A2(new_n11797_), .B(new_n11783_), .ZN(new_n11994_));
  OAI22_X1   g11737(.A1(new_n2846_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n2841_), .ZN(new_n11995_));
  OAI21_X1   g11738(.A1(new_n3247_), .A2(new_n3015_), .B(new_n11995_), .ZN(new_n11996_));
  AOI21_X1   g11739(.A1(new_n3565_), .A2(new_n2848_), .B(new_n11996_), .ZN(new_n11997_));
  INV_X1     g11740(.I(new_n11997_), .ZN(new_n11998_));
  NOR2_X1    g11741(.A1(new_n11753_), .A2(new_n11757_), .ZN(new_n11999_));
  XOR2_X1    g11742(.A1(new_n11606_), .A2(new_n3288_), .Z(new_n12000_));
  INV_X1     g11743(.I(new_n12000_), .ZN(new_n12001_));
  XOR2_X1    g11744(.A1(new_n11760_), .A2(new_n12001_), .Z(new_n12002_));
  OAI21_X1   g11745(.A1(new_n11999_), .A2(new_n12000_), .B(new_n12002_), .ZN(new_n12003_));
  AOI21_X1   g11746(.A1(new_n11754_), .A2(new_n11756_), .B(new_n11764_), .ZN(new_n12004_));
  INV_X1     g11747(.I(new_n12004_), .ZN(new_n12005_));
  NAND2_X1   g11748(.A1(new_n11730_), .A2(new_n11733_), .ZN(new_n12006_));
  NAND2_X1   g11749(.A1(new_n12006_), .A2(new_n11727_), .ZN(new_n12007_));
  NOR2_X1    g11750(.A1(new_n12006_), .A2(new_n11727_), .ZN(new_n12008_));
  XOR2_X1    g11751(.A1(new_n11613_), .A2(new_n4198_), .Z(new_n12009_));
  OAI21_X1   g11752(.A1(new_n12008_), .A2(new_n12009_), .B(new_n12007_), .ZN(new_n12010_));
  INV_X1     g11753(.I(new_n12010_), .ZN(new_n12011_));
  AOI21_X1   g11754(.A1(new_n11721_), .A2(new_n11719_), .B(new_n11728_), .ZN(new_n12012_));
  INV_X1     g11755(.I(new_n12012_), .ZN(new_n12013_));
  AOI21_X1   g11756(.A1(new_n11700_), .A2(new_n11698_), .B(new_n11713_), .ZN(new_n12014_));
  INV_X1     g11757(.I(new_n12014_), .ZN(new_n12015_));
  OAI22_X1   g11758(.A1(new_n4711_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n4706_), .ZN(new_n12016_));
  NAND2_X1   g11759(.A1(new_n5814_), .A2(\b[24] ), .ZN(new_n12017_));
  AOI21_X1   g11760(.A1(new_n12016_), .A2(new_n12017_), .B(new_n4714_), .ZN(new_n12018_));
  NAND2_X1   g11761(.A1(new_n1926_), .A2(new_n12018_), .ZN(new_n12019_));
  XOR2_X1    g11762(.A1(new_n12019_), .A2(\a[47] ), .Z(new_n12020_));
  INV_X1     g11763(.I(new_n12020_), .ZN(new_n12021_));
  OAI22_X1   g11764(.A1(new_n5228_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n5225_), .ZN(new_n12022_));
  NAND2_X1   g11765(.A1(new_n5387_), .A2(\b[21] ), .ZN(new_n12023_));
  AOI21_X1   g11766(.A1(new_n12022_), .A2(new_n12023_), .B(new_n5231_), .ZN(new_n12024_));
  NAND2_X1   g11767(.A1(new_n1604_), .A2(new_n12024_), .ZN(new_n12025_));
  XOR2_X1    g11768(.A1(new_n12025_), .A2(\a[50] ), .Z(new_n12026_));
  INV_X1     g11769(.I(new_n12026_), .ZN(new_n12027_));
  OAI22_X1   g11770(.A1(new_n5786_), .A2(new_n1305_), .B1(new_n1222_), .B2(new_n5792_), .ZN(new_n12028_));
  NAND2_X1   g11771(.A1(new_n6745_), .A2(\b[18] ), .ZN(new_n12029_));
  AOI21_X1   g11772(.A1(new_n12029_), .A2(new_n12028_), .B(new_n5796_), .ZN(new_n12030_));
  NAND2_X1   g11773(.A1(new_n1304_), .A2(new_n12030_), .ZN(new_n12031_));
  XOR2_X1    g11774(.A1(new_n12031_), .A2(\a[53] ), .Z(new_n12032_));
  INV_X1     g11775(.I(new_n11639_), .ZN(new_n12033_));
  OAI21_X1   g11776(.A1(new_n12033_), .A2(new_n11643_), .B(new_n11637_), .ZN(new_n12034_));
  OAI21_X1   g11777(.A1(new_n11639_), .A2(new_n11646_), .B(new_n12034_), .ZN(new_n12035_));
  NOR3_X1    g11778(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n450_), .ZN(new_n12036_));
  NOR2_X1    g11779(.A1(new_n9364_), .A2(new_n450_), .ZN(new_n12037_));
  NOR3_X1    g11780(.A1(new_n12037_), .A2(new_n495_), .A3(new_n8985_), .ZN(new_n12038_));
  NOR2_X1    g11781(.A1(new_n12038_), .A2(new_n12036_), .ZN(new_n12039_));
  NOR2_X1    g11782(.A1(new_n11646_), .A2(new_n12039_), .ZN(new_n12040_));
  INV_X1     g11783(.I(new_n12039_), .ZN(new_n12041_));
  NOR2_X1    g11784(.A1(new_n12041_), .A2(new_n11643_), .ZN(new_n12042_));
  OAI21_X1   g11785(.A1(new_n12040_), .A2(new_n12042_), .B(new_n12035_), .ZN(new_n12043_));
  XOR2_X1    g11786(.A1(new_n11643_), .A2(new_n12039_), .Z(new_n12044_));
  OAI21_X1   g11787(.A1(new_n12035_), .A2(new_n12044_), .B(new_n12043_), .ZN(new_n12045_));
  INV_X1     g11788(.I(new_n12045_), .ZN(new_n12046_));
  OAI22_X1   g11789(.A1(new_n848_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n795_), .ZN(new_n12047_));
  NAND2_X1   g11790(.A1(new_n8628_), .A2(\b[12] ), .ZN(new_n12048_));
  AOI21_X1   g11791(.A1(new_n12048_), .A2(new_n12047_), .B(new_n7354_), .ZN(new_n12049_));
  NAND2_X1   g11792(.A1(new_n847_), .A2(new_n12049_), .ZN(new_n12050_));
  XOR2_X1    g11793(.A1(new_n12050_), .A2(\a[59] ), .Z(new_n12051_));
  OAI22_X1   g11794(.A1(new_n659_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n617_), .ZN(new_n12052_));
  NAND2_X1   g11795(.A1(new_n9644_), .A2(\b[9] ), .ZN(new_n12053_));
  AOI21_X1   g11796(.A1(new_n12053_), .A2(new_n12052_), .B(new_n8321_), .ZN(new_n12054_));
  NAND2_X1   g11797(.A1(new_n663_), .A2(new_n12054_), .ZN(new_n12055_));
  XOR2_X1    g11798(.A1(new_n12055_), .A2(\a[62] ), .Z(new_n12056_));
  XNOR2_X1   g11799(.A1(new_n12051_), .A2(new_n12056_), .ZN(new_n12057_));
  NOR2_X1    g11800(.A1(new_n12046_), .A2(new_n12057_), .ZN(new_n12058_));
  NOR2_X1    g11801(.A1(new_n12051_), .A2(new_n12056_), .ZN(new_n12059_));
  INV_X1     g11802(.I(new_n12059_), .ZN(new_n12060_));
  NAND2_X1   g11803(.A1(new_n12051_), .A2(new_n12056_), .ZN(new_n12061_));
  AOI21_X1   g11804(.A1(new_n12060_), .A2(new_n12061_), .B(new_n12045_), .ZN(new_n12062_));
  NOR2_X1    g11805(.A1(new_n12058_), .A2(new_n12062_), .ZN(new_n12063_));
  OAI22_X1   g11806(.A1(new_n6721_), .A2(new_n992_), .B1(new_n6723_), .B2(new_n1044_), .ZN(new_n12064_));
  NAND2_X1   g11807(.A1(new_n7617_), .A2(\b[15] ), .ZN(new_n12065_));
  AOI21_X1   g11808(.A1(new_n12065_), .A2(new_n12064_), .B(new_n6731_), .ZN(new_n12066_));
  NAND2_X1   g11809(.A1(new_n1047_), .A2(new_n12066_), .ZN(new_n12067_));
  XOR2_X1    g11810(.A1(new_n12067_), .A2(new_n6516_), .Z(new_n12068_));
  INV_X1     g11811(.I(new_n11655_), .ZN(new_n12069_));
  AOI21_X1   g11812(.A1(new_n11657_), .A2(new_n11656_), .B(new_n11632_), .ZN(new_n12070_));
  NOR2_X1    g11813(.A1(new_n12069_), .A2(new_n12070_), .ZN(new_n12071_));
  XOR2_X1    g11814(.A1(new_n12068_), .A2(new_n12071_), .Z(new_n12072_));
  NOR2_X1    g11815(.A1(new_n12072_), .A2(new_n12063_), .ZN(new_n12073_));
  INV_X1     g11816(.I(new_n12063_), .ZN(new_n12074_));
  XOR2_X1    g11817(.A1(new_n12067_), .A2(\a[56] ), .Z(new_n12075_));
  NOR2_X1    g11818(.A1(new_n12075_), .A2(new_n12071_), .ZN(new_n12076_));
  INV_X1     g11819(.I(new_n12076_), .ZN(new_n12077_));
  NAND2_X1   g11820(.A1(new_n12075_), .A2(new_n12071_), .ZN(new_n12078_));
  AOI21_X1   g11821(.A1(new_n12077_), .A2(new_n12078_), .B(new_n12074_), .ZN(new_n12079_));
  NOR2_X1    g11822(.A1(new_n12073_), .A2(new_n12079_), .ZN(new_n12080_));
  AOI21_X1   g11823(.A1(new_n11664_), .A2(new_n11665_), .B(new_n11630_), .ZN(new_n12081_));
  NOR2_X1    g11824(.A1(new_n12081_), .A2(new_n11666_), .ZN(new_n12082_));
  INV_X1     g11825(.I(new_n12082_), .ZN(new_n12083_));
  XOR2_X1    g11826(.A1(new_n12080_), .A2(new_n12083_), .Z(new_n12084_));
  NOR2_X1    g11827(.A1(new_n12084_), .A2(new_n12032_), .ZN(new_n12085_));
  INV_X1     g11828(.I(new_n12032_), .ZN(new_n12086_));
  NOR2_X1    g11829(.A1(new_n12080_), .A2(new_n12082_), .ZN(new_n12087_));
  INV_X1     g11830(.I(new_n12087_), .ZN(new_n12088_));
  NAND2_X1   g11831(.A1(new_n12080_), .A2(new_n12082_), .ZN(new_n12089_));
  AOI21_X1   g11832(.A1(new_n12088_), .A2(new_n12089_), .B(new_n12086_), .ZN(new_n12090_));
  NOR2_X1    g11833(.A1(new_n12085_), .A2(new_n12090_), .ZN(new_n12091_));
  AOI21_X1   g11834(.A1(new_n11687_), .A2(new_n11685_), .B(new_n11683_), .ZN(new_n12092_));
  NOR2_X1    g11835(.A1(new_n12091_), .A2(new_n12092_), .ZN(new_n12093_));
  NAND2_X1   g11836(.A1(new_n12091_), .A2(new_n12092_), .ZN(new_n12094_));
  INV_X1     g11837(.I(new_n12094_), .ZN(new_n12095_));
  OAI21_X1   g11838(.A1(new_n12095_), .A2(new_n12093_), .B(new_n12027_), .ZN(new_n12096_));
  INV_X1     g11839(.I(new_n12092_), .ZN(new_n12097_));
  NAND2_X1   g11840(.A1(new_n12091_), .A2(new_n12097_), .ZN(new_n12098_));
  OAI21_X1   g11841(.A1(new_n12085_), .A2(new_n12090_), .B(new_n12092_), .ZN(new_n12099_));
  AOI21_X1   g11842(.A1(new_n12098_), .A2(new_n12099_), .B(new_n12027_), .ZN(new_n12100_));
  INV_X1     g11843(.I(new_n12100_), .ZN(new_n12101_));
  AOI21_X1   g11844(.A1(new_n12101_), .A2(new_n12096_), .B(new_n12021_), .ZN(new_n12102_));
  INV_X1     g11845(.I(new_n12093_), .ZN(new_n12103_));
  AOI21_X1   g11846(.A1(new_n12103_), .A2(new_n12094_), .B(new_n12026_), .ZN(new_n12104_));
  NOR3_X1    g11847(.A1(new_n12104_), .A2(new_n12100_), .A3(new_n12020_), .ZN(new_n12105_));
  OAI21_X1   g11848(.A1(new_n12102_), .A2(new_n12105_), .B(new_n12015_), .ZN(new_n12106_));
  AOI21_X1   g11849(.A1(new_n12101_), .A2(new_n12096_), .B(new_n12020_), .ZN(new_n12107_));
  NOR3_X1    g11850(.A1(new_n12104_), .A2(new_n12100_), .A3(new_n12021_), .ZN(new_n12108_));
  OAI21_X1   g11851(.A1(new_n12107_), .A2(new_n12108_), .B(new_n12014_), .ZN(new_n12109_));
  OAI22_X1   g11852(.A1(new_n4208_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n4203_), .ZN(new_n12110_));
  NAND2_X1   g11853(.A1(new_n5244_), .A2(\b[27] ), .ZN(new_n12111_));
  AOI21_X1   g11854(.A1(new_n12110_), .A2(new_n12111_), .B(new_n4211_), .ZN(new_n12112_));
  NAND2_X1   g11855(.A1(new_n2276_), .A2(new_n12112_), .ZN(new_n12113_));
  XOR2_X1    g11856(.A1(new_n12113_), .A2(\a[44] ), .Z(new_n12114_));
  AOI21_X1   g11857(.A1(new_n12106_), .A2(new_n12109_), .B(new_n12114_), .ZN(new_n12115_));
  OAI21_X1   g11858(.A1(new_n12104_), .A2(new_n12100_), .B(new_n12020_), .ZN(new_n12116_));
  NAND3_X1   g11859(.A1(new_n12101_), .A2(new_n12096_), .A3(new_n12021_), .ZN(new_n12117_));
  AOI21_X1   g11860(.A1(new_n12117_), .A2(new_n12116_), .B(new_n12014_), .ZN(new_n12118_));
  OAI21_X1   g11861(.A1(new_n12104_), .A2(new_n12100_), .B(new_n12021_), .ZN(new_n12119_));
  NAND3_X1   g11862(.A1(new_n12101_), .A2(new_n12096_), .A3(new_n12020_), .ZN(new_n12120_));
  AOI21_X1   g11863(.A1(new_n12120_), .A2(new_n12119_), .B(new_n12015_), .ZN(new_n12121_));
  INV_X1     g11864(.I(new_n12114_), .ZN(new_n12122_));
  NOR3_X1    g11865(.A1(new_n12118_), .A2(new_n12121_), .A3(new_n12122_), .ZN(new_n12123_));
  OAI21_X1   g11866(.A1(new_n12115_), .A2(new_n12123_), .B(new_n12013_), .ZN(new_n12124_));
  NOR3_X1    g11867(.A1(new_n12118_), .A2(new_n12121_), .A3(new_n12114_), .ZN(new_n12125_));
  AOI21_X1   g11868(.A1(new_n12106_), .A2(new_n12109_), .B(new_n12122_), .ZN(new_n12126_));
  OAI21_X1   g11869(.A1(new_n12126_), .A2(new_n12125_), .B(new_n12012_), .ZN(new_n12127_));
  OAI22_X1   g11870(.A1(new_n3736_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n3731_), .ZN(new_n12128_));
  NAND2_X1   g11871(.A1(new_n4730_), .A2(\b[30] ), .ZN(new_n12129_));
  AOI21_X1   g11872(.A1(new_n12128_), .A2(new_n12129_), .B(new_n3739_), .ZN(new_n12130_));
  NAND2_X1   g11873(.A1(new_n2659_), .A2(new_n12130_), .ZN(new_n12131_));
  XOR2_X1    g11874(.A1(new_n12131_), .A2(\a[41] ), .Z(new_n12132_));
  INV_X1     g11875(.I(new_n12132_), .ZN(new_n12133_));
  NAND3_X1   g11876(.A1(new_n12124_), .A2(new_n12127_), .A3(new_n12133_), .ZN(new_n12134_));
  OAI21_X1   g11877(.A1(new_n12118_), .A2(new_n12121_), .B(new_n12122_), .ZN(new_n12135_));
  NAND3_X1   g11878(.A1(new_n12106_), .A2(new_n12109_), .A3(new_n12114_), .ZN(new_n12136_));
  AOI21_X1   g11879(.A1(new_n12135_), .A2(new_n12136_), .B(new_n12012_), .ZN(new_n12137_));
  NAND3_X1   g11880(.A1(new_n12106_), .A2(new_n12109_), .A3(new_n12122_), .ZN(new_n12138_));
  OAI21_X1   g11881(.A1(new_n12118_), .A2(new_n12121_), .B(new_n12114_), .ZN(new_n12139_));
  AOI21_X1   g11882(.A1(new_n12139_), .A2(new_n12138_), .B(new_n12013_), .ZN(new_n12140_));
  OAI21_X1   g11883(.A1(new_n12137_), .A2(new_n12140_), .B(new_n12132_), .ZN(new_n12141_));
  AOI21_X1   g11884(.A1(new_n12141_), .A2(new_n12134_), .B(new_n12011_), .ZN(new_n12142_));
  OAI21_X1   g11885(.A1(new_n12137_), .A2(new_n12140_), .B(new_n12133_), .ZN(new_n12143_));
  NAND3_X1   g11886(.A1(new_n12124_), .A2(new_n12127_), .A3(new_n12132_), .ZN(new_n12144_));
  AOI21_X1   g11887(.A1(new_n12143_), .A2(new_n12144_), .B(new_n12010_), .ZN(new_n12145_));
  OAI22_X1   g11888(.A1(new_n3298_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n3293_), .ZN(new_n12146_));
  NAND2_X1   g11889(.A1(new_n4227_), .A2(\b[33] ), .ZN(new_n12147_));
  AOI21_X1   g11890(.A1(new_n12146_), .A2(new_n12147_), .B(new_n3301_), .ZN(new_n12148_));
  NAND2_X1   g11891(.A1(new_n3101_), .A2(new_n12148_), .ZN(new_n12149_));
  XOR2_X1    g11892(.A1(new_n12149_), .A2(\a[38] ), .Z(new_n12150_));
  NOR3_X1    g11893(.A1(new_n12142_), .A2(new_n12145_), .A3(new_n12150_), .ZN(new_n12151_));
  NOR3_X1    g11894(.A1(new_n12137_), .A2(new_n12140_), .A3(new_n12132_), .ZN(new_n12152_));
  AOI21_X1   g11895(.A1(new_n12124_), .A2(new_n12127_), .B(new_n12133_), .ZN(new_n12153_));
  OAI21_X1   g11896(.A1(new_n12153_), .A2(new_n12152_), .B(new_n12010_), .ZN(new_n12154_));
  AOI21_X1   g11897(.A1(new_n12124_), .A2(new_n12127_), .B(new_n12132_), .ZN(new_n12155_));
  NOR3_X1    g11898(.A1(new_n12137_), .A2(new_n12140_), .A3(new_n12133_), .ZN(new_n12156_));
  OAI21_X1   g11899(.A1(new_n12155_), .A2(new_n12156_), .B(new_n12011_), .ZN(new_n12157_));
  INV_X1     g11900(.I(new_n12150_), .ZN(new_n12158_));
  AOI21_X1   g11901(.A1(new_n12157_), .A2(new_n12154_), .B(new_n12158_), .ZN(new_n12159_));
  OAI21_X1   g11902(.A1(new_n12159_), .A2(new_n12151_), .B(new_n12005_), .ZN(new_n12160_));
  AOI21_X1   g11903(.A1(new_n12157_), .A2(new_n12154_), .B(new_n12150_), .ZN(new_n12161_));
  NOR3_X1    g11904(.A1(new_n12142_), .A2(new_n12145_), .A3(new_n12158_), .ZN(new_n12162_));
  OAI21_X1   g11905(.A1(new_n12161_), .A2(new_n12162_), .B(new_n12004_), .ZN(new_n12163_));
  NAND2_X1   g11906(.A1(new_n12160_), .A2(new_n12163_), .ZN(new_n12164_));
  NAND2_X1   g11907(.A1(new_n12164_), .A2(new_n12003_), .ZN(new_n12165_));
  INV_X1     g11908(.I(new_n12003_), .ZN(new_n12166_));
  NAND3_X1   g11909(.A1(new_n12157_), .A2(new_n12154_), .A3(new_n12158_), .ZN(new_n12167_));
  OAI21_X1   g11910(.A1(new_n12142_), .A2(new_n12145_), .B(new_n12150_), .ZN(new_n12168_));
  AOI21_X1   g11911(.A1(new_n12168_), .A2(new_n12167_), .B(new_n12004_), .ZN(new_n12169_));
  OAI21_X1   g11912(.A1(new_n12142_), .A2(new_n12145_), .B(new_n12158_), .ZN(new_n12170_));
  NAND3_X1   g11913(.A1(new_n12157_), .A2(new_n12154_), .A3(new_n12150_), .ZN(new_n12171_));
  AOI21_X1   g11914(.A1(new_n12170_), .A2(new_n12171_), .B(new_n12005_), .ZN(new_n12172_));
  NOR2_X1    g11915(.A1(new_n12169_), .A2(new_n12172_), .ZN(new_n12173_));
  NAND2_X1   g11916(.A1(new_n12173_), .A2(new_n12166_), .ZN(new_n12174_));
  AOI21_X1   g11917(.A1(new_n12165_), .A2(new_n12174_), .B(\a[35] ), .ZN(new_n12175_));
  NOR2_X1    g11918(.A1(new_n12173_), .A2(new_n12166_), .ZN(new_n12176_));
  NOR2_X1    g11919(.A1(new_n12164_), .A2(new_n12003_), .ZN(new_n12177_));
  NOR3_X1    g11920(.A1(new_n12177_), .A2(new_n12176_), .A3(new_n2836_), .ZN(new_n12178_));
  OAI21_X1   g11921(.A1(new_n12175_), .A2(new_n12178_), .B(new_n11998_), .ZN(new_n12179_));
  OAI21_X1   g11922(.A1(new_n12177_), .A2(new_n12176_), .B(new_n2836_), .ZN(new_n12180_));
  NAND3_X1   g11923(.A1(new_n12165_), .A2(new_n12174_), .A3(\a[35] ), .ZN(new_n12181_));
  NAND3_X1   g11924(.A1(new_n12180_), .A2(new_n12181_), .A3(new_n11997_), .ZN(new_n12182_));
  OAI22_X1   g11925(.A1(new_n2452_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n2447_), .ZN(new_n12183_));
  NAND2_X1   g11926(.A1(new_n3312_), .A2(\b[39] ), .ZN(new_n12184_));
  AOI21_X1   g11927(.A1(new_n12183_), .A2(new_n12184_), .B(new_n2455_), .ZN(new_n12185_));
  NAND2_X1   g11928(.A1(new_n3996_), .A2(new_n12185_), .ZN(new_n12186_));
  XOR2_X1    g11929(.A1(new_n12186_), .A2(\a[32] ), .Z(new_n12187_));
  INV_X1     g11930(.I(new_n12187_), .ZN(new_n12188_));
  NAND3_X1   g11931(.A1(new_n12179_), .A2(new_n12182_), .A3(new_n12188_), .ZN(new_n12189_));
  AOI21_X1   g11932(.A1(new_n12180_), .A2(new_n12181_), .B(new_n11997_), .ZN(new_n12190_));
  NOR3_X1    g11933(.A1(new_n12175_), .A2(new_n12178_), .A3(new_n11998_), .ZN(new_n12191_));
  OAI21_X1   g11934(.A1(new_n12191_), .A2(new_n12190_), .B(new_n12187_), .ZN(new_n12192_));
  AOI21_X1   g11935(.A1(new_n12192_), .A2(new_n12189_), .B(new_n11994_), .ZN(new_n12193_));
  INV_X1     g11936(.I(new_n11994_), .ZN(new_n12194_));
  OAI21_X1   g11937(.A1(new_n12191_), .A2(new_n12190_), .B(new_n12188_), .ZN(new_n12195_));
  NAND3_X1   g11938(.A1(new_n12179_), .A2(new_n12182_), .A3(new_n12187_), .ZN(new_n12196_));
  AOI21_X1   g11939(.A1(new_n12195_), .A2(new_n12196_), .B(new_n12194_), .ZN(new_n12197_));
  OAI22_X1   g11940(.A1(new_n2084_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n2079_), .ZN(new_n12198_));
  NAND2_X1   g11941(.A1(new_n2864_), .A2(\b[42] ), .ZN(new_n12199_));
  AOI21_X1   g11942(.A1(new_n12198_), .A2(new_n12199_), .B(new_n2087_), .ZN(new_n12200_));
  NAND2_X1   g11943(.A1(new_n4500_), .A2(new_n12200_), .ZN(new_n12201_));
  XOR2_X1    g11944(.A1(new_n12201_), .A2(\a[29] ), .Z(new_n12202_));
  INV_X1     g11945(.I(new_n12202_), .ZN(new_n12203_));
  OAI21_X1   g11946(.A1(new_n12193_), .A2(new_n12197_), .B(new_n12203_), .ZN(new_n12204_));
  NOR3_X1    g11947(.A1(new_n12193_), .A2(new_n12197_), .A3(new_n12203_), .ZN(new_n12205_));
  INV_X1     g11948(.I(new_n12205_), .ZN(new_n12206_));
  AOI21_X1   g11949(.A1(new_n12206_), .A2(new_n12204_), .B(new_n11993_), .ZN(new_n12207_));
  INV_X1     g11950(.I(new_n11993_), .ZN(new_n12208_));
  NOR3_X1    g11951(.A1(new_n12193_), .A2(new_n12197_), .A3(new_n12202_), .ZN(new_n12209_));
  INV_X1     g11952(.I(new_n12209_), .ZN(new_n12210_));
  OAI21_X1   g11953(.A1(new_n12193_), .A2(new_n12197_), .B(new_n12202_), .ZN(new_n12211_));
  AOI21_X1   g11954(.A1(new_n12210_), .A2(new_n12211_), .B(new_n12208_), .ZN(new_n12212_));
  OAI22_X1   g11955(.A1(new_n1760_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n1755_), .ZN(new_n12213_));
  NAND2_X1   g11956(.A1(new_n2470_), .A2(\b[45] ), .ZN(new_n12214_));
  AOI21_X1   g11957(.A1(new_n12213_), .A2(new_n12214_), .B(new_n1763_), .ZN(new_n12215_));
  NAND2_X1   g11958(.A1(new_n5004_), .A2(new_n12215_), .ZN(new_n12216_));
  XOR2_X1    g11959(.A1(new_n12216_), .A2(\a[26] ), .Z(new_n12217_));
  INV_X1     g11960(.I(new_n12217_), .ZN(new_n12218_));
  OAI21_X1   g11961(.A1(new_n12207_), .A2(new_n12212_), .B(new_n12218_), .ZN(new_n12219_));
  INV_X1     g11962(.I(new_n12204_), .ZN(new_n12220_));
  OAI21_X1   g11963(.A1(new_n12220_), .A2(new_n12205_), .B(new_n12208_), .ZN(new_n12221_));
  INV_X1     g11964(.I(new_n12211_), .ZN(new_n12222_));
  OAI21_X1   g11965(.A1(new_n12222_), .A2(new_n12209_), .B(new_n11993_), .ZN(new_n12223_));
  NAND3_X1   g11966(.A1(new_n12221_), .A2(new_n12223_), .A3(new_n12217_), .ZN(new_n12224_));
  AOI21_X1   g11967(.A1(new_n12219_), .A2(new_n12224_), .B(new_n11991_), .ZN(new_n12225_));
  INV_X1     g11968(.I(new_n11991_), .ZN(new_n12226_));
  NAND3_X1   g11969(.A1(new_n12221_), .A2(new_n12223_), .A3(new_n12218_), .ZN(new_n12227_));
  OAI21_X1   g11970(.A1(new_n12207_), .A2(new_n12212_), .B(new_n12217_), .ZN(new_n12228_));
  AOI21_X1   g11971(.A1(new_n12228_), .A2(new_n12227_), .B(new_n12226_), .ZN(new_n12229_));
  OAI22_X1   g11972(.A1(new_n1444_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n1439_), .ZN(new_n12230_));
  NAND2_X1   g11973(.A1(new_n2098_), .A2(\b[48] ), .ZN(new_n12231_));
  AOI21_X1   g11974(.A1(new_n12230_), .A2(new_n12231_), .B(new_n1447_), .ZN(new_n12232_));
  NAND2_X1   g11975(.A1(new_n5537_), .A2(new_n12232_), .ZN(new_n12233_));
  XOR2_X1    g11976(.A1(new_n12233_), .A2(\a[23] ), .Z(new_n12234_));
  NOR3_X1    g11977(.A1(new_n12225_), .A2(new_n12229_), .A3(new_n12234_), .ZN(new_n12235_));
  AOI21_X1   g11978(.A1(new_n12221_), .A2(new_n12223_), .B(new_n12217_), .ZN(new_n12236_));
  NOR3_X1    g11979(.A1(new_n12207_), .A2(new_n12212_), .A3(new_n12218_), .ZN(new_n12237_));
  OAI21_X1   g11980(.A1(new_n12236_), .A2(new_n12237_), .B(new_n12226_), .ZN(new_n12238_));
  NOR3_X1    g11981(.A1(new_n12207_), .A2(new_n12212_), .A3(new_n12217_), .ZN(new_n12239_));
  AOI21_X1   g11982(.A1(new_n12221_), .A2(new_n12223_), .B(new_n12218_), .ZN(new_n12240_));
  OAI21_X1   g11983(.A1(new_n12240_), .A2(new_n12239_), .B(new_n11991_), .ZN(new_n12241_));
  INV_X1     g11984(.I(new_n12234_), .ZN(new_n12242_));
  AOI21_X1   g11985(.A1(new_n12238_), .A2(new_n12241_), .B(new_n12242_), .ZN(new_n12243_));
  OAI21_X1   g11986(.A1(new_n12243_), .A2(new_n12235_), .B(new_n11990_), .ZN(new_n12244_));
  AOI21_X1   g11987(.A1(new_n12238_), .A2(new_n12241_), .B(new_n12234_), .ZN(new_n12245_));
  NOR3_X1    g11988(.A1(new_n12225_), .A2(new_n12229_), .A3(new_n12242_), .ZN(new_n12246_));
  OAI21_X1   g11989(.A1(new_n12245_), .A2(new_n12246_), .B(new_n11989_), .ZN(new_n12247_));
  OAI22_X1   g11990(.A1(new_n1168_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n1163_), .ZN(new_n12248_));
  NAND2_X1   g11991(.A1(new_n1774_), .A2(\b[51] ), .ZN(new_n12249_));
  AOI21_X1   g11992(.A1(new_n12248_), .A2(new_n12249_), .B(new_n1171_), .ZN(new_n12250_));
  NAND2_X1   g11993(.A1(new_n6219_), .A2(new_n12250_), .ZN(new_n12251_));
  XOR2_X1    g11994(.A1(new_n12251_), .A2(\a[20] ), .Z(new_n12252_));
  INV_X1     g11995(.I(new_n12252_), .ZN(new_n12253_));
  NAND3_X1   g11996(.A1(new_n12244_), .A2(new_n12247_), .A3(new_n12253_), .ZN(new_n12254_));
  NAND3_X1   g11997(.A1(new_n12238_), .A2(new_n12241_), .A3(new_n12242_), .ZN(new_n12255_));
  OAI21_X1   g11998(.A1(new_n12225_), .A2(new_n12229_), .B(new_n12234_), .ZN(new_n12256_));
  AOI21_X1   g11999(.A1(new_n12256_), .A2(new_n12255_), .B(new_n11989_), .ZN(new_n12257_));
  OAI21_X1   g12000(.A1(new_n12225_), .A2(new_n12229_), .B(new_n12242_), .ZN(new_n12258_));
  NAND3_X1   g12001(.A1(new_n12238_), .A2(new_n12241_), .A3(new_n12234_), .ZN(new_n12259_));
  AOI21_X1   g12002(.A1(new_n12258_), .A2(new_n12259_), .B(new_n11990_), .ZN(new_n12260_));
  OAI21_X1   g12003(.A1(new_n12257_), .A2(new_n12260_), .B(new_n12252_), .ZN(new_n12261_));
  AOI21_X1   g12004(.A1(new_n12261_), .A2(new_n12254_), .B(new_n11988_), .ZN(new_n12262_));
  INV_X1     g12005(.I(new_n11988_), .ZN(new_n12263_));
  OAI21_X1   g12006(.A1(new_n12257_), .A2(new_n12260_), .B(new_n12253_), .ZN(new_n12264_));
  NAND3_X1   g12007(.A1(new_n12244_), .A2(new_n12247_), .A3(new_n12252_), .ZN(new_n12265_));
  AOI21_X1   g12008(.A1(new_n12264_), .A2(new_n12265_), .B(new_n12263_), .ZN(new_n12266_));
  OAI22_X1   g12009(.A1(new_n940_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n935_), .ZN(new_n12267_));
  NAND2_X1   g12010(.A1(new_n1458_), .A2(\b[54] ), .ZN(new_n12268_));
  AOI21_X1   g12011(.A1(new_n12267_), .A2(new_n12268_), .B(new_n943_), .ZN(new_n12269_));
  NAND2_X1   g12012(.A1(new_n6994_), .A2(new_n12269_), .ZN(new_n12270_));
  XOR2_X1    g12013(.A1(new_n12270_), .A2(\a[17] ), .Z(new_n12271_));
  INV_X1     g12014(.I(new_n12271_), .ZN(new_n12272_));
  OAI21_X1   g12015(.A1(new_n12262_), .A2(new_n12266_), .B(new_n12272_), .ZN(new_n12273_));
  NOR3_X1    g12016(.A1(new_n12257_), .A2(new_n12260_), .A3(new_n12252_), .ZN(new_n12274_));
  AOI21_X1   g12017(.A1(new_n12244_), .A2(new_n12247_), .B(new_n12253_), .ZN(new_n12275_));
  OAI21_X1   g12018(.A1(new_n12275_), .A2(new_n12274_), .B(new_n12263_), .ZN(new_n12276_));
  AOI21_X1   g12019(.A1(new_n12244_), .A2(new_n12247_), .B(new_n12252_), .ZN(new_n12277_));
  NOR3_X1    g12020(.A1(new_n12257_), .A2(new_n12260_), .A3(new_n12253_), .ZN(new_n12278_));
  OAI21_X1   g12021(.A1(new_n12277_), .A2(new_n12278_), .B(new_n11988_), .ZN(new_n12279_));
  NAND3_X1   g12022(.A1(new_n12276_), .A2(new_n12279_), .A3(new_n12271_), .ZN(new_n12280_));
  AOI21_X1   g12023(.A1(new_n12273_), .A2(new_n12280_), .B(new_n11987_), .ZN(new_n12281_));
  INV_X1     g12024(.I(new_n11987_), .ZN(new_n12282_));
  NAND3_X1   g12025(.A1(new_n12276_), .A2(new_n12279_), .A3(new_n12272_), .ZN(new_n12283_));
  OAI21_X1   g12026(.A1(new_n12262_), .A2(new_n12266_), .B(new_n12271_), .ZN(new_n12284_));
  AOI21_X1   g12027(.A1(new_n12284_), .A2(new_n12283_), .B(new_n12282_), .ZN(new_n12285_));
  OAI22_X1   g12028(.A1(new_n757_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n752_), .ZN(new_n12286_));
  NAND2_X1   g12029(.A1(new_n1182_), .A2(\b[57] ), .ZN(new_n12287_));
  AOI21_X1   g12030(.A1(new_n12286_), .A2(new_n12287_), .B(new_n760_), .ZN(new_n12288_));
  NAND2_X1   g12031(.A1(new_n7895_), .A2(new_n12288_), .ZN(new_n12289_));
  XOR2_X1    g12032(.A1(new_n12289_), .A2(\a[14] ), .Z(new_n12290_));
  INV_X1     g12033(.I(new_n12290_), .ZN(new_n12291_));
  OAI21_X1   g12034(.A1(new_n12281_), .A2(new_n12285_), .B(new_n12291_), .ZN(new_n12292_));
  AOI21_X1   g12035(.A1(new_n12276_), .A2(new_n12279_), .B(new_n12271_), .ZN(new_n12293_));
  NOR3_X1    g12036(.A1(new_n12262_), .A2(new_n12266_), .A3(new_n12272_), .ZN(new_n12294_));
  OAI21_X1   g12037(.A1(new_n12293_), .A2(new_n12294_), .B(new_n12282_), .ZN(new_n12295_));
  NOR3_X1    g12038(.A1(new_n12262_), .A2(new_n12266_), .A3(new_n12271_), .ZN(new_n12296_));
  AOI21_X1   g12039(.A1(new_n12276_), .A2(new_n12279_), .B(new_n12272_), .ZN(new_n12297_));
  OAI21_X1   g12040(.A1(new_n12297_), .A2(new_n12296_), .B(new_n11987_), .ZN(new_n12298_));
  NAND3_X1   g12041(.A1(new_n12295_), .A2(new_n12298_), .A3(new_n12290_), .ZN(new_n12299_));
  NAND2_X1   g12042(.A1(new_n12292_), .A2(new_n12299_), .ZN(new_n12300_));
  NAND3_X1   g12043(.A1(new_n12295_), .A2(new_n12298_), .A3(new_n12291_), .ZN(new_n12301_));
  OAI21_X1   g12044(.A1(new_n12281_), .A2(new_n12285_), .B(new_n12290_), .ZN(new_n12302_));
  NAND2_X1   g12045(.A1(new_n12302_), .A2(new_n12301_), .ZN(new_n12303_));
  MUX2_X1    g12046(.I0(new_n12303_), .I1(new_n12300_), .S(new_n11986_), .Z(new_n12304_));
  NAND2_X1   g12047(.A1(new_n11914_), .A2(new_n11588_), .ZN(new_n12305_));
  NAND2_X1   g12048(.A1(new_n12305_), .A2(new_n11910_), .ZN(new_n12306_));
  OAI22_X1   g12049(.A1(new_n582_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n577_), .ZN(new_n12307_));
  NAND2_X1   g12050(.A1(new_n960_), .A2(\b[60] ), .ZN(new_n12308_));
  AOI21_X1   g12051(.A1(new_n12307_), .A2(new_n12308_), .B(new_n585_), .ZN(new_n12309_));
  NAND2_X1   g12052(.A1(new_n8935_), .A2(new_n12309_), .ZN(new_n12310_));
  XOR2_X1    g12053(.A1(new_n12310_), .A2(new_n572_), .Z(new_n12311_));
  XOR2_X1    g12054(.A1(new_n12306_), .A2(new_n12311_), .Z(new_n12312_));
  NAND2_X1   g12055(.A1(new_n12304_), .A2(new_n12312_), .ZN(new_n12313_));
  NAND2_X1   g12056(.A1(new_n12306_), .A2(new_n12311_), .ZN(new_n12314_));
  OR2_X2     g12057(.A1(new_n12306_), .A2(new_n12311_), .Z(new_n12315_));
  AND2_X2    g12058(.A1(new_n12315_), .A2(new_n12314_), .Z(new_n12316_));
  OAI21_X1   g12059(.A1(new_n12304_), .A2(new_n12316_), .B(new_n12313_), .ZN(new_n12317_));
  XNOR2_X1   g12060(.A1(new_n12317_), .A2(new_n11984_), .ZN(new_n12318_));
  NAND2_X1   g12061(.A1(new_n12318_), .A2(new_n429_), .ZN(new_n12319_));
  XOR2_X1    g12062(.A1(new_n12317_), .A2(new_n11984_), .Z(new_n12320_));
  NAND2_X1   g12063(.A1(new_n12320_), .A2(\a[8] ), .ZN(new_n12321_));
  AOI21_X1   g12064(.A1(new_n12319_), .A2(new_n12321_), .B(new_n11982_), .ZN(new_n12322_));
  NOR2_X1    g12065(.A1(new_n12320_), .A2(\a[8] ), .ZN(new_n12323_));
  NOR2_X1    g12066(.A1(new_n12318_), .A2(new_n429_), .ZN(new_n12324_));
  NOR3_X1    g12067(.A1(new_n12324_), .A2(new_n12323_), .A3(new_n11981_), .ZN(new_n12325_));
  NOR2_X1    g12068(.A1(new_n12325_), .A2(new_n12322_), .ZN(new_n12326_));
  XOR2_X1    g12069(.A1(new_n12326_), .A2(new_n11980_), .Z(new_n12327_));
  OAI21_X1   g12070(.A1(new_n12324_), .A2(new_n12323_), .B(new_n11981_), .ZN(new_n12328_));
  NAND3_X1   g12071(.A1(new_n12319_), .A2(new_n12321_), .A3(new_n11982_), .ZN(new_n12329_));
  AOI21_X1   g12072(.A1(new_n12328_), .A2(new_n12329_), .B(new_n11979_), .ZN(new_n12330_));
  NOR3_X1    g12073(.A1(new_n12325_), .A2(new_n12322_), .A3(new_n11980_), .ZN(new_n12331_));
  OAI21_X1   g12074(.A1(new_n12330_), .A2(new_n12331_), .B(new_n11977_), .ZN(new_n12332_));
  OAI21_X1   g12075(.A1(new_n11977_), .A2(new_n12327_), .B(new_n12332_), .ZN(\f[71] ));
  XOR2_X1    g12076(.A1(new_n11981_), .A2(new_n429_), .Z(new_n12334_));
  XOR2_X1    g12077(.A1(new_n11984_), .A2(new_n12334_), .Z(new_n12335_));
  AOI21_X1   g12078(.A1(new_n12317_), .A2(new_n12334_), .B(new_n12335_), .ZN(new_n12336_));
  NAND2_X1   g12079(.A1(new_n12304_), .A2(new_n12315_), .ZN(new_n12337_));
  NAND2_X1   g12080(.A1(new_n12337_), .A2(new_n12314_), .ZN(new_n12338_));
  NAND2_X1   g12081(.A1(new_n12299_), .A2(new_n11986_), .ZN(new_n12339_));
  AND2_X2    g12082(.A1(new_n12339_), .A2(new_n12292_), .Z(new_n12340_));
  AOI21_X1   g12083(.A1(new_n12282_), .A2(new_n12280_), .B(new_n12293_), .ZN(new_n12341_));
  INV_X1     g12084(.I(new_n12341_), .ZN(new_n12342_));
  AOI21_X1   g12085(.A1(new_n12263_), .A2(new_n12261_), .B(new_n12274_), .ZN(new_n12343_));
  AOI21_X1   g12086(.A1(new_n11990_), .A2(new_n12259_), .B(new_n12245_), .ZN(new_n12344_));
  AOI21_X1   g12087(.A1(new_n12226_), .A2(new_n12224_), .B(new_n12236_), .ZN(new_n12345_));
  INV_X1     g12088(.I(new_n12189_), .ZN(new_n12346_));
  AOI21_X1   g12089(.A1(new_n12194_), .A2(new_n12192_), .B(new_n12346_), .ZN(new_n12347_));
  NAND2_X1   g12090(.A1(new_n12164_), .A2(new_n12166_), .ZN(new_n12348_));
  XOR2_X1    g12091(.A1(new_n11997_), .A2(\a[35] ), .Z(new_n12349_));
  OAI21_X1   g12092(.A1(new_n12164_), .A2(new_n12166_), .B(new_n12349_), .ZN(new_n12350_));
  NAND2_X1   g12093(.A1(new_n12350_), .A2(new_n12348_), .ZN(new_n12351_));
  INV_X1     g12094(.I(new_n12351_), .ZN(new_n12352_));
  AOI21_X1   g12095(.A1(new_n12005_), .A2(new_n12168_), .B(new_n12151_), .ZN(new_n12353_));
  INV_X1     g12096(.I(new_n12353_), .ZN(new_n12354_));
  AOI21_X1   g12097(.A1(new_n12010_), .A2(new_n12144_), .B(new_n12155_), .ZN(new_n12355_));
  AOI21_X1   g12098(.A1(new_n12013_), .A2(new_n12136_), .B(new_n12115_), .ZN(new_n12356_));
  AOI21_X1   g12099(.A1(new_n12015_), .A2(new_n12116_), .B(new_n12105_), .ZN(new_n12357_));
  NAND2_X1   g12100(.A1(new_n12099_), .A2(new_n12027_), .ZN(new_n12358_));
  AND2_X2    g12101(.A1(new_n12358_), .A2(new_n12098_), .Z(new_n12359_));
  INV_X1     g12102(.I(new_n12359_), .ZN(new_n12360_));
  OAI22_X1   g12103(.A1(new_n5228_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n5225_), .ZN(new_n12361_));
  NAND2_X1   g12104(.A1(new_n5387_), .A2(\b[22] ), .ZN(new_n12362_));
  AOI21_X1   g12105(.A1(new_n12361_), .A2(new_n12362_), .B(new_n5231_), .ZN(new_n12363_));
  NAND2_X1   g12106(.A1(new_n1708_), .A2(new_n12363_), .ZN(new_n12364_));
  XOR2_X1    g12107(.A1(new_n12364_), .A2(\a[50] ), .Z(new_n12365_));
  INV_X1     g12108(.I(new_n12365_), .ZN(new_n12366_));
  AOI21_X1   g12109(.A1(new_n12086_), .A2(new_n12089_), .B(new_n12087_), .ZN(new_n12367_));
  AOI21_X1   g12110(.A1(new_n12045_), .A2(new_n12061_), .B(new_n12059_), .ZN(new_n12368_));
  INV_X1     g12111(.I(new_n12040_), .ZN(new_n12369_));
  AOI21_X1   g12112(.A1(new_n12035_), .A2(new_n12369_), .B(new_n12042_), .ZN(new_n12370_));
  OAI22_X1   g12113(.A1(new_n717_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n659_), .ZN(new_n12371_));
  NAND2_X1   g12114(.A1(new_n9644_), .A2(\b[10] ), .ZN(new_n12372_));
  AOI21_X1   g12115(.A1(new_n12372_), .A2(new_n12371_), .B(new_n8321_), .ZN(new_n12373_));
  NAND2_X1   g12116(.A1(new_n716_), .A2(new_n12373_), .ZN(new_n12374_));
  XOR2_X1    g12117(.A1(new_n12374_), .A2(new_n8309_), .Z(new_n12375_));
  NOR2_X1    g12118(.A1(new_n8985_), .A2(new_n510_), .ZN(new_n12376_));
  NOR2_X1    g12119(.A1(new_n9364_), .A2(new_n495_), .ZN(new_n12377_));
  XNOR2_X1   g12120(.A1(new_n12376_), .A2(new_n12377_), .ZN(new_n12378_));
  XOR2_X1    g12121(.A1(new_n12378_), .A2(\a[8] ), .Z(new_n12379_));
  NOR2_X1    g12122(.A1(new_n12379_), .A2(new_n12039_), .ZN(new_n12380_));
  NOR2_X1    g12123(.A1(new_n12378_), .A2(new_n429_), .ZN(new_n12381_));
  INV_X1     g12124(.I(new_n12381_), .ZN(new_n12382_));
  NAND2_X1   g12125(.A1(new_n12378_), .A2(new_n429_), .ZN(new_n12383_));
  AOI21_X1   g12126(.A1(new_n12382_), .A2(new_n12383_), .B(new_n12041_), .ZN(new_n12384_));
  NOR2_X1    g12127(.A1(new_n12380_), .A2(new_n12384_), .ZN(new_n12385_));
  NOR2_X1    g12128(.A1(new_n12375_), .A2(new_n12385_), .ZN(new_n12386_));
  NAND2_X1   g12129(.A1(new_n12375_), .A2(new_n12385_), .ZN(new_n12387_));
  INV_X1     g12130(.I(new_n12387_), .ZN(new_n12388_));
  NOR2_X1    g12131(.A1(new_n12388_), .A2(new_n12386_), .ZN(new_n12389_));
  XOR2_X1    g12132(.A1(new_n12375_), .A2(new_n12385_), .Z(new_n12390_));
  NAND2_X1   g12133(.A1(new_n12390_), .A2(new_n12370_), .ZN(new_n12391_));
  OAI21_X1   g12134(.A1(new_n12370_), .A2(new_n12389_), .B(new_n12391_), .ZN(new_n12392_));
  OAI22_X1   g12135(.A1(new_n904_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n848_), .ZN(new_n12393_));
  NAND2_X1   g12136(.A1(new_n8628_), .A2(\b[13] ), .ZN(new_n12394_));
  AOI21_X1   g12137(.A1(new_n12394_), .A2(new_n12393_), .B(new_n7354_), .ZN(new_n12395_));
  NAND2_X1   g12138(.A1(new_n907_), .A2(new_n12395_), .ZN(new_n12396_));
  XOR2_X1    g12139(.A1(new_n12396_), .A2(new_n7343_), .Z(new_n12397_));
  XNOR2_X1   g12140(.A1(new_n12392_), .A2(new_n12397_), .ZN(new_n12398_));
  NOR2_X1    g12141(.A1(new_n12398_), .A2(new_n12368_), .ZN(new_n12399_));
  INV_X1     g12142(.I(new_n12368_), .ZN(new_n12400_));
  NAND2_X1   g12143(.A1(new_n12392_), .A2(new_n12397_), .ZN(new_n12401_));
  NOR2_X1    g12144(.A1(new_n12392_), .A2(new_n12397_), .ZN(new_n12402_));
  INV_X1     g12145(.I(new_n12402_), .ZN(new_n12403_));
  AOI21_X1   g12146(.A1(new_n12403_), .A2(new_n12401_), .B(new_n12400_), .ZN(new_n12404_));
  NOR2_X1    g12147(.A1(new_n12399_), .A2(new_n12404_), .ZN(new_n12405_));
  OAI22_X1   g12148(.A1(new_n6721_), .A2(new_n1044_), .B1(new_n6723_), .B2(new_n1124_), .ZN(new_n12406_));
  NAND2_X1   g12149(.A1(new_n7617_), .A2(\b[16] ), .ZN(new_n12407_));
  AOI21_X1   g12150(.A1(new_n12407_), .A2(new_n12406_), .B(new_n6731_), .ZN(new_n12408_));
  NAND2_X1   g12151(.A1(new_n1123_), .A2(new_n12408_), .ZN(new_n12409_));
  XOR2_X1    g12152(.A1(new_n12409_), .A2(\a[56] ), .Z(new_n12410_));
  INV_X1     g12153(.I(new_n12410_), .ZN(new_n12411_));
  AOI21_X1   g12154(.A1(new_n12075_), .A2(new_n12071_), .B(new_n12074_), .ZN(new_n12412_));
  OAI21_X1   g12155(.A1(new_n12412_), .A2(new_n12076_), .B(new_n12411_), .ZN(new_n12413_));
  NOR2_X1    g12156(.A1(new_n12412_), .A2(new_n12076_), .ZN(new_n12414_));
  NAND2_X1   g12157(.A1(new_n12414_), .A2(new_n12410_), .ZN(new_n12415_));
  AOI21_X1   g12158(.A1(new_n12415_), .A2(new_n12413_), .B(new_n12405_), .ZN(new_n12416_));
  XOR2_X1    g12159(.A1(new_n12414_), .A2(new_n12411_), .Z(new_n12417_));
  NOR3_X1    g12160(.A1(new_n12417_), .A2(new_n12399_), .A3(new_n12404_), .ZN(new_n12418_));
  NOR2_X1    g12161(.A1(new_n12418_), .A2(new_n12416_), .ZN(new_n12419_));
  OAI22_X1   g12162(.A1(new_n5786_), .A2(new_n1393_), .B1(new_n1305_), .B2(new_n5792_), .ZN(new_n12420_));
  NAND2_X1   g12163(.A1(new_n6745_), .A2(\b[19] ), .ZN(new_n12421_));
  AOI21_X1   g12164(.A1(new_n12421_), .A2(new_n12420_), .B(new_n5796_), .ZN(new_n12422_));
  NAND2_X1   g12165(.A1(new_n1396_), .A2(new_n12422_), .ZN(new_n12423_));
  XOR2_X1    g12166(.A1(new_n12423_), .A2(\a[53] ), .Z(new_n12424_));
  XOR2_X1    g12167(.A1(new_n12419_), .A2(new_n12424_), .Z(new_n12425_));
  NOR2_X1    g12168(.A1(new_n12425_), .A2(new_n12367_), .ZN(new_n12426_));
  INV_X1     g12169(.I(new_n12367_), .ZN(new_n12427_));
  INV_X1     g12170(.I(new_n12424_), .ZN(new_n12428_));
  NAND2_X1   g12171(.A1(new_n12419_), .A2(new_n12428_), .ZN(new_n12429_));
  INV_X1     g12172(.I(new_n12419_), .ZN(new_n12430_));
  NAND2_X1   g12173(.A1(new_n12430_), .A2(new_n12424_), .ZN(new_n12431_));
  AOI21_X1   g12174(.A1(new_n12431_), .A2(new_n12429_), .B(new_n12427_), .ZN(new_n12432_));
  NOR2_X1    g12175(.A1(new_n12426_), .A2(new_n12432_), .ZN(new_n12433_));
  NOR2_X1    g12176(.A1(new_n12433_), .A2(new_n12366_), .ZN(new_n12434_));
  NAND2_X1   g12177(.A1(new_n12433_), .A2(new_n12366_), .ZN(new_n12435_));
  INV_X1     g12178(.I(new_n12435_), .ZN(new_n12436_));
  OAI21_X1   g12179(.A1(new_n12436_), .A2(new_n12434_), .B(new_n12360_), .ZN(new_n12437_));
  NOR2_X1    g12180(.A1(new_n12433_), .A2(new_n12365_), .ZN(new_n12438_));
  NAND2_X1   g12181(.A1(new_n12433_), .A2(new_n12365_), .ZN(new_n12439_));
  INV_X1     g12182(.I(new_n12439_), .ZN(new_n12440_));
  OAI21_X1   g12183(.A1(new_n12440_), .A2(new_n12438_), .B(new_n12359_), .ZN(new_n12441_));
  OAI22_X1   g12184(.A1(new_n4711_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n4706_), .ZN(new_n12442_));
  NAND2_X1   g12185(.A1(new_n5814_), .A2(\b[25] ), .ZN(new_n12443_));
  AOI21_X1   g12186(.A1(new_n12442_), .A2(new_n12443_), .B(new_n4714_), .ZN(new_n12444_));
  NAND2_X1   g12187(.A1(new_n2042_), .A2(new_n12444_), .ZN(new_n12445_));
  XOR2_X1    g12188(.A1(new_n12445_), .A2(\a[47] ), .Z(new_n12446_));
  INV_X1     g12189(.I(new_n12446_), .ZN(new_n12447_));
  NAND3_X1   g12190(.A1(new_n12437_), .A2(new_n12441_), .A3(new_n12447_), .ZN(new_n12448_));
  NAND2_X1   g12191(.A1(new_n12437_), .A2(new_n12441_), .ZN(new_n12449_));
  NAND2_X1   g12192(.A1(new_n12449_), .A2(new_n12446_), .ZN(new_n12450_));
  AOI21_X1   g12193(.A1(new_n12450_), .A2(new_n12448_), .B(new_n12357_), .ZN(new_n12451_));
  INV_X1     g12194(.I(new_n12357_), .ZN(new_n12452_));
  AOI21_X1   g12195(.A1(new_n12437_), .A2(new_n12441_), .B(new_n12446_), .ZN(new_n12453_));
  INV_X1     g12196(.I(new_n12453_), .ZN(new_n12454_));
  NAND3_X1   g12197(.A1(new_n12437_), .A2(new_n12441_), .A3(new_n12446_), .ZN(new_n12455_));
  AOI21_X1   g12198(.A1(new_n12454_), .A2(new_n12455_), .B(new_n12452_), .ZN(new_n12456_));
  OAI22_X1   g12199(.A1(new_n4208_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n4203_), .ZN(new_n12457_));
  NAND2_X1   g12200(.A1(new_n5244_), .A2(\b[28] ), .ZN(new_n12458_));
  AOI21_X1   g12201(.A1(new_n12457_), .A2(new_n12458_), .B(new_n4211_), .ZN(new_n12459_));
  NAND2_X1   g12202(.A1(new_n2404_), .A2(new_n12459_), .ZN(new_n12460_));
  XOR2_X1    g12203(.A1(new_n12460_), .A2(\a[44] ), .Z(new_n12461_));
  NOR3_X1    g12204(.A1(new_n12456_), .A2(new_n12451_), .A3(new_n12461_), .ZN(new_n12462_));
  INV_X1     g12205(.I(new_n12462_), .ZN(new_n12463_));
  OAI21_X1   g12206(.A1(new_n12456_), .A2(new_n12451_), .B(new_n12461_), .ZN(new_n12464_));
  AOI21_X1   g12207(.A1(new_n12463_), .A2(new_n12464_), .B(new_n12356_), .ZN(new_n12465_));
  INV_X1     g12208(.I(new_n12356_), .ZN(new_n12466_));
  INV_X1     g12209(.I(new_n12461_), .ZN(new_n12467_));
  OAI21_X1   g12210(.A1(new_n12456_), .A2(new_n12451_), .B(new_n12467_), .ZN(new_n12468_));
  NOR3_X1    g12211(.A1(new_n12456_), .A2(new_n12451_), .A3(new_n12467_), .ZN(new_n12469_));
  INV_X1     g12212(.I(new_n12469_), .ZN(new_n12470_));
  AOI21_X1   g12213(.A1(new_n12470_), .A2(new_n12468_), .B(new_n12466_), .ZN(new_n12471_));
  OAI22_X1   g12214(.A1(new_n3736_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n3731_), .ZN(new_n12472_));
  NAND2_X1   g12215(.A1(new_n4730_), .A2(\b[31] ), .ZN(new_n12473_));
  AOI21_X1   g12216(.A1(new_n12472_), .A2(new_n12473_), .B(new_n3739_), .ZN(new_n12474_));
  NAND2_X1   g12217(.A1(new_n2797_), .A2(new_n12474_), .ZN(new_n12475_));
  XOR2_X1    g12218(.A1(new_n12475_), .A2(\a[41] ), .Z(new_n12476_));
  INV_X1     g12219(.I(new_n12476_), .ZN(new_n12477_));
  OAI21_X1   g12220(.A1(new_n12465_), .A2(new_n12471_), .B(new_n12477_), .ZN(new_n12478_));
  INV_X1     g12221(.I(new_n12464_), .ZN(new_n12479_));
  OAI21_X1   g12222(.A1(new_n12479_), .A2(new_n12462_), .B(new_n12466_), .ZN(new_n12480_));
  INV_X1     g12223(.I(new_n12468_), .ZN(new_n12481_));
  OAI21_X1   g12224(.A1(new_n12481_), .A2(new_n12469_), .B(new_n12356_), .ZN(new_n12482_));
  NAND3_X1   g12225(.A1(new_n12480_), .A2(new_n12482_), .A3(new_n12476_), .ZN(new_n12483_));
  AOI21_X1   g12226(.A1(new_n12478_), .A2(new_n12483_), .B(new_n12355_), .ZN(new_n12484_));
  INV_X1     g12227(.I(new_n12355_), .ZN(new_n12485_));
  NAND3_X1   g12228(.A1(new_n12480_), .A2(new_n12482_), .A3(new_n12477_), .ZN(new_n12486_));
  OAI21_X1   g12229(.A1(new_n12465_), .A2(new_n12471_), .B(new_n12476_), .ZN(new_n12487_));
  AOI21_X1   g12230(.A1(new_n12487_), .A2(new_n12486_), .B(new_n12485_), .ZN(new_n12488_));
  OAI22_X1   g12231(.A1(new_n3298_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n3293_), .ZN(new_n12489_));
  NAND2_X1   g12232(.A1(new_n4227_), .A2(\b[34] ), .ZN(new_n12490_));
  AOI21_X1   g12233(.A1(new_n12489_), .A2(new_n12490_), .B(new_n3301_), .ZN(new_n12491_));
  NAND2_X1   g12234(.A1(new_n3246_), .A2(new_n12491_), .ZN(new_n12492_));
  XOR2_X1    g12235(.A1(new_n12492_), .A2(\a[38] ), .Z(new_n12493_));
  NOR3_X1    g12236(.A1(new_n12484_), .A2(new_n12488_), .A3(new_n12493_), .ZN(new_n12494_));
  AOI21_X1   g12237(.A1(new_n12480_), .A2(new_n12482_), .B(new_n12476_), .ZN(new_n12495_));
  NOR3_X1    g12238(.A1(new_n12465_), .A2(new_n12471_), .A3(new_n12477_), .ZN(new_n12496_));
  OAI21_X1   g12239(.A1(new_n12495_), .A2(new_n12496_), .B(new_n12485_), .ZN(new_n12497_));
  NOR3_X1    g12240(.A1(new_n12465_), .A2(new_n12471_), .A3(new_n12476_), .ZN(new_n12498_));
  AOI21_X1   g12241(.A1(new_n12480_), .A2(new_n12482_), .B(new_n12477_), .ZN(new_n12499_));
  OAI21_X1   g12242(.A1(new_n12499_), .A2(new_n12498_), .B(new_n12355_), .ZN(new_n12500_));
  INV_X1     g12243(.I(new_n12493_), .ZN(new_n12501_));
  AOI21_X1   g12244(.A1(new_n12497_), .A2(new_n12500_), .B(new_n12501_), .ZN(new_n12502_));
  OAI21_X1   g12245(.A1(new_n12502_), .A2(new_n12494_), .B(new_n12354_), .ZN(new_n12503_));
  AOI21_X1   g12246(.A1(new_n12497_), .A2(new_n12500_), .B(new_n12493_), .ZN(new_n12504_));
  NOR3_X1    g12247(.A1(new_n12484_), .A2(new_n12488_), .A3(new_n12501_), .ZN(new_n12505_));
  OAI21_X1   g12248(.A1(new_n12504_), .A2(new_n12505_), .B(new_n12353_), .ZN(new_n12506_));
  OAI22_X1   g12249(.A1(new_n2846_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n2841_), .ZN(new_n12507_));
  NAND2_X1   g12250(.A1(new_n3755_), .A2(\b[37] ), .ZN(new_n12508_));
  AOI21_X1   g12251(.A1(new_n12507_), .A2(new_n12508_), .B(new_n2849_), .ZN(new_n12509_));
  NAND2_X1   g12252(.A1(new_n3700_), .A2(new_n12509_), .ZN(new_n12510_));
  XOR2_X1    g12253(.A1(new_n12510_), .A2(\a[35] ), .Z(new_n12511_));
  INV_X1     g12254(.I(new_n12511_), .ZN(new_n12512_));
  NAND3_X1   g12255(.A1(new_n12503_), .A2(new_n12506_), .A3(new_n12512_), .ZN(new_n12513_));
  NAND3_X1   g12256(.A1(new_n12497_), .A2(new_n12500_), .A3(new_n12501_), .ZN(new_n12514_));
  OAI21_X1   g12257(.A1(new_n12484_), .A2(new_n12488_), .B(new_n12493_), .ZN(new_n12515_));
  AOI21_X1   g12258(.A1(new_n12515_), .A2(new_n12514_), .B(new_n12353_), .ZN(new_n12516_));
  OAI21_X1   g12259(.A1(new_n12484_), .A2(new_n12488_), .B(new_n12501_), .ZN(new_n12517_));
  NAND3_X1   g12260(.A1(new_n12497_), .A2(new_n12500_), .A3(new_n12493_), .ZN(new_n12518_));
  AOI21_X1   g12261(.A1(new_n12517_), .A2(new_n12518_), .B(new_n12354_), .ZN(new_n12519_));
  OAI21_X1   g12262(.A1(new_n12516_), .A2(new_n12519_), .B(new_n12511_), .ZN(new_n12520_));
  AOI21_X1   g12263(.A1(new_n12520_), .A2(new_n12513_), .B(new_n12352_), .ZN(new_n12521_));
  OAI21_X1   g12264(.A1(new_n12516_), .A2(new_n12519_), .B(new_n12512_), .ZN(new_n12522_));
  NAND3_X1   g12265(.A1(new_n12503_), .A2(new_n12506_), .A3(new_n12511_), .ZN(new_n12523_));
  AOI21_X1   g12266(.A1(new_n12522_), .A2(new_n12523_), .B(new_n12351_), .ZN(new_n12524_));
  OAI22_X1   g12267(.A1(new_n2452_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n2447_), .ZN(new_n12525_));
  NAND2_X1   g12268(.A1(new_n3312_), .A2(\b[40] ), .ZN(new_n12526_));
  AOI21_X1   g12269(.A1(new_n12525_), .A2(new_n12526_), .B(new_n2455_), .ZN(new_n12527_));
  NAND2_X1   g12270(.A1(new_n4017_), .A2(new_n12527_), .ZN(new_n12528_));
  XOR2_X1    g12271(.A1(new_n12528_), .A2(\a[32] ), .Z(new_n12529_));
  INV_X1     g12272(.I(new_n12529_), .ZN(new_n12530_));
  OAI21_X1   g12273(.A1(new_n12521_), .A2(new_n12524_), .B(new_n12530_), .ZN(new_n12531_));
  INV_X1     g12274(.I(new_n12531_), .ZN(new_n12532_));
  NOR3_X1    g12275(.A1(new_n12521_), .A2(new_n12524_), .A3(new_n12530_), .ZN(new_n12533_));
  NOR2_X1    g12276(.A1(new_n12532_), .A2(new_n12533_), .ZN(new_n12534_));
  NOR3_X1    g12277(.A1(new_n12521_), .A2(new_n12524_), .A3(new_n12529_), .ZN(new_n12535_));
  NOR3_X1    g12278(.A1(new_n12516_), .A2(new_n12519_), .A3(new_n12511_), .ZN(new_n12536_));
  AOI21_X1   g12279(.A1(new_n12503_), .A2(new_n12506_), .B(new_n12512_), .ZN(new_n12537_));
  OAI21_X1   g12280(.A1(new_n12537_), .A2(new_n12536_), .B(new_n12351_), .ZN(new_n12538_));
  AOI21_X1   g12281(.A1(new_n12503_), .A2(new_n12506_), .B(new_n12511_), .ZN(new_n12539_));
  NOR3_X1    g12282(.A1(new_n12516_), .A2(new_n12519_), .A3(new_n12512_), .ZN(new_n12540_));
  OAI21_X1   g12283(.A1(new_n12539_), .A2(new_n12540_), .B(new_n12352_), .ZN(new_n12541_));
  AOI21_X1   g12284(.A1(new_n12538_), .A2(new_n12541_), .B(new_n12530_), .ZN(new_n12542_));
  OAI21_X1   g12285(.A1(new_n12535_), .A2(new_n12542_), .B(new_n12347_), .ZN(new_n12543_));
  OAI21_X1   g12286(.A1(new_n12534_), .A2(new_n12347_), .B(new_n12543_), .ZN(new_n12544_));
  OAI22_X1   g12287(.A1(new_n2084_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n2079_), .ZN(new_n12545_));
  NAND2_X1   g12288(.A1(new_n2864_), .A2(\b[43] ), .ZN(new_n12546_));
  AOI21_X1   g12289(.A1(new_n12545_), .A2(new_n12546_), .B(new_n2087_), .ZN(new_n12547_));
  NAND2_X1   g12290(.A1(new_n4513_), .A2(new_n12547_), .ZN(new_n12548_));
  XOR2_X1    g12291(.A1(new_n12548_), .A2(\a[29] ), .Z(new_n12549_));
  INV_X1     g12292(.I(new_n12549_), .ZN(new_n12550_));
  NOR2_X1    g12293(.A1(new_n12208_), .A2(new_n12203_), .ZN(new_n12551_));
  INV_X1     g12294(.I(new_n12551_), .ZN(new_n12552_));
  NOR2_X1    g12295(.A1(new_n12193_), .A2(new_n12197_), .ZN(new_n12553_));
  XOR2_X1    g12296(.A1(new_n11993_), .A2(new_n12203_), .Z(new_n12554_));
  INV_X1     g12297(.I(new_n12554_), .ZN(new_n12555_));
  NAND2_X1   g12298(.A1(new_n12553_), .A2(new_n12555_), .ZN(new_n12556_));
  AOI21_X1   g12299(.A1(new_n12556_), .A2(new_n12552_), .B(new_n12550_), .ZN(new_n12557_));
  INV_X1     g12300(.I(new_n12557_), .ZN(new_n12558_));
  NAND3_X1   g12301(.A1(new_n12556_), .A2(new_n12552_), .A3(new_n12550_), .ZN(new_n12559_));
  AOI21_X1   g12302(.A1(new_n12558_), .A2(new_n12559_), .B(new_n12544_), .ZN(new_n12560_));
  NAND3_X1   g12303(.A1(new_n12558_), .A2(new_n12544_), .A3(new_n12559_), .ZN(new_n12561_));
  INV_X1     g12304(.I(new_n12561_), .ZN(new_n12562_));
  OAI22_X1   g12305(.A1(new_n1760_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n1755_), .ZN(new_n12563_));
  NAND2_X1   g12306(.A1(new_n2470_), .A2(\b[46] ), .ZN(new_n12564_));
  AOI21_X1   g12307(.A1(new_n12563_), .A2(new_n12564_), .B(new_n1763_), .ZN(new_n12565_));
  NAND2_X1   g12308(.A1(new_n5177_), .A2(new_n12565_), .ZN(new_n12566_));
  XOR2_X1    g12309(.A1(new_n12566_), .A2(\a[26] ), .Z(new_n12567_));
  INV_X1     g12310(.I(new_n12567_), .ZN(new_n12568_));
  OAI21_X1   g12311(.A1(new_n12562_), .A2(new_n12560_), .B(new_n12568_), .ZN(new_n12569_));
  INV_X1     g12312(.I(new_n12560_), .ZN(new_n12570_));
  NAND3_X1   g12313(.A1(new_n12570_), .A2(new_n12561_), .A3(new_n12567_), .ZN(new_n12571_));
  AOI21_X1   g12314(.A1(new_n12571_), .A2(new_n12569_), .B(new_n12345_), .ZN(new_n12572_));
  INV_X1     g12315(.I(new_n12345_), .ZN(new_n12573_));
  NAND3_X1   g12316(.A1(new_n12570_), .A2(new_n12561_), .A3(new_n12568_), .ZN(new_n12574_));
  OAI21_X1   g12317(.A1(new_n12562_), .A2(new_n12560_), .B(new_n12567_), .ZN(new_n12575_));
  AOI21_X1   g12318(.A1(new_n12574_), .A2(new_n12575_), .B(new_n12573_), .ZN(new_n12576_));
  OAI22_X1   g12319(.A1(new_n1444_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n1439_), .ZN(new_n12577_));
  NAND2_X1   g12320(.A1(new_n2098_), .A2(\b[49] ), .ZN(new_n12578_));
  AOI21_X1   g12321(.A1(new_n12577_), .A2(new_n12578_), .B(new_n1447_), .ZN(new_n12579_));
  NAND2_X1   g12322(.A1(new_n5741_), .A2(new_n12579_), .ZN(new_n12580_));
  XOR2_X1    g12323(.A1(new_n12580_), .A2(\a[23] ), .Z(new_n12581_));
  INV_X1     g12324(.I(new_n12581_), .ZN(new_n12582_));
  OAI21_X1   g12325(.A1(new_n12572_), .A2(new_n12576_), .B(new_n12582_), .ZN(new_n12583_));
  AOI21_X1   g12326(.A1(new_n12570_), .A2(new_n12561_), .B(new_n12567_), .ZN(new_n12584_));
  NOR3_X1    g12327(.A1(new_n12562_), .A2(new_n12560_), .A3(new_n12568_), .ZN(new_n12585_));
  OAI21_X1   g12328(.A1(new_n12584_), .A2(new_n12585_), .B(new_n12573_), .ZN(new_n12586_));
  NOR3_X1    g12329(.A1(new_n12562_), .A2(new_n12560_), .A3(new_n12567_), .ZN(new_n12587_));
  AOI21_X1   g12330(.A1(new_n12570_), .A2(new_n12561_), .B(new_n12568_), .ZN(new_n12588_));
  OAI21_X1   g12331(.A1(new_n12588_), .A2(new_n12587_), .B(new_n12345_), .ZN(new_n12589_));
  NAND3_X1   g12332(.A1(new_n12586_), .A2(new_n12589_), .A3(new_n12581_), .ZN(new_n12590_));
  AOI21_X1   g12333(.A1(new_n12583_), .A2(new_n12590_), .B(new_n12344_), .ZN(new_n12591_));
  INV_X1     g12334(.I(new_n12344_), .ZN(new_n12592_));
  NAND3_X1   g12335(.A1(new_n12586_), .A2(new_n12589_), .A3(new_n12582_), .ZN(new_n12593_));
  OAI21_X1   g12336(.A1(new_n12572_), .A2(new_n12576_), .B(new_n12581_), .ZN(new_n12594_));
  AOI21_X1   g12337(.A1(new_n12594_), .A2(new_n12593_), .B(new_n12592_), .ZN(new_n12595_));
  OAI22_X1   g12338(.A1(new_n1168_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n1163_), .ZN(new_n12596_));
  NAND2_X1   g12339(.A1(new_n1774_), .A2(\b[52] ), .ZN(new_n12597_));
  AOI21_X1   g12340(.A1(new_n12596_), .A2(new_n12597_), .B(new_n1171_), .ZN(new_n12598_));
  NAND2_X1   g12341(.A1(new_n6237_), .A2(new_n12598_), .ZN(new_n12599_));
  XOR2_X1    g12342(.A1(new_n12599_), .A2(\a[20] ), .Z(new_n12600_));
  INV_X1     g12343(.I(new_n12600_), .ZN(new_n12601_));
  OAI21_X1   g12344(.A1(new_n12591_), .A2(new_n12595_), .B(new_n12601_), .ZN(new_n12602_));
  AOI21_X1   g12345(.A1(new_n12586_), .A2(new_n12589_), .B(new_n12581_), .ZN(new_n12603_));
  NOR3_X1    g12346(.A1(new_n12572_), .A2(new_n12576_), .A3(new_n12582_), .ZN(new_n12604_));
  OAI21_X1   g12347(.A1(new_n12603_), .A2(new_n12604_), .B(new_n12592_), .ZN(new_n12605_));
  NOR3_X1    g12348(.A1(new_n12572_), .A2(new_n12576_), .A3(new_n12581_), .ZN(new_n12606_));
  AOI21_X1   g12349(.A1(new_n12586_), .A2(new_n12589_), .B(new_n12582_), .ZN(new_n12607_));
  OAI21_X1   g12350(.A1(new_n12607_), .A2(new_n12606_), .B(new_n12344_), .ZN(new_n12608_));
  NAND3_X1   g12351(.A1(new_n12605_), .A2(new_n12608_), .A3(new_n12600_), .ZN(new_n12609_));
  AOI21_X1   g12352(.A1(new_n12602_), .A2(new_n12609_), .B(new_n12343_), .ZN(new_n12610_));
  INV_X1     g12353(.I(new_n12343_), .ZN(new_n12611_));
  NAND3_X1   g12354(.A1(new_n12605_), .A2(new_n12608_), .A3(new_n12601_), .ZN(new_n12612_));
  OAI21_X1   g12355(.A1(new_n12591_), .A2(new_n12595_), .B(new_n12600_), .ZN(new_n12613_));
  AOI21_X1   g12356(.A1(new_n12613_), .A2(new_n12612_), .B(new_n12611_), .ZN(new_n12614_));
  OAI22_X1   g12357(.A1(new_n940_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n935_), .ZN(new_n12615_));
  NAND2_X1   g12358(.A1(new_n1458_), .A2(\b[55] ), .ZN(new_n12616_));
  AOI21_X1   g12359(.A1(new_n12615_), .A2(new_n12616_), .B(new_n943_), .ZN(new_n12617_));
  NAND2_X1   g12360(.A1(new_n7308_), .A2(new_n12617_), .ZN(new_n12618_));
  XOR2_X1    g12361(.A1(new_n12618_), .A2(\a[17] ), .Z(new_n12619_));
  NOR3_X1    g12362(.A1(new_n12610_), .A2(new_n12614_), .A3(new_n12619_), .ZN(new_n12620_));
  AOI21_X1   g12363(.A1(new_n12605_), .A2(new_n12608_), .B(new_n12600_), .ZN(new_n12621_));
  NOR3_X1    g12364(.A1(new_n12591_), .A2(new_n12595_), .A3(new_n12601_), .ZN(new_n12622_));
  OAI21_X1   g12365(.A1(new_n12621_), .A2(new_n12622_), .B(new_n12611_), .ZN(new_n12623_));
  NOR3_X1    g12366(.A1(new_n12591_), .A2(new_n12595_), .A3(new_n12600_), .ZN(new_n12624_));
  AOI21_X1   g12367(.A1(new_n12605_), .A2(new_n12608_), .B(new_n12601_), .ZN(new_n12625_));
  OAI21_X1   g12368(.A1(new_n12625_), .A2(new_n12624_), .B(new_n12343_), .ZN(new_n12626_));
  INV_X1     g12369(.I(new_n12619_), .ZN(new_n12627_));
  AOI21_X1   g12370(.A1(new_n12623_), .A2(new_n12626_), .B(new_n12627_), .ZN(new_n12628_));
  OAI21_X1   g12371(.A1(new_n12628_), .A2(new_n12620_), .B(new_n12342_), .ZN(new_n12629_));
  AOI21_X1   g12372(.A1(new_n12623_), .A2(new_n12626_), .B(new_n12619_), .ZN(new_n12630_));
  NOR3_X1    g12373(.A1(new_n12610_), .A2(new_n12614_), .A3(new_n12627_), .ZN(new_n12631_));
  OAI21_X1   g12374(.A1(new_n12630_), .A2(new_n12631_), .B(new_n12341_), .ZN(new_n12632_));
  OAI22_X1   g12375(.A1(new_n757_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n752_), .ZN(new_n12633_));
  NAND2_X1   g12376(.A1(new_n1182_), .A2(\b[58] ), .ZN(new_n12634_));
  AOI21_X1   g12377(.A1(new_n12633_), .A2(new_n12634_), .B(new_n760_), .ZN(new_n12635_));
  NAND2_X1   g12378(.A1(new_n7929_), .A2(new_n12635_), .ZN(new_n12636_));
  XOR2_X1    g12379(.A1(new_n12636_), .A2(\a[14] ), .Z(new_n12637_));
  INV_X1     g12380(.I(new_n12637_), .ZN(new_n12638_));
  NAND3_X1   g12381(.A1(new_n12629_), .A2(new_n12632_), .A3(new_n12638_), .ZN(new_n12639_));
  NAND3_X1   g12382(.A1(new_n12623_), .A2(new_n12626_), .A3(new_n12627_), .ZN(new_n12640_));
  OAI21_X1   g12383(.A1(new_n12610_), .A2(new_n12614_), .B(new_n12619_), .ZN(new_n12641_));
  AOI21_X1   g12384(.A1(new_n12641_), .A2(new_n12640_), .B(new_n12341_), .ZN(new_n12642_));
  OAI21_X1   g12385(.A1(new_n12610_), .A2(new_n12614_), .B(new_n12627_), .ZN(new_n12643_));
  NAND3_X1   g12386(.A1(new_n12623_), .A2(new_n12626_), .A3(new_n12619_), .ZN(new_n12644_));
  AOI21_X1   g12387(.A1(new_n12643_), .A2(new_n12644_), .B(new_n12342_), .ZN(new_n12645_));
  OAI21_X1   g12388(.A1(new_n12642_), .A2(new_n12645_), .B(new_n12637_), .ZN(new_n12646_));
  AOI21_X1   g12389(.A1(new_n12646_), .A2(new_n12639_), .B(new_n12340_), .ZN(new_n12647_));
  NAND2_X1   g12390(.A1(new_n12339_), .A2(new_n12292_), .ZN(new_n12648_));
  OAI21_X1   g12391(.A1(new_n12642_), .A2(new_n12645_), .B(new_n12638_), .ZN(new_n12649_));
  NAND3_X1   g12392(.A1(new_n12629_), .A2(new_n12632_), .A3(new_n12637_), .ZN(new_n12650_));
  AOI21_X1   g12393(.A1(new_n12649_), .A2(new_n12650_), .B(new_n12648_), .ZN(new_n12651_));
  NOR2_X1    g12394(.A1(new_n12647_), .A2(new_n12651_), .ZN(new_n12652_));
  OAI22_X1   g12395(.A1(new_n582_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n577_), .ZN(new_n12653_));
  NAND2_X1   g12396(.A1(new_n960_), .A2(\b[61] ), .ZN(new_n12654_));
  AOI21_X1   g12397(.A1(new_n12653_), .A2(new_n12654_), .B(new_n585_), .ZN(new_n12655_));
  NAND2_X1   g12398(.A1(new_n8963_), .A2(new_n12655_), .ZN(new_n12656_));
  XOR2_X1    g12399(.A1(new_n12656_), .A2(\a[11] ), .Z(new_n12657_));
  NOR2_X1    g12400(.A1(new_n12652_), .A2(new_n12657_), .ZN(new_n12658_));
  INV_X1     g12401(.I(new_n12657_), .ZN(new_n12659_));
  NOR3_X1    g12402(.A1(new_n12647_), .A2(new_n12651_), .A3(new_n12659_), .ZN(new_n12660_));
  OAI21_X1   g12403(.A1(new_n12658_), .A2(new_n12660_), .B(new_n12338_), .ZN(new_n12661_));
  XOR2_X1    g12404(.A1(new_n12652_), .A2(new_n12659_), .Z(new_n12662_));
  OAI21_X1   g12405(.A1(new_n12662_), .A2(new_n12338_), .B(new_n12661_), .ZN(new_n12663_));
  XNOR2_X1   g12406(.A1(new_n12663_), .A2(new_n12336_), .ZN(new_n12664_));
  XOR2_X1    g12407(.A1(new_n11977_), .A2(new_n11980_), .Z(new_n12665_));
  NAND2_X1   g12408(.A1(new_n12665_), .A2(new_n12326_), .ZN(new_n12666_));
  XNOR2_X1   g12409(.A1(new_n12666_), .A2(new_n12664_), .ZN(new_n12667_));
  NOR2_X1    g12410(.A1(new_n11977_), .A2(new_n11980_), .ZN(new_n12668_));
  XOR2_X1    g12411(.A1(new_n12667_), .A2(new_n12668_), .Z(\f[72] ));
  INV_X1     g12412(.I(new_n12660_), .ZN(new_n12670_));
  AOI21_X1   g12413(.A1(new_n12338_), .A2(new_n12670_), .B(new_n12658_), .ZN(new_n12671_));
  NAND2_X1   g12414(.A1(new_n12646_), .A2(new_n12648_), .ZN(new_n12672_));
  AND2_X2    g12415(.A1(new_n12672_), .A2(new_n12639_), .Z(new_n12673_));
  AOI21_X1   g12416(.A1(new_n12342_), .A2(new_n12644_), .B(new_n12630_), .ZN(new_n12674_));
  INV_X1     g12417(.I(new_n12674_), .ZN(new_n12675_));
  AOI21_X1   g12418(.A1(new_n12611_), .A2(new_n12609_), .B(new_n12621_), .ZN(new_n12676_));
  AOI21_X1   g12419(.A1(new_n12592_), .A2(new_n12590_), .B(new_n12603_), .ZN(new_n12677_));
  OAI22_X1   g12420(.A1(new_n1444_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n1439_), .ZN(new_n12678_));
  OAI21_X1   g12421(.A1(new_n5538_), .A2(new_n1548_), .B(new_n12678_), .ZN(new_n12679_));
  AOI21_X1   g12422(.A1(new_n5954_), .A2(new_n1446_), .B(new_n12679_), .ZN(new_n12680_));
  INV_X1     g12423(.I(new_n12680_), .ZN(new_n12681_));
  AOI21_X1   g12424(.A1(new_n12573_), .A2(new_n12571_), .B(new_n12584_), .ZN(new_n12682_));
  NAND2_X1   g12425(.A1(new_n12556_), .A2(new_n12552_), .ZN(new_n12683_));
  INV_X1     g12426(.I(new_n12683_), .ZN(new_n12684_));
  XOR2_X1    g12427(.A1(new_n12544_), .A2(new_n12550_), .Z(new_n12685_));
  OAI21_X1   g12428(.A1(new_n12549_), .A2(new_n12684_), .B(new_n12685_), .ZN(new_n12686_));
  OAI22_X1   g12429(.A1(new_n2084_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n2079_), .ZN(new_n12687_));
  OAI21_X1   g12430(.A1(new_n4501_), .A2(new_n2214_), .B(new_n12687_), .ZN(new_n12688_));
  AOI21_X1   g12431(.A1(new_n4833_), .A2(new_n2086_), .B(new_n12688_), .ZN(new_n12689_));
  INV_X1     g12432(.I(new_n12689_), .ZN(new_n12690_));
  NOR2_X1    g12433(.A1(new_n12347_), .A2(new_n12533_), .ZN(new_n12691_));
  AOI21_X1   g12434(.A1(new_n12351_), .A2(new_n12520_), .B(new_n12536_), .ZN(new_n12692_));
  AOI21_X1   g12435(.A1(new_n12354_), .A2(new_n12518_), .B(new_n12504_), .ZN(new_n12693_));
  AOI21_X1   g12436(.A1(new_n12485_), .A2(new_n12483_), .B(new_n12495_), .ZN(new_n12694_));
  INV_X1     g12437(.I(new_n12694_), .ZN(new_n12695_));
  AOI21_X1   g12438(.A1(new_n12466_), .A2(new_n12464_), .B(new_n12462_), .ZN(new_n12696_));
  INV_X1     g12439(.I(new_n12696_), .ZN(new_n12697_));
  OAI22_X1   g12440(.A1(new_n3736_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n3731_), .ZN(new_n12698_));
  NAND2_X1   g12441(.A1(new_n4730_), .A2(\b[32] ), .ZN(new_n12699_));
  AOI21_X1   g12442(.A1(new_n12698_), .A2(new_n12699_), .B(new_n3739_), .ZN(new_n12700_));
  NAND2_X1   g12443(.A1(new_n2963_), .A2(new_n12700_), .ZN(new_n12701_));
  XOR2_X1    g12444(.A1(new_n12701_), .A2(\a[41] ), .Z(new_n12702_));
  OAI22_X1   g12445(.A1(new_n4711_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n4706_), .ZN(new_n12703_));
  NAND2_X1   g12446(.A1(new_n5814_), .A2(\b[26] ), .ZN(new_n12704_));
  AOI21_X1   g12447(.A1(new_n12703_), .A2(new_n12704_), .B(new_n4714_), .ZN(new_n12705_));
  NAND2_X1   g12448(.A1(new_n2174_), .A2(new_n12705_), .ZN(new_n12706_));
  XOR2_X1    g12449(.A1(new_n12706_), .A2(\a[47] ), .Z(new_n12707_));
  OAI22_X1   g12450(.A1(new_n5786_), .A2(new_n1518_), .B1(new_n1393_), .B2(new_n5792_), .ZN(new_n12708_));
  NAND2_X1   g12451(.A1(new_n6745_), .A2(\b[20] ), .ZN(new_n12709_));
  AOI21_X1   g12452(.A1(new_n12709_), .A2(new_n12708_), .B(new_n5796_), .ZN(new_n12710_));
  NAND2_X1   g12453(.A1(new_n1517_), .A2(new_n12710_), .ZN(new_n12711_));
  XOR2_X1    g12454(.A1(new_n12711_), .A2(\a[53] ), .Z(new_n12712_));
  OAI21_X1   g12455(.A1(new_n12370_), .A2(new_n12386_), .B(new_n12387_), .ZN(new_n12713_));
  INV_X1     g12456(.I(new_n12713_), .ZN(new_n12714_));
  OAI22_X1   g12457(.A1(new_n992_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n904_), .ZN(new_n12715_));
  NAND2_X1   g12458(.A1(new_n8628_), .A2(\b[14] ), .ZN(new_n12716_));
  AOI21_X1   g12459(.A1(new_n12716_), .A2(new_n12715_), .B(new_n7354_), .ZN(new_n12717_));
  NAND2_X1   g12460(.A1(new_n991_), .A2(new_n12717_), .ZN(new_n12718_));
  XOR2_X1    g12461(.A1(new_n12718_), .A2(\a[59] ), .Z(new_n12719_));
  OAI22_X1   g12462(.A1(new_n795_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n717_), .ZN(new_n12720_));
  NAND2_X1   g12463(.A1(new_n9644_), .A2(\b[11] ), .ZN(new_n12721_));
  AOI21_X1   g12464(.A1(new_n12721_), .A2(new_n12720_), .B(new_n8321_), .ZN(new_n12722_));
  NAND2_X1   g12465(.A1(new_n799_), .A2(new_n12722_), .ZN(new_n12723_));
  XOR2_X1    g12466(.A1(new_n12723_), .A2(new_n8309_), .Z(new_n12724_));
  NAND2_X1   g12467(.A1(new_n12383_), .A2(new_n12041_), .ZN(new_n12725_));
  NAND2_X1   g12468(.A1(new_n12725_), .A2(new_n12382_), .ZN(new_n12726_));
  NOR3_X1    g12469(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n510_), .ZN(new_n12727_));
  NOR2_X1    g12470(.A1(new_n9364_), .A2(new_n510_), .ZN(new_n12728_));
  NOR3_X1    g12471(.A1(new_n12728_), .A2(new_n617_), .A3(new_n8985_), .ZN(new_n12729_));
  NOR2_X1    g12472(.A1(new_n12729_), .A2(new_n12727_), .ZN(new_n12730_));
  NOR2_X1    g12473(.A1(new_n12726_), .A2(new_n12730_), .ZN(new_n12731_));
  INV_X1     g12474(.I(new_n12731_), .ZN(new_n12732_));
  NAND2_X1   g12475(.A1(new_n12726_), .A2(new_n12730_), .ZN(new_n12733_));
  NAND2_X1   g12476(.A1(new_n12732_), .A2(new_n12733_), .ZN(new_n12734_));
  INV_X1     g12477(.I(new_n12730_), .ZN(new_n12735_));
  XOR2_X1    g12478(.A1(new_n12726_), .A2(new_n12735_), .Z(new_n12736_));
  NOR2_X1    g12479(.A1(new_n12724_), .A2(new_n12736_), .ZN(new_n12737_));
  AOI21_X1   g12480(.A1(new_n12724_), .A2(new_n12734_), .B(new_n12737_), .ZN(new_n12738_));
  NOR2_X1    g12481(.A1(new_n12738_), .A2(new_n12719_), .ZN(new_n12739_));
  INV_X1     g12482(.I(new_n12739_), .ZN(new_n12740_));
  NAND2_X1   g12483(.A1(new_n12738_), .A2(new_n12719_), .ZN(new_n12741_));
  AOI21_X1   g12484(.A1(new_n12740_), .A2(new_n12741_), .B(new_n12714_), .ZN(new_n12742_));
  XNOR2_X1   g12485(.A1(new_n12738_), .A2(new_n12719_), .ZN(new_n12743_));
  NOR2_X1    g12486(.A1(new_n12743_), .A2(new_n12713_), .ZN(new_n12744_));
  NOR2_X1    g12487(.A1(new_n12744_), .A2(new_n12742_), .ZN(new_n12745_));
  OAI21_X1   g12488(.A1(new_n12368_), .A2(new_n12402_), .B(new_n12401_), .ZN(new_n12746_));
  INV_X1     g12489(.I(new_n12746_), .ZN(new_n12747_));
  OAI22_X1   g12490(.A1(new_n6721_), .A2(new_n1124_), .B1(new_n6723_), .B2(new_n1222_), .ZN(new_n12748_));
  NAND2_X1   g12491(.A1(new_n7617_), .A2(\b[17] ), .ZN(new_n12749_));
  AOI21_X1   g12492(.A1(new_n12749_), .A2(new_n12748_), .B(new_n6731_), .ZN(new_n12750_));
  NAND2_X1   g12493(.A1(new_n1225_), .A2(new_n12750_), .ZN(new_n12751_));
  XOR2_X1    g12494(.A1(new_n12751_), .A2(\a[56] ), .Z(new_n12752_));
  NOR2_X1    g12495(.A1(new_n12752_), .A2(new_n12747_), .ZN(new_n12753_));
  INV_X1     g12496(.I(new_n12753_), .ZN(new_n12754_));
  NAND2_X1   g12497(.A1(new_n12752_), .A2(new_n12747_), .ZN(new_n12755_));
  AOI21_X1   g12498(.A1(new_n12754_), .A2(new_n12755_), .B(new_n12745_), .ZN(new_n12756_));
  XOR2_X1    g12499(.A1(new_n12752_), .A2(new_n12747_), .Z(new_n12757_));
  AOI21_X1   g12500(.A1(new_n12745_), .A2(new_n12757_), .B(new_n12756_), .ZN(new_n12758_));
  NAND2_X1   g12501(.A1(new_n12415_), .A2(new_n12405_), .ZN(new_n12759_));
  NAND2_X1   g12502(.A1(new_n12759_), .A2(new_n12413_), .ZN(new_n12760_));
  INV_X1     g12503(.I(new_n12760_), .ZN(new_n12761_));
  NOR2_X1    g12504(.A1(new_n12758_), .A2(new_n12761_), .ZN(new_n12762_));
  INV_X1     g12505(.I(new_n12762_), .ZN(new_n12763_));
  NAND2_X1   g12506(.A1(new_n12758_), .A2(new_n12761_), .ZN(new_n12764_));
  AOI21_X1   g12507(.A1(new_n12763_), .A2(new_n12764_), .B(new_n12712_), .ZN(new_n12765_));
  INV_X1     g12508(.I(new_n12712_), .ZN(new_n12766_));
  XOR2_X1    g12509(.A1(new_n12758_), .A2(new_n12760_), .Z(new_n12767_));
  NOR2_X1    g12510(.A1(new_n12767_), .A2(new_n12766_), .ZN(new_n12768_));
  NOR2_X1    g12511(.A1(new_n12768_), .A2(new_n12765_), .ZN(new_n12769_));
  INV_X1     g12512(.I(new_n12429_), .ZN(new_n12770_));
  AOI21_X1   g12513(.A1(new_n12430_), .A2(new_n12424_), .B(new_n12367_), .ZN(new_n12771_));
  NOR2_X1    g12514(.A1(new_n12771_), .A2(new_n12770_), .ZN(new_n12772_));
  OAI22_X1   g12515(.A1(new_n5228_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n5225_), .ZN(new_n12773_));
  NAND2_X1   g12516(.A1(new_n5387_), .A2(\b[23] ), .ZN(new_n12774_));
  AOI21_X1   g12517(.A1(new_n12773_), .A2(new_n12774_), .B(new_n5231_), .ZN(new_n12775_));
  NAND2_X1   g12518(.A1(new_n1828_), .A2(new_n12775_), .ZN(new_n12776_));
  XOR2_X1    g12519(.A1(new_n12776_), .A2(\a[50] ), .Z(new_n12777_));
  NOR2_X1    g12520(.A1(new_n12772_), .A2(new_n12777_), .ZN(new_n12778_));
  INV_X1     g12521(.I(new_n12778_), .ZN(new_n12779_));
  NAND2_X1   g12522(.A1(new_n12772_), .A2(new_n12777_), .ZN(new_n12780_));
  AOI21_X1   g12523(.A1(new_n12779_), .A2(new_n12780_), .B(new_n12769_), .ZN(new_n12781_));
  XNOR2_X1   g12524(.A1(new_n12772_), .A2(new_n12777_), .ZN(new_n12782_));
  NOR3_X1    g12525(.A1(new_n12782_), .A2(new_n12765_), .A3(new_n12768_), .ZN(new_n12783_));
  NOR2_X1    g12526(.A1(new_n12783_), .A2(new_n12781_), .ZN(new_n12784_));
  OAI21_X1   g12527(.A1(new_n12359_), .A2(new_n12434_), .B(new_n12435_), .ZN(new_n12785_));
  INV_X1     g12528(.I(new_n12785_), .ZN(new_n12786_));
  NOR2_X1    g12529(.A1(new_n12784_), .A2(new_n12786_), .ZN(new_n12787_));
  INV_X1     g12530(.I(new_n12787_), .ZN(new_n12788_));
  NAND2_X1   g12531(.A1(new_n12784_), .A2(new_n12786_), .ZN(new_n12789_));
  AOI21_X1   g12532(.A1(new_n12788_), .A2(new_n12789_), .B(new_n12707_), .ZN(new_n12790_));
  INV_X1     g12533(.I(new_n12707_), .ZN(new_n12791_));
  XOR2_X1    g12534(.A1(new_n12784_), .A2(new_n12785_), .Z(new_n12792_));
  NOR2_X1    g12535(.A1(new_n12792_), .A2(new_n12791_), .ZN(new_n12793_));
  NOR2_X1    g12536(.A1(new_n12793_), .A2(new_n12790_), .ZN(new_n12794_));
  AOI21_X1   g12537(.A1(new_n12452_), .A2(new_n12455_), .B(new_n12453_), .ZN(new_n12795_));
  OAI22_X1   g12538(.A1(new_n4208_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n4203_), .ZN(new_n12796_));
  NAND2_X1   g12539(.A1(new_n5244_), .A2(\b[29] ), .ZN(new_n12797_));
  AOI21_X1   g12540(.A1(new_n12796_), .A2(new_n12797_), .B(new_n4211_), .ZN(new_n12798_));
  NAND2_X1   g12541(.A1(new_n2546_), .A2(new_n12798_), .ZN(new_n12799_));
  XOR2_X1    g12542(.A1(new_n12799_), .A2(\a[44] ), .Z(new_n12800_));
  INV_X1     g12543(.I(new_n12800_), .ZN(new_n12801_));
  XOR2_X1    g12544(.A1(new_n12795_), .A2(new_n12801_), .Z(new_n12802_));
  NOR2_X1    g12545(.A1(new_n12802_), .A2(new_n12794_), .ZN(new_n12803_));
  INV_X1     g12546(.I(new_n12803_), .ZN(new_n12804_));
  NOR2_X1    g12547(.A1(new_n12795_), .A2(new_n12800_), .ZN(new_n12805_));
  NAND2_X1   g12548(.A1(new_n12795_), .A2(new_n12800_), .ZN(new_n12806_));
  INV_X1     g12549(.I(new_n12806_), .ZN(new_n12807_));
  OAI21_X1   g12550(.A1(new_n12805_), .A2(new_n12807_), .B(new_n12794_), .ZN(new_n12808_));
  AOI21_X1   g12551(.A1(new_n12804_), .A2(new_n12808_), .B(new_n12702_), .ZN(new_n12809_));
  INV_X1     g12552(.I(new_n12702_), .ZN(new_n12810_));
  INV_X1     g12553(.I(new_n12808_), .ZN(new_n12811_));
  NOR3_X1    g12554(.A1(new_n12811_), .A2(new_n12803_), .A3(new_n12810_), .ZN(new_n12812_));
  OAI21_X1   g12555(.A1(new_n12809_), .A2(new_n12812_), .B(new_n12697_), .ZN(new_n12813_));
  AOI21_X1   g12556(.A1(new_n12804_), .A2(new_n12808_), .B(new_n12810_), .ZN(new_n12814_));
  NOR3_X1    g12557(.A1(new_n12811_), .A2(new_n12803_), .A3(new_n12702_), .ZN(new_n12815_));
  OAI21_X1   g12558(.A1(new_n12814_), .A2(new_n12815_), .B(new_n12696_), .ZN(new_n12816_));
  OAI22_X1   g12559(.A1(new_n3298_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n3293_), .ZN(new_n12817_));
  NAND2_X1   g12560(.A1(new_n4227_), .A2(\b[35] ), .ZN(new_n12818_));
  AOI21_X1   g12561(.A1(new_n12817_), .A2(new_n12818_), .B(new_n3301_), .ZN(new_n12819_));
  NAND2_X1   g12562(.A1(new_n3411_), .A2(new_n12819_), .ZN(new_n12820_));
  XOR2_X1    g12563(.A1(new_n12820_), .A2(\a[38] ), .Z(new_n12821_));
  AOI21_X1   g12564(.A1(new_n12813_), .A2(new_n12816_), .B(new_n12821_), .ZN(new_n12822_));
  OAI21_X1   g12565(.A1(new_n12811_), .A2(new_n12803_), .B(new_n12810_), .ZN(new_n12823_));
  NAND3_X1   g12566(.A1(new_n12804_), .A2(new_n12702_), .A3(new_n12808_), .ZN(new_n12824_));
  AOI21_X1   g12567(.A1(new_n12823_), .A2(new_n12824_), .B(new_n12696_), .ZN(new_n12825_));
  OAI21_X1   g12568(.A1(new_n12811_), .A2(new_n12803_), .B(new_n12702_), .ZN(new_n12826_));
  NAND3_X1   g12569(.A1(new_n12804_), .A2(new_n12810_), .A3(new_n12808_), .ZN(new_n12827_));
  AOI21_X1   g12570(.A1(new_n12826_), .A2(new_n12827_), .B(new_n12697_), .ZN(new_n12828_));
  INV_X1     g12571(.I(new_n12821_), .ZN(new_n12829_));
  NOR3_X1    g12572(.A1(new_n12825_), .A2(new_n12828_), .A3(new_n12829_), .ZN(new_n12830_));
  OAI21_X1   g12573(.A1(new_n12822_), .A2(new_n12830_), .B(new_n12695_), .ZN(new_n12831_));
  NOR3_X1    g12574(.A1(new_n12825_), .A2(new_n12828_), .A3(new_n12821_), .ZN(new_n12832_));
  AOI21_X1   g12575(.A1(new_n12813_), .A2(new_n12816_), .B(new_n12829_), .ZN(new_n12833_));
  OAI21_X1   g12576(.A1(new_n12833_), .A2(new_n12832_), .B(new_n12694_), .ZN(new_n12834_));
  OAI22_X1   g12577(.A1(new_n2846_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n2841_), .ZN(new_n12835_));
  NAND2_X1   g12578(.A1(new_n3755_), .A2(\b[38] ), .ZN(new_n12836_));
  AOI21_X1   g12579(.A1(new_n12835_), .A2(new_n12836_), .B(new_n2849_), .ZN(new_n12837_));
  NAND2_X1   g12580(.A1(new_n3844_), .A2(new_n12837_), .ZN(new_n12838_));
  XOR2_X1    g12581(.A1(new_n12838_), .A2(\a[35] ), .Z(new_n12839_));
  INV_X1     g12582(.I(new_n12839_), .ZN(new_n12840_));
  NAND3_X1   g12583(.A1(new_n12831_), .A2(new_n12834_), .A3(new_n12840_), .ZN(new_n12841_));
  OAI21_X1   g12584(.A1(new_n12825_), .A2(new_n12828_), .B(new_n12829_), .ZN(new_n12842_));
  NAND3_X1   g12585(.A1(new_n12813_), .A2(new_n12816_), .A3(new_n12821_), .ZN(new_n12843_));
  AOI21_X1   g12586(.A1(new_n12842_), .A2(new_n12843_), .B(new_n12694_), .ZN(new_n12844_));
  NAND3_X1   g12587(.A1(new_n12813_), .A2(new_n12816_), .A3(new_n12829_), .ZN(new_n12845_));
  OAI21_X1   g12588(.A1(new_n12825_), .A2(new_n12828_), .B(new_n12821_), .ZN(new_n12846_));
  AOI21_X1   g12589(.A1(new_n12846_), .A2(new_n12845_), .B(new_n12695_), .ZN(new_n12847_));
  OAI21_X1   g12590(.A1(new_n12844_), .A2(new_n12847_), .B(new_n12839_), .ZN(new_n12848_));
  AOI21_X1   g12591(.A1(new_n12848_), .A2(new_n12841_), .B(new_n12693_), .ZN(new_n12849_));
  INV_X1     g12592(.I(new_n12693_), .ZN(new_n12850_));
  OAI21_X1   g12593(.A1(new_n12844_), .A2(new_n12847_), .B(new_n12840_), .ZN(new_n12851_));
  NAND3_X1   g12594(.A1(new_n12831_), .A2(new_n12834_), .A3(new_n12839_), .ZN(new_n12852_));
  AOI21_X1   g12595(.A1(new_n12851_), .A2(new_n12852_), .B(new_n12850_), .ZN(new_n12853_));
  OAI22_X1   g12596(.A1(new_n2452_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n2447_), .ZN(new_n12854_));
  NAND2_X1   g12597(.A1(new_n3312_), .A2(\b[41] ), .ZN(new_n12855_));
  AOI21_X1   g12598(.A1(new_n12854_), .A2(new_n12855_), .B(new_n2455_), .ZN(new_n12856_));
  NAND2_X1   g12599(.A1(new_n4320_), .A2(new_n12856_), .ZN(new_n12857_));
  XOR2_X1    g12600(.A1(new_n12857_), .A2(\a[32] ), .Z(new_n12858_));
  INV_X1     g12601(.I(new_n12858_), .ZN(new_n12859_));
  OAI21_X1   g12602(.A1(new_n12849_), .A2(new_n12853_), .B(new_n12859_), .ZN(new_n12860_));
  NOR3_X1    g12603(.A1(new_n12844_), .A2(new_n12847_), .A3(new_n12839_), .ZN(new_n12861_));
  AOI21_X1   g12604(.A1(new_n12831_), .A2(new_n12834_), .B(new_n12840_), .ZN(new_n12862_));
  OAI21_X1   g12605(.A1(new_n12862_), .A2(new_n12861_), .B(new_n12850_), .ZN(new_n12863_));
  AOI21_X1   g12606(.A1(new_n12831_), .A2(new_n12834_), .B(new_n12839_), .ZN(new_n12864_));
  NOR3_X1    g12607(.A1(new_n12844_), .A2(new_n12847_), .A3(new_n12840_), .ZN(new_n12865_));
  OAI21_X1   g12608(.A1(new_n12864_), .A2(new_n12865_), .B(new_n12693_), .ZN(new_n12866_));
  NAND3_X1   g12609(.A1(new_n12863_), .A2(new_n12866_), .A3(new_n12858_), .ZN(new_n12867_));
  AOI21_X1   g12610(.A1(new_n12860_), .A2(new_n12867_), .B(new_n12692_), .ZN(new_n12868_));
  INV_X1     g12611(.I(new_n12692_), .ZN(new_n12869_));
  NAND3_X1   g12612(.A1(new_n12863_), .A2(new_n12866_), .A3(new_n12859_), .ZN(new_n12870_));
  OAI21_X1   g12613(.A1(new_n12849_), .A2(new_n12853_), .B(new_n12858_), .ZN(new_n12871_));
  AOI21_X1   g12614(.A1(new_n12871_), .A2(new_n12870_), .B(new_n12869_), .ZN(new_n12872_));
  NOR2_X1    g12615(.A1(new_n12868_), .A2(new_n12872_), .ZN(new_n12873_));
  NOR3_X1    g12616(.A1(new_n12873_), .A2(new_n12532_), .A3(new_n12691_), .ZN(new_n12874_));
  INV_X1     g12617(.I(new_n12691_), .ZN(new_n12875_));
  AOI21_X1   g12618(.A1(new_n12863_), .A2(new_n12866_), .B(new_n12858_), .ZN(new_n12876_));
  NOR3_X1    g12619(.A1(new_n12849_), .A2(new_n12853_), .A3(new_n12859_), .ZN(new_n12877_));
  OAI21_X1   g12620(.A1(new_n12876_), .A2(new_n12877_), .B(new_n12869_), .ZN(new_n12878_));
  NOR3_X1    g12621(.A1(new_n12849_), .A2(new_n12853_), .A3(new_n12858_), .ZN(new_n12879_));
  AOI21_X1   g12622(.A1(new_n12863_), .A2(new_n12866_), .B(new_n12859_), .ZN(new_n12880_));
  OAI21_X1   g12623(.A1(new_n12880_), .A2(new_n12879_), .B(new_n12692_), .ZN(new_n12881_));
  NAND2_X1   g12624(.A1(new_n12878_), .A2(new_n12881_), .ZN(new_n12882_));
  AOI21_X1   g12625(.A1(new_n12875_), .A2(new_n12531_), .B(new_n12882_), .ZN(new_n12883_));
  OAI21_X1   g12626(.A1(new_n12883_), .A2(new_n12874_), .B(new_n2074_), .ZN(new_n12884_));
  NAND3_X1   g12627(.A1(new_n12882_), .A2(new_n12531_), .A3(new_n12875_), .ZN(new_n12885_));
  OAI21_X1   g12628(.A1(new_n12532_), .A2(new_n12691_), .B(new_n12873_), .ZN(new_n12886_));
  NAND3_X1   g12629(.A1(new_n12886_), .A2(\a[29] ), .A3(new_n12885_), .ZN(new_n12887_));
  AOI21_X1   g12630(.A1(new_n12884_), .A2(new_n12887_), .B(new_n12690_), .ZN(new_n12888_));
  AOI21_X1   g12631(.A1(new_n12886_), .A2(new_n12885_), .B(\a[29] ), .ZN(new_n12889_));
  NOR3_X1    g12632(.A1(new_n12883_), .A2(new_n12874_), .A3(new_n2074_), .ZN(new_n12890_));
  NOR3_X1    g12633(.A1(new_n12890_), .A2(new_n12889_), .A3(new_n12689_), .ZN(new_n12891_));
  OAI22_X1   g12634(.A1(new_n1760_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n1755_), .ZN(new_n12892_));
  NAND2_X1   g12635(.A1(new_n2470_), .A2(\b[47] ), .ZN(new_n12893_));
  AOI21_X1   g12636(.A1(new_n12892_), .A2(new_n12893_), .B(new_n1763_), .ZN(new_n12894_));
  NAND2_X1   g12637(.A1(new_n5196_), .A2(new_n12894_), .ZN(new_n12895_));
  XOR2_X1    g12638(.A1(new_n12895_), .A2(\a[26] ), .Z(new_n12896_));
  INV_X1     g12639(.I(new_n12896_), .ZN(new_n12897_));
  OAI21_X1   g12640(.A1(new_n12891_), .A2(new_n12888_), .B(new_n12897_), .ZN(new_n12898_));
  OAI21_X1   g12641(.A1(new_n12890_), .A2(new_n12889_), .B(new_n12689_), .ZN(new_n12899_));
  NAND3_X1   g12642(.A1(new_n12884_), .A2(new_n12887_), .A3(new_n12690_), .ZN(new_n12900_));
  NAND3_X1   g12643(.A1(new_n12899_), .A2(new_n12900_), .A3(new_n12896_), .ZN(new_n12901_));
  AOI21_X1   g12644(.A1(new_n12898_), .A2(new_n12901_), .B(new_n12686_), .ZN(new_n12902_));
  INV_X1     g12645(.I(new_n12686_), .ZN(new_n12903_));
  NAND3_X1   g12646(.A1(new_n12899_), .A2(new_n12900_), .A3(new_n12897_), .ZN(new_n12904_));
  OAI21_X1   g12647(.A1(new_n12891_), .A2(new_n12888_), .B(new_n12896_), .ZN(new_n12905_));
  AOI21_X1   g12648(.A1(new_n12905_), .A2(new_n12904_), .B(new_n12903_), .ZN(new_n12906_));
  OR2_X2     g12649(.A1(new_n12902_), .A2(new_n12906_), .Z(new_n12907_));
  NAND2_X1   g12650(.A1(new_n12907_), .A2(new_n12682_), .ZN(new_n12908_));
  INV_X1     g12651(.I(new_n12682_), .ZN(new_n12909_));
  NOR2_X1    g12652(.A1(new_n12902_), .A2(new_n12906_), .ZN(new_n12910_));
  NAND2_X1   g12653(.A1(new_n12910_), .A2(new_n12909_), .ZN(new_n12911_));
  AOI21_X1   g12654(.A1(new_n12908_), .A2(new_n12911_), .B(\a[23] ), .ZN(new_n12912_));
  NOR2_X1    g12655(.A1(new_n12910_), .A2(new_n12909_), .ZN(new_n12913_));
  INV_X1     g12656(.I(new_n12911_), .ZN(new_n12914_));
  NOR3_X1    g12657(.A1(new_n12914_), .A2(new_n12913_), .A3(new_n1434_), .ZN(new_n12915_));
  OAI21_X1   g12658(.A1(new_n12915_), .A2(new_n12912_), .B(new_n12681_), .ZN(new_n12916_));
  OAI21_X1   g12659(.A1(new_n12914_), .A2(new_n12913_), .B(new_n1434_), .ZN(new_n12917_));
  NAND3_X1   g12660(.A1(new_n12908_), .A2(new_n12911_), .A3(\a[23] ), .ZN(new_n12918_));
  NAND3_X1   g12661(.A1(new_n12917_), .A2(new_n12918_), .A3(new_n12680_), .ZN(new_n12919_));
  OAI22_X1   g12662(.A1(new_n1168_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n1163_), .ZN(new_n12920_));
  NAND2_X1   g12663(.A1(new_n1774_), .A2(\b[53] ), .ZN(new_n12921_));
  AOI21_X1   g12664(.A1(new_n12920_), .A2(new_n12921_), .B(new_n1171_), .ZN(new_n12922_));
  NAND2_X1   g12665(.A1(new_n6471_), .A2(new_n12922_), .ZN(new_n12923_));
  XOR2_X1    g12666(.A1(new_n12923_), .A2(\a[20] ), .Z(new_n12924_));
  INV_X1     g12667(.I(new_n12924_), .ZN(new_n12925_));
  NAND3_X1   g12668(.A1(new_n12916_), .A2(new_n12919_), .A3(new_n12925_), .ZN(new_n12926_));
  AOI21_X1   g12669(.A1(new_n12917_), .A2(new_n12918_), .B(new_n12680_), .ZN(new_n12927_));
  NOR3_X1    g12670(.A1(new_n12915_), .A2(new_n12912_), .A3(new_n12681_), .ZN(new_n12928_));
  OAI21_X1   g12671(.A1(new_n12928_), .A2(new_n12927_), .B(new_n12924_), .ZN(new_n12929_));
  AOI21_X1   g12672(.A1(new_n12929_), .A2(new_n12926_), .B(new_n12677_), .ZN(new_n12930_));
  INV_X1     g12673(.I(new_n12677_), .ZN(new_n12931_));
  OAI21_X1   g12674(.A1(new_n12928_), .A2(new_n12927_), .B(new_n12925_), .ZN(new_n12932_));
  NAND3_X1   g12675(.A1(new_n12916_), .A2(new_n12919_), .A3(new_n12924_), .ZN(new_n12933_));
  AOI21_X1   g12676(.A1(new_n12932_), .A2(new_n12933_), .B(new_n12931_), .ZN(new_n12934_));
  OAI22_X1   g12677(.A1(new_n940_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n935_), .ZN(new_n12935_));
  NAND2_X1   g12678(.A1(new_n1458_), .A2(\b[56] ), .ZN(new_n12936_));
  AOI21_X1   g12679(.A1(new_n12935_), .A2(new_n12936_), .B(new_n943_), .ZN(new_n12937_));
  NAND2_X1   g12680(.A1(new_n7559_), .A2(new_n12937_), .ZN(new_n12938_));
  XOR2_X1    g12681(.A1(new_n12938_), .A2(\a[17] ), .Z(new_n12939_));
  INV_X1     g12682(.I(new_n12939_), .ZN(new_n12940_));
  OAI21_X1   g12683(.A1(new_n12930_), .A2(new_n12934_), .B(new_n12940_), .ZN(new_n12941_));
  NOR3_X1    g12684(.A1(new_n12928_), .A2(new_n12927_), .A3(new_n12924_), .ZN(new_n12942_));
  AOI21_X1   g12685(.A1(new_n12916_), .A2(new_n12919_), .B(new_n12925_), .ZN(new_n12943_));
  OAI21_X1   g12686(.A1(new_n12942_), .A2(new_n12943_), .B(new_n12931_), .ZN(new_n12944_));
  AOI21_X1   g12687(.A1(new_n12916_), .A2(new_n12919_), .B(new_n12924_), .ZN(new_n12945_));
  NOR3_X1    g12688(.A1(new_n12928_), .A2(new_n12927_), .A3(new_n12925_), .ZN(new_n12946_));
  OAI21_X1   g12689(.A1(new_n12946_), .A2(new_n12945_), .B(new_n12677_), .ZN(new_n12947_));
  NAND3_X1   g12690(.A1(new_n12944_), .A2(new_n12947_), .A3(new_n12939_), .ZN(new_n12948_));
  AOI21_X1   g12691(.A1(new_n12941_), .A2(new_n12948_), .B(new_n12676_), .ZN(new_n12949_));
  INV_X1     g12692(.I(new_n12676_), .ZN(new_n12950_));
  NAND3_X1   g12693(.A1(new_n12944_), .A2(new_n12947_), .A3(new_n12940_), .ZN(new_n12951_));
  OAI21_X1   g12694(.A1(new_n12930_), .A2(new_n12934_), .B(new_n12939_), .ZN(new_n12952_));
  AOI21_X1   g12695(.A1(new_n12952_), .A2(new_n12951_), .B(new_n12950_), .ZN(new_n12953_));
  OAI22_X1   g12696(.A1(new_n757_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n752_), .ZN(new_n12954_));
  NAND2_X1   g12697(.A1(new_n1182_), .A2(\b[59] ), .ZN(new_n12955_));
  AOI21_X1   g12698(.A1(new_n12954_), .A2(new_n12955_), .B(new_n760_), .ZN(new_n12956_));
  NAND2_X1   g12699(.A1(new_n8550_), .A2(new_n12956_), .ZN(new_n12957_));
  XOR2_X1    g12700(.A1(new_n12957_), .A2(\a[14] ), .Z(new_n12958_));
  INV_X1     g12701(.I(new_n12958_), .ZN(new_n12959_));
  OAI21_X1   g12702(.A1(new_n12949_), .A2(new_n12953_), .B(new_n12959_), .ZN(new_n12960_));
  INV_X1     g12703(.I(new_n12960_), .ZN(new_n12961_));
  NOR3_X1    g12704(.A1(new_n12949_), .A2(new_n12953_), .A3(new_n12959_), .ZN(new_n12962_));
  OAI21_X1   g12705(.A1(new_n12961_), .A2(new_n12962_), .B(new_n12675_), .ZN(new_n12963_));
  NOR3_X1    g12706(.A1(new_n12949_), .A2(new_n12953_), .A3(new_n12958_), .ZN(new_n12964_));
  AOI21_X1   g12707(.A1(new_n12944_), .A2(new_n12947_), .B(new_n12939_), .ZN(new_n12965_));
  NOR3_X1    g12708(.A1(new_n12930_), .A2(new_n12934_), .A3(new_n12940_), .ZN(new_n12966_));
  OAI21_X1   g12709(.A1(new_n12965_), .A2(new_n12966_), .B(new_n12950_), .ZN(new_n12967_));
  INV_X1     g12710(.I(new_n12953_), .ZN(new_n12968_));
  AOI21_X1   g12711(.A1(new_n12968_), .A2(new_n12967_), .B(new_n12959_), .ZN(new_n12969_));
  OAI21_X1   g12712(.A1(new_n12969_), .A2(new_n12964_), .B(new_n12674_), .ZN(new_n12970_));
  NOR2_X1    g12713(.A1(new_n635_), .A2(new_n8932_), .ZN(new_n12971_));
  NOR2_X1    g12714(.A1(new_n577_), .A2(new_n8956_), .ZN(new_n12972_));
  NOR4_X1    g12715(.A1(new_n9323_), .A2(new_n585_), .A3(new_n12971_), .A4(new_n12972_), .ZN(new_n12973_));
  XOR2_X1    g12716(.A1(new_n12973_), .A2(new_n572_), .Z(new_n12974_));
  INV_X1     g12717(.I(new_n12974_), .ZN(new_n12975_));
  NAND3_X1   g12718(.A1(new_n12963_), .A2(new_n12970_), .A3(new_n12975_), .ZN(new_n12976_));
  INV_X1     g12719(.I(new_n12962_), .ZN(new_n12977_));
  AOI21_X1   g12720(.A1(new_n12977_), .A2(new_n12960_), .B(new_n12674_), .ZN(new_n12978_));
  INV_X1     g12721(.I(new_n12964_), .ZN(new_n12979_));
  OAI21_X1   g12722(.A1(new_n12949_), .A2(new_n12953_), .B(new_n12958_), .ZN(new_n12980_));
  AOI21_X1   g12723(.A1(new_n12979_), .A2(new_n12980_), .B(new_n12675_), .ZN(new_n12981_));
  OAI21_X1   g12724(.A1(new_n12978_), .A2(new_n12981_), .B(new_n12974_), .ZN(new_n12982_));
  AOI21_X1   g12725(.A1(new_n12982_), .A2(new_n12976_), .B(new_n12673_), .ZN(new_n12983_));
  INV_X1     g12726(.I(new_n12673_), .ZN(new_n12984_));
  OAI21_X1   g12727(.A1(new_n12978_), .A2(new_n12981_), .B(new_n12975_), .ZN(new_n12985_));
  NAND3_X1   g12728(.A1(new_n12963_), .A2(new_n12970_), .A3(new_n12974_), .ZN(new_n12986_));
  AOI21_X1   g12729(.A1(new_n12985_), .A2(new_n12986_), .B(new_n12984_), .ZN(new_n12987_));
  OR2_X2     g12730(.A1(new_n12983_), .A2(new_n12987_), .Z(new_n12988_));
  INV_X1     g12731(.I(new_n11971_), .ZN(new_n12989_));
  NOR2_X1    g12732(.A1(new_n11583_), .A2(new_n11571_), .ZN(new_n12990_));
  INV_X1     g12733(.I(new_n11974_), .ZN(new_n12991_));
  AOI21_X1   g12734(.A1(new_n11972_), .A2(new_n12991_), .B(new_n11966_), .ZN(new_n12992_));
  OAI21_X1   g12735(.A1(new_n11581_), .A2(new_n12990_), .B(new_n12992_), .ZN(new_n12993_));
  NAND3_X1   g12736(.A1(new_n12993_), .A2(new_n12989_), .A3(new_n12330_), .ZN(new_n12994_));
  NOR2_X1    g12737(.A1(new_n12663_), .A2(new_n12336_), .ZN(new_n12995_));
  NOR3_X1    g12738(.A1(new_n12330_), .A2(new_n12664_), .A3(new_n12995_), .ZN(new_n12996_));
  AOI21_X1   g12739(.A1(new_n12994_), .A2(new_n12996_), .B(new_n12988_), .ZN(new_n12997_));
  NOR2_X1    g12740(.A1(new_n12983_), .A2(new_n12987_), .ZN(new_n12998_));
  OAI21_X1   g12741(.A1(new_n12325_), .A2(new_n12322_), .B(new_n11980_), .ZN(new_n12999_));
  NOR3_X1    g12742(.A1(new_n11976_), .A2(new_n11971_), .A3(new_n12999_), .ZN(new_n13000_));
  XOR2_X1    g12743(.A1(new_n12663_), .A2(new_n12336_), .Z(new_n13001_));
  NAND2_X1   g12744(.A1(new_n12999_), .A2(new_n13001_), .ZN(new_n13002_));
  NOR3_X1    g12745(.A1(new_n13000_), .A2(new_n12998_), .A3(new_n13002_), .ZN(new_n13003_));
  NOR2_X1    g12746(.A1(new_n12997_), .A2(new_n13003_), .ZN(new_n13004_));
  XOR2_X1    g12747(.A1(new_n13004_), .A2(new_n12671_), .Z(\f[73] ));
  NOR2_X1    g12748(.A1(new_n13000_), .A2(new_n13002_), .ZN(new_n13006_));
  OAI22_X1   g12749(.A1(new_n12997_), .A2(new_n13003_), .B1(new_n13006_), .B2(new_n12671_), .ZN(new_n13007_));
  NAND2_X1   g12750(.A1(new_n12986_), .A2(new_n12984_), .ZN(new_n13008_));
  NAND2_X1   g12751(.A1(new_n13008_), .A2(new_n12985_), .ZN(new_n13009_));
  INV_X1     g12752(.I(new_n13009_), .ZN(new_n13010_));
  AOI22_X1   g12753(.A1(new_n10814_), .A2(new_n584_), .B1(\b[63] ), .B2(new_n960_), .ZN(new_n13011_));
  OAI21_X1   g12754(.A1(new_n12674_), .A2(new_n12962_), .B(new_n12960_), .ZN(new_n13012_));
  INV_X1     g12755(.I(new_n13012_), .ZN(new_n13013_));
  OAI22_X1   g12756(.A1(new_n757_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n752_), .ZN(new_n13014_));
  OAI21_X1   g12757(.A1(new_n7930_), .A2(new_n823_), .B(new_n13014_), .ZN(new_n13015_));
  AOI21_X1   g12758(.A1(new_n8935_), .A2(new_n759_), .B(new_n13015_), .ZN(new_n13016_));
  INV_X1     g12759(.I(new_n13016_), .ZN(new_n13017_));
  OAI21_X1   g12760(.A1(new_n12676_), .A2(new_n12966_), .B(new_n12941_), .ZN(new_n13018_));
  AOI21_X1   g12761(.A1(new_n12931_), .A2(new_n12929_), .B(new_n12942_), .ZN(new_n13019_));
  INV_X1     g12762(.I(new_n13019_), .ZN(new_n13020_));
  OAI22_X1   g12763(.A1(new_n1168_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n1163_), .ZN(new_n13021_));
  OAI21_X1   g12764(.A1(new_n6238_), .A2(new_n1255_), .B(new_n13021_), .ZN(new_n13022_));
  AOI21_X1   g12765(.A1(new_n6994_), .A2(new_n1170_), .B(new_n13022_), .ZN(new_n13023_));
  NOR2_X1    g12766(.A1(new_n12910_), .A2(new_n12682_), .ZN(new_n13024_));
  XOR2_X1    g12767(.A1(new_n12680_), .A2(new_n1434_), .Z(new_n13025_));
  AOI21_X1   g12768(.A1(new_n12910_), .A2(new_n12682_), .B(new_n13025_), .ZN(new_n13026_));
  NOR2_X1    g12769(.A1(new_n13026_), .A2(new_n13024_), .ZN(new_n13027_));
  NAND2_X1   g12770(.A1(new_n12901_), .A2(new_n12903_), .ZN(new_n13028_));
  OAI22_X1   g12771(.A1(new_n1760_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n1755_), .ZN(new_n13029_));
  OAI21_X1   g12772(.A1(new_n5178_), .A2(new_n1857_), .B(new_n13029_), .ZN(new_n13030_));
  AOI21_X1   g12773(.A1(new_n5537_), .A2(new_n1762_), .B(new_n13030_), .ZN(new_n13031_));
  INV_X1     g12774(.I(new_n13031_), .ZN(new_n13032_));
  AOI21_X1   g12775(.A1(new_n12875_), .A2(new_n12531_), .B(new_n12873_), .ZN(new_n13033_));
  INV_X1     g12776(.I(new_n13033_), .ZN(new_n13034_));
  XOR2_X1    g12777(.A1(new_n12689_), .A2(\a[29] ), .Z(new_n13035_));
  INV_X1     g12778(.I(new_n13035_), .ZN(new_n13036_));
  NAND4_X1   g12779(.A1(new_n12873_), .A2(new_n12531_), .A3(new_n12875_), .A4(new_n13036_), .ZN(new_n13037_));
  NAND2_X1   g12780(.A1(new_n13034_), .A2(new_n13037_), .ZN(new_n13038_));
  AOI21_X1   g12781(.A1(new_n12869_), .A2(new_n12867_), .B(new_n12876_), .ZN(new_n13039_));
  INV_X1     g12782(.I(new_n13039_), .ZN(new_n13040_));
  OAI22_X1   g12783(.A1(new_n2452_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n2447_), .ZN(new_n13041_));
  OAI21_X1   g12784(.A1(new_n4018_), .A2(new_n2602_), .B(new_n13041_), .ZN(new_n13042_));
  AOI21_X1   g12785(.A1(new_n4500_), .A2(new_n2454_), .B(new_n13042_), .ZN(new_n13043_));
  INV_X1     g12786(.I(new_n13043_), .ZN(new_n13044_));
  OAI21_X1   g12787(.A1(new_n12693_), .A2(new_n12862_), .B(new_n12841_), .ZN(new_n13045_));
  AOI21_X1   g12788(.A1(new_n12695_), .A2(new_n12846_), .B(new_n12832_), .ZN(new_n13046_));
  INV_X1     g12789(.I(new_n13046_), .ZN(new_n13047_));
  OAI22_X1   g12790(.A1(new_n2846_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n2841_), .ZN(new_n13048_));
  NAND2_X1   g12791(.A1(new_n3755_), .A2(\b[39] ), .ZN(new_n13049_));
  AOI21_X1   g12792(.A1(new_n13048_), .A2(new_n13049_), .B(new_n2849_), .ZN(new_n13050_));
  NAND2_X1   g12793(.A1(new_n3996_), .A2(new_n13050_), .ZN(new_n13051_));
  XOR2_X1    g12794(.A1(new_n13051_), .A2(\a[35] ), .Z(new_n13052_));
  INV_X1     g12795(.I(new_n13052_), .ZN(new_n13053_));
  AOI21_X1   g12796(.A1(new_n12697_), .A2(new_n12826_), .B(new_n12815_), .ZN(new_n13054_));
  INV_X1     g12797(.I(new_n13054_), .ZN(new_n13055_));
  OAI22_X1   g12798(.A1(new_n3298_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n3293_), .ZN(new_n13056_));
  NAND2_X1   g12799(.A1(new_n4227_), .A2(\b[36] ), .ZN(new_n13057_));
  AOI21_X1   g12800(.A1(new_n13056_), .A2(new_n13057_), .B(new_n3301_), .ZN(new_n13058_));
  NAND2_X1   g12801(.A1(new_n3565_), .A2(new_n13058_), .ZN(new_n13059_));
  XOR2_X1    g12802(.A1(new_n13059_), .A2(\a[38] ), .Z(new_n13060_));
  INV_X1     g12803(.I(new_n13060_), .ZN(new_n13061_));
  OAI22_X1   g12804(.A1(new_n4208_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n4203_), .ZN(new_n13062_));
  NAND2_X1   g12805(.A1(new_n5244_), .A2(\b[30] ), .ZN(new_n13063_));
  AOI21_X1   g12806(.A1(new_n13062_), .A2(new_n13063_), .B(new_n4211_), .ZN(new_n13064_));
  NAND2_X1   g12807(.A1(new_n2659_), .A2(new_n13064_), .ZN(new_n13065_));
  XOR2_X1    g12808(.A1(new_n13065_), .A2(\a[44] ), .Z(new_n13066_));
  OAI22_X1   g12809(.A1(new_n5228_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n5225_), .ZN(new_n13067_));
  NAND2_X1   g12810(.A1(new_n5387_), .A2(\b[24] ), .ZN(new_n13068_));
  AOI21_X1   g12811(.A1(new_n13067_), .A2(new_n13068_), .B(new_n5231_), .ZN(new_n13069_));
  NAND2_X1   g12812(.A1(new_n1926_), .A2(new_n13069_), .ZN(new_n13070_));
  XOR2_X1    g12813(.A1(new_n13070_), .A2(\a[50] ), .Z(new_n13071_));
  AOI21_X1   g12814(.A1(new_n12766_), .A2(new_n12764_), .B(new_n12762_), .ZN(new_n13072_));
  OAI22_X1   g12815(.A1(new_n5786_), .A2(new_n1601_), .B1(new_n1518_), .B2(new_n5792_), .ZN(new_n13073_));
  NAND2_X1   g12816(.A1(new_n6745_), .A2(\b[21] ), .ZN(new_n13074_));
  AOI21_X1   g12817(.A1(new_n13074_), .A2(new_n13073_), .B(new_n5796_), .ZN(new_n13075_));
  NAND2_X1   g12818(.A1(new_n1604_), .A2(new_n13075_), .ZN(new_n13076_));
  XOR2_X1    g12819(.A1(new_n13076_), .A2(\a[53] ), .Z(new_n13077_));
  OAI22_X1   g12820(.A1(new_n6721_), .A2(new_n1222_), .B1(new_n6723_), .B2(new_n1305_), .ZN(new_n13078_));
  NAND2_X1   g12821(.A1(new_n7617_), .A2(\b[18] ), .ZN(new_n13079_));
  AOI21_X1   g12822(.A1(new_n13079_), .A2(new_n13078_), .B(new_n6731_), .ZN(new_n13080_));
  NAND2_X1   g12823(.A1(new_n1304_), .A2(new_n13080_), .ZN(new_n13081_));
  XOR2_X1    g12824(.A1(new_n13081_), .A2(\a[56] ), .Z(new_n13082_));
  NAND2_X1   g12825(.A1(new_n12724_), .A2(new_n12732_), .ZN(new_n13083_));
  NAND2_X1   g12826(.A1(new_n13083_), .A2(new_n12733_), .ZN(new_n13084_));
  NOR3_X1    g12827(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n617_), .ZN(new_n13085_));
  NOR2_X1    g12828(.A1(new_n9364_), .A2(new_n617_), .ZN(new_n13086_));
  NOR3_X1    g12829(.A1(new_n13086_), .A2(new_n659_), .A3(new_n8985_), .ZN(new_n13087_));
  NOR2_X1    g12830(.A1(new_n13087_), .A2(new_n13085_), .ZN(new_n13088_));
  NOR2_X1    g12831(.A1(new_n12735_), .A2(new_n13088_), .ZN(new_n13089_));
  INV_X1     g12832(.I(new_n13088_), .ZN(new_n13090_));
  NOR2_X1    g12833(.A1(new_n13090_), .A2(new_n12730_), .ZN(new_n13091_));
  NOR2_X1    g12834(.A1(new_n13089_), .A2(new_n13091_), .ZN(new_n13092_));
  INV_X1     g12835(.I(new_n13092_), .ZN(new_n13093_));
  NAND2_X1   g12836(.A1(new_n13084_), .A2(new_n13093_), .ZN(new_n13094_));
  XOR2_X1    g12837(.A1(new_n12730_), .A2(new_n13088_), .Z(new_n13095_));
  OAI21_X1   g12838(.A1(new_n13084_), .A2(new_n13095_), .B(new_n13094_), .ZN(new_n13096_));
  INV_X1     g12839(.I(new_n13096_), .ZN(new_n13097_));
  OAI22_X1   g12840(.A1(new_n1044_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n992_), .ZN(new_n13098_));
  NAND2_X1   g12841(.A1(new_n8628_), .A2(\b[15] ), .ZN(new_n13099_));
  AOI21_X1   g12842(.A1(new_n13099_), .A2(new_n13098_), .B(new_n7354_), .ZN(new_n13100_));
  NAND2_X1   g12843(.A1(new_n1047_), .A2(new_n13100_), .ZN(new_n13101_));
  XOR2_X1    g12844(.A1(new_n13101_), .A2(new_n7343_), .Z(new_n13102_));
  OAI22_X1   g12845(.A1(new_n848_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n795_), .ZN(new_n13103_));
  NAND2_X1   g12846(.A1(new_n9644_), .A2(\b[12] ), .ZN(new_n13104_));
  AOI21_X1   g12847(.A1(new_n13104_), .A2(new_n13103_), .B(new_n8321_), .ZN(new_n13105_));
  NAND2_X1   g12848(.A1(new_n847_), .A2(new_n13105_), .ZN(new_n13106_));
  XOR2_X1    g12849(.A1(new_n13106_), .A2(\a[62] ), .Z(new_n13107_));
  INV_X1     g12850(.I(new_n13107_), .ZN(new_n13108_));
  NAND2_X1   g12851(.A1(new_n13102_), .A2(new_n13108_), .ZN(new_n13109_));
  XOR2_X1    g12852(.A1(new_n13101_), .A2(\a[59] ), .Z(new_n13110_));
  NAND2_X1   g12853(.A1(new_n13110_), .A2(new_n13107_), .ZN(new_n13111_));
  AOI21_X1   g12854(.A1(new_n13109_), .A2(new_n13111_), .B(new_n13097_), .ZN(new_n13112_));
  XOR2_X1    g12855(.A1(new_n13102_), .A2(new_n13107_), .Z(new_n13113_));
  NOR2_X1    g12856(.A1(new_n13113_), .A2(new_n13096_), .ZN(new_n13114_));
  NOR2_X1    g12857(.A1(new_n13114_), .A2(new_n13112_), .ZN(new_n13115_));
  AOI21_X1   g12858(.A1(new_n12713_), .A2(new_n12741_), .B(new_n12739_), .ZN(new_n13116_));
  INV_X1     g12859(.I(new_n13116_), .ZN(new_n13117_));
  XOR2_X1    g12860(.A1(new_n13115_), .A2(new_n13117_), .Z(new_n13118_));
  NOR2_X1    g12861(.A1(new_n13118_), .A2(new_n13082_), .ZN(new_n13119_));
  INV_X1     g12862(.I(new_n13082_), .ZN(new_n13120_));
  OAI21_X1   g12863(.A1(new_n13114_), .A2(new_n13112_), .B(new_n13117_), .ZN(new_n13121_));
  NAND2_X1   g12864(.A1(new_n13115_), .A2(new_n13116_), .ZN(new_n13122_));
  AOI21_X1   g12865(.A1(new_n13122_), .A2(new_n13121_), .B(new_n13120_), .ZN(new_n13123_));
  NOR2_X1    g12866(.A1(new_n13119_), .A2(new_n13123_), .ZN(new_n13124_));
  INV_X1     g12867(.I(new_n12745_), .ZN(new_n13125_));
  AOI21_X1   g12868(.A1(new_n13125_), .A2(new_n12755_), .B(new_n12753_), .ZN(new_n13126_));
  XOR2_X1    g12869(.A1(new_n13124_), .A2(new_n13126_), .Z(new_n13127_));
  NOR2_X1    g12870(.A1(new_n13127_), .A2(new_n13077_), .ZN(new_n13128_));
  INV_X1     g12871(.I(new_n13077_), .ZN(new_n13129_));
  INV_X1     g12872(.I(new_n13126_), .ZN(new_n13130_));
  NAND2_X1   g12873(.A1(new_n13124_), .A2(new_n13130_), .ZN(new_n13131_));
  OAI21_X1   g12874(.A1(new_n13119_), .A2(new_n13123_), .B(new_n13126_), .ZN(new_n13132_));
  AOI21_X1   g12875(.A1(new_n13131_), .A2(new_n13132_), .B(new_n13129_), .ZN(new_n13133_));
  NOR2_X1    g12876(.A1(new_n13128_), .A2(new_n13133_), .ZN(new_n13134_));
  XOR2_X1    g12877(.A1(new_n13134_), .A2(new_n13072_), .Z(new_n13135_));
  NOR2_X1    g12878(.A1(new_n13135_), .A2(new_n13071_), .ZN(new_n13136_));
  INV_X1     g12879(.I(new_n13071_), .ZN(new_n13137_));
  OAI21_X1   g12880(.A1(new_n13128_), .A2(new_n13133_), .B(new_n13072_), .ZN(new_n13138_));
  INV_X1     g12881(.I(new_n13072_), .ZN(new_n13139_));
  NAND2_X1   g12882(.A1(new_n13134_), .A2(new_n13139_), .ZN(new_n13140_));
  AOI21_X1   g12883(.A1(new_n13140_), .A2(new_n13138_), .B(new_n13137_), .ZN(new_n13141_));
  NOR2_X1    g12884(.A1(new_n13136_), .A2(new_n13141_), .ZN(new_n13142_));
  OAI22_X1   g12885(.A1(new_n4711_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n4706_), .ZN(new_n13143_));
  NAND2_X1   g12886(.A1(new_n5814_), .A2(\b[27] ), .ZN(new_n13144_));
  AOI21_X1   g12887(.A1(new_n13143_), .A2(new_n13144_), .B(new_n4714_), .ZN(new_n13145_));
  NAND2_X1   g12888(.A1(new_n2276_), .A2(new_n13145_), .ZN(new_n13146_));
  XOR2_X1    g12889(.A1(new_n13146_), .A2(\a[47] ), .Z(new_n13147_));
  INV_X1     g12890(.I(new_n13147_), .ZN(new_n13148_));
  AOI21_X1   g12891(.A1(new_n12772_), .A2(new_n12777_), .B(new_n12769_), .ZN(new_n13149_));
  NOR2_X1    g12892(.A1(new_n13149_), .A2(new_n12778_), .ZN(new_n13150_));
  XOR2_X1    g12893(.A1(new_n13150_), .A2(new_n13148_), .Z(new_n13151_));
  NOR2_X1    g12894(.A1(new_n13142_), .A2(new_n13151_), .ZN(new_n13152_));
  INV_X1     g12895(.I(new_n13152_), .ZN(new_n13153_));
  NOR2_X1    g12896(.A1(new_n13150_), .A2(new_n13147_), .ZN(new_n13154_));
  NOR3_X1    g12897(.A1(new_n13148_), .A2(new_n13149_), .A3(new_n12778_), .ZN(new_n13155_));
  OAI21_X1   g12898(.A1(new_n13154_), .A2(new_n13155_), .B(new_n13142_), .ZN(new_n13156_));
  AOI21_X1   g12899(.A1(new_n12791_), .A2(new_n12789_), .B(new_n12787_), .ZN(new_n13157_));
  INV_X1     g12900(.I(new_n13157_), .ZN(new_n13158_));
  NAND3_X1   g12901(.A1(new_n13153_), .A2(new_n13156_), .A3(new_n13158_), .ZN(new_n13159_));
  INV_X1     g12902(.I(new_n13142_), .ZN(new_n13160_));
  NOR2_X1    g12903(.A1(new_n13154_), .A2(new_n13155_), .ZN(new_n13161_));
  NOR2_X1    g12904(.A1(new_n13160_), .A2(new_n13161_), .ZN(new_n13162_));
  OAI21_X1   g12905(.A1(new_n13162_), .A2(new_n13152_), .B(new_n13157_), .ZN(new_n13163_));
  AOI21_X1   g12906(.A1(new_n13163_), .A2(new_n13159_), .B(new_n13066_), .ZN(new_n13164_));
  INV_X1     g12907(.I(new_n13066_), .ZN(new_n13165_));
  OAI21_X1   g12908(.A1(new_n13162_), .A2(new_n13152_), .B(new_n13158_), .ZN(new_n13166_));
  NAND3_X1   g12909(.A1(new_n13153_), .A2(new_n13156_), .A3(new_n13157_), .ZN(new_n13167_));
  AOI21_X1   g12910(.A1(new_n13166_), .A2(new_n13167_), .B(new_n13165_), .ZN(new_n13168_));
  OAI22_X1   g12911(.A1(new_n3736_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n3731_), .ZN(new_n13169_));
  NAND2_X1   g12912(.A1(new_n4730_), .A2(\b[33] ), .ZN(new_n13170_));
  AOI21_X1   g12913(.A1(new_n13169_), .A2(new_n13170_), .B(new_n3739_), .ZN(new_n13171_));
  NAND2_X1   g12914(.A1(new_n3101_), .A2(new_n13171_), .ZN(new_n13172_));
  XOR2_X1    g12915(.A1(new_n13172_), .A2(\a[41] ), .Z(new_n13173_));
  INV_X1     g12916(.I(new_n12805_), .ZN(new_n13174_));
  OAI21_X1   g12917(.A1(new_n12793_), .A2(new_n12790_), .B(new_n12806_), .ZN(new_n13175_));
  NAND2_X1   g12918(.A1(new_n13175_), .A2(new_n13174_), .ZN(new_n13176_));
  NAND2_X1   g12919(.A1(new_n13176_), .A2(new_n13173_), .ZN(new_n13177_));
  INV_X1     g12920(.I(new_n13177_), .ZN(new_n13178_));
  NOR2_X1    g12921(.A1(new_n13176_), .A2(new_n13173_), .ZN(new_n13179_));
  OAI22_X1   g12922(.A1(new_n13178_), .A2(new_n13179_), .B1(new_n13164_), .B2(new_n13168_), .ZN(new_n13180_));
  NOR2_X1    g12923(.A1(new_n13164_), .A2(new_n13168_), .ZN(new_n13181_));
  INV_X1     g12924(.I(new_n13173_), .ZN(new_n13182_));
  NAND2_X1   g12925(.A1(new_n13176_), .A2(new_n13182_), .ZN(new_n13183_));
  INV_X1     g12926(.I(new_n13183_), .ZN(new_n13184_));
  NOR2_X1    g12927(.A1(new_n13176_), .A2(new_n13182_), .ZN(new_n13185_));
  OAI21_X1   g12928(.A1(new_n13184_), .A2(new_n13185_), .B(new_n13181_), .ZN(new_n13186_));
  AOI21_X1   g12929(.A1(new_n13186_), .A2(new_n13180_), .B(new_n13061_), .ZN(new_n13187_));
  INV_X1     g12930(.I(new_n13180_), .ZN(new_n13188_));
  NOR2_X1    g12931(.A1(new_n13184_), .A2(new_n13185_), .ZN(new_n13189_));
  NOR3_X1    g12932(.A1(new_n13189_), .A2(new_n13164_), .A3(new_n13168_), .ZN(new_n13190_));
  NOR3_X1    g12933(.A1(new_n13190_), .A2(new_n13188_), .A3(new_n13060_), .ZN(new_n13191_));
  OAI21_X1   g12934(.A1(new_n13191_), .A2(new_n13187_), .B(new_n13055_), .ZN(new_n13192_));
  AOI21_X1   g12935(.A1(new_n13186_), .A2(new_n13180_), .B(new_n13060_), .ZN(new_n13193_));
  NOR3_X1    g12936(.A1(new_n13190_), .A2(new_n13188_), .A3(new_n13061_), .ZN(new_n13194_));
  OAI21_X1   g12937(.A1(new_n13194_), .A2(new_n13193_), .B(new_n13054_), .ZN(new_n13195_));
  AOI21_X1   g12938(.A1(new_n13192_), .A2(new_n13195_), .B(new_n13053_), .ZN(new_n13196_));
  OAI21_X1   g12939(.A1(new_n13190_), .A2(new_n13188_), .B(new_n13060_), .ZN(new_n13197_));
  NAND3_X1   g12940(.A1(new_n13186_), .A2(new_n13061_), .A3(new_n13180_), .ZN(new_n13198_));
  AOI21_X1   g12941(.A1(new_n13197_), .A2(new_n13198_), .B(new_n13054_), .ZN(new_n13199_));
  OAI21_X1   g12942(.A1(new_n13190_), .A2(new_n13188_), .B(new_n13061_), .ZN(new_n13200_));
  NAND3_X1   g12943(.A1(new_n13186_), .A2(new_n13060_), .A3(new_n13180_), .ZN(new_n13201_));
  AOI21_X1   g12944(.A1(new_n13200_), .A2(new_n13201_), .B(new_n13055_), .ZN(new_n13202_));
  NOR3_X1    g12945(.A1(new_n13199_), .A2(new_n13202_), .A3(new_n13052_), .ZN(new_n13203_));
  OAI21_X1   g12946(.A1(new_n13196_), .A2(new_n13203_), .B(new_n13047_), .ZN(new_n13204_));
  AOI21_X1   g12947(.A1(new_n13192_), .A2(new_n13195_), .B(new_n13052_), .ZN(new_n13205_));
  NOR3_X1    g12948(.A1(new_n13199_), .A2(new_n13202_), .A3(new_n13053_), .ZN(new_n13206_));
  OAI21_X1   g12949(.A1(new_n13205_), .A2(new_n13206_), .B(new_n13046_), .ZN(new_n13207_));
  AOI21_X1   g12950(.A1(new_n13204_), .A2(new_n13207_), .B(new_n13045_), .ZN(new_n13208_));
  AOI21_X1   g12951(.A1(new_n12850_), .A2(new_n12848_), .B(new_n12861_), .ZN(new_n13209_));
  OAI21_X1   g12952(.A1(new_n13199_), .A2(new_n13202_), .B(new_n13052_), .ZN(new_n13210_));
  NAND3_X1   g12953(.A1(new_n13192_), .A2(new_n13195_), .A3(new_n13053_), .ZN(new_n13211_));
  AOI21_X1   g12954(.A1(new_n13210_), .A2(new_n13211_), .B(new_n13046_), .ZN(new_n13212_));
  OAI21_X1   g12955(.A1(new_n13199_), .A2(new_n13202_), .B(new_n13053_), .ZN(new_n13213_));
  NAND3_X1   g12956(.A1(new_n13192_), .A2(new_n13195_), .A3(new_n13052_), .ZN(new_n13214_));
  AOI21_X1   g12957(.A1(new_n13213_), .A2(new_n13214_), .B(new_n13047_), .ZN(new_n13215_));
  NOR3_X1    g12958(.A1(new_n13212_), .A2(new_n13215_), .A3(new_n13209_), .ZN(new_n13216_));
  OAI21_X1   g12959(.A1(new_n13208_), .A2(new_n13216_), .B(new_n2442_), .ZN(new_n13217_));
  OAI21_X1   g12960(.A1(new_n13212_), .A2(new_n13215_), .B(new_n13209_), .ZN(new_n13218_));
  NAND3_X1   g12961(.A1(new_n13204_), .A2(new_n13207_), .A3(new_n13045_), .ZN(new_n13219_));
  NAND3_X1   g12962(.A1(new_n13218_), .A2(new_n13219_), .A3(\a[32] ), .ZN(new_n13220_));
  AOI21_X1   g12963(.A1(new_n13217_), .A2(new_n13220_), .B(new_n13044_), .ZN(new_n13221_));
  AOI21_X1   g12964(.A1(new_n13218_), .A2(new_n13219_), .B(\a[32] ), .ZN(new_n13222_));
  NOR3_X1    g12965(.A1(new_n13208_), .A2(new_n13216_), .A3(new_n2442_), .ZN(new_n13223_));
  NOR3_X1    g12966(.A1(new_n13223_), .A2(new_n13222_), .A3(new_n13043_), .ZN(new_n13224_));
  OAI22_X1   g12967(.A1(new_n2084_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n2079_), .ZN(new_n13225_));
  NAND2_X1   g12968(.A1(new_n2864_), .A2(\b[45] ), .ZN(new_n13226_));
  AOI21_X1   g12969(.A1(new_n13225_), .A2(new_n13226_), .B(new_n2087_), .ZN(new_n13227_));
  NAND2_X1   g12970(.A1(new_n5004_), .A2(new_n13227_), .ZN(new_n13228_));
  XOR2_X1    g12971(.A1(new_n13228_), .A2(\a[29] ), .Z(new_n13229_));
  NOR3_X1    g12972(.A1(new_n13224_), .A2(new_n13221_), .A3(new_n13229_), .ZN(new_n13230_));
  OAI21_X1   g12973(.A1(new_n13223_), .A2(new_n13222_), .B(new_n13043_), .ZN(new_n13231_));
  NAND3_X1   g12974(.A1(new_n13217_), .A2(new_n13220_), .A3(new_n13044_), .ZN(new_n13232_));
  INV_X1     g12975(.I(new_n13229_), .ZN(new_n13233_));
  AOI21_X1   g12976(.A1(new_n13231_), .A2(new_n13232_), .B(new_n13233_), .ZN(new_n13234_));
  OAI21_X1   g12977(.A1(new_n13230_), .A2(new_n13234_), .B(new_n13040_), .ZN(new_n13235_));
  AOI21_X1   g12978(.A1(new_n13231_), .A2(new_n13232_), .B(new_n13229_), .ZN(new_n13236_));
  NOR3_X1    g12979(.A1(new_n13224_), .A2(new_n13221_), .A3(new_n13233_), .ZN(new_n13237_));
  OAI21_X1   g12980(.A1(new_n13237_), .A2(new_n13236_), .B(new_n13039_), .ZN(new_n13238_));
  AOI21_X1   g12981(.A1(new_n13235_), .A2(new_n13238_), .B(new_n13038_), .ZN(new_n13239_));
  INV_X1     g12982(.I(new_n13037_), .ZN(new_n13240_));
  NOR2_X1    g12983(.A1(new_n13240_), .A2(new_n13033_), .ZN(new_n13241_));
  NAND3_X1   g12984(.A1(new_n13231_), .A2(new_n13232_), .A3(new_n13233_), .ZN(new_n13242_));
  OAI21_X1   g12985(.A1(new_n13224_), .A2(new_n13221_), .B(new_n13229_), .ZN(new_n13243_));
  AOI21_X1   g12986(.A1(new_n13243_), .A2(new_n13242_), .B(new_n13039_), .ZN(new_n13244_));
  OAI21_X1   g12987(.A1(new_n13224_), .A2(new_n13221_), .B(new_n13233_), .ZN(new_n13245_));
  NAND3_X1   g12988(.A1(new_n13231_), .A2(new_n13232_), .A3(new_n13229_), .ZN(new_n13246_));
  AOI21_X1   g12989(.A1(new_n13245_), .A2(new_n13246_), .B(new_n13040_), .ZN(new_n13247_));
  NOR3_X1    g12990(.A1(new_n13241_), .A2(new_n13244_), .A3(new_n13247_), .ZN(new_n13248_));
  OAI21_X1   g12991(.A1(new_n13239_), .A2(new_n13248_), .B(new_n1750_), .ZN(new_n13249_));
  OAI21_X1   g12992(.A1(new_n13244_), .A2(new_n13247_), .B(new_n13241_), .ZN(new_n13250_));
  NAND3_X1   g12993(.A1(new_n13038_), .A2(new_n13235_), .A3(new_n13238_), .ZN(new_n13251_));
  NAND3_X1   g12994(.A1(new_n13251_), .A2(new_n13250_), .A3(\a[26] ), .ZN(new_n13252_));
  AOI21_X1   g12995(.A1(new_n13249_), .A2(new_n13252_), .B(new_n13032_), .ZN(new_n13253_));
  AOI21_X1   g12996(.A1(new_n13251_), .A2(new_n13250_), .B(\a[26] ), .ZN(new_n13254_));
  NOR3_X1    g12997(.A1(new_n13239_), .A2(new_n13248_), .A3(new_n1750_), .ZN(new_n13255_));
  NOR3_X1    g12998(.A1(new_n13254_), .A2(new_n13255_), .A3(new_n13031_), .ZN(new_n13256_));
  OAI22_X1   g12999(.A1(new_n1444_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n1439_), .ZN(new_n13257_));
  NAND2_X1   g13000(.A1(new_n2098_), .A2(\b[51] ), .ZN(new_n13258_));
  AOI21_X1   g13001(.A1(new_n13257_), .A2(new_n13258_), .B(new_n1447_), .ZN(new_n13259_));
  NAND2_X1   g13002(.A1(new_n6219_), .A2(new_n13259_), .ZN(new_n13260_));
  XOR2_X1    g13003(.A1(new_n13260_), .A2(\a[23] ), .Z(new_n13261_));
  INV_X1     g13004(.I(new_n13261_), .ZN(new_n13262_));
  OAI21_X1   g13005(.A1(new_n13256_), .A2(new_n13253_), .B(new_n13262_), .ZN(new_n13263_));
  OAI21_X1   g13006(.A1(new_n13254_), .A2(new_n13255_), .B(new_n13031_), .ZN(new_n13264_));
  NAND3_X1   g13007(.A1(new_n13249_), .A2(new_n13252_), .A3(new_n13032_), .ZN(new_n13265_));
  NAND3_X1   g13008(.A1(new_n13264_), .A2(new_n13265_), .A3(new_n13261_), .ZN(new_n13266_));
  AOI22_X1   g13009(.A1(new_n13263_), .A2(new_n13266_), .B1(new_n12898_), .B2(new_n13028_), .ZN(new_n13267_));
  NAND2_X1   g13010(.A1(new_n13028_), .A2(new_n12898_), .ZN(new_n13268_));
  NAND3_X1   g13011(.A1(new_n13264_), .A2(new_n13265_), .A3(new_n13262_), .ZN(new_n13269_));
  OAI21_X1   g13012(.A1(new_n13256_), .A2(new_n13253_), .B(new_n13261_), .ZN(new_n13270_));
  AOI21_X1   g13013(.A1(new_n13270_), .A2(new_n13269_), .B(new_n13268_), .ZN(new_n13271_));
  OAI21_X1   g13014(.A1(new_n13267_), .A2(new_n13271_), .B(new_n13027_), .ZN(new_n13272_));
  INV_X1     g13015(.I(new_n13272_), .ZN(new_n13273_));
  NOR3_X1    g13016(.A1(new_n13267_), .A2(new_n13027_), .A3(new_n13271_), .ZN(new_n13274_));
  OAI21_X1   g13017(.A1(new_n13273_), .A2(new_n13274_), .B(new_n1158_), .ZN(new_n13275_));
  INV_X1     g13018(.I(new_n13274_), .ZN(new_n13276_));
  NAND3_X1   g13019(.A1(new_n13276_), .A2(new_n13272_), .A3(\a[20] ), .ZN(new_n13277_));
  AOI21_X1   g13020(.A1(new_n13275_), .A2(new_n13277_), .B(new_n13023_), .ZN(new_n13278_));
  INV_X1     g13021(.I(new_n13023_), .ZN(new_n13279_));
  AOI21_X1   g13022(.A1(new_n13276_), .A2(new_n13272_), .B(\a[20] ), .ZN(new_n13280_));
  NOR3_X1    g13023(.A1(new_n13273_), .A2(new_n1158_), .A3(new_n13274_), .ZN(new_n13281_));
  NOR3_X1    g13024(.A1(new_n13281_), .A2(new_n13280_), .A3(new_n13279_), .ZN(new_n13282_));
  OAI22_X1   g13025(.A1(new_n940_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n935_), .ZN(new_n13283_));
  NAND2_X1   g13026(.A1(new_n1458_), .A2(\b[57] ), .ZN(new_n13284_));
  AOI21_X1   g13027(.A1(new_n13283_), .A2(new_n13284_), .B(new_n943_), .ZN(new_n13285_));
  NAND2_X1   g13028(.A1(new_n7895_), .A2(new_n13285_), .ZN(new_n13286_));
  XOR2_X1    g13029(.A1(new_n13286_), .A2(\a[17] ), .Z(new_n13287_));
  NOR3_X1    g13030(.A1(new_n13282_), .A2(new_n13278_), .A3(new_n13287_), .ZN(new_n13288_));
  OAI21_X1   g13031(.A1(new_n13281_), .A2(new_n13280_), .B(new_n13279_), .ZN(new_n13289_));
  NAND3_X1   g13032(.A1(new_n13275_), .A2(new_n13277_), .A3(new_n13023_), .ZN(new_n13290_));
  INV_X1     g13033(.I(new_n13287_), .ZN(new_n13291_));
  AOI21_X1   g13034(.A1(new_n13289_), .A2(new_n13290_), .B(new_n13291_), .ZN(new_n13292_));
  OAI21_X1   g13035(.A1(new_n13288_), .A2(new_n13292_), .B(new_n13020_), .ZN(new_n13293_));
  AOI21_X1   g13036(.A1(new_n13289_), .A2(new_n13290_), .B(new_n13287_), .ZN(new_n13294_));
  NOR3_X1    g13037(.A1(new_n13282_), .A2(new_n13278_), .A3(new_n13291_), .ZN(new_n13295_));
  OAI21_X1   g13038(.A1(new_n13295_), .A2(new_n13294_), .B(new_n13019_), .ZN(new_n13296_));
  AOI21_X1   g13039(.A1(new_n13293_), .A2(new_n13296_), .B(new_n13018_), .ZN(new_n13297_));
  AOI21_X1   g13040(.A1(new_n12950_), .A2(new_n12948_), .B(new_n12965_), .ZN(new_n13298_));
  NAND3_X1   g13041(.A1(new_n13289_), .A2(new_n13290_), .A3(new_n13291_), .ZN(new_n13299_));
  OAI21_X1   g13042(.A1(new_n13282_), .A2(new_n13278_), .B(new_n13287_), .ZN(new_n13300_));
  AOI21_X1   g13043(.A1(new_n13300_), .A2(new_n13299_), .B(new_n13019_), .ZN(new_n13301_));
  OAI21_X1   g13044(.A1(new_n13282_), .A2(new_n13278_), .B(new_n13291_), .ZN(new_n13302_));
  NAND3_X1   g13045(.A1(new_n13289_), .A2(new_n13290_), .A3(new_n13287_), .ZN(new_n13303_));
  AOI21_X1   g13046(.A1(new_n13302_), .A2(new_n13303_), .B(new_n13020_), .ZN(new_n13304_));
  NOR3_X1    g13047(.A1(new_n13298_), .A2(new_n13301_), .A3(new_n13304_), .ZN(new_n13305_));
  OAI21_X1   g13048(.A1(new_n13297_), .A2(new_n13305_), .B(new_n747_), .ZN(new_n13306_));
  OAI21_X1   g13049(.A1(new_n13301_), .A2(new_n13304_), .B(new_n13298_), .ZN(new_n13307_));
  NAND3_X1   g13050(.A1(new_n13018_), .A2(new_n13293_), .A3(new_n13296_), .ZN(new_n13308_));
  NAND3_X1   g13051(.A1(new_n13307_), .A2(new_n13308_), .A3(\a[14] ), .ZN(new_n13309_));
  AOI21_X1   g13052(.A1(new_n13306_), .A2(new_n13309_), .B(new_n13017_), .ZN(new_n13310_));
  AOI21_X1   g13053(.A1(new_n13307_), .A2(new_n13308_), .B(\a[14] ), .ZN(new_n13311_));
  NOR3_X1    g13054(.A1(new_n13297_), .A2(new_n13305_), .A3(new_n747_), .ZN(new_n13312_));
  NOR3_X1    g13055(.A1(new_n13311_), .A2(new_n13312_), .A3(new_n13016_), .ZN(new_n13313_));
  OAI21_X1   g13056(.A1(new_n13310_), .A2(new_n13313_), .B(new_n13013_), .ZN(new_n13314_));
  OAI21_X1   g13057(.A1(new_n13311_), .A2(new_n13312_), .B(new_n13016_), .ZN(new_n13315_));
  NAND3_X1   g13058(.A1(new_n13306_), .A2(new_n13309_), .A3(new_n13017_), .ZN(new_n13316_));
  NAND3_X1   g13059(.A1(new_n13315_), .A2(new_n13316_), .A3(new_n13012_), .ZN(new_n13317_));
  AOI21_X1   g13060(.A1(new_n13314_), .A2(new_n13317_), .B(\a[11] ), .ZN(new_n13318_));
  AOI21_X1   g13061(.A1(new_n13315_), .A2(new_n13316_), .B(new_n13012_), .ZN(new_n13319_));
  NOR3_X1    g13062(.A1(new_n13310_), .A2(new_n13313_), .A3(new_n13013_), .ZN(new_n13320_));
  NOR3_X1    g13063(.A1(new_n13320_), .A2(new_n13319_), .A3(new_n572_), .ZN(new_n13321_));
  OAI21_X1   g13064(.A1(new_n13321_), .A2(new_n13318_), .B(new_n13011_), .ZN(new_n13322_));
  INV_X1     g13065(.I(new_n13011_), .ZN(new_n13323_));
  OAI21_X1   g13066(.A1(new_n13320_), .A2(new_n13319_), .B(new_n572_), .ZN(new_n13324_));
  NAND3_X1   g13067(.A1(new_n13314_), .A2(new_n13317_), .A3(\a[11] ), .ZN(new_n13325_));
  NAND3_X1   g13068(.A1(new_n13324_), .A2(new_n13325_), .A3(new_n13323_), .ZN(new_n13326_));
  NAND2_X1   g13069(.A1(new_n13322_), .A2(new_n13326_), .ZN(new_n13327_));
  XOR2_X1    g13070(.A1(new_n13327_), .A2(new_n13010_), .Z(new_n13328_));
  AOI21_X1   g13071(.A1(new_n13322_), .A2(new_n13326_), .B(new_n13010_), .ZN(new_n13329_));
  NAND3_X1   g13072(.A1(new_n13322_), .A2(new_n13326_), .A3(new_n13010_), .ZN(new_n13330_));
  INV_X1     g13073(.I(new_n13330_), .ZN(new_n13331_));
  OAI21_X1   g13074(.A1(new_n13329_), .A2(new_n13331_), .B(new_n13007_), .ZN(new_n13332_));
  OAI21_X1   g13075(.A1(new_n13007_), .A2(new_n13328_), .B(new_n13332_), .ZN(\f[74] ));
  OAI21_X1   g13076(.A1(new_n13310_), .A2(new_n13313_), .B(new_n13012_), .ZN(new_n13334_));
  INV_X1     g13077(.I(new_n13334_), .ZN(new_n13335_));
  NOR3_X1    g13078(.A1(new_n13310_), .A2(new_n13313_), .A3(new_n13012_), .ZN(new_n13336_));
  XOR2_X1    g13079(.A1(new_n13011_), .A2(\a[11] ), .Z(new_n13337_));
  NOR2_X1    g13080(.A1(new_n13336_), .A2(new_n13337_), .ZN(new_n13338_));
  XOR2_X1    g13081(.A1(new_n13016_), .A2(\a[14] ), .Z(new_n13339_));
  NOR3_X1    g13082(.A1(new_n13301_), .A2(new_n13304_), .A3(new_n13339_), .ZN(new_n13340_));
  INV_X1     g13083(.I(new_n13339_), .ZN(new_n13341_));
  AOI21_X1   g13084(.A1(new_n13293_), .A2(new_n13296_), .B(new_n13341_), .ZN(new_n13342_));
  OAI22_X1   g13085(.A1(new_n13342_), .A2(new_n13340_), .B1(new_n13298_), .B2(new_n13339_), .ZN(new_n13343_));
  NOR2_X1    g13086(.A1(new_n13295_), .A2(new_n13019_), .ZN(new_n13344_));
  NOR2_X1    g13087(.A1(new_n13344_), .A2(new_n13294_), .ZN(new_n13345_));
  NOR2_X1    g13088(.A1(new_n13267_), .A2(new_n13271_), .ZN(new_n13346_));
  NOR2_X1    g13089(.A1(new_n13346_), .A2(new_n13027_), .ZN(new_n13347_));
  XOR2_X1    g13090(.A1(new_n13023_), .A2(new_n1158_), .Z(new_n13348_));
  AOI21_X1   g13091(.A1(new_n13346_), .A2(new_n13027_), .B(new_n13348_), .ZN(new_n13349_));
  NOR2_X1    g13092(.A1(new_n13349_), .A2(new_n13347_), .ZN(new_n13350_));
  NAND2_X1   g13093(.A1(new_n13266_), .A2(new_n13268_), .ZN(new_n13351_));
  NAND2_X1   g13094(.A1(new_n13351_), .A2(new_n13263_), .ZN(new_n13352_));
  XOR2_X1    g13095(.A1(new_n13031_), .A2(\a[26] ), .Z(new_n13353_));
  NOR3_X1    g13096(.A1(new_n13244_), .A2(new_n13247_), .A3(new_n13353_), .ZN(new_n13354_));
  INV_X1     g13097(.I(new_n13353_), .ZN(new_n13355_));
  AOI21_X1   g13098(.A1(new_n13235_), .A2(new_n13238_), .B(new_n13355_), .ZN(new_n13356_));
  OAI22_X1   g13099(.A1(new_n13356_), .A2(new_n13354_), .B1(new_n13241_), .B2(new_n13353_), .ZN(new_n13357_));
  AOI21_X1   g13100(.A1(new_n13040_), .A2(new_n13246_), .B(new_n13236_), .ZN(new_n13358_));
  INV_X1     g13101(.I(new_n13358_), .ZN(new_n13359_));
  OAI21_X1   g13102(.A1(new_n13212_), .A2(new_n13215_), .B(new_n13045_), .ZN(new_n13360_));
  XOR2_X1    g13103(.A1(new_n13043_), .A2(new_n2442_), .Z(new_n13361_));
  NAND4_X1   g13104(.A1(new_n13204_), .A2(new_n13207_), .A3(new_n13209_), .A4(new_n13361_), .ZN(new_n13362_));
  NAND2_X1   g13105(.A1(new_n13362_), .A2(new_n13360_), .ZN(new_n13363_));
  INV_X1     g13106(.I(new_n13363_), .ZN(new_n13364_));
  AOI21_X1   g13107(.A1(new_n13047_), .A2(new_n13210_), .B(new_n13203_), .ZN(new_n13365_));
  AOI21_X1   g13108(.A1(new_n13055_), .A2(new_n13201_), .B(new_n13193_), .ZN(new_n13366_));
  INV_X1     g13109(.I(new_n13366_), .ZN(new_n13367_));
  INV_X1     g13110(.I(new_n13185_), .ZN(new_n13368_));
  AOI21_X1   g13111(.A1(new_n13181_), .A2(new_n13368_), .B(new_n13184_), .ZN(new_n13369_));
  INV_X1     g13112(.I(new_n13369_), .ZN(new_n13370_));
  INV_X1     g13113(.I(new_n13166_), .ZN(new_n13371_));
  AOI21_X1   g13114(.A1(new_n13165_), .A2(new_n13167_), .B(new_n13371_), .ZN(new_n13372_));
  INV_X1     g13115(.I(new_n13154_), .ZN(new_n13373_));
  OAI21_X1   g13116(.A1(new_n13160_), .A2(new_n13155_), .B(new_n13373_), .ZN(new_n13374_));
  INV_X1     g13117(.I(new_n13374_), .ZN(new_n13375_));
  NAND2_X1   g13118(.A1(new_n13138_), .A2(new_n13137_), .ZN(new_n13376_));
  NAND2_X1   g13119(.A1(new_n13376_), .A2(new_n13140_), .ZN(new_n13377_));
  NAND2_X1   g13120(.A1(new_n13132_), .A2(new_n13129_), .ZN(new_n13378_));
  OAI22_X1   g13121(.A1(new_n5786_), .A2(new_n1709_), .B1(new_n1601_), .B2(new_n5792_), .ZN(new_n13379_));
  NAND2_X1   g13122(.A1(new_n6745_), .A2(\b[22] ), .ZN(new_n13380_));
  AOI21_X1   g13123(.A1(new_n13380_), .A2(new_n13379_), .B(new_n5796_), .ZN(new_n13381_));
  NAND2_X1   g13124(.A1(new_n1708_), .A2(new_n13381_), .ZN(new_n13382_));
  XOR2_X1    g13125(.A1(new_n13382_), .A2(\a[53] ), .Z(new_n13383_));
  NAND2_X1   g13126(.A1(new_n13122_), .A2(new_n13120_), .ZN(new_n13384_));
  NAND2_X1   g13127(.A1(new_n13384_), .A2(new_n13121_), .ZN(new_n13385_));
  INV_X1     g13128(.I(new_n13385_), .ZN(new_n13386_));
  INV_X1     g13129(.I(new_n13089_), .ZN(new_n13387_));
  OAI21_X1   g13130(.A1(new_n12730_), .A2(new_n13090_), .B(new_n13084_), .ZN(new_n13388_));
  NAND2_X1   g13131(.A1(new_n13388_), .A2(new_n13387_), .ZN(new_n13389_));
  OAI22_X1   g13132(.A1(new_n904_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n848_), .ZN(new_n13390_));
  NAND2_X1   g13133(.A1(new_n9644_), .A2(\b[13] ), .ZN(new_n13391_));
  AOI21_X1   g13134(.A1(new_n13391_), .A2(new_n13390_), .B(new_n8321_), .ZN(new_n13392_));
  NAND2_X1   g13135(.A1(new_n907_), .A2(new_n13392_), .ZN(new_n13393_));
  XOR2_X1    g13136(.A1(new_n13393_), .A2(\a[62] ), .Z(new_n13394_));
  NOR2_X1    g13137(.A1(new_n8985_), .A2(new_n717_), .ZN(new_n13395_));
  NOR2_X1    g13138(.A1(new_n9364_), .A2(new_n659_), .ZN(new_n13396_));
  XNOR2_X1   g13139(.A1(new_n13395_), .A2(new_n13396_), .ZN(new_n13397_));
  XOR2_X1    g13140(.A1(new_n13397_), .A2(\a[11] ), .Z(new_n13398_));
  NOR2_X1    g13141(.A1(new_n13398_), .A2(new_n12730_), .ZN(new_n13399_));
  NOR2_X1    g13142(.A1(new_n13397_), .A2(new_n572_), .ZN(new_n13400_));
  INV_X1     g13143(.I(new_n13400_), .ZN(new_n13401_));
  NAND2_X1   g13144(.A1(new_n13397_), .A2(new_n572_), .ZN(new_n13402_));
  AOI21_X1   g13145(.A1(new_n13401_), .A2(new_n13402_), .B(new_n12735_), .ZN(new_n13403_));
  NOR2_X1    g13146(.A1(new_n13399_), .A2(new_n13403_), .ZN(new_n13404_));
  INV_X1     g13147(.I(new_n13404_), .ZN(new_n13405_));
  NAND2_X1   g13148(.A1(new_n13394_), .A2(new_n13405_), .ZN(new_n13406_));
  INV_X1     g13149(.I(new_n13406_), .ZN(new_n13407_));
  NOR2_X1    g13150(.A1(new_n13394_), .A2(new_n13405_), .ZN(new_n13408_));
  OAI21_X1   g13151(.A1(new_n13407_), .A2(new_n13408_), .B(new_n13389_), .ZN(new_n13409_));
  INV_X1     g13152(.I(new_n13389_), .ZN(new_n13410_));
  XOR2_X1    g13153(.A1(new_n13394_), .A2(new_n13405_), .Z(new_n13411_));
  NAND2_X1   g13154(.A1(new_n13410_), .A2(new_n13411_), .ZN(new_n13412_));
  NAND2_X1   g13155(.A1(new_n13412_), .A2(new_n13409_), .ZN(new_n13413_));
  OAI22_X1   g13156(.A1(new_n1124_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1044_), .ZN(new_n13414_));
  NAND2_X1   g13157(.A1(new_n8628_), .A2(\b[16] ), .ZN(new_n13415_));
  AOI21_X1   g13158(.A1(new_n13415_), .A2(new_n13414_), .B(new_n7354_), .ZN(new_n13416_));
  NAND2_X1   g13159(.A1(new_n1123_), .A2(new_n13416_), .ZN(new_n13417_));
  XOR2_X1    g13160(.A1(new_n13417_), .A2(\a[59] ), .Z(new_n13418_));
  INV_X1     g13161(.I(new_n13418_), .ZN(new_n13419_));
  NAND2_X1   g13162(.A1(new_n13111_), .A2(new_n13096_), .ZN(new_n13420_));
  NAND2_X1   g13163(.A1(new_n13420_), .A2(new_n13109_), .ZN(new_n13421_));
  XOR2_X1    g13164(.A1(new_n13421_), .A2(new_n13419_), .Z(new_n13422_));
  NAND2_X1   g13165(.A1(new_n13422_), .A2(new_n13413_), .ZN(new_n13423_));
  INV_X1     g13166(.I(new_n13413_), .ZN(new_n13424_));
  AOI21_X1   g13167(.A1(new_n13420_), .A2(new_n13109_), .B(new_n13418_), .ZN(new_n13425_));
  NOR2_X1    g13168(.A1(new_n13421_), .A2(new_n13419_), .ZN(new_n13426_));
  OAI21_X1   g13169(.A1(new_n13425_), .A2(new_n13426_), .B(new_n13424_), .ZN(new_n13427_));
  NAND2_X1   g13170(.A1(new_n13423_), .A2(new_n13427_), .ZN(new_n13428_));
  OAI22_X1   g13171(.A1(new_n6721_), .A2(new_n1305_), .B1(new_n6723_), .B2(new_n1393_), .ZN(new_n13429_));
  NAND2_X1   g13172(.A1(new_n7617_), .A2(\b[19] ), .ZN(new_n13430_));
  AOI21_X1   g13173(.A1(new_n13430_), .A2(new_n13429_), .B(new_n6731_), .ZN(new_n13431_));
  NAND2_X1   g13174(.A1(new_n1396_), .A2(new_n13431_), .ZN(new_n13432_));
  XOR2_X1    g13175(.A1(new_n13432_), .A2(\a[56] ), .Z(new_n13433_));
  INV_X1     g13176(.I(new_n13433_), .ZN(new_n13434_));
  XOR2_X1    g13177(.A1(new_n13428_), .A2(new_n13434_), .Z(new_n13435_));
  NOR2_X1    g13178(.A1(new_n13428_), .A2(new_n13433_), .ZN(new_n13436_));
  INV_X1     g13179(.I(new_n13428_), .ZN(new_n13437_));
  NOR2_X1    g13180(.A1(new_n13437_), .A2(new_n13434_), .ZN(new_n13438_));
  OAI21_X1   g13181(.A1(new_n13438_), .A2(new_n13436_), .B(new_n13386_), .ZN(new_n13439_));
  OAI21_X1   g13182(.A1(new_n13386_), .A2(new_n13435_), .B(new_n13439_), .ZN(new_n13440_));
  NAND2_X1   g13183(.A1(new_n13440_), .A2(new_n13383_), .ZN(new_n13441_));
  OR2_X2     g13184(.A1(new_n13440_), .A2(new_n13383_), .Z(new_n13442_));
  AOI22_X1   g13185(.A1(new_n13442_), .A2(new_n13441_), .B1(new_n13131_), .B2(new_n13378_), .ZN(new_n13443_));
  NAND2_X1   g13186(.A1(new_n13378_), .A2(new_n13131_), .ZN(new_n13444_));
  XNOR2_X1   g13187(.A1(new_n13440_), .A2(new_n13383_), .ZN(new_n13445_));
  NOR2_X1    g13188(.A1(new_n13445_), .A2(new_n13444_), .ZN(new_n13446_));
  NOR2_X1    g13189(.A1(new_n13446_), .A2(new_n13443_), .ZN(new_n13447_));
  OAI22_X1   g13190(.A1(new_n5228_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n5225_), .ZN(new_n13448_));
  NAND2_X1   g13191(.A1(new_n5387_), .A2(\b[25] ), .ZN(new_n13449_));
  AOI21_X1   g13192(.A1(new_n13448_), .A2(new_n13449_), .B(new_n5231_), .ZN(new_n13450_));
  NAND2_X1   g13193(.A1(new_n2042_), .A2(new_n13450_), .ZN(new_n13451_));
  XOR2_X1    g13194(.A1(new_n13451_), .A2(\a[50] ), .Z(new_n13452_));
  XOR2_X1    g13195(.A1(new_n13447_), .A2(new_n13452_), .Z(new_n13453_));
  NAND2_X1   g13196(.A1(new_n13453_), .A2(new_n13377_), .ZN(new_n13454_));
  INV_X1     g13197(.I(new_n13377_), .ZN(new_n13455_));
  NOR2_X1    g13198(.A1(new_n13447_), .A2(new_n13452_), .ZN(new_n13456_));
  NAND2_X1   g13199(.A1(new_n13447_), .A2(new_n13452_), .ZN(new_n13457_));
  INV_X1     g13200(.I(new_n13457_), .ZN(new_n13458_));
  OAI21_X1   g13201(.A1(new_n13458_), .A2(new_n13456_), .B(new_n13455_), .ZN(new_n13459_));
  OAI22_X1   g13202(.A1(new_n4711_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n4706_), .ZN(new_n13460_));
  NAND2_X1   g13203(.A1(new_n5814_), .A2(\b[28] ), .ZN(new_n13461_));
  AOI21_X1   g13204(.A1(new_n13460_), .A2(new_n13461_), .B(new_n4714_), .ZN(new_n13462_));
  NAND2_X1   g13205(.A1(new_n2404_), .A2(new_n13462_), .ZN(new_n13463_));
  XOR2_X1    g13206(.A1(new_n13463_), .A2(\a[47] ), .Z(new_n13464_));
  INV_X1     g13207(.I(new_n13464_), .ZN(new_n13465_));
  NAND3_X1   g13208(.A1(new_n13454_), .A2(new_n13459_), .A3(new_n13465_), .ZN(new_n13466_));
  AOI21_X1   g13209(.A1(new_n13454_), .A2(new_n13459_), .B(new_n13465_), .ZN(new_n13467_));
  INV_X1     g13210(.I(new_n13467_), .ZN(new_n13468_));
  AOI21_X1   g13211(.A1(new_n13468_), .A2(new_n13466_), .B(new_n13375_), .ZN(new_n13469_));
  INV_X1     g13212(.I(new_n13469_), .ZN(new_n13470_));
  NAND2_X1   g13213(.A1(new_n13454_), .A2(new_n13459_), .ZN(new_n13471_));
  NAND2_X1   g13214(.A1(new_n13471_), .A2(new_n13465_), .ZN(new_n13472_));
  INV_X1     g13215(.I(new_n13472_), .ZN(new_n13473_));
  NOR2_X1    g13216(.A1(new_n13471_), .A2(new_n13465_), .ZN(new_n13474_));
  OAI21_X1   g13217(.A1(new_n13473_), .A2(new_n13474_), .B(new_n13375_), .ZN(new_n13475_));
  OAI22_X1   g13218(.A1(new_n4208_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n4203_), .ZN(new_n13476_));
  NAND2_X1   g13219(.A1(new_n5244_), .A2(\b[31] ), .ZN(new_n13477_));
  AOI21_X1   g13220(.A1(new_n13476_), .A2(new_n13477_), .B(new_n4211_), .ZN(new_n13478_));
  NAND2_X1   g13221(.A1(new_n2797_), .A2(new_n13478_), .ZN(new_n13479_));
  XOR2_X1    g13222(.A1(new_n13479_), .A2(\a[44] ), .Z(new_n13480_));
  AOI21_X1   g13223(.A1(new_n13470_), .A2(new_n13475_), .B(new_n13480_), .ZN(new_n13481_));
  INV_X1     g13224(.I(new_n13481_), .ZN(new_n13482_));
  NAND3_X1   g13225(.A1(new_n13470_), .A2(new_n13475_), .A3(new_n13480_), .ZN(new_n13483_));
  AOI21_X1   g13226(.A1(new_n13482_), .A2(new_n13483_), .B(new_n13372_), .ZN(new_n13484_));
  INV_X1     g13227(.I(new_n13372_), .ZN(new_n13485_));
  INV_X1     g13228(.I(new_n13480_), .ZN(new_n13486_));
  NAND3_X1   g13229(.A1(new_n13470_), .A2(new_n13475_), .A3(new_n13486_), .ZN(new_n13487_));
  AOI21_X1   g13230(.A1(new_n13470_), .A2(new_n13475_), .B(new_n13486_), .ZN(new_n13488_));
  INV_X1     g13231(.I(new_n13488_), .ZN(new_n13489_));
  AOI21_X1   g13232(.A1(new_n13489_), .A2(new_n13487_), .B(new_n13485_), .ZN(new_n13490_));
  OAI22_X1   g13233(.A1(new_n3736_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n3731_), .ZN(new_n13491_));
  NAND2_X1   g13234(.A1(new_n4730_), .A2(\b[34] ), .ZN(new_n13492_));
  AOI21_X1   g13235(.A1(new_n13491_), .A2(new_n13492_), .B(new_n3739_), .ZN(new_n13493_));
  NAND2_X1   g13236(.A1(new_n3246_), .A2(new_n13493_), .ZN(new_n13494_));
  XOR2_X1    g13237(.A1(new_n13494_), .A2(\a[41] ), .Z(new_n13495_));
  NOR3_X1    g13238(.A1(new_n13484_), .A2(new_n13490_), .A3(new_n13495_), .ZN(new_n13496_));
  INV_X1     g13239(.I(new_n13483_), .ZN(new_n13497_));
  OAI21_X1   g13240(.A1(new_n13497_), .A2(new_n13481_), .B(new_n13485_), .ZN(new_n13498_));
  INV_X1     g13241(.I(new_n13487_), .ZN(new_n13499_));
  OAI21_X1   g13242(.A1(new_n13499_), .A2(new_n13488_), .B(new_n13372_), .ZN(new_n13500_));
  INV_X1     g13243(.I(new_n13495_), .ZN(new_n13501_));
  AOI21_X1   g13244(.A1(new_n13498_), .A2(new_n13500_), .B(new_n13501_), .ZN(new_n13502_));
  OAI21_X1   g13245(.A1(new_n13496_), .A2(new_n13502_), .B(new_n13370_), .ZN(new_n13503_));
  AOI21_X1   g13246(.A1(new_n13498_), .A2(new_n13500_), .B(new_n13495_), .ZN(new_n13504_));
  NOR3_X1    g13247(.A1(new_n13484_), .A2(new_n13490_), .A3(new_n13501_), .ZN(new_n13505_));
  OAI21_X1   g13248(.A1(new_n13505_), .A2(new_n13504_), .B(new_n13369_), .ZN(new_n13506_));
  OAI22_X1   g13249(.A1(new_n3298_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n3293_), .ZN(new_n13507_));
  NAND2_X1   g13250(.A1(new_n4227_), .A2(\b[37] ), .ZN(new_n13508_));
  AOI21_X1   g13251(.A1(new_n13507_), .A2(new_n13508_), .B(new_n3301_), .ZN(new_n13509_));
  NAND2_X1   g13252(.A1(new_n3700_), .A2(new_n13509_), .ZN(new_n13510_));
  XOR2_X1    g13253(.A1(new_n13510_), .A2(\a[38] ), .Z(new_n13511_));
  INV_X1     g13254(.I(new_n13511_), .ZN(new_n13512_));
  NAND3_X1   g13255(.A1(new_n13503_), .A2(new_n13506_), .A3(new_n13512_), .ZN(new_n13513_));
  INV_X1     g13256(.I(new_n13513_), .ZN(new_n13514_));
  AOI21_X1   g13257(.A1(new_n13503_), .A2(new_n13506_), .B(new_n13512_), .ZN(new_n13515_));
  OAI21_X1   g13258(.A1(new_n13514_), .A2(new_n13515_), .B(new_n13367_), .ZN(new_n13516_));
  AOI21_X1   g13259(.A1(new_n13503_), .A2(new_n13506_), .B(new_n13511_), .ZN(new_n13517_));
  NAND3_X1   g13260(.A1(new_n13498_), .A2(new_n13500_), .A3(new_n13501_), .ZN(new_n13518_));
  INV_X1     g13261(.I(new_n13502_), .ZN(new_n13519_));
  AOI21_X1   g13262(.A1(new_n13519_), .A2(new_n13518_), .B(new_n13369_), .ZN(new_n13520_));
  OAI21_X1   g13263(.A1(new_n13484_), .A2(new_n13490_), .B(new_n13501_), .ZN(new_n13521_));
  NAND3_X1   g13264(.A1(new_n13498_), .A2(new_n13500_), .A3(new_n13495_), .ZN(new_n13522_));
  AOI21_X1   g13265(.A1(new_n13521_), .A2(new_n13522_), .B(new_n13370_), .ZN(new_n13523_));
  NOR3_X1    g13266(.A1(new_n13520_), .A2(new_n13523_), .A3(new_n13512_), .ZN(new_n13524_));
  OAI21_X1   g13267(.A1(new_n13524_), .A2(new_n13517_), .B(new_n13366_), .ZN(new_n13525_));
  OAI22_X1   g13268(.A1(new_n2846_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n2841_), .ZN(new_n13526_));
  NAND2_X1   g13269(.A1(new_n3755_), .A2(\b[40] ), .ZN(new_n13527_));
  AOI21_X1   g13270(.A1(new_n13526_), .A2(new_n13527_), .B(new_n2849_), .ZN(new_n13528_));
  NAND2_X1   g13271(.A1(new_n4017_), .A2(new_n13528_), .ZN(new_n13529_));
  XOR2_X1    g13272(.A1(new_n13529_), .A2(\a[35] ), .Z(new_n13530_));
  INV_X1     g13273(.I(new_n13530_), .ZN(new_n13531_));
  NAND3_X1   g13274(.A1(new_n13516_), .A2(new_n13525_), .A3(new_n13531_), .ZN(new_n13532_));
  OAI21_X1   g13275(.A1(new_n13520_), .A2(new_n13523_), .B(new_n13511_), .ZN(new_n13533_));
  AOI21_X1   g13276(.A1(new_n13533_), .A2(new_n13513_), .B(new_n13366_), .ZN(new_n13534_));
  OAI21_X1   g13277(.A1(new_n13520_), .A2(new_n13523_), .B(new_n13512_), .ZN(new_n13535_));
  NAND3_X1   g13278(.A1(new_n13503_), .A2(new_n13506_), .A3(new_n13511_), .ZN(new_n13536_));
  AOI21_X1   g13279(.A1(new_n13535_), .A2(new_n13536_), .B(new_n13367_), .ZN(new_n13537_));
  OAI21_X1   g13280(.A1(new_n13534_), .A2(new_n13537_), .B(new_n13530_), .ZN(new_n13538_));
  AOI21_X1   g13281(.A1(new_n13532_), .A2(new_n13538_), .B(new_n13365_), .ZN(new_n13539_));
  INV_X1     g13282(.I(new_n13365_), .ZN(new_n13540_));
  OAI21_X1   g13283(.A1(new_n13534_), .A2(new_n13537_), .B(new_n13531_), .ZN(new_n13541_));
  NAND3_X1   g13284(.A1(new_n13516_), .A2(new_n13525_), .A3(new_n13530_), .ZN(new_n13542_));
  AOI21_X1   g13285(.A1(new_n13542_), .A2(new_n13541_), .B(new_n13540_), .ZN(new_n13543_));
  OAI22_X1   g13286(.A1(new_n2452_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n2447_), .ZN(new_n13544_));
  NAND2_X1   g13287(.A1(new_n3312_), .A2(\b[43] ), .ZN(new_n13545_));
  AOI21_X1   g13288(.A1(new_n13544_), .A2(new_n13545_), .B(new_n2455_), .ZN(new_n13546_));
  NAND2_X1   g13289(.A1(new_n4513_), .A2(new_n13546_), .ZN(new_n13547_));
  XOR2_X1    g13290(.A1(new_n13547_), .A2(\a[32] ), .Z(new_n13548_));
  INV_X1     g13291(.I(new_n13548_), .ZN(new_n13549_));
  OAI21_X1   g13292(.A1(new_n13539_), .A2(new_n13543_), .B(new_n13549_), .ZN(new_n13550_));
  NOR3_X1    g13293(.A1(new_n13534_), .A2(new_n13537_), .A3(new_n13530_), .ZN(new_n13551_));
  AOI21_X1   g13294(.A1(new_n13516_), .A2(new_n13525_), .B(new_n13531_), .ZN(new_n13552_));
  OAI21_X1   g13295(.A1(new_n13552_), .A2(new_n13551_), .B(new_n13540_), .ZN(new_n13553_));
  AOI21_X1   g13296(.A1(new_n13516_), .A2(new_n13525_), .B(new_n13530_), .ZN(new_n13554_));
  NOR3_X1    g13297(.A1(new_n13534_), .A2(new_n13537_), .A3(new_n13531_), .ZN(new_n13555_));
  OAI21_X1   g13298(.A1(new_n13554_), .A2(new_n13555_), .B(new_n13365_), .ZN(new_n13556_));
  NAND3_X1   g13299(.A1(new_n13553_), .A2(new_n13556_), .A3(new_n13548_), .ZN(new_n13557_));
  AOI21_X1   g13300(.A1(new_n13550_), .A2(new_n13557_), .B(new_n13364_), .ZN(new_n13558_));
  NAND3_X1   g13301(.A1(new_n13553_), .A2(new_n13556_), .A3(new_n13549_), .ZN(new_n13559_));
  OAI21_X1   g13302(.A1(new_n13539_), .A2(new_n13543_), .B(new_n13548_), .ZN(new_n13560_));
  AOI21_X1   g13303(.A1(new_n13560_), .A2(new_n13559_), .B(new_n13363_), .ZN(new_n13561_));
  OAI22_X1   g13304(.A1(new_n2084_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n2079_), .ZN(new_n13562_));
  NAND2_X1   g13305(.A1(new_n2864_), .A2(\b[46] ), .ZN(new_n13563_));
  AOI21_X1   g13306(.A1(new_n13562_), .A2(new_n13563_), .B(new_n2087_), .ZN(new_n13564_));
  NAND2_X1   g13307(.A1(new_n5177_), .A2(new_n13564_), .ZN(new_n13565_));
  XOR2_X1    g13308(.A1(new_n13565_), .A2(\a[29] ), .Z(new_n13566_));
  NOR3_X1    g13309(.A1(new_n13558_), .A2(new_n13561_), .A3(new_n13566_), .ZN(new_n13567_));
  AOI21_X1   g13310(.A1(new_n13553_), .A2(new_n13556_), .B(new_n13548_), .ZN(new_n13568_));
  NOR3_X1    g13311(.A1(new_n13539_), .A2(new_n13543_), .A3(new_n13549_), .ZN(new_n13569_));
  OAI21_X1   g13312(.A1(new_n13568_), .A2(new_n13569_), .B(new_n13363_), .ZN(new_n13570_));
  NOR3_X1    g13313(.A1(new_n13539_), .A2(new_n13543_), .A3(new_n13548_), .ZN(new_n13571_));
  AOI21_X1   g13314(.A1(new_n13553_), .A2(new_n13556_), .B(new_n13549_), .ZN(new_n13572_));
  OAI21_X1   g13315(.A1(new_n13572_), .A2(new_n13571_), .B(new_n13364_), .ZN(new_n13573_));
  INV_X1     g13316(.I(new_n13566_), .ZN(new_n13574_));
  AOI21_X1   g13317(.A1(new_n13570_), .A2(new_n13573_), .B(new_n13574_), .ZN(new_n13575_));
  OAI21_X1   g13318(.A1(new_n13575_), .A2(new_n13567_), .B(new_n13359_), .ZN(new_n13576_));
  AOI21_X1   g13319(.A1(new_n13570_), .A2(new_n13573_), .B(new_n13566_), .ZN(new_n13577_));
  NOR3_X1    g13320(.A1(new_n13558_), .A2(new_n13561_), .A3(new_n13574_), .ZN(new_n13578_));
  OAI21_X1   g13321(.A1(new_n13577_), .A2(new_n13578_), .B(new_n13358_), .ZN(new_n13579_));
  OAI22_X1   g13322(.A1(new_n1760_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n1755_), .ZN(new_n13580_));
  NAND2_X1   g13323(.A1(new_n2470_), .A2(\b[49] ), .ZN(new_n13581_));
  AOI21_X1   g13324(.A1(new_n13580_), .A2(new_n13581_), .B(new_n1763_), .ZN(new_n13582_));
  NAND2_X1   g13325(.A1(new_n5741_), .A2(new_n13582_), .ZN(new_n13583_));
  XOR2_X1    g13326(.A1(new_n13583_), .A2(\a[26] ), .Z(new_n13584_));
  INV_X1     g13327(.I(new_n13584_), .ZN(new_n13585_));
  NAND3_X1   g13328(.A1(new_n13576_), .A2(new_n13579_), .A3(new_n13585_), .ZN(new_n13586_));
  NAND3_X1   g13329(.A1(new_n13570_), .A2(new_n13573_), .A3(new_n13574_), .ZN(new_n13587_));
  OAI21_X1   g13330(.A1(new_n13558_), .A2(new_n13561_), .B(new_n13566_), .ZN(new_n13588_));
  AOI21_X1   g13331(.A1(new_n13588_), .A2(new_n13587_), .B(new_n13358_), .ZN(new_n13589_));
  OAI21_X1   g13332(.A1(new_n13558_), .A2(new_n13561_), .B(new_n13574_), .ZN(new_n13590_));
  NAND3_X1   g13333(.A1(new_n13570_), .A2(new_n13573_), .A3(new_n13566_), .ZN(new_n13591_));
  AOI21_X1   g13334(.A1(new_n13590_), .A2(new_n13591_), .B(new_n13359_), .ZN(new_n13592_));
  OAI21_X1   g13335(.A1(new_n13589_), .A2(new_n13592_), .B(new_n13584_), .ZN(new_n13593_));
  AOI21_X1   g13336(.A1(new_n13593_), .A2(new_n13586_), .B(new_n13357_), .ZN(new_n13594_));
  INV_X1     g13337(.I(new_n13357_), .ZN(new_n13595_));
  OAI21_X1   g13338(.A1(new_n13589_), .A2(new_n13592_), .B(new_n13585_), .ZN(new_n13596_));
  NAND3_X1   g13339(.A1(new_n13576_), .A2(new_n13579_), .A3(new_n13584_), .ZN(new_n13597_));
  AOI21_X1   g13340(.A1(new_n13596_), .A2(new_n13597_), .B(new_n13595_), .ZN(new_n13598_));
  OAI22_X1   g13341(.A1(new_n1444_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n1439_), .ZN(new_n13599_));
  NAND2_X1   g13342(.A1(new_n2098_), .A2(\b[52] ), .ZN(new_n13600_));
  AOI21_X1   g13343(.A1(new_n13599_), .A2(new_n13600_), .B(new_n1447_), .ZN(new_n13601_));
  NAND2_X1   g13344(.A1(new_n6237_), .A2(new_n13601_), .ZN(new_n13602_));
  XOR2_X1    g13345(.A1(new_n13602_), .A2(\a[23] ), .Z(new_n13603_));
  NOR3_X1    g13346(.A1(new_n13594_), .A2(new_n13598_), .A3(new_n13603_), .ZN(new_n13604_));
  NOR3_X1    g13347(.A1(new_n13589_), .A2(new_n13592_), .A3(new_n13584_), .ZN(new_n13605_));
  AOI21_X1   g13348(.A1(new_n13576_), .A2(new_n13579_), .B(new_n13585_), .ZN(new_n13606_));
  OAI21_X1   g13349(.A1(new_n13606_), .A2(new_n13605_), .B(new_n13595_), .ZN(new_n13607_));
  AOI21_X1   g13350(.A1(new_n13576_), .A2(new_n13579_), .B(new_n13584_), .ZN(new_n13608_));
  NOR3_X1    g13351(.A1(new_n13589_), .A2(new_n13592_), .A3(new_n13585_), .ZN(new_n13609_));
  OAI21_X1   g13352(.A1(new_n13608_), .A2(new_n13609_), .B(new_n13357_), .ZN(new_n13610_));
  INV_X1     g13353(.I(new_n13603_), .ZN(new_n13611_));
  AOI21_X1   g13354(.A1(new_n13607_), .A2(new_n13610_), .B(new_n13611_), .ZN(new_n13612_));
  OAI21_X1   g13355(.A1(new_n13612_), .A2(new_n13604_), .B(new_n13352_), .ZN(new_n13613_));
  INV_X1     g13356(.I(new_n13352_), .ZN(new_n13614_));
  AOI21_X1   g13357(.A1(new_n13607_), .A2(new_n13610_), .B(new_n13603_), .ZN(new_n13615_));
  NOR3_X1    g13358(.A1(new_n13594_), .A2(new_n13598_), .A3(new_n13611_), .ZN(new_n13616_));
  OAI21_X1   g13359(.A1(new_n13615_), .A2(new_n13616_), .B(new_n13614_), .ZN(new_n13617_));
  OAI22_X1   g13360(.A1(new_n1168_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n1163_), .ZN(new_n13618_));
  NAND2_X1   g13361(.A1(new_n1774_), .A2(\b[55] ), .ZN(new_n13619_));
  AOI21_X1   g13362(.A1(new_n13618_), .A2(new_n13619_), .B(new_n1171_), .ZN(new_n13620_));
  NAND2_X1   g13363(.A1(new_n7308_), .A2(new_n13620_), .ZN(new_n13621_));
  XOR2_X1    g13364(.A1(new_n13621_), .A2(\a[20] ), .Z(new_n13622_));
  INV_X1     g13365(.I(new_n13622_), .ZN(new_n13623_));
  NAND3_X1   g13366(.A1(new_n13617_), .A2(new_n13613_), .A3(new_n13623_), .ZN(new_n13624_));
  NAND3_X1   g13367(.A1(new_n13607_), .A2(new_n13610_), .A3(new_n13611_), .ZN(new_n13625_));
  OAI21_X1   g13368(.A1(new_n13594_), .A2(new_n13598_), .B(new_n13603_), .ZN(new_n13626_));
  AOI21_X1   g13369(.A1(new_n13625_), .A2(new_n13626_), .B(new_n13614_), .ZN(new_n13627_));
  OAI21_X1   g13370(.A1(new_n13594_), .A2(new_n13598_), .B(new_n13611_), .ZN(new_n13628_));
  NAND3_X1   g13371(.A1(new_n13607_), .A2(new_n13610_), .A3(new_n13603_), .ZN(new_n13629_));
  AOI21_X1   g13372(.A1(new_n13628_), .A2(new_n13629_), .B(new_n13352_), .ZN(new_n13630_));
  OAI21_X1   g13373(.A1(new_n13627_), .A2(new_n13630_), .B(new_n13622_), .ZN(new_n13631_));
  AOI21_X1   g13374(.A1(new_n13631_), .A2(new_n13624_), .B(new_n13350_), .ZN(new_n13632_));
  INV_X1     g13375(.I(new_n13632_), .ZN(new_n13633_));
  INV_X1     g13376(.I(new_n13350_), .ZN(new_n13634_));
  OAI21_X1   g13377(.A1(new_n13627_), .A2(new_n13630_), .B(new_n13623_), .ZN(new_n13635_));
  NAND3_X1   g13378(.A1(new_n13617_), .A2(new_n13613_), .A3(new_n13622_), .ZN(new_n13636_));
  AOI21_X1   g13379(.A1(new_n13635_), .A2(new_n13636_), .B(new_n13634_), .ZN(new_n13637_));
  INV_X1     g13380(.I(new_n13637_), .ZN(new_n13638_));
  OAI22_X1   g13381(.A1(new_n940_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n935_), .ZN(new_n13639_));
  NAND2_X1   g13382(.A1(new_n1458_), .A2(\b[58] ), .ZN(new_n13640_));
  AOI21_X1   g13383(.A1(new_n13639_), .A2(new_n13640_), .B(new_n943_), .ZN(new_n13641_));
  NAND2_X1   g13384(.A1(new_n7929_), .A2(new_n13641_), .ZN(new_n13642_));
  XOR2_X1    g13385(.A1(new_n13642_), .A2(\a[17] ), .Z(new_n13643_));
  INV_X1     g13386(.I(new_n13643_), .ZN(new_n13644_));
  NAND3_X1   g13387(.A1(new_n13638_), .A2(new_n13633_), .A3(new_n13644_), .ZN(new_n13645_));
  OAI21_X1   g13388(.A1(new_n13637_), .A2(new_n13632_), .B(new_n13643_), .ZN(new_n13646_));
  AOI21_X1   g13389(.A1(new_n13645_), .A2(new_n13646_), .B(new_n13345_), .ZN(new_n13647_));
  INV_X1     g13390(.I(new_n13345_), .ZN(new_n13648_));
  AOI21_X1   g13391(.A1(new_n13638_), .A2(new_n13633_), .B(new_n13643_), .ZN(new_n13649_));
  NOR3_X1    g13392(.A1(new_n13637_), .A2(new_n13632_), .A3(new_n13644_), .ZN(new_n13650_));
  NOR2_X1    g13393(.A1(new_n13649_), .A2(new_n13650_), .ZN(new_n13651_));
  NOR2_X1    g13394(.A1(new_n13648_), .A2(new_n13651_), .ZN(new_n13652_));
  OAI22_X1   g13395(.A1(new_n757_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n752_), .ZN(new_n13653_));
  NAND2_X1   g13396(.A1(new_n1182_), .A2(\b[61] ), .ZN(new_n13654_));
  AOI21_X1   g13397(.A1(new_n13653_), .A2(new_n13654_), .B(new_n760_), .ZN(new_n13655_));
  NAND2_X1   g13398(.A1(new_n8963_), .A2(new_n13655_), .ZN(new_n13656_));
  XOR2_X1    g13399(.A1(new_n13656_), .A2(\a[14] ), .Z(new_n13657_));
  INV_X1     g13400(.I(new_n13657_), .ZN(new_n13658_));
  OAI21_X1   g13401(.A1(new_n13652_), .A2(new_n13647_), .B(new_n13658_), .ZN(new_n13659_));
  NAND2_X1   g13402(.A1(new_n13645_), .A2(new_n13646_), .ZN(new_n13660_));
  NAND2_X1   g13403(.A1(new_n13648_), .A2(new_n13660_), .ZN(new_n13661_));
  OAI21_X1   g13404(.A1(new_n13649_), .A2(new_n13650_), .B(new_n13345_), .ZN(new_n13662_));
  NAND3_X1   g13405(.A1(new_n13661_), .A2(new_n13662_), .A3(new_n13657_), .ZN(new_n13663_));
  AOI21_X1   g13406(.A1(new_n13659_), .A2(new_n13663_), .B(new_n13343_), .ZN(new_n13664_));
  INV_X1     g13407(.I(new_n13343_), .ZN(new_n13665_));
  NAND3_X1   g13408(.A1(new_n13661_), .A2(new_n13662_), .A3(new_n13658_), .ZN(new_n13666_));
  OAI21_X1   g13409(.A1(new_n13652_), .A2(new_n13647_), .B(new_n13657_), .ZN(new_n13667_));
  AOI21_X1   g13410(.A1(new_n13666_), .A2(new_n13667_), .B(new_n13665_), .ZN(new_n13668_));
  OAI22_X1   g13411(.A1(new_n13338_), .A2(new_n13335_), .B1(new_n13664_), .B2(new_n13668_), .ZN(new_n13669_));
  NAND3_X1   g13412(.A1(new_n13315_), .A2(new_n13316_), .A3(new_n13013_), .ZN(new_n13670_));
  INV_X1     g13413(.I(new_n13337_), .ZN(new_n13671_));
  NAND2_X1   g13414(.A1(new_n13670_), .A2(new_n13671_), .ZN(new_n13672_));
  NOR2_X1    g13415(.A1(new_n13668_), .A2(new_n13664_), .ZN(new_n13673_));
  NAND3_X1   g13416(.A1(new_n13672_), .A2(new_n13673_), .A3(new_n13334_), .ZN(new_n13674_));
  NAND2_X1   g13417(.A1(new_n13669_), .A2(new_n13674_), .ZN(new_n13675_));
  INV_X1     g13418(.I(new_n12671_), .ZN(new_n13676_));
  NAND2_X1   g13419(.A1(new_n12994_), .A2(new_n12996_), .ZN(new_n13677_));
  OAI21_X1   g13420(.A1(new_n13000_), .A2(new_n13002_), .B(new_n12998_), .ZN(new_n13678_));
  NAND3_X1   g13421(.A1(new_n12994_), .A2(new_n12988_), .A3(new_n12996_), .ZN(new_n13679_));
  AOI22_X1   g13422(.A1(new_n13678_), .A2(new_n13679_), .B1(new_n13677_), .B2(new_n13676_), .ZN(new_n13680_));
  NAND2_X1   g13423(.A1(new_n13680_), .A2(new_n13009_), .ZN(new_n13681_));
  XOR2_X1    g13424(.A1(new_n13681_), .A2(new_n13675_), .Z(new_n13682_));
  XOR2_X1    g13425(.A1(new_n13680_), .A2(new_n13009_), .Z(new_n13683_));
  NAND2_X1   g13426(.A1(new_n13683_), .A2(new_n13327_), .ZN(new_n13684_));
  XOR2_X1    g13427(.A1(new_n13682_), .A2(new_n13684_), .Z(\f[75] ));
  NAND2_X1   g13428(.A1(new_n13665_), .A2(new_n13663_), .ZN(new_n13686_));
  AND2_X2    g13429(.A1(new_n13686_), .A2(new_n13659_), .Z(new_n13687_));
  INV_X1     g13430(.I(new_n13645_), .ZN(new_n13688_));
  AOI21_X1   g13431(.A1(new_n13648_), .A2(new_n13646_), .B(new_n13688_), .ZN(new_n13689_));
  INV_X1     g13432(.I(new_n13689_), .ZN(new_n13690_));
  INV_X1     g13433(.I(new_n13635_), .ZN(new_n13691_));
  AOI21_X1   g13434(.A1(new_n13634_), .A2(new_n13636_), .B(new_n13691_), .ZN(new_n13692_));
  OAI22_X1   g13435(.A1(new_n1168_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n1163_), .ZN(new_n13693_));
  OAI21_X1   g13436(.A1(new_n6995_), .A2(new_n1255_), .B(new_n13693_), .ZN(new_n13694_));
  AOI21_X1   g13437(.A1(new_n7559_), .A2(new_n1170_), .B(new_n13694_), .ZN(new_n13695_));
  INV_X1     g13438(.I(new_n13695_), .ZN(new_n13696_));
  AOI21_X1   g13439(.A1(new_n13352_), .A2(new_n13626_), .B(new_n13604_), .ZN(new_n13697_));
  INV_X1     g13440(.I(new_n13697_), .ZN(new_n13698_));
  AOI21_X1   g13441(.A1(new_n13595_), .A2(new_n13597_), .B(new_n13608_), .ZN(new_n13699_));
  INV_X1     g13442(.I(new_n13699_), .ZN(new_n13700_));
  AOI21_X1   g13443(.A1(new_n13359_), .A2(new_n13588_), .B(new_n13567_), .ZN(new_n13701_));
  INV_X1     g13444(.I(new_n13701_), .ZN(new_n13702_));
  AOI21_X1   g13445(.A1(new_n13363_), .A2(new_n13560_), .B(new_n13571_), .ZN(new_n13703_));
  INV_X1     g13446(.I(new_n13703_), .ZN(new_n13704_));
  AOI21_X1   g13447(.A1(new_n13367_), .A2(new_n13533_), .B(new_n13514_), .ZN(new_n13705_));
  INV_X1     g13448(.I(new_n13705_), .ZN(new_n13706_));
  OAI22_X1   g13449(.A1(new_n3298_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n3293_), .ZN(new_n13707_));
  NAND2_X1   g13450(.A1(new_n4227_), .A2(\b[38] ), .ZN(new_n13708_));
  AOI21_X1   g13451(.A1(new_n13707_), .A2(new_n13708_), .B(new_n3301_), .ZN(new_n13709_));
  NAND2_X1   g13452(.A1(new_n3844_), .A2(new_n13709_), .ZN(new_n13710_));
  XOR2_X1    g13453(.A1(new_n13710_), .A2(\a[38] ), .Z(new_n13711_));
  AOI21_X1   g13454(.A1(new_n13370_), .A2(new_n13522_), .B(new_n13504_), .ZN(new_n13712_));
  OAI22_X1   g13455(.A1(new_n3736_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n3731_), .ZN(new_n13713_));
  NAND2_X1   g13456(.A1(new_n4730_), .A2(\b[35] ), .ZN(new_n13714_));
  AOI21_X1   g13457(.A1(new_n13713_), .A2(new_n13714_), .B(new_n3739_), .ZN(new_n13715_));
  NAND2_X1   g13458(.A1(new_n3411_), .A2(new_n13715_), .ZN(new_n13716_));
  XOR2_X1    g13459(.A1(new_n13716_), .A2(\a[41] ), .Z(new_n13717_));
  AOI21_X1   g13460(.A1(new_n13485_), .A2(new_n13483_), .B(new_n13481_), .ZN(new_n13718_));
  OAI22_X1   g13461(.A1(new_n4208_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n4203_), .ZN(new_n13719_));
  NAND2_X1   g13462(.A1(new_n5244_), .A2(\b[32] ), .ZN(new_n13720_));
  AOI21_X1   g13463(.A1(new_n13719_), .A2(new_n13720_), .B(new_n4211_), .ZN(new_n13721_));
  NAND2_X1   g13464(.A1(new_n2963_), .A2(new_n13721_), .ZN(new_n13722_));
  XOR2_X1    g13465(.A1(new_n13722_), .A2(\a[44] ), .Z(new_n13723_));
  OAI21_X1   g13466(.A1(new_n13375_), .A2(new_n13467_), .B(new_n13466_), .ZN(new_n13724_));
  OAI22_X1   g13467(.A1(new_n4711_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n4706_), .ZN(new_n13725_));
  NAND2_X1   g13468(.A1(new_n5814_), .A2(\b[29] ), .ZN(new_n13726_));
  AOI21_X1   g13469(.A1(new_n13725_), .A2(new_n13726_), .B(new_n4714_), .ZN(new_n13727_));
  NAND2_X1   g13470(.A1(new_n2546_), .A2(new_n13727_), .ZN(new_n13728_));
  XOR2_X1    g13471(.A1(new_n13728_), .A2(\a[47] ), .Z(new_n13729_));
  INV_X1     g13472(.I(new_n13729_), .ZN(new_n13730_));
  AOI21_X1   g13473(.A1(new_n13377_), .A2(new_n13457_), .B(new_n13456_), .ZN(new_n13731_));
  OAI22_X1   g13474(.A1(new_n5228_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n5225_), .ZN(new_n13732_));
  NAND2_X1   g13475(.A1(new_n5387_), .A2(\b[26] ), .ZN(new_n13733_));
  AOI21_X1   g13476(.A1(new_n13732_), .A2(new_n13733_), .B(new_n5231_), .ZN(new_n13734_));
  NAND2_X1   g13477(.A1(new_n2174_), .A2(new_n13734_), .ZN(new_n13735_));
  XOR2_X1    g13478(.A1(new_n13735_), .A2(\a[50] ), .Z(new_n13736_));
  INV_X1     g13479(.I(new_n13736_), .ZN(new_n13737_));
  OAI22_X1   g13480(.A1(new_n6721_), .A2(new_n1393_), .B1(new_n6723_), .B2(new_n1518_), .ZN(new_n13738_));
  NAND2_X1   g13481(.A1(new_n7617_), .A2(\b[20] ), .ZN(new_n13739_));
  AOI21_X1   g13482(.A1(new_n13739_), .A2(new_n13738_), .B(new_n6731_), .ZN(new_n13740_));
  NAND2_X1   g13483(.A1(new_n1517_), .A2(new_n13740_), .ZN(new_n13741_));
  XOR2_X1    g13484(.A1(new_n13741_), .A2(\a[56] ), .Z(new_n13742_));
  OAI22_X1   g13485(.A1(new_n992_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n904_), .ZN(new_n13743_));
  NAND2_X1   g13486(.A1(new_n9644_), .A2(\b[14] ), .ZN(new_n13744_));
  AOI21_X1   g13487(.A1(new_n13744_), .A2(new_n13743_), .B(new_n8321_), .ZN(new_n13745_));
  NAND2_X1   g13488(.A1(new_n991_), .A2(new_n13745_), .ZN(new_n13746_));
  XOR2_X1    g13489(.A1(new_n13746_), .A2(\a[62] ), .Z(new_n13747_));
  NAND2_X1   g13490(.A1(new_n13402_), .A2(new_n12735_), .ZN(new_n13748_));
  NAND2_X1   g13491(.A1(new_n13748_), .A2(new_n13401_), .ZN(new_n13749_));
  NOR3_X1    g13492(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n717_), .ZN(new_n13750_));
  NOR2_X1    g13493(.A1(new_n9364_), .A2(new_n717_), .ZN(new_n13751_));
  NOR3_X1    g13494(.A1(new_n13751_), .A2(new_n795_), .A3(new_n8985_), .ZN(new_n13752_));
  NOR2_X1    g13495(.A1(new_n13752_), .A2(new_n13750_), .ZN(new_n13753_));
  NOR2_X1    g13496(.A1(new_n13749_), .A2(new_n13753_), .ZN(new_n13754_));
  INV_X1     g13497(.I(new_n13754_), .ZN(new_n13755_));
  NAND2_X1   g13498(.A1(new_n13749_), .A2(new_n13753_), .ZN(new_n13756_));
  AOI21_X1   g13499(.A1(new_n13755_), .A2(new_n13756_), .B(new_n13747_), .ZN(new_n13757_));
  INV_X1     g13500(.I(new_n13753_), .ZN(new_n13758_));
  XOR2_X1    g13501(.A1(new_n13749_), .A2(new_n13758_), .Z(new_n13759_));
  INV_X1     g13502(.I(new_n13759_), .ZN(new_n13760_));
  AOI21_X1   g13503(.A1(new_n13747_), .A2(new_n13760_), .B(new_n13757_), .ZN(new_n13761_));
  INV_X1     g13504(.I(new_n13761_), .ZN(new_n13762_));
  AOI21_X1   g13505(.A1(new_n13389_), .A2(new_n13406_), .B(new_n13408_), .ZN(new_n13763_));
  OAI22_X1   g13506(.A1(new_n1222_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1124_), .ZN(new_n13764_));
  NAND2_X1   g13507(.A1(new_n8628_), .A2(\b[17] ), .ZN(new_n13765_));
  AOI21_X1   g13508(.A1(new_n13765_), .A2(new_n13764_), .B(new_n7354_), .ZN(new_n13766_));
  NAND2_X1   g13509(.A1(new_n1225_), .A2(new_n13766_), .ZN(new_n13767_));
  XOR2_X1    g13510(.A1(new_n13767_), .A2(\a[59] ), .Z(new_n13768_));
  NOR2_X1    g13511(.A1(new_n13768_), .A2(new_n13763_), .ZN(new_n13769_));
  AND2_X2    g13512(.A1(new_n13768_), .A2(new_n13763_), .Z(new_n13770_));
  OAI21_X1   g13513(.A1(new_n13770_), .A2(new_n13769_), .B(new_n13762_), .ZN(new_n13771_));
  XOR2_X1    g13514(.A1(new_n13768_), .A2(new_n13763_), .Z(new_n13772_));
  NAND2_X1   g13515(.A1(new_n13772_), .A2(new_n13761_), .ZN(new_n13773_));
  NAND2_X1   g13516(.A1(new_n13773_), .A2(new_n13771_), .ZN(new_n13774_));
  INV_X1     g13517(.I(new_n13774_), .ZN(new_n13775_));
  NOR2_X1    g13518(.A1(new_n13424_), .A2(new_n13426_), .ZN(new_n13776_));
  NOR2_X1    g13519(.A1(new_n13776_), .A2(new_n13425_), .ZN(new_n13777_));
  NOR2_X1    g13520(.A1(new_n13775_), .A2(new_n13777_), .ZN(new_n13778_));
  INV_X1     g13521(.I(new_n13778_), .ZN(new_n13779_));
  NAND2_X1   g13522(.A1(new_n13775_), .A2(new_n13777_), .ZN(new_n13780_));
  AOI21_X1   g13523(.A1(new_n13779_), .A2(new_n13780_), .B(new_n13742_), .ZN(new_n13781_));
  INV_X1     g13524(.I(new_n13742_), .ZN(new_n13782_));
  XOR2_X1    g13525(.A1(new_n13774_), .A2(new_n13777_), .Z(new_n13783_));
  NOR2_X1    g13526(.A1(new_n13783_), .A2(new_n13782_), .ZN(new_n13784_));
  NAND2_X1   g13527(.A1(new_n13437_), .A2(new_n13434_), .ZN(new_n13785_));
  OAI21_X1   g13528(.A1(new_n13386_), .A2(new_n13438_), .B(new_n13785_), .ZN(new_n13786_));
  OAI22_X1   g13529(.A1(new_n5786_), .A2(new_n1825_), .B1(new_n1709_), .B2(new_n5792_), .ZN(new_n13787_));
  NAND2_X1   g13530(.A1(new_n6745_), .A2(\b[23] ), .ZN(new_n13788_));
  AOI21_X1   g13531(.A1(new_n13788_), .A2(new_n13787_), .B(new_n5796_), .ZN(new_n13789_));
  NAND2_X1   g13532(.A1(new_n1828_), .A2(new_n13789_), .ZN(new_n13790_));
  XOR2_X1    g13533(.A1(new_n13790_), .A2(new_n5783_), .Z(new_n13791_));
  AND2_X2    g13534(.A1(new_n13786_), .A2(new_n13791_), .Z(new_n13792_));
  NOR2_X1    g13535(.A1(new_n13786_), .A2(new_n13791_), .ZN(new_n13793_));
  OAI22_X1   g13536(.A1(new_n13792_), .A2(new_n13793_), .B1(new_n13781_), .B2(new_n13784_), .ZN(new_n13794_));
  NOR2_X1    g13537(.A1(new_n13781_), .A2(new_n13784_), .ZN(new_n13795_));
  XOR2_X1    g13538(.A1(new_n13786_), .A2(new_n13791_), .Z(new_n13796_));
  NAND2_X1   g13539(.A1(new_n13796_), .A2(new_n13795_), .ZN(new_n13797_));
  NAND2_X1   g13540(.A1(new_n13797_), .A2(new_n13794_), .ZN(new_n13798_));
  NAND2_X1   g13541(.A1(new_n13441_), .A2(new_n13444_), .ZN(new_n13799_));
  NAND2_X1   g13542(.A1(new_n13799_), .A2(new_n13442_), .ZN(new_n13800_));
  XOR2_X1    g13543(.A1(new_n13798_), .A2(new_n13800_), .Z(new_n13801_));
  NAND2_X1   g13544(.A1(new_n13801_), .A2(new_n13737_), .ZN(new_n13802_));
  AOI22_X1   g13545(.A1(new_n13797_), .A2(new_n13794_), .B1(new_n13799_), .B2(new_n13442_), .ZN(new_n13803_));
  NOR2_X1    g13546(.A1(new_n13798_), .A2(new_n13800_), .ZN(new_n13804_));
  OAI21_X1   g13547(.A1(new_n13804_), .A2(new_n13803_), .B(new_n13736_), .ZN(new_n13805_));
  NAND2_X1   g13548(.A1(new_n13802_), .A2(new_n13805_), .ZN(new_n13806_));
  XOR2_X1    g13549(.A1(new_n13806_), .A2(new_n13731_), .Z(new_n13807_));
  NAND2_X1   g13550(.A1(new_n13807_), .A2(new_n13730_), .ZN(new_n13808_));
  INV_X1     g13551(.I(new_n13731_), .ZN(new_n13809_));
  INV_X1     g13552(.I(new_n13806_), .ZN(new_n13810_));
  NOR2_X1    g13553(.A1(new_n13810_), .A2(new_n13809_), .ZN(new_n13811_));
  NOR2_X1    g13554(.A1(new_n13806_), .A2(new_n13731_), .ZN(new_n13812_));
  OAI21_X1   g13555(.A1(new_n13811_), .A2(new_n13812_), .B(new_n13729_), .ZN(new_n13813_));
  NAND2_X1   g13556(.A1(new_n13808_), .A2(new_n13813_), .ZN(new_n13814_));
  XOR2_X1    g13557(.A1(new_n13814_), .A2(new_n13724_), .Z(new_n13815_));
  NOR2_X1    g13558(.A1(new_n13815_), .A2(new_n13723_), .ZN(new_n13816_));
  INV_X1     g13559(.I(new_n13723_), .ZN(new_n13817_));
  INV_X1     g13560(.I(new_n13724_), .ZN(new_n13818_));
  NAND2_X1   g13561(.A1(new_n13814_), .A2(new_n13818_), .ZN(new_n13819_));
  NAND3_X1   g13562(.A1(new_n13808_), .A2(new_n13724_), .A3(new_n13813_), .ZN(new_n13820_));
  AOI21_X1   g13563(.A1(new_n13819_), .A2(new_n13820_), .B(new_n13817_), .ZN(new_n13821_));
  NOR2_X1    g13564(.A1(new_n13816_), .A2(new_n13821_), .ZN(new_n13822_));
  XOR2_X1    g13565(.A1(new_n13822_), .A2(new_n13718_), .Z(new_n13823_));
  NOR2_X1    g13566(.A1(new_n13823_), .A2(new_n13717_), .ZN(new_n13824_));
  INV_X1     g13567(.I(new_n13717_), .ZN(new_n13825_));
  OAI21_X1   g13568(.A1(new_n13816_), .A2(new_n13821_), .B(new_n13718_), .ZN(new_n13826_));
  INV_X1     g13569(.I(new_n13718_), .ZN(new_n13827_));
  NAND2_X1   g13570(.A1(new_n13822_), .A2(new_n13827_), .ZN(new_n13828_));
  AOI21_X1   g13571(.A1(new_n13828_), .A2(new_n13826_), .B(new_n13825_), .ZN(new_n13829_));
  NOR2_X1    g13572(.A1(new_n13824_), .A2(new_n13829_), .ZN(new_n13830_));
  XOR2_X1    g13573(.A1(new_n13830_), .A2(new_n13712_), .Z(new_n13831_));
  NOR2_X1    g13574(.A1(new_n13831_), .A2(new_n13711_), .ZN(new_n13832_));
  INV_X1     g13575(.I(new_n13711_), .ZN(new_n13833_));
  OAI21_X1   g13576(.A1(new_n13824_), .A2(new_n13829_), .B(new_n13712_), .ZN(new_n13834_));
  INV_X1     g13577(.I(new_n13712_), .ZN(new_n13835_));
  NAND2_X1   g13578(.A1(new_n13830_), .A2(new_n13835_), .ZN(new_n13836_));
  AOI21_X1   g13579(.A1(new_n13836_), .A2(new_n13834_), .B(new_n13833_), .ZN(new_n13837_));
  NOR2_X1    g13580(.A1(new_n13832_), .A2(new_n13837_), .ZN(new_n13838_));
  OAI22_X1   g13581(.A1(new_n2846_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n2841_), .ZN(new_n13839_));
  NAND2_X1   g13582(.A1(new_n3755_), .A2(\b[41] ), .ZN(new_n13840_));
  AOI21_X1   g13583(.A1(new_n13839_), .A2(new_n13840_), .B(new_n2849_), .ZN(new_n13841_));
  NAND2_X1   g13584(.A1(new_n4320_), .A2(new_n13841_), .ZN(new_n13842_));
  XOR2_X1    g13585(.A1(new_n13842_), .A2(\a[35] ), .Z(new_n13843_));
  INV_X1     g13586(.I(new_n13843_), .ZN(new_n13844_));
  NAND2_X1   g13587(.A1(new_n13838_), .A2(new_n13844_), .ZN(new_n13845_));
  INV_X1     g13588(.I(new_n13845_), .ZN(new_n13846_));
  NOR2_X1    g13589(.A1(new_n13838_), .A2(new_n13844_), .ZN(new_n13847_));
  OAI21_X1   g13590(.A1(new_n13846_), .A2(new_n13847_), .B(new_n13706_), .ZN(new_n13848_));
  INV_X1     g13591(.I(new_n13848_), .ZN(new_n13849_));
  XOR2_X1    g13592(.A1(new_n13838_), .A2(new_n13843_), .Z(new_n13850_));
  NOR2_X1    g13593(.A1(new_n13850_), .A2(new_n13706_), .ZN(new_n13851_));
  NOR2_X1    g13594(.A1(new_n13849_), .A2(new_n13851_), .ZN(new_n13852_));
  NOR2_X1    g13595(.A1(new_n13555_), .A2(new_n13365_), .ZN(new_n13853_));
  NOR2_X1    g13596(.A1(new_n13853_), .A2(new_n13554_), .ZN(new_n13854_));
  INV_X1     g13597(.I(new_n13854_), .ZN(new_n13855_));
  OAI22_X1   g13598(.A1(new_n2452_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n2447_), .ZN(new_n13856_));
  OAI21_X1   g13599(.A1(new_n4501_), .A2(new_n2602_), .B(new_n13856_), .ZN(new_n13857_));
  AOI21_X1   g13600(.A1(new_n4833_), .A2(new_n2454_), .B(new_n13857_), .ZN(new_n13858_));
  NOR2_X1    g13601(.A1(new_n13855_), .A2(new_n13858_), .ZN(new_n13859_));
  INV_X1     g13602(.I(new_n13858_), .ZN(new_n13860_));
  NOR2_X1    g13603(.A1(new_n13854_), .A2(new_n13860_), .ZN(new_n13861_));
  OAI21_X1   g13604(.A1(new_n13859_), .A2(new_n13861_), .B(new_n2442_), .ZN(new_n13862_));
  INV_X1     g13605(.I(new_n13862_), .ZN(new_n13863_));
  NOR3_X1    g13606(.A1(new_n13859_), .A2(new_n13861_), .A3(new_n2442_), .ZN(new_n13864_));
  OAI21_X1   g13607(.A1(new_n13863_), .A2(new_n13864_), .B(new_n13852_), .ZN(new_n13865_));
  OAI21_X1   g13608(.A1(new_n13850_), .A2(new_n13706_), .B(new_n13848_), .ZN(new_n13866_));
  INV_X1     g13609(.I(new_n13864_), .ZN(new_n13867_));
  NAND3_X1   g13610(.A1(new_n13866_), .A2(new_n13862_), .A3(new_n13867_), .ZN(new_n13868_));
  OAI22_X1   g13611(.A1(new_n2084_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n2079_), .ZN(new_n13869_));
  NAND2_X1   g13612(.A1(new_n2864_), .A2(\b[47] ), .ZN(new_n13870_));
  AOI21_X1   g13613(.A1(new_n13869_), .A2(new_n13870_), .B(new_n2087_), .ZN(new_n13871_));
  NAND2_X1   g13614(.A1(new_n5196_), .A2(new_n13871_), .ZN(new_n13872_));
  XOR2_X1    g13615(.A1(new_n13872_), .A2(\a[29] ), .Z(new_n13873_));
  AOI21_X1   g13616(.A1(new_n13865_), .A2(new_n13868_), .B(new_n13873_), .ZN(new_n13874_));
  AOI21_X1   g13617(.A1(new_n13862_), .A2(new_n13867_), .B(new_n13866_), .ZN(new_n13875_));
  NOR3_X1    g13618(.A1(new_n13852_), .A2(new_n13863_), .A3(new_n13864_), .ZN(new_n13876_));
  INV_X1     g13619(.I(new_n13873_), .ZN(new_n13877_));
  NOR3_X1    g13620(.A1(new_n13876_), .A2(new_n13875_), .A3(new_n13877_), .ZN(new_n13878_));
  OAI21_X1   g13621(.A1(new_n13874_), .A2(new_n13878_), .B(new_n13704_), .ZN(new_n13879_));
  NOR3_X1    g13622(.A1(new_n13876_), .A2(new_n13875_), .A3(new_n13873_), .ZN(new_n13880_));
  AOI21_X1   g13623(.A1(new_n13865_), .A2(new_n13868_), .B(new_n13877_), .ZN(new_n13881_));
  OAI21_X1   g13624(.A1(new_n13881_), .A2(new_n13880_), .B(new_n13703_), .ZN(new_n13882_));
  OAI22_X1   g13625(.A1(new_n1760_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n1755_), .ZN(new_n13883_));
  NAND2_X1   g13626(.A1(new_n2470_), .A2(\b[50] ), .ZN(new_n13884_));
  AOI21_X1   g13627(.A1(new_n13883_), .A2(new_n13884_), .B(new_n1763_), .ZN(new_n13885_));
  NAND2_X1   g13628(.A1(new_n5954_), .A2(new_n13885_), .ZN(new_n13886_));
  XOR2_X1    g13629(.A1(new_n13886_), .A2(\a[26] ), .Z(new_n13887_));
  AOI21_X1   g13630(.A1(new_n13879_), .A2(new_n13882_), .B(new_n13887_), .ZN(new_n13888_));
  OAI21_X1   g13631(.A1(new_n13876_), .A2(new_n13875_), .B(new_n13877_), .ZN(new_n13889_));
  NAND3_X1   g13632(.A1(new_n13865_), .A2(new_n13868_), .A3(new_n13873_), .ZN(new_n13890_));
  AOI21_X1   g13633(.A1(new_n13890_), .A2(new_n13889_), .B(new_n13703_), .ZN(new_n13891_));
  NAND3_X1   g13634(.A1(new_n13865_), .A2(new_n13868_), .A3(new_n13877_), .ZN(new_n13892_));
  OAI21_X1   g13635(.A1(new_n13876_), .A2(new_n13875_), .B(new_n13873_), .ZN(new_n13893_));
  AOI21_X1   g13636(.A1(new_n13892_), .A2(new_n13893_), .B(new_n13704_), .ZN(new_n13894_));
  INV_X1     g13637(.I(new_n13887_), .ZN(new_n13895_));
  NOR3_X1    g13638(.A1(new_n13891_), .A2(new_n13894_), .A3(new_n13895_), .ZN(new_n13896_));
  OAI21_X1   g13639(.A1(new_n13888_), .A2(new_n13896_), .B(new_n13702_), .ZN(new_n13897_));
  NOR3_X1    g13640(.A1(new_n13891_), .A2(new_n13894_), .A3(new_n13887_), .ZN(new_n13898_));
  AOI21_X1   g13641(.A1(new_n13879_), .A2(new_n13882_), .B(new_n13895_), .ZN(new_n13899_));
  OAI21_X1   g13642(.A1(new_n13899_), .A2(new_n13898_), .B(new_n13701_), .ZN(new_n13900_));
  OAI22_X1   g13643(.A1(new_n1444_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n1439_), .ZN(new_n13901_));
  NAND2_X1   g13644(.A1(new_n2098_), .A2(\b[53] ), .ZN(new_n13902_));
  AOI21_X1   g13645(.A1(new_n13901_), .A2(new_n13902_), .B(new_n1447_), .ZN(new_n13903_));
  NAND2_X1   g13646(.A1(new_n6471_), .A2(new_n13903_), .ZN(new_n13904_));
  XOR2_X1    g13647(.A1(new_n13904_), .A2(\a[23] ), .Z(new_n13905_));
  AOI21_X1   g13648(.A1(new_n13897_), .A2(new_n13900_), .B(new_n13905_), .ZN(new_n13906_));
  OAI21_X1   g13649(.A1(new_n13891_), .A2(new_n13894_), .B(new_n13895_), .ZN(new_n13907_));
  NAND3_X1   g13650(.A1(new_n13879_), .A2(new_n13882_), .A3(new_n13887_), .ZN(new_n13908_));
  AOI21_X1   g13651(.A1(new_n13907_), .A2(new_n13908_), .B(new_n13701_), .ZN(new_n13909_));
  NAND3_X1   g13652(.A1(new_n13879_), .A2(new_n13882_), .A3(new_n13895_), .ZN(new_n13910_));
  OAI21_X1   g13653(.A1(new_n13891_), .A2(new_n13894_), .B(new_n13887_), .ZN(new_n13911_));
  AOI21_X1   g13654(.A1(new_n13911_), .A2(new_n13910_), .B(new_n13702_), .ZN(new_n13912_));
  INV_X1     g13655(.I(new_n13905_), .ZN(new_n13913_));
  NOR3_X1    g13656(.A1(new_n13909_), .A2(new_n13912_), .A3(new_n13913_), .ZN(new_n13914_));
  OAI21_X1   g13657(.A1(new_n13906_), .A2(new_n13914_), .B(new_n13700_), .ZN(new_n13915_));
  NOR3_X1    g13658(.A1(new_n13909_), .A2(new_n13912_), .A3(new_n13905_), .ZN(new_n13916_));
  AOI21_X1   g13659(.A1(new_n13897_), .A2(new_n13900_), .B(new_n13913_), .ZN(new_n13917_));
  OAI21_X1   g13660(.A1(new_n13917_), .A2(new_n13916_), .B(new_n13699_), .ZN(new_n13918_));
  AOI21_X1   g13661(.A1(new_n13915_), .A2(new_n13918_), .B(new_n13698_), .ZN(new_n13919_));
  OAI21_X1   g13662(.A1(new_n13909_), .A2(new_n13912_), .B(new_n13913_), .ZN(new_n13920_));
  NAND3_X1   g13663(.A1(new_n13897_), .A2(new_n13900_), .A3(new_n13905_), .ZN(new_n13921_));
  AOI21_X1   g13664(.A1(new_n13920_), .A2(new_n13921_), .B(new_n13699_), .ZN(new_n13922_));
  NAND3_X1   g13665(.A1(new_n13897_), .A2(new_n13900_), .A3(new_n13913_), .ZN(new_n13923_));
  OAI21_X1   g13666(.A1(new_n13909_), .A2(new_n13912_), .B(new_n13905_), .ZN(new_n13924_));
  AOI21_X1   g13667(.A1(new_n13924_), .A2(new_n13923_), .B(new_n13700_), .ZN(new_n13925_));
  NOR3_X1    g13668(.A1(new_n13922_), .A2(new_n13925_), .A3(new_n13697_), .ZN(new_n13926_));
  OAI21_X1   g13669(.A1(new_n13919_), .A2(new_n13926_), .B(new_n1158_), .ZN(new_n13927_));
  OAI21_X1   g13670(.A1(new_n13922_), .A2(new_n13925_), .B(new_n13697_), .ZN(new_n13928_));
  NAND3_X1   g13671(.A1(new_n13915_), .A2(new_n13918_), .A3(new_n13698_), .ZN(new_n13929_));
  NAND3_X1   g13672(.A1(new_n13928_), .A2(new_n13929_), .A3(\a[20] ), .ZN(new_n13930_));
  AOI21_X1   g13673(.A1(new_n13927_), .A2(new_n13930_), .B(new_n13696_), .ZN(new_n13931_));
  AOI21_X1   g13674(.A1(new_n13928_), .A2(new_n13929_), .B(\a[20] ), .ZN(new_n13932_));
  NOR3_X1    g13675(.A1(new_n13919_), .A2(new_n13926_), .A3(new_n1158_), .ZN(new_n13933_));
  NOR3_X1    g13676(.A1(new_n13933_), .A2(new_n13932_), .A3(new_n13695_), .ZN(new_n13934_));
  OAI22_X1   g13677(.A1(new_n940_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n935_), .ZN(new_n13935_));
  NAND2_X1   g13678(.A1(new_n1458_), .A2(\b[59] ), .ZN(new_n13936_));
  AOI21_X1   g13679(.A1(new_n13935_), .A2(new_n13936_), .B(new_n943_), .ZN(new_n13937_));
  NAND2_X1   g13680(.A1(new_n8550_), .A2(new_n13937_), .ZN(new_n13938_));
  XOR2_X1    g13681(.A1(new_n13938_), .A2(\a[17] ), .Z(new_n13939_));
  INV_X1     g13682(.I(new_n13939_), .ZN(new_n13940_));
  OAI21_X1   g13683(.A1(new_n13934_), .A2(new_n13931_), .B(new_n13940_), .ZN(new_n13941_));
  OAI21_X1   g13684(.A1(new_n13933_), .A2(new_n13932_), .B(new_n13695_), .ZN(new_n13942_));
  NAND3_X1   g13685(.A1(new_n13927_), .A2(new_n13930_), .A3(new_n13696_), .ZN(new_n13943_));
  NAND3_X1   g13686(.A1(new_n13942_), .A2(new_n13943_), .A3(new_n13939_), .ZN(new_n13944_));
  AOI21_X1   g13687(.A1(new_n13941_), .A2(new_n13944_), .B(new_n13692_), .ZN(new_n13945_));
  INV_X1     g13688(.I(new_n13692_), .ZN(new_n13946_));
  NAND3_X1   g13689(.A1(new_n13942_), .A2(new_n13943_), .A3(new_n13940_), .ZN(new_n13947_));
  OAI21_X1   g13690(.A1(new_n13934_), .A2(new_n13931_), .B(new_n13939_), .ZN(new_n13948_));
  AOI21_X1   g13691(.A1(new_n13948_), .A2(new_n13947_), .B(new_n13946_), .ZN(new_n13949_));
  NOR2_X1    g13692(.A1(new_n823_), .A2(new_n8932_), .ZN(new_n13950_));
  NOR2_X1    g13693(.A1(new_n752_), .A2(new_n8956_), .ZN(new_n13951_));
  NOR4_X1    g13694(.A1(new_n9323_), .A2(new_n760_), .A3(new_n13950_), .A4(new_n13951_), .ZN(new_n13952_));
  XOR2_X1    g13695(.A1(new_n13952_), .A2(new_n747_), .Z(new_n13953_));
  NOR3_X1    g13696(.A1(new_n13945_), .A2(new_n13949_), .A3(new_n13953_), .ZN(new_n13954_));
  AOI21_X1   g13697(.A1(new_n13942_), .A2(new_n13943_), .B(new_n13939_), .ZN(new_n13955_));
  NOR3_X1    g13698(.A1(new_n13934_), .A2(new_n13931_), .A3(new_n13940_), .ZN(new_n13956_));
  OAI21_X1   g13699(.A1(new_n13956_), .A2(new_n13955_), .B(new_n13946_), .ZN(new_n13957_));
  NOR3_X1    g13700(.A1(new_n13934_), .A2(new_n13931_), .A3(new_n13939_), .ZN(new_n13958_));
  AOI21_X1   g13701(.A1(new_n13942_), .A2(new_n13943_), .B(new_n13940_), .ZN(new_n13959_));
  OAI21_X1   g13702(.A1(new_n13958_), .A2(new_n13959_), .B(new_n13692_), .ZN(new_n13960_));
  INV_X1     g13703(.I(new_n13953_), .ZN(new_n13961_));
  AOI21_X1   g13704(.A1(new_n13957_), .A2(new_n13960_), .B(new_n13961_), .ZN(new_n13962_));
  OAI21_X1   g13705(.A1(new_n13962_), .A2(new_n13954_), .B(new_n13690_), .ZN(new_n13963_));
  AOI21_X1   g13706(.A1(new_n13957_), .A2(new_n13960_), .B(new_n13953_), .ZN(new_n13964_));
  NOR3_X1    g13707(.A1(new_n13945_), .A2(new_n13949_), .A3(new_n13961_), .ZN(new_n13965_));
  OAI21_X1   g13708(.A1(new_n13964_), .A2(new_n13965_), .B(new_n13689_), .ZN(new_n13966_));
  NAND2_X1   g13709(.A1(new_n13963_), .A2(new_n13966_), .ZN(new_n13967_));
  NAND2_X1   g13710(.A1(new_n13680_), .A2(new_n13330_), .ZN(new_n13968_));
  NAND2_X1   g13711(.A1(new_n13669_), .A2(new_n13674_), .ZN(new_n13969_));
  NOR2_X1    g13712(.A1(new_n13329_), .A2(new_n13969_), .ZN(new_n13970_));
  AOI21_X1   g13713(.A1(new_n13968_), .A2(new_n13970_), .B(new_n13967_), .ZN(new_n13971_));
  INV_X1     g13714(.I(new_n13967_), .ZN(new_n13972_));
  OAI21_X1   g13715(.A1(new_n13007_), .A2(new_n13331_), .B(new_n13970_), .ZN(new_n13973_));
  NOR2_X1    g13716(.A1(new_n13973_), .A2(new_n13972_), .ZN(new_n13974_));
  OAI21_X1   g13717(.A1(new_n13974_), .A2(new_n13971_), .B(new_n13687_), .ZN(new_n13975_));
  INV_X1     g13718(.I(new_n13687_), .ZN(new_n13976_));
  NAND2_X1   g13719(.A1(new_n13973_), .A2(new_n13972_), .ZN(new_n13977_));
  NAND3_X1   g13720(.A1(new_n13968_), .A2(new_n13967_), .A3(new_n13970_), .ZN(new_n13978_));
  NAND3_X1   g13721(.A1(new_n13977_), .A2(new_n13978_), .A3(new_n13976_), .ZN(new_n13979_));
  NAND2_X1   g13722(.A1(new_n13975_), .A2(new_n13979_), .ZN(\f[76] ));
  AOI22_X1   g13723(.A1(new_n13977_), .A2(new_n13978_), .B1(new_n13976_), .B2(new_n13973_), .ZN(new_n13981_));
  NOR2_X1    g13724(.A1(new_n13965_), .A2(new_n13689_), .ZN(new_n13982_));
  NOR2_X1    g13725(.A1(new_n13982_), .A2(new_n13964_), .ZN(new_n13983_));
  AOI22_X1   g13726(.A1(new_n10814_), .A2(new_n759_), .B1(\b[63] ), .B2(new_n1182_), .ZN(new_n13984_));
  AOI21_X1   g13727(.A1(new_n13946_), .A2(new_n13944_), .B(new_n13955_), .ZN(new_n13985_));
  OAI22_X1   g13728(.A1(new_n940_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n935_), .ZN(new_n13986_));
  OAI21_X1   g13729(.A1(new_n7930_), .A2(new_n1020_), .B(new_n13986_), .ZN(new_n13987_));
  AOI21_X1   g13730(.A1(new_n8935_), .A2(new_n942_), .B(new_n13987_), .ZN(new_n13988_));
  INV_X1     g13731(.I(new_n13988_), .ZN(new_n13989_));
  AOI21_X1   g13732(.A1(new_n13915_), .A2(new_n13918_), .B(new_n13697_), .ZN(new_n13990_));
  XOR2_X1    g13733(.A1(new_n13695_), .A2(\a[20] ), .Z(new_n13991_));
  NOR4_X1    g13734(.A1(new_n13922_), .A2(new_n13925_), .A3(new_n13698_), .A4(new_n13991_), .ZN(new_n13992_));
  NOR2_X1    g13735(.A1(new_n13992_), .A2(new_n13990_), .ZN(new_n13993_));
  INV_X1     g13736(.I(new_n13993_), .ZN(new_n13994_));
  AOI21_X1   g13737(.A1(new_n13700_), .A2(new_n13921_), .B(new_n13906_), .ZN(new_n13995_));
  INV_X1     g13738(.I(new_n13995_), .ZN(new_n13996_));
  OAI22_X1   g13739(.A1(new_n1444_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n1439_), .ZN(new_n13997_));
  OAI21_X1   g13740(.A1(new_n6238_), .A2(new_n1548_), .B(new_n13997_), .ZN(new_n13998_));
  AOI21_X1   g13741(.A1(new_n6994_), .A2(new_n1446_), .B(new_n13998_), .ZN(new_n13999_));
  INV_X1     g13742(.I(new_n13999_), .ZN(new_n14000_));
  AOI21_X1   g13743(.A1(new_n13702_), .A2(new_n13908_), .B(new_n13888_), .ZN(new_n14001_));
  AOI21_X1   g13744(.A1(new_n13704_), .A2(new_n13890_), .B(new_n13874_), .ZN(new_n14002_));
  OAI22_X1   g13745(.A1(new_n1760_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n1755_), .ZN(new_n14003_));
  NAND2_X1   g13746(.A1(new_n2470_), .A2(\b[51] ), .ZN(new_n14004_));
  AOI21_X1   g13747(.A1(new_n14003_), .A2(new_n14004_), .B(new_n1763_), .ZN(new_n14005_));
  NAND2_X1   g13748(.A1(new_n6219_), .A2(new_n14005_), .ZN(new_n14006_));
  XOR2_X1    g13749(.A1(new_n14006_), .A2(\a[26] ), .Z(new_n14007_));
  INV_X1     g13750(.I(new_n14007_), .ZN(new_n14008_));
  OAI22_X1   g13751(.A1(new_n2452_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n2447_), .ZN(new_n14009_));
  NAND2_X1   g13752(.A1(new_n3312_), .A2(\b[45] ), .ZN(new_n14010_));
  AOI21_X1   g13753(.A1(new_n14009_), .A2(new_n14010_), .B(new_n2455_), .ZN(new_n14011_));
  NAND2_X1   g13754(.A1(new_n5004_), .A2(new_n14011_), .ZN(new_n14012_));
  XOR2_X1    g13755(.A1(new_n14012_), .A2(\a[32] ), .Z(new_n14013_));
  INV_X1     g13756(.I(new_n14013_), .ZN(new_n14014_));
  OAI22_X1   g13757(.A1(new_n2846_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n2841_), .ZN(new_n14015_));
  NAND2_X1   g13758(.A1(new_n3755_), .A2(\b[42] ), .ZN(new_n14016_));
  AOI21_X1   g13759(.A1(new_n14015_), .A2(new_n14016_), .B(new_n2849_), .ZN(new_n14017_));
  NAND2_X1   g13760(.A1(new_n4500_), .A2(new_n14017_), .ZN(new_n14018_));
  XOR2_X1    g13761(.A1(new_n14018_), .A2(\a[35] ), .Z(new_n14019_));
  INV_X1     g13762(.I(new_n14019_), .ZN(new_n14020_));
  NAND2_X1   g13763(.A1(new_n13834_), .A2(new_n13833_), .ZN(new_n14021_));
  NAND2_X1   g13764(.A1(new_n14021_), .A2(new_n13836_), .ZN(new_n14022_));
  OAI22_X1   g13765(.A1(new_n3298_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n3293_), .ZN(new_n14023_));
  NAND2_X1   g13766(.A1(new_n4227_), .A2(\b[39] ), .ZN(new_n14024_));
  AOI21_X1   g13767(.A1(new_n14023_), .A2(new_n14024_), .B(new_n3301_), .ZN(new_n14025_));
  NAND2_X1   g13768(.A1(new_n3996_), .A2(new_n14025_), .ZN(new_n14026_));
  XOR2_X1    g13769(.A1(new_n14026_), .A2(\a[38] ), .Z(new_n14027_));
  INV_X1     g13770(.I(new_n14027_), .ZN(new_n14028_));
  OAI22_X1   g13771(.A1(new_n3736_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n3731_), .ZN(new_n14029_));
  NAND2_X1   g13772(.A1(new_n4730_), .A2(\b[36] ), .ZN(new_n14030_));
  AOI21_X1   g13773(.A1(new_n14029_), .A2(new_n14030_), .B(new_n3739_), .ZN(new_n14031_));
  NAND2_X1   g13774(.A1(new_n3565_), .A2(new_n14031_), .ZN(new_n14032_));
  XOR2_X1    g13775(.A1(new_n14032_), .A2(\a[41] ), .Z(new_n14033_));
  INV_X1     g13776(.I(new_n14033_), .ZN(new_n14034_));
  OAI22_X1   g13777(.A1(new_n4711_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n4706_), .ZN(new_n14035_));
  NAND2_X1   g13778(.A1(new_n5814_), .A2(\b[30] ), .ZN(new_n14036_));
  AOI21_X1   g13779(.A1(new_n14035_), .A2(new_n14036_), .B(new_n4714_), .ZN(new_n14037_));
  NAND2_X1   g13780(.A1(new_n2659_), .A2(new_n14037_), .ZN(new_n14038_));
  XOR2_X1    g13781(.A1(new_n14038_), .A2(\a[47] ), .Z(new_n14039_));
  INV_X1     g13782(.I(new_n14039_), .ZN(new_n14040_));
  OAI22_X1   g13783(.A1(new_n5786_), .A2(new_n1927_), .B1(new_n1825_), .B2(new_n5792_), .ZN(new_n14041_));
  NAND2_X1   g13784(.A1(new_n6745_), .A2(\b[24] ), .ZN(new_n14042_));
  AOI21_X1   g13785(.A1(new_n14042_), .A2(new_n14041_), .B(new_n5796_), .ZN(new_n14043_));
  NAND2_X1   g13786(.A1(new_n1926_), .A2(new_n14043_), .ZN(new_n14044_));
  XOR2_X1    g13787(.A1(new_n14044_), .A2(\a[53] ), .Z(new_n14045_));
  AOI21_X1   g13788(.A1(new_n13775_), .A2(new_n13777_), .B(new_n13742_), .ZN(new_n14046_));
  NOR2_X1    g13789(.A1(new_n14046_), .A2(new_n13778_), .ZN(new_n14047_));
  OAI22_X1   g13790(.A1(new_n1305_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1222_), .ZN(new_n14048_));
  NAND2_X1   g13791(.A1(new_n8628_), .A2(\b[18] ), .ZN(new_n14049_));
  AOI21_X1   g13792(.A1(new_n14049_), .A2(new_n14048_), .B(new_n7354_), .ZN(new_n14050_));
  NAND2_X1   g13793(.A1(new_n1304_), .A2(new_n14050_), .ZN(new_n14051_));
  XOR2_X1    g13794(.A1(new_n14051_), .A2(\a[59] ), .Z(new_n14052_));
  OAI21_X1   g13795(.A1(new_n13747_), .A2(new_n13754_), .B(new_n13756_), .ZN(new_n14053_));
  OAI22_X1   g13796(.A1(new_n1044_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n992_), .ZN(new_n14054_));
  NAND2_X1   g13797(.A1(new_n9644_), .A2(\b[15] ), .ZN(new_n14055_));
  AOI21_X1   g13798(.A1(new_n14055_), .A2(new_n14054_), .B(new_n8321_), .ZN(new_n14056_));
  NAND2_X1   g13799(.A1(new_n1047_), .A2(new_n14056_), .ZN(new_n14057_));
  XOR2_X1    g13800(.A1(new_n14057_), .A2(\a[62] ), .Z(new_n14058_));
  NOR2_X1    g13801(.A1(new_n8985_), .A2(new_n848_), .ZN(new_n14059_));
  NOR2_X1    g13802(.A1(new_n9364_), .A2(new_n795_), .ZN(new_n14060_));
  XNOR2_X1   g13803(.A1(new_n14059_), .A2(new_n14060_), .ZN(new_n14061_));
  XOR2_X1    g13804(.A1(new_n14061_), .A2(new_n13753_), .Z(new_n14062_));
  NOR2_X1    g13805(.A1(new_n14058_), .A2(new_n14062_), .ZN(new_n14063_));
  XOR2_X1    g13806(.A1(new_n14057_), .A2(new_n8309_), .Z(new_n14064_));
  NOR2_X1    g13807(.A1(new_n13758_), .A2(new_n14061_), .ZN(new_n14065_));
  INV_X1     g13808(.I(new_n14065_), .ZN(new_n14066_));
  NAND2_X1   g13809(.A1(new_n13758_), .A2(new_n14061_), .ZN(new_n14067_));
  AOI21_X1   g13810(.A1(new_n14066_), .A2(new_n14067_), .B(new_n14064_), .ZN(new_n14068_));
  NOR2_X1    g13811(.A1(new_n14068_), .A2(new_n14063_), .ZN(new_n14069_));
  OR2_X2     g13812(.A1(new_n14069_), .A2(new_n14053_), .Z(new_n14070_));
  NAND2_X1   g13813(.A1(new_n14069_), .A2(new_n14053_), .ZN(new_n14071_));
  AOI21_X1   g13814(.A1(new_n14070_), .A2(new_n14071_), .B(new_n14052_), .ZN(new_n14072_));
  XOR2_X1    g13815(.A1(new_n14069_), .A2(new_n14053_), .Z(new_n14073_));
  AND2_X2    g13816(.A1(new_n14073_), .A2(new_n14052_), .Z(new_n14074_));
  NOR2_X1    g13817(.A1(new_n14074_), .A2(new_n14072_), .ZN(new_n14075_));
  OAI22_X1   g13818(.A1(new_n6721_), .A2(new_n1518_), .B1(new_n6723_), .B2(new_n1601_), .ZN(new_n14076_));
  NAND2_X1   g13819(.A1(new_n7617_), .A2(\b[21] ), .ZN(new_n14077_));
  AOI21_X1   g13820(.A1(new_n14077_), .A2(new_n14076_), .B(new_n6731_), .ZN(new_n14078_));
  NAND2_X1   g13821(.A1(new_n1604_), .A2(new_n14078_), .ZN(new_n14079_));
  XOR2_X1    g13822(.A1(new_n14079_), .A2(\a[56] ), .Z(new_n14080_));
  NOR2_X1    g13823(.A1(new_n13770_), .A2(new_n13761_), .ZN(new_n14081_));
  NOR2_X1    g13824(.A1(new_n14081_), .A2(new_n13769_), .ZN(new_n14082_));
  XNOR2_X1   g13825(.A1(new_n14080_), .A2(new_n14082_), .ZN(new_n14083_));
  NOR2_X1    g13826(.A1(new_n14083_), .A2(new_n14075_), .ZN(new_n14084_));
  INV_X1     g13827(.I(new_n14075_), .ZN(new_n14085_));
  NOR2_X1    g13828(.A1(new_n14080_), .A2(new_n14082_), .ZN(new_n14086_));
  INV_X1     g13829(.I(new_n14086_), .ZN(new_n14087_));
  NAND2_X1   g13830(.A1(new_n14080_), .A2(new_n14082_), .ZN(new_n14088_));
  AOI21_X1   g13831(.A1(new_n14087_), .A2(new_n14088_), .B(new_n14085_), .ZN(new_n14089_));
  NOR2_X1    g13832(.A1(new_n14089_), .A2(new_n14084_), .ZN(new_n14090_));
  XOR2_X1    g13833(.A1(new_n14090_), .A2(new_n14047_), .Z(new_n14091_));
  NOR2_X1    g13834(.A1(new_n14091_), .A2(new_n14045_), .ZN(new_n14092_));
  INV_X1     g13835(.I(new_n14045_), .ZN(new_n14093_));
  OAI21_X1   g13836(.A1(new_n14089_), .A2(new_n14084_), .B(new_n14047_), .ZN(new_n14094_));
  OAI21_X1   g13837(.A1(new_n13778_), .A2(new_n14046_), .B(new_n14090_), .ZN(new_n14095_));
  AOI21_X1   g13838(.A1(new_n14095_), .A2(new_n14094_), .B(new_n14093_), .ZN(new_n14096_));
  NOR2_X1    g13839(.A1(new_n14092_), .A2(new_n14096_), .ZN(new_n14097_));
  OAI22_X1   g13840(.A1(new_n5228_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n5225_), .ZN(new_n14098_));
  NAND2_X1   g13841(.A1(new_n5387_), .A2(\b[27] ), .ZN(new_n14099_));
  AOI21_X1   g13842(.A1(new_n14098_), .A2(new_n14099_), .B(new_n5231_), .ZN(new_n14100_));
  NAND2_X1   g13843(.A1(new_n2276_), .A2(new_n14100_), .ZN(new_n14101_));
  XOR2_X1    g13844(.A1(new_n14101_), .A2(\a[50] ), .Z(new_n14102_));
  INV_X1     g13845(.I(new_n14102_), .ZN(new_n14103_));
  NOR2_X1    g13846(.A1(new_n13793_), .A2(new_n13795_), .ZN(new_n14104_));
  NOR2_X1    g13847(.A1(new_n14104_), .A2(new_n13792_), .ZN(new_n14105_));
  XOR2_X1    g13848(.A1(new_n14105_), .A2(new_n14103_), .Z(new_n14106_));
  NOR2_X1    g13849(.A1(new_n14106_), .A2(new_n14097_), .ZN(new_n14107_));
  OAI21_X1   g13850(.A1(new_n13792_), .A2(new_n14104_), .B(new_n14103_), .ZN(new_n14108_));
  NAND2_X1   g13851(.A1(new_n14105_), .A2(new_n14102_), .ZN(new_n14109_));
  NAND2_X1   g13852(.A1(new_n14109_), .A2(new_n14108_), .ZN(new_n14110_));
  AOI21_X1   g13853(.A1(new_n14097_), .A2(new_n14110_), .B(new_n14107_), .ZN(new_n14111_));
  NOR2_X1    g13854(.A1(new_n13804_), .A2(new_n13736_), .ZN(new_n14112_));
  NOR2_X1    g13855(.A1(new_n14112_), .A2(new_n13803_), .ZN(new_n14113_));
  NOR2_X1    g13856(.A1(new_n14111_), .A2(new_n14113_), .ZN(new_n14114_));
  INV_X1     g13857(.I(new_n14114_), .ZN(new_n14115_));
  NAND2_X1   g13858(.A1(new_n14111_), .A2(new_n14113_), .ZN(new_n14116_));
  NAND2_X1   g13859(.A1(new_n14115_), .A2(new_n14116_), .ZN(new_n14117_));
  NAND2_X1   g13860(.A1(new_n14117_), .A2(new_n14040_), .ZN(new_n14118_));
  XNOR2_X1   g13861(.A1(new_n14111_), .A2(new_n14113_), .ZN(new_n14119_));
  OAI21_X1   g13862(.A1(new_n14040_), .A2(new_n14119_), .B(new_n14118_), .ZN(new_n14120_));
  OAI22_X1   g13863(.A1(new_n4208_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n4203_), .ZN(new_n14121_));
  NAND2_X1   g13864(.A1(new_n5244_), .A2(\b[33] ), .ZN(new_n14122_));
  AOI21_X1   g13865(.A1(new_n14121_), .A2(new_n14122_), .B(new_n4211_), .ZN(new_n14123_));
  NAND2_X1   g13866(.A1(new_n3101_), .A2(new_n14123_), .ZN(new_n14124_));
  XOR2_X1    g13867(.A1(new_n14124_), .A2(\a[44] ), .Z(new_n14125_));
  INV_X1     g13868(.I(new_n14125_), .ZN(new_n14126_));
  INV_X1     g13869(.I(new_n13812_), .ZN(new_n14127_));
  OAI21_X1   g13870(.A1(new_n13729_), .A2(new_n13811_), .B(new_n14127_), .ZN(new_n14128_));
  AND2_X2    g13871(.A1(new_n14128_), .A2(new_n14126_), .Z(new_n14129_));
  NOR2_X1    g13872(.A1(new_n14128_), .A2(new_n14126_), .ZN(new_n14130_));
  OAI21_X1   g13873(.A1(new_n14129_), .A2(new_n14130_), .B(new_n14120_), .ZN(new_n14131_));
  XOR2_X1    g13874(.A1(new_n14128_), .A2(new_n14125_), .Z(new_n14132_));
  OAI21_X1   g13875(.A1(new_n14120_), .A2(new_n14132_), .B(new_n14131_), .ZN(new_n14133_));
  NAND2_X1   g13876(.A1(new_n13819_), .A2(new_n13817_), .ZN(new_n14134_));
  NAND2_X1   g13877(.A1(new_n14134_), .A2(new_n13820_), .ZN(new_n14135_));
  XOR2_X1    g13878(.A1(new_n14133_), .A2(new_n14135_), .Z(new_n14136_));
  NAND2_X1   g13879(.A1(new_n14133_), .A2(new_n14135_), .ZN(new_n14137_));
  OR2_X2     g13880(.A1(new_n14133_), .A2(new_n14135_), .Z(new_n14138_));
  AOI21_X1   g13881(.A1(new_n14138_), .A2(new_n14137_), .B(new_n14034_), .ZN(new_n14139_));
  AOI21_X1   g13882(.A1(new_n14034_), .A2(new_n14136_), .B(new_n14139_), .ZN(new_n14140_));
  NAND2_X1   g13883(.A1(new_n13826_), .A2(new_n13825_), .ZN(new_n14141_));
  NAND2_X1   g13884(.A1(new_n14141_), .A2(new_n13828_), .ZN(new_n14142_));
  XOR2_X1    g13885(.A1(new_n14140_), .A2(new_n14142_), .Z(new_n14143_));
  NAND2_X1   g13886(.A1(new_n14140_), .A2(new_n14142_), .ZN(new_n14144_));
  OR2_X2     g13887(.A1(new_n14140_), .A2(new_n14142_), .Z(new_n14145_));
  AOI21_X1   g13888(.A1(new_n14145_), .A2(new_n14144_), .B(new_n14028_), .ZN(new_n14146_));
  AOI21_X1   g13889(.A1(new_n14028_), .A2(new_n14143_), .B(new_n14146_), .ZN(new_n14147_));
  NOR2_X1    g13890(.A1(new_n14147_), .A2(new_n14022_), .ZN(new_n14148_));
  AND2_X2    g13891(.A1(new_n14147_), .A2(new_n14022_), .Z(new_n14149_));
  OAI21_X1   g13892(.A1(new_n14149_), .A2(new_n14148_), .B(new_n14020_), .ZN(new_n14150_));
  XNOR2_X1   g13893(.A1(new_n14147_), .A2(new_n14022_), .ZN(new_n14151_));
  OAI21_X1   g13894(.A1(new_n14020_), .A2(new_n14151_), .B(new_n14150_), .ZN(new_n14152_));
  OAI21_X1   g13895(.A1(new_n13705_), .A2(new_n13847_), .B(new_n13845_), .ZN(new_n14153_));
  AND2_X2    g13896(.A1(new_n14152_), .A2(new_n14153_), .Z(new_n14154_));
  NOR2_X1    g13897(.A1(new_n14152_), .A2(new_n14153_), .ZN(new_n14155_));
  OAI21_X1   g13898(.A1(new_n14154_), .A2(new_n14155_), .B(new_n14014_), .ZN(new_n14156_));
  XNOR2_X1   g13899(.A1(new_n14152_), .A2(new_n14153_), .ZN(new_n14157_));
  OAI21_X1   g13900(.A1(new_n14014_), .A2(new_n14157_), .B(new_n14156_), .ZN(new_n14158_));
  NOR2_X1    g13901(.A1(new_n13852_), .A2(new_n13854_), .ZN(new_n14159_));
  XOR2_X1    g13902(.A1(new_n13858_), .A2(\a[32] ), .Z(new_n14160_));
  NOR3_X1    g13903(.A1(new_n13866_), .A2(new_n13855_), .A3(new_n14160_), .ZN(new_n14161_));
  OAI22_X1   g13904(.A1(new_n2084_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n2079_), .ZN(new_n14162_));
  OAI21_X1   g13905(.A1(new_n5178_), .A2(new_n2214_), .B(new_n14162_), .ZN(new_n14163_));
  AOI21_X1   g13906(.A1(new_n5537_), .A2(new_n2086_), .B(new_n14163_), .ZN(new_n14164_));
  NOR3_X1    g13907(.A1(new_n14159_), .A2(new_n14161_), .A3(new_n14164_), .ZN(new_n14165_));
  NAND2_X1   g13908(.A1(new_n13866_), .A2(new_n13855_), .ZN(new_n14166_));
  INV_X1     g13909(.I(new_n14160_), .ZN(new_n14167_));
  NAND3_X1   g13910(.A1(new_n13852_), .A2(new_n13854_), .A3(new_n14167_), .ZN(new_n14168_));
  INV_X1     g13911(.I(new_n14164_), .ZN(new_n14169_));
  AOI21_X1   g13912(.A1(new_n14168_), .A2(new_n14166_), .B(new_n14169_), .ZN(new_n14170_));
  OAI21_X1   g13913(.A1(new_n14170_), .A2(new_n14165_), .B(new_n2074_), .ZN(new_n14171_));
  NAND3_X1   g13914(.A1(new_n14168_), .A2(new_n14166_), .A3(new_n14169_), .ZN(new_n14172_));
  OAI21_X1   g13915(.A1(new_n14159_), .A2(new_n14161_), .B(new_n14164_), .ZN(new_n14173_));
  NAND3_X1   g13916(.A1(new_n14172_), .A2(new_n14173_), .A3(\a[29] ), .ZN(new_n14174_));
  AOI21_X1   g13917(.A1(new_n14171_), .A2(new_n14174_), .B(new_n14158_), .ZN(new_n14175_));
  INV_X1     g13918(.I(new_n14158_), .ZN(new_n14176_));
  AOI21_X1   g13919(.A1(new_n14172_), .A2(new_n14173_), .B(\a[29] ), .ZN(new_n14177_));
  NOR3_X1    g13920(.A1(new_n14170_), .A2(new_n14165_), .A3(new_n2074_), .ZN(new_n14178_));
  NOR3_X1    g13921(.A1(new_n14177_), .A2(new_n14178_), .A3(new_n14176_), .ZN(new_n14179_));
  OAI21_X1   g13922(.A1(new_n14179_), .A2(new_n14175_), .B(new_n14008_), .ZN(new_n14180_));
  OAI21_X1   g13923(.A1(new_n14177_), .A2(new_n14178_), .B(new_n14176_), .ZN(new_n14181_));
  NAND3_X1   g13924(.A1(new_n14171_), .A2(new_n14174_), .A3(new_n14158_), .ZN(new_n14182_));
  NAND3_X1   g13925(.A1(new_n14181_), .A2(new_n14182_), .A3(new_n14007_), .ZN(new_n14183_));
  AOI21_X1   g13926(.A1(new_n14180_), .A2(new_n14183_), .B(new_n14002_), .ZN(new_n14184_));
  INV_X1     g13927(.I(new_n14002_), .ZN(new_n14185_));
  OAI21_X1   g13928(.A1(new_n14179_), .A2(new_n14175_), .B(new_n14007_), .ZN(new_n14186_));
  NAND3_X1   g13929(.A1(new_n14181_), .A2(new_n14182_), .A3(new_n14008_), .ZN(new_n14187_));
  AOI21_X1   g13930(.A1(new_n14186_), .A2(new_n14187_), .B(new_n14185_), .ZN(new_n14188_));
  OAI21_X1   g13931(.A1(new_n14184_), .A2(new_n14188_), .B(new_n14001_), .ZN(new_n14189_));
  INV_X1     g13932(.I(new_n14001_), .ZN(new_n14190_));
  AOI21_X1   g13933(.A1(new_n14181_), .A2(new_n14182_), .B(new_n14007_), .ZN(new_n14191_));
  NOR3_X1    g13934(.A1(new_n14179_), .A2(new_n14175_), .A3(new_n14008_), .ZN(new_n14192_));
  OAI21_X1   g13935(.A1(new_n14192_), .A2(new_n14191_), .B(new_n14185_), .ZN(new_n14193_));
  AOI21_X1   g13936(.A1(new_n14181_), .A2(new_n14182_), .B(new_n14008_), .ZN(new_n14194_));
  NOR3_X1    g13937(.A1(new_n14179_), .A2(new_n14175_), .A3(new_n14007_), .ZN(new_n14195_));
  OAI21_X1   g13938(.A1(new_n14195_), .A2(new_n14194_), .B(new_n14002_), .ZN(new_n14196_));
  NAND3_X1   g13939(.A1(new_n14193_), .A2(new_n14196_), .A3(new_n14190_), .ZN(new_n14197_));
  AOI21_X1   g13940(.A1(new_n14197_), .A2(new_n14189_), .B(\a[23] ), .ZN(new_n14198_));
  AOI21_X1   g13941(.A1(new_n14193_), .A2(new_n14196_), .B(new_n14190_), .ZN(new_n14199_));
  NOR3_X1    g13942(.A1(new_n14184_), .A2(new_n14188_), .A3(new_n14001_), .ZN(new_n14200_));
  NOR3_X1    g13943(.A1(new_n14199_), .A2(new_n14200_), .A3(new_n1434_), .ZN(new_n14201_));
  OAI21_X1   g13944(.A1(new_n14198_), .A2(new_n14201_), .B(new_n14000_), .ZN(new_n14202_));
  OAI21_X1   g13945(.A1(new_n14199_), .A2(new_n14200_), .B(new_n1434_), .ZN(new_n14203_));
  NAND3_X1   g13946(.A1(new_n14197_), .A2(new_n14189_), .A3(\a[23] ), .ZN(new_n14204_));
  NAND3_X1   g13947(.A1(new_n14203_), .A2(new_n14204_), .A3(new_n13999_), .ZN(new_n14205_));
  OAI22_X1   g13948(.A1(new_n1168_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n1163_), .ZN(new_n14206_));
  NAND2_X1   g13949(.A1(new_n1774_), .A2(\b[57] ), .ZN(new_n14207_));
  AOI21_X1   g13950(.A1(new_n14206_), .A2(new_n14207_), .B(new_n1171_), .ZN(new_n14208_));
  NAND2_X1   g13951(.A1(new_n7895_), .A2(new_n14208_), .ZN(new_n14209_));
  XOR2_X1    g13952(.A1(new_n14209_), .A2(\a[20] ), .Z(new_n14210_));
  INV_X1     g13953(.I(new_n14210_), .ZN(new_n14211_));
  NAND3_X1   g13954(.A1(new_n14202_), .A2(new_n14205_), .A3(new_n14211_), .ZN(new_n14212_));
  INV_X1     g13955(.I(new_n14212_), .ZN(new_n14213_));
  AOI21_X1   g13956(.A1(new_n14202_), .A2(new_n14205_), .B(new_n14211_), .ZN(new_n14214_));
  OAI21_X1   g13957(.A1(new_n14213_), .A2(new_n14214_), .B(new_n13996_), .ZN(new_n14215_));
  AOI21_X1   g13958(.A1(new_n14202_), .A2(new_n14205_), .B(new_n14210_), .ZN(new_n14216_));
  NAND3_X1   g13959(.A1(new_n14202_), .A2(new_n14205_), .A3(new_n14210_), .ZN(new_n14217_));
  INV_X1     g13960(.I(new_n14217_), .ZN(new_n14218_));
  OAI21_X1   g13961(.A1(new_n14218_), .A2(new_n14216_), .B(new_n13995_), .ZN(new_n14219_));
  AOI21_X1   g13962(.A1(new_n14215_), .A2(new_n14219_), .B(new_n13994_), .ZN(new_n14220_));
  INV_X1     g13963(.I(new_n14214_), .ZN(new_n14221_));
  AOI21_X1   g13964(.A1(new_n14221_), .A2(new_n14212_), .B(new_n13995_), .ZN(new_n14222_));
  INV_X1     g13965(.I(new_n14216_), .ZN(new_n14223_));
  AOI21_X1   g13966(.A1(new_n14223_), .A2(new_n14217_), .B(new_n13996_), .ZN(new_n14224_));
  NOR3_X1    g13967(.A1(new_n14222_), .A2(new_n14224_), .A3(new_n13993_), .ZN(new_n14225_));
  OAI21_X1   g13968(.A1(new_n14225_), .A2(new_n14220_), .B(new_n930_), .ZN(new_n14226_));
  OAI21_X1   g13969(.A1(new_n14222_), .A2(new_n14224_), .B(new_n13993_), .ZN(new_n14227_));
  NAND3_X1   g13970(.A1(new_n14215_), .A2(new_n14219_), .A3(new_n13994_), .ZN(new_n14228_));
  NAND3_X1   g13971(.A1(new_n14227_), .A2(new_n14228_), .A3(\a[17] ), .ZN(new_n14229_));
  AOI21_X1   g13972(.A1(new_n14226_), .A2(new_n14229_), .B(new_n13989_), .ZN(new_n14230_));
  AOI21_X1   g13973(.A1(new_n14227_), .A2(new_n14228_), .B(\a[17] ), .ZN(new_n14231_));
  NOR3_X1    g13974(.A1(new_n14225_), .A2(new_n14220_), .A3(new_n930_), .ZN(new_n14232_));
  NOR3_X1    g13975(.A1(new_n14232_), .A2(new_n14231_), .A3(new_n13988_), .ZN(new_n14233_));
  OAI21_X1   g13976(.A1(new_n14233_), .A2(new_n14230_), .B(new_n13985_), .ZN(new_n14234_));
  INV_X1     g13977(.I(new_n13985_), .ZN(new_n14235_));
  OAI21_X1   g13978(.A1(new_n14232_), .A2(new_n14231_), .B(new_n13988_), .ZN(new_n14236_));
  NAND3_X1   g13979(.A1(new_n14226_), .A2(new_n14229_), .A3(new_n13989_), .ZN(new_n14237_));
  NAND3_X1   g13980(.A1(new_n14236_), .A2(new_n14237_), .A3(new_n14235_), .ZN(new_n14238_));
  AOI21_X1   g13981(.A1(new_n14234_), .A2(new_n14238_), .B(\a[14] ), .ZN(new_n14239_));
  AOI21_X1   g13982(.A1(new_n14236_), .A2(new_n14237_), .B(new_n14235_), .ZN(new_n14240_));
  NOR3_X1    g13983(.A1(new_n14233_), .A2(new_n14230_), .A3(new_n13985_), .ZN(new_n14241_));
  NOR3_X1    g13984(.A1(new_n14241_), .A2(new_n14240_), .A3(new_n747_), .ZN(new_n14242_));
  OAI21_X1   g13985(.A1(new_n14242_), .A2(new_n14239_), .B(new_n13984_), .ZN(new_n14243_));
  INV_X1     g13986(.I(new_n13984_), .ZN(new_n14244_));
  OAI21_X1   g13987(.A1(new_n14241_), .A2(new_n14240_), .B(new_n747_), .ZN(new_n14245_));
  NAND3_X1   g13988(.A1(new_n14234_), .A2(new_n14238_), .A3(\a[14] ), .ZN(new_n14246_));
  NAND3_X1   g13989(.A1(new_n14245_), .A2(new_n14246_), .A3(new_n14244_), .ZN(new_n14247_));
  NAND2_X1   g13990(.A1(new_n14243_), .A2(new_n14247_), .ZN(new_n14248_));
  XOR2_X1    g13991(.A1(new_n14248_), .A2(new_n13983_), .Z(new_n14249_));
  NAND2_X1   g13992(.A1(new_n14249_), .A2(new_n13981_), .ZN(new_n14250_));
  XOR2_X1    g13993(.A1(new_n14248_), .A2(new_n13983_), .Z(new_n14251_));
  OAI21_X1   g13994(.A1(new_n13981_), .A2(new_n14251_), .B(new_n14250_), .ZN(\f[77] ));
  NAND2_X1   g13995(.A1(new_n14236_), .A2(new_n14237_), .ZN(new_n14253_));
  XOR2_X1    g13996(.A1(new_n13984_), .A2(\a[14] ), .Z(new_n14254_));
  INV_X1     g13997(.I(new_n14254_), .ZN(new_n14255_));
  XNOR2_X1   g13998(.A1(new_n13985_), .A2(new_n14254_), .ZN(new_n14256_));
  AOI21_X1   g13999(.A1(new_n14253_), .A2(new_n14255_), .B(new_n14256_), .ZN(new_n14257_));
  AOI21_X1   g14000(.A1(new_n14215_), .A2(new_n14219_), .B(new_n13993_), .ZN(new_n14258_));
  XOR2_X1    g14001(.A1(new_n13988_), .A2(new_n930_), .Z(new_n14259_));
  NAND2_X1   g14002(.A1(new_n13993_), .A2(new_n14259_), .ZN(new_n14260_));
  NOR3_X1    g14003(.A1(new_n14222_), .A2(new_n14224_), .A3(new_n14260_), .ZN(new_n14261_));
  NOR2_X1    g14004(.A1(new_n14261_), .A2(new_n14258_), .ZN(new_n14262_));
  AOI21_X1   g14005(.A1(new_n13996_), .A2(new_n14221_), .B(new_n14213_), .ZN(new_n14263_));
  INV_X1     g14006(.I(new_n14263_), .ZN(new_n14264_));
  OAI21_X1   g14007(.A1(new_n14184_), .A2(new_n14188_), .B(new_n14190_), .ZN(new_n14265_));
  NAND2_X1   g14008(.A1(new_n14193_), .A2(new_n14196_), .ZN(new_n14266_));
  NOR2_X1    g14009(.A1(new_n13999_), .A2(new_n1434_), .ZN(new_n14267_));
  NOR2_X1    g14010(.A1(new_n14000_), .A2(\a[23] ), .ZN(new_n14268_));
  OAI22_X1   g14011(.A1(new_n14266_), .A2(new_n14190_), .B1(new_n14267_), .B2(new_n14268_), .ZN(new_n14269_));
  NAND2_X1   g14012(.A1(new_n14269_), .A2(new_n14265_), .ZN(new_n14270_));
  INV_X1     g14013(.I(new_n14270_), .ZN(new_n14271_));
  AOI21_X1   g14014(.A1(new_n14185_), .A2(new_n14183_), .B(new_n14191_), .ZN(new_n14272_));
  INV_X1     g14015(.I(new_n14272_), .ZN(new_n14273_));
  OAI22_X1   g14016(.A1(new_n1760_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n1755_), .ZN(new_n14274_));
  NAND2_X1   g14017(.A1(new_n2470_), .A2(\b[52] ), .ZN(new_n14275_));
  AOI21_X1   g14018(.A1(new_n14274_), .A2(new_n14275_), .B(new_n1763_), .ZN(new_n14276_));
  NAND2_X1   g14019(.A1(new_n6237_), .A2(new_n14276_), .ZN(new_n14277_));
  XOR2_X1    g14020(.A1(new_n14277_), .A2(\a[26] ), .Z(new_n14278_));
  INV_X1     g14021(.I(new_n14278_), .ZN(new_n14279_));
  NAND2_X1   g14022(.A1(new_n14168_), .A2(new_n14166_), .ZN(new_n14280_));
  NAND2_X1   g14023(.A1(new_n14158_), .A2(new_n14280_), .ZN(new_n14281_));
  XOR2_X1    g14024(.A1(new_n14164_), .A2(\a[29] ), .Z(new_n14282_));
  OR2_X2     g14025(.A1(new_n14158_), .A2(new_n14282_), .Z(new_n14283_));
  OAI21_X1   g14026(.A1(new_n14283_), .A2(new_n14280_), .B(new_n14281_), .ZN(new_n14284_));
  INV_X1     g14027(.I(new_n14284_), .ZN(new_n14285_));
  OAI22_X1   g14028(.A1(new_n2084_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n2079_), .ZN(new_n14286_));
  NAND2_X1   g14029(.A1(new_n2864_), .A2(\b[49] ), .ZN(new_n14287_));
  AOI21_X1   g14030(.A1(new_n14286_), .A2(new_n14287_), .B(new_n2087_), .ZN(new_n14288_));
  NAND2_X1   g14031(.A1(new_n5741_), .A2(new_n14288_), .ZN(new_n14289_));
  XOR2_X1    g14032(.A1(new_n14289_), .A2(\a[29] ), .Z(new_n14290_));
  INV_X1     g14033(.I(new_n14290_), .ZN(new_n14291_));
  NOR2_X1    g14034(.A1(new_n14148_), .A2(new_n14019_), .ZN(new_n14292_));
  NOR2_X1    g14035(.A1(new_n14292_), .A2(new_n14149_), .ZN(new_n14293_));
  INV_X1     g14036(.I(new_n14293_), .ZN(new_n14294_));
  NAND2_X1   g14037(.A1(new_n14145_), .A2(new_n14028_), .ZN(new_n14295_));
  NAND2_X1   g14038(.A1(new_n14138_), .A2(new_n14034_), .ZN(new_n14296_));
  NAND2_X1   g14039(.A1(new_n14296_), .A2(new_n14137_), .ZN(new_n14297_));
  INV_X1     g14040(.I(new_n14130_), .ZN(new_n14298_));
  AOI21_X1   g14041(.A1(new_n14298_), .A2(new_n14120_), .B(new_n14129_), .ZN(new_n14299_));
  INV_X1     g14042(.I(new_n14299_), .ZN(new_n14300_));
  AOI21_X1   g14043(.A1(new_n14040_), .A2(new_n14116_), .B(new_n14114_), .ZN(new_n14301_));
  NAND2_X1   g14044(.A1(new_n14094_), .A2(new_n14093_), .ZN(new_n14302_));
  NAND2_X1   g14045(.A1(new_n14095_), .A2(new_n14302_), .ZN(new_n14303_));
  INV_X1     g14046(.I(new_n14303_), .ZN(new_n14304_));
  AOI21_X1   g14047(.A1(new_n14085_), .A2(new_n14088_), .B(new_n14086_), .ZN(new_n14305_));
  INV_X1     g14048(.I(new_n14305_), .ZN(new_n14306_));
  INV_X1     g14049(.I(new_n14052_), .ZN(new_n14307_));
  NAND2_X1   g14050(.A1(new_n14070_), .A2(new_n14307_), .ZN(new_n14308_));
  NAND2_X1   g14051(.A1(new_n14308_), .A2(new_n14071_), .ZN(new_n14309_));
  OAI22_X1   g14052(.A1(new_n1124_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1044_), .ZN(new_n14310_));
  NAND2_X1   g14053(.A1(new_n9644_), .A2(\b[16] ), .ZN(new_n14311_));
  AOI21_X1   g14054(.A1(new_n14311_), .A2(new_n14310_), .B(new_n8321_), .ZN(new_n14312_));
  NAND2_X1   g14055(.A1(new_n1123_), .A2(new_n14312_), .ZN(new_n14313_));
  XOR2_X1    g14056(.A1(new_n14313_), .A2(\a[62] ), .Z(new_n14314_));
  INV_X1     g14057(.I(new_n14314_), .ZN(new_n14315_));
  AOI21_X1   g14058(.A1(new_n13758_), .A2(new_n14061_), .B(new_n14058_), .ZN(new_n14316_));
  NOR2_X1    g14059(.A1(new_n14316_), .A2(new_n14065_), .ZN(new_n14317_));
  NOR2_X1    g14060(.A1(new_n8985_), .A2(new_n904_), .ZN(new_n14318_));
  NOR2_X1    g14061(.A1(new_n9364_), .A2(new_n848_), .ZN(new_n14319_));
  XNOR2_X1   g14062(.A1(new_n14318_), .A2(new_n14319_), .ZN(new_n14320_));
  NOR2_X1    g14063(.A1(new_n14320_), .A2(new_n747_), .ZN(new_n14321_));
  INV_X1     g14064(.I(new_n14321_), .ZN(new_n14322_));
  NAND2_X1   g14065(.A1(new_n14320_), .A2(new_n747_), .ZN(new_n14323_));
  AOI21_X1   g14066(.A1(new_n14322_), .A2(new_n14323_), .B(new_n13753_), .ZN(new_n14324_));
  XOR2_X1    g14067(.A1(new_n14320_), .A2(\a[14] ), .Z(new_n14325_));
  NOR2_X1    g14068(.A1(new_n14325_), .A2(new_n13758_), .ZN(new_n14326_));
  NOR2_X1    g14069(.A1(new_n14326_), .A2(new_n14324_), .ZN(new_n14327_));
  XOR2_X1    g14070(.A1(new_n14317_), .A2(new_n14327_), .Z(new_n14328_));
  NAND2_X1   g14071(.A1(new_n14328_), .A2(new_n14315_), .ZN(new_n14329_));
  NOR2_X1    g14072(.A1(new_n14317_), .A2(new_n14327_), .ZN(new_n14330_));
  NOR4_X1    g14073(.A1(new_n14316_), .A2(new_n14065_), .A3(new_n14324_), .A4(new_n14326_), .ZN(new_n14331_));
  OAI21_X1   g14074(.A1(new_n14330_), .A2(new_n14331_), .B(new_n14314_), .ZN(new_n14332_));
  NAND2_X1   g14075(.A1(new_n14329_), .A2(new_n14332_), .ZN(new_n14333_));
  OAI22_X1   g14076(.A1(new_n1393_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1305_), .ZN(new_n14334_));
  NAND2_X1   g14077(.A1(new_n8628_), .A2(\b[19] ), .ZN(new_n14335_));
  AOI21_X1   g14078(.A1(new_n14335_), .A2(new_n14334_), .B(new_n7354_), .ZN(new_n14336_));
  NAND2_X1   g14079(.A1(new_n1396_), .A2(new_n14336_), .ZN(new_n14337_));
  XOR2_X1    g14080(.A1(new_n14337_), .A2(\a[59] ), .Z(new_n14338_));
  XOR2_X1    g14081(.A1(new_n14333_), .A2(new_n14338_), .Z(new_n14339_));
  NAND2_X1   g14082(.A1(new_n14339_), .A2(new_n14309_), .ZN(new_n14340_));
  INV_X1     g14083(.I(new_n14309_), .ZN(new_n14341_));
  NOR2_X1    g14084(.A1(new_n14333_), .A2(new_n14338_), .ZN(new_n14342_));
  AND2_X2    g14085(.A1(new_n14333_), .A2(new_n14338_), .Z(new_n14343_));
  OAI21_X1   g14086(.A1(new_n14343_), .A2(new_n14342_), .B(new_n14341_), .ZN(new_n14344_));
  NAND2_X1   g14087(.A1(new_n14340_), .A2(new_n14344_), .ZN(new_n14345_));
  OAI22_X1   g14088(.A1(new_n6721_), .A2(new_n1601_), .B1(new_n6723_), .B2(new_n1709_), .ZN(new_n14346_));
  NAND2_X1   g14089(.A1(new_n7617_), .A2(\b[22] ), .ZN(new_n14347_));
  AOI21_X1   g14090(.A1(new_n14347_), .A2(new_n14346_), .B(new_n6731_), .ZN(new_n14348_));
  NAND2_X1   g14091(.A1(new_n1708_), .A2(new_n14348_), .ZN(new_n14349_));
  XOR2_X1    g14092(.A1(new_n14349_), .A2(\a[56] ), .Z(new_n14350_));
  NOR2_X1    g14093(.A1(new_n14345_), .A2(new_n14350_), .ZN(new_n14351_));
  NAND2_X1   g14094(.A1(new_n14345_), .A2(new_n14350_), .ZN(new_n14352_));
  INV_X1     g14095(.I(new_n14352_), .ZN(new_n14353_));
  OAI21_X1   g14096(.A1(new_n14353_), .A2(new_n14351_), .B(new_n14306_), .ZN(new_n14354_));
  XNOR2_X1   g14097(.A1(new_n14345_), .A2(new_n14350_), .ZN(new_n14355_));
  OAI21_X1   g14098(.A1(new_n14306_), .A2(new_n14355_), .B(new_n14354_), .ZN(new_n14356_));
  OAI22_X1   g14099(.A1(new_n5786_), .A2(new_n2039_), .B1(new_n1927_), .B2(new_n5792_), .ZN(new_n14357_));
  NAND2_X1   g14100(.A1(new_n6745_), .A2(\b[25] ), .ZN(new_n14358_));
  AOI21_X1   g14101(.A1(new_n14358_), .A2(new_n14357_), .B(new_n5796_), .ZN(new_n14359_));
  NAND2_X1   g14102(.A1(new_n2042_), .A2(new_n14359_), .ZN(new_n14360_));
  XOR2_X1    g14103(.A1(new_n14360_), .A2(\a[53] ), .Z(new_n14361_));
  XOR2_X1    g14104(.A1(new_n14356_), .A2(new_n14361_), .Z(new_n14362_));
  INV_X1     g14105(.I(new_n14361_), .ZN(new_n14363_));
  AND2_X2    g14106(.A1(new_n14356_), .A2(new_n14363_), .Z(new_n14364_));
  NOR2_X1    g14107(.A1(new_n14356_), .A2(new_n14363_), .ZN(new_n14365_));
  OAI21_X1   g14108(.A1(new_n14364_), .A2(new_n14365_), .B(new_n14304_), .ZN(new_n14366_));
  OAI21_X1   g14109(.A1(new_n14362_), .A2(new_n14304_), .B(new_n14366_), .ZN(new_n14367_));
  OAI22_X1   g14110(.A1(new_n5228_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n5225_), .ZN(new_n14368_));
  NAND2_X1   g14111(.A1(new_n5387_), .A2(\b[28] ), .ZN(new_n14369_));
  AOI21_X1   g14112(.A1(new_n14368_), .A2(new_n14369_), .B(new_n5231_), .ZN(new_n14370_));
  NAND2_X1   g14113(.A1(new_n2404_), .A2(new_n14370_), .ZN(new_n14371_));
  XOR2_X1    g14114(.A1(new_n14371_), .A2(\a[50] ), .Z(new_n14372_));
  NAND2_X1   g14115(.A1(new_n14097_), .A2(new_n14109_), .ZN(new_n14373_));
  AOI21_X1   g14116(.A1(new_n14373_), .A2(new_n14108_), .B(new_n14372_), .ZN(new_n14374_));
  INV_X1     g14117(.I(new_n14372_), .ZN(new_n14375_));
  NAND2_X1   g14118(.A1(new_n14373_), .A2(new_n14108_), .ZN(new_n14376_));
  NOR2_X1    g14119(.A1(new_n14376_), .A2(new_n14375_), .ZN(new_n14377_));
  OAI21_X1   g14120(.A1(new_n14374_), .A2(new_n14377_), .B(new_n14367_), .ZN(new_n14378_));
  XOR2_X1    g14121(.A1(new_n14376_), .A2(new_n14372_), .Z(new_n14379_));
  OR2_X2     g14122(.A1(new_n14367_), .A2(new_n14379_), .Z(new_n14380_));
  OAI22_X1   g14123(.A1(new_n4711_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n4706_), .ZN(new_n14381_));
  NAND2_X1   g14124(.A1(new_n5814_), .A2(\b[31] ), .ZN(new_n14382_));
  AOI21_X1   g14125(.A1(new_n14381_), .A2(new_n14382_), .B(new_n4714_), .ZN(new_n14383_));
  NAND2_X1   g14126(.A1(new_n2797_), .A2(new_n14383_), .ZN(new_n14384_));
  XOR2_X1    g14127(.A1(new_n14384_), .A2(\a[47] ), .Z(new_n14385_));
  INV_X1     g14128(.I(new_n14385_), .ZN(new_n14386_));
  NAND3_X1   g14129(.A1(new_n14380_), .A2(new_n14378_), .A3(new_n14386_), .ZN(new_n14387_));
  NAND2_X1   g14130(.A1(new_n14380_), .A2(new_n14378_), .ZN(new_n14388_));
  NAND2_X1   g14131(.A1(new_n14388_), .A2(new_n14385_), .ZN(new_n14389_));
  AOI21_X1   g14132(.A1(new_n14389_), .A2(new_n14387_), .B(new_n14301_), .ZN(new_n14390_));
  INV_X1     g14133(.I(new_n14301_), .ZN(new_n14391_));
  XOR2_X1    g14134(.A1(new_n14388_), .A2(new_n14386_), .Z(new_n14392_));
  NOR2_X1    g14135(.A1(new_n14392_), .A2(new_n14391_), .ZN(new_n14393_));
  NOR2_X1    g14136(.A1(new_n14393_), .A2(new_n14390_), .ZN(new_n14394_));
  OAI22_X1   g14137(.A1(new_n4208_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n4203_), .ZN(new_n14395_));
  NAND2_X1   g14138(.A1(new_n5244_), .A2(\b[34] ), .ZN(new_n14396_));
  AOI21_X1   g14139(.A1(new_n14395_), .A2(new_n14396_), .B(new_n4211_), .ZN(new_n14397_));
  NAND2_X1   g14140(.A1(new_n3246_), .A2(new_n14397_), .ZN(new_n14398_));
  XOR2_X1    g14141(.A1(new_n14398_), .A2(\a[44] ), .Z(new_n14399_));
  XOR2_X1    g14142(.A1(new_n14394_), .A2(new_n14399_), .Z(new_n14400_));
  NAND2_X1   g14143(.A1(new_n14400_), .A2(new_n14300_), .ZN(new_n14401_));
  NOR2_X1    g14144(.A1(new_n14394_), .A2(new_n14399_), .ZN(new_n14402_));
  AND2_X2    g14145(.A1(new_n14394_), .A2(new_n14399_), .Z(new_n14403_));
  OAI21_X1   g14146(.A1(new_n14403_), .A2(new_n14402_), .B(new_n14299_), .ZN(new_n14404_));
  NAND2_X1   g14147(.A1(new_n14401_), .A2(new_n14404_), .ZN(new_n14405_));
  OAI22_X1   g14148(.A1(new_n3736_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n3731_), .ZN(new_n14406_));
  NAND2_X1   g14149(.A1(new_n4730_), .A2(\b[37] ), .ZN(new_n14407_));
  AOI21_X1   g14150(.A1(new_n14406_), .A2(new_n14407_), .B(new_n3739_), .ZN(new_n14408_));
  NAND2_X1   g14151(.A1(new_n3700_), .A2(new_n14408_), .ZN(new_n14409_));
  XOR2_X1    g14152(.A1(new_n14409_), .A2(\a[41] ), .Z(new_n14410_));
  NOR2_X1    g14153(.A1(new_n14405_), .A2(new_n14410_), .ZN(new_n14411_));
  INV_X1     g14154(.I(new_n14410_), .ZN(new_n14412_));
  AOI21_X1   g14155(.A1(new_n14401_), .A2(new_n14404_), .B(new_n14412_), .ZN(new_n14413_));
  OAI21_X1   g14156(.A1(new_n14411_), .A2(new_n14413_), .B(new_n14297_), .ZN(new_n14414_));
  XOR2_X1    g14157(.A1(new_n14405_), .A2(new_n14412_), .Z(new_n14415_));
  OAI21_X1   g14158(.A1(new_n14415_), .A2(new_n14297_), .B(new_n14414_), .ZN(new_n14416_));
  OAI22_X1   g14159(.A1(new_n3298_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n3293_), .ZN(new_n14417_));
  NAND2_X1   g14160(.A1(new_n4227_), .A2(\b[40] ), .ZN(new_n14418_));
  AOI21_X1   g14161(.A1(new_n14417_), .A2(new_n14418_), .B(new_n3301_), .ZN(new_n14419_));
  NAND2_X1   g14162(.A1(new_n4017_), .A2(new_n14419_), .ZN(new_n14420_));
  XOR2_X1    g14163(.A1(new_n14420_), .A2(\a[38] ), .Z(new_n14421_));
  XOR2_X1    g14164(.A1(new_n14416_), .A2(new_n14421_), .Z(new_n14422_));
  AOI21_X1   g14165(.A1(new_n14144_), .A2(new_n14295_), .B(new_n14422_), .ZN(new_n14423_));
  NAND2_X1   g14166(.A1(new_n14295_), .A2(new_n14144_), .ZN(new_n14424_));
  INV_X1     g14167(.I(new_n14421_), .ZN(new_n14425_));
  NAND2_X1   g14168(.A1(new_n14416_), .A2(new_n14425_), .ZN(new_n14426_));
  OR2_X2     g14169(.A1(new_n14416_), .A2(new_n14425_), .Z(new_n14427_));
  AOI21_X1   g14170(.A1(new_n14427_), .A2(new_n14426_), .B(new_n14424_), .ZN(new_n14428_));
  NOR2_X1    g14171(.A1(new_n14423_), .A2(new_n14428_), .ZN(new_n14429_));
  OAI22_X1   g14172(.A1(new_n2846_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n2841_), .ZN(new_n14430_));
  NAND2_X1   g14173(.A1(new_n3755_), .A2(\b[43] ), .ZN(new_n14431_));
  AOI21_X1   g14174(.A1(new_n14430_), .A2(new_n14431_), .B(new_n2849_), .ZN(new_n14432_));
  NAND2_X1   g14175(.A1(new_n4513_), .A2(new_n14432_), .ZN(new_n14433_));
  XOR2_X1    g14176(.A1(new_n14433_), .A2(\a[35] ), .Z(new_n14434_));
  INV_X1     g14177(.I(new_n14434_), .ZN(new_n14435_));
  XOR2_X1    g14178(.A1(new_n14429_), .A2(new_n14435_), .Z(new_n14436_));
  NAND2_X1   g14179(.A1(new_n14436_), .A2(new_n14294_), .ZN(new_n14437_));
  NAND2_X1   g14180(.A1(new_n14429_), .A2(new_n14435_), .ZN(new_n14438_));
  OAI21_X1   g14181(.A1(new_n14423_), .A2(new_n14428_), .B(new_n14434_), .ZN(new_n14439_));
  NAND2_X1   g14182(.A1(new_n14438_), .A2(new_n14439_), .ZN(new_n14440_));
  NAND2_X1   g14183(.A1(new_n14440_), .A2(new_n14293_), .ZN(new_n14441_));
  NAND2_X1   g14184(.A1(new_n14437_), .A2(new_n14441_), .ZN(new_n14442_));
  NOR2_X1    g14185(.A1(new_n14155_), .A2(new_n14013_), .ZN(new_n14443_));
  NOR2_X1    g14186(.A1(new_n14443_), .A2(new_n14154_), .ZN(new_n14444_));
  OAI22_X1   g14187(.A1(new_n2452_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n2447_), .ZN(new_n14445_));
  NAND2_X1   g14188(.A1(new_n3312_), .A2(\b[46] ), .ZN(new_n14446_));
  AOI21_X1   g14189(.A1(new_n14445_), .A2(new_n14446_), .B(new_n2455_), .ZN(new_n14447_));
  NAND2_X1   g14190(.A1(new_n5177_), .A2(new_n14447_), .ZN(new_n14448_));
  XOR2_X1    g14191(.A1(new_n14448_), .A2(\a[32] ), .Z(new_n14449_));
  NOR2_X1    g14192(.A1(new_n14444_), .A2(new_n14449_), .ZN(new_n14450_));
  AND2_X2    g14193(.A1(new_n14444_), .A2(new_n14449_), .Z(new_n14451_));
  OAI21_X1   g14194(.A1(new_n14451_), .A2(new_n14450_), .B(new_n14442_), .ZN(new_n14452_));
  XOR2_X1    g14195(.A1(new_n14444_), .A2(new_n14449_), .Z(new_n14453_));
  NAND3_X1   g14196(.A1(new_n14453_), .A2(new_n14437_), .A3(new_n14441_), .ZN(new_n14454_));
  AOI21_X1   g14197(.A1(new_n14454_), .A2(new_n14452_), .B(new_n14291_), .ZN(new_n14455_));
  INV_X1     g14198(.I(new_n14455_), .ZN(new_n14456_));
  NAND3_X1   g14199(.A1(new_n14454_), .A2(new_n14452_), .A3(new_n14291_), .ZN(new_n14457_));
  AOI21_X1   g14200(.A1(new_n14456_), .A2(new_n14457_), .B(new_n14285_), .ZN(new_n14458_));
  INV_X1     g14201(.I(new_n14458_), .ZN(new_n14459_));
  NAND2_X1   g14202(.A1(new_n14454_), .A2(new_n14452_), .ZN(new_n14460_));
  NAND2_X1   g14203(.A1(new_n14460_), .A2(new_n14291_), .ZN(new_n14461_));
  NAND3_X1   g14204(.A1(new_n14454_), .A2(new_n14452_), .A3(new_n14290_), .ZN(new_n14462_));
  AOI21_X1   g14205(.A1(new_n14461_), .A2(new_n14462_), .B(new_n14284_), .ZN(new_n14463_));
  INV_X1     g14206(.I(new_n14463_), .ZN(new_n14464_));
  AOI21_X1   g14207(.A1(new_n14464_), .A2(new_n14459_), .B(new_n14279_), .ZN(new_n14465_));
  NOR3_X1    g14208(.A1(new_n14458_), .A2(new_n14463_), .A3(new_n14278_), .ZN(new_n14466_));
  OAI21_X1   g14209(.A1(new_n14465_), .A2(new_n14466_), .B(new_n14273_), .ZN(new_n14467_));
  OAI21_X1   g14210(.A1(new_n14458_), .A2(new_n14463_), .B(new_n14279_), .ZN(new_n14468_));
  INV_X1     g14211(.I(new_n14468_), .ZN(new_n14469_));
  NOR3_X1    g14212(.A1(new_n14458_), .A2(new_n14463_), .A3(new_n14279_), .ZN(new_n14470_));
  OAI21_X1   g14213(.A1(new_n14469_), .A2(new_n14470_), .B(new_n14272_), .ZN(new_n14471_));
  OAI22_X1   g14214(.A1(new_n1444_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n1439_), .ZN(new_n14472_));
  NAND2_X1   g14215(.A1(new_n2098_), .A2(\b[55] ), .ZN(new_n14473_));
  AOI21_X1   g14216(.A1(new_n14472_), .A2(new_n14473_), .B(new_n1447_), .ZN(new_n14474_));
  NAND2_X1   g14217(.A1(new_n7308_), .A2(new_n14474_), .ZN(new_n14475_));
  XOR2_X1    g14218(.A1(new_n14475_), .A2(\a[23] ), .Z(new_n14476_));
  INV_X1     g14219(.I(new_n14476_), .ZN(new_n14477_));
  NAND3_X1   g14220(.A1(new_n14467_), .A2(new_n14471_), .A3(new_n14477_), .ZN(new_n14478_));
  AOI21_X1   g14221(.A1(new_n14467_), .A2(new_n14471_), .B(new_n14477_), .ZN(new_n14479_));
  INV_X1     g14222(.I(new_n14479_), .ZN(new_n14480_));
  AOI21_X1   g14223(.A1(new_n14480_), .A2(new_n14478_), .B(new_n14271_), .ZN(new_n14481_));
  INV_X1     g14224(.I(new_n14467_), .ZN(new_n14482_));
  INV_X1     g14225(.I(new_n14470_), .ZN(new_n14483_));
  AOI21_X1   g14226(.A1(new_n14483_), .A2(new_n14468_), .B(new_n14273_), .ZN(new_n14484_));
  OAI21_X1   g14227(.A1(new_n14482_), .A2(new_n14484_), .B(new_n14477_), .ZN(new_n14485_));
  NAND3_X1   g14228(.A1(new_n14467_), .A2(new_n14471_), .A3(new_n14476_), .ZN(new_n14486_));
  AOI21_X1   g14229(.A1(new_n14485_), .A2(new_n14486_), .B(new_n14270_), .ZN(new_n14487_));
  OAI22_X1   g14230(.A1(new_n1168_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n1163_), .ZN(new_n14488_));
  NAND2_X1   g14231(.A1(new_n1774_), .A2(\b[58] ), .ZN(new_n14489_));
  AOI21_X1   g14232(.A1(new_n14488_), .A2(new_n14489_), .B(new_n1171_), .ZN(new_n14490_));
  NAND2_X1   g14233(.A1(new_n7929_), .A2(new_n14490_), .ZN(new_n14491_));
  XOR2_X1    g14234(.A1(new_n14491_), .A2(\a[20] ), .Z(new_n14492_));
  NOR3_X1    g14235(.A1(new_n14481_), .A2(new_n14487_), .A3(new_n14492_), .ZN(new_n14493_));
  INV_X1     g14236(.I(new_n14478_), .ZN(new_n14494_));
  OAI21_X1   g14237(.A1(new_n14494_), .A2(new_n14479_), .B(new_n14270_), .ZN(new_n14495_));
  AOI21_X1   g14238(.A1(new_n14467_), .A2(new_n14471_), .B(new_n14476_), .ZN(new_n14496_));
  NOR3_X1    g14239(.A1(new_n14482_), .A2(new_n14484_), .A3(new_n14477_), .ZN(new_n14497_));
  OAI21_X1   g14240(.A1(new_n14497_), .A2(new_n14496_), .B(new_n14271_), .ZN(new_n14498_));
  INV_X1     g14241(.I(new_n14492_), .ZN(new_n14499_));
  AOI21_X1   g14242(.A1(new_n14495_), .A2(new_n14498_), .B(new_n14499_), .ZN(new_n14500_));
  OAI21_X1   g14243(.A1(new_n14500_), .A2(new_n14493_), .B(new_n14264_), .ZN(new_n14501_));
  AOI21_X1   g14244(.A1(new_n14495_), .A2(new_n14498_), .B(new_n14492_), .ZN(new_n14502_));
  NOR3_X1    g14245(.A1(new_n14481_), .A2(new_n14487_), .A3(new_n14499_), .ZN(new_n14503_));
  OAI21_X1   g14246(.A1(new_n14502_), .A2(new_n14503_), .B(new_n14263_), .ZN(new_n14504_));
  OAI22_X1   g14247(.A1(new_n940_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n935_), .ZN(new_n14505_));
  NAND2_X1   g14248(.A1(new_n1458_), .A2(\b[61] ), .ZN(new_n14506_));
  AOI21_X1   g14249(.A1(new_n14505_), .A2(new_n14506_), .B(new_n943_), .ZN(new_n14507_));
  NAND2_X1   g14250(.A1(new_n8963_), .A2(new_n14507_), .ZN(new_n14508_));
  XOR2_X1    g14251(.A1(new_n14508_), .A2(\a[17] ), .Z(new_n14509_));
  INV_X1     g14252(.I(new_n14509_), .ZN(new_n14510_));
  NAND3_X1   g14253(.A1(new_n14501_), .A2(new_n14504_), .A3(new_n14510_), .ZN(new_n14511_));
  NAND3_X1   g14254(.A1(new_n14495_), .A2(new_n14498_), .A3(new_n14499_), .ZN(new_n14512_));
  OAI21_X1   g14255(.A1(new_n14481_), .A2(new_n14487_), .B(new_n14492_), .ZN(new_n14513_));
  AOI21_X1   g14256(.A1(new_n14513_), .A2(new_n14512_), .B(new_n14263_), .ZN(new_n14514_));
  OAI21_X1   g14257(.A1(new_n14481_), .A2(new_n14487_), .B(new_n14499_), .ZN(new_n14515_));
  NAND3_X1   g14258(.A1(new_n14495_), .A2(new_n14498_), .A3(new_n14492_), .ZN(new_n14516_));
  AOI21_X1   g14259(.A1(new_n14515_), .A2(new_n14516_), .B(new_n14264_), .ZN(new_n14517_));
  OAI21_X1   g14260(.A1(new_n14517_), .A2(new_n14514_), .B(new_n14509_), .ZN(new_n14518_));
  AOI21_X1   g14261(.A1(new_n14518_), .A2(new_n14511_), .B(new_n14262_), .ZN(new_n14519_));
  INV_X1     g14262(.I(new_n14262_), .ZN(new_n14520_));
  OAI21_X1   g14263(.A1(new_n14517_), .A2(new_n14514_), .B(new_n14510_), .ZN(new_n14521_));
  NAND3_X1   g14264(.A1(new_n14501_), .A2(new_n14504_), .A3(new_n14509_), .ZN(new_n14522_));
  AOI21_X1   g14265(.A1(new_n14521_), .A2(new_n14522_), .B(new_n14520_), .ZN(new_n14523_));
  NOR2_X1    g14266(.A1(new_n14519_), .A2(new_n14523_), .ZN(new_n14524_));
  XNOR2_X1   g14267(.A1(new_n14524_), .A2(new_n14257_), .ZN(new_n14525_));
  NOR2_X1    g14268(.A1(new_n13973_), .A2(new_n13972_), .ZN(new_n14526_));
  INV_X1     g14269(.I(new_n14526_), .ZN(new_n14527_));
  INV_X1     g14270(.I(new_n13983_), .ZN(new_n14528_));
  NAND3_X1   g14271(.A1(new_n13975_), .A2(new_n14527_), .A3(new_n14528_), .ZN(new_n14529_));
  NAND2_X1   g14272(.A1(new_n13981_), .A2(new_n13983_), .ZN(new_n14530_));
  AOI21_X1   g14273(.A1(new_n14530_), .A2(new_n14529_), .B(new_n14248_), .ZN(new_n14531_));
  XOR2_X1    g14274(.A1(new_n14531_), .A2(new_n14525_), .Z(new_n14532_));
  INV_X1     g14275(.I(new_n13981_), .ZN(new_n14533_));
  NOR2_X1    g14276(.A1(new_n14533_), .A2(new_n13983_), .ZN(new_n14534_));
  XOR2_X1    g14277(.A1(new_n14532_), .A2(new_n14534_), .Z(\f[78] ));
  NAND2_X1   g14278(.A1(new_n14518_), .A2(new_n14520_), .ZN(new_n14536_));
  NAND2_X1   g14279(.A1(new_n14536_), .A2(new_n14511_), .ZN(new_n14537_));
  INV_X1     g14280(.I(new_n14537_), .ZN(new_n14538_));
  AOI21_X1   g14281(.A1(new_n14264_), .A2(new_n14516_), .B(new_n14502_), .ZN(new_n14539_));
  INV_X1     g14282(.I(new_n14539_), .ZN(new_n14540_));
  AOI21_X1   g14283(.A1(new_n14270_), .A2(new_n14480_), .B(new_n14494_), .ZN(new_n14541_));
  OAI22_X1   g14284(.A1(new_n1760_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n1755_), .ZN(new_n14542_));
  NAND2_X1   g14285(.A1(new_n2470_), .A2(\b[53] ), .ZN(new_n14543_));
  AOI21_X1   g14286(.A1(new_n14542_), .A2(new_n14543_), .B(new_n1763_), .ZN(new_n14544_));
  NAND2_X1   g14287(.A1(new_n6471_), .A2(new_n14544_), .ZN(new_n14545_));
  XOR2_X1    g14288(.A1(new_n14545_), .A2(\a[26] ), .Z(new_n14546_));
  OAI21_X1   g14289(.A1(new_n14285_), .A2(new_n14455_), .B(new_n14457_), .ZN(new_n14547_));
  INV_X1     g14290(.I(new_n14547_), .ZN(new_n14548_));
  OAI22_X1   g14291(.A1(new_n2452_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n2447_), .ZN(new_n14549_));
  NAND2_X1   g14292(.A1(new_n3312_), .A2(\b[47] ), .ZN(new_n14550_));
  AOI21_X1   g14293(.A1(new_n14549_), .A2(new_n14550_), .B(new_n2455_), .ZN(new_n14551_));
  NAND2_X1   g14294(.A1(new_n5196_), .A2(new_n14551_), .ZN(new_n14552_));
  XOR2_X1    g14295(.A1(new_n14552_), .A2(\a[32] ), .Z(new_n14553_));
  INV_X1     g14296(.I(new_n14553_), .ZN(new_n14554_));
  NAND2_X1   g14297(.A1(new_n14439_), .A2(new_n14294_), .ZN(new_n14555_));
  NAND2_X1   g14298(.A1(new_n14555_), .A2(new_n14438_), .ZN(new_n14556_));
  OAI22_X1   g14299(.A1(new_n2846_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n2841_), .ZN(new_n14557_));
  NAND2_X1   g14300(.A1(new_n3755_), .A2(\b[44] ), .ZN(new_n14558_));
  AOI21_X1   g14301(.A1(new_n14557_), .A2(new_n14558_), .B(new_n2849_), .ZN(new_n14559_));
  NAND2_X1   g14302(.A1(new_n4833_), .A2(new_n14559_), .ZN(new_n14560_));
  XOR2_X1    g14303(.A1(new_n14560_), .A2(\a[35] ), .Z(new_n14561_));
  INV_X1     g14304(.I(new_n14561_), .ZN(new_n14562_));
  INV_X1     g14305(.I(new_n14413_), .ZN(new_n14563_));
  AOI21_X1   g14306(.A1(new_n14297_), .A2(new_n14563_), .B(new_n14411_), .ZN(new_n14564_));
  OAI22_X1   g14307(.A1(new_n3736_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n3731_), .ZN(new_n14565_));
  NAND2_X1   g14308(.A1(new_n4730_), .A2(\b[38] ), .ZN(new_n14566_));
  AOI21_X1   g14309(.A1(new_n14565_), .A2(new_n14566_), .B(new_n3739_), .ZN(new_n14567_));
  NAND2_X1   g14310(.A1(new_n3844_), .A2(new_n14567_), .ZN(new_n14568_));
  XOR2_X1    g14311(.A1(new_n14568_), .A2(\a[41] ), .Z(new_n14569_));
  INV_X1     g14312(.I(new_n14569_), .ZN(new_n14570_));
  NOR2_X1    g14313(.A1(new_n14403_), .A2(new_n14299_), .ZN(new_n14571_));
  NOR2_X1    g14314(.A1(new_n14571_), .A2(new_n14402_), .ZN(new_n14572_));
  OAI22_X1   g14315(.A1(new_n4208_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n4203_), .ZN(new_n14573_));
  NAND2_X1   g14316(.A1(new_n5244_), .A2(\b[35] ), .ZN(new_n14574_));
  AOI21_X1   g14317(.A1(new_n14573_), .A2(new_n14574_), .B(new_n4211_), .ZN(new_n14575_));
  NAND2_X1   g14318(.A1(new_n3411_), .A2(new_n14575_), .ZN(new_n14576_));
  XOR2_X1    g14319(.A1(new_n14576_), .A2(\a[44] ), .Z(new_n14577_));
  INV_X1     g14320(.I(new_n14577_), .ZN(new_n14578_));
  NAND2_X1   g14321(.A1(new_n14389_), .A2(new_n14391_), .ZN(new_n14579_));
  NAND2_X1   g14322(.A1(new_n14579_), .A2(new_n14387_), .ZN(new_n14580_));
  OAI22_X1   g14323(.A1(new_n4711_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n4706_), .ZN(new_n14581_));
  NAND2_X1   g14324(.A1(new_n5814_), .A2(\b[32] ), .ZN(new_n14582_));
  AOI21_X1   g14325(.A1(new_n14581_), .A2(new_n14582_), .B(new_n4714_), .ZN(new_n14583_));
  NAND2_X1   g14326(.A1(new_n2963_), .A2(new_n14583_), .ZN(new_n14584_));
  XOR2_X1    g14327(.A1(new_n14584_), .A2(\a[47] ), .Z(new_n14585_));
  OAI22_X1   g14328(.A1(new_n5786_), .A2(new_n2175_), .B1(new_n2039_), .B2(new_n5792_), .ZN(new_n14586_));
  NAND2_X1   g14329(.A1(new_n6745_), .A2(\b[26] ), .ZN(new_n14587_));
  AOI21_X1   g14330(.A1(new_n14587_), .A2(new_n14586_), .B(new_n5796_), .ZN(new_n14588_));
  NAND2_X1   g14331(.A1(new_n2174_), .A2(new_n14588_), .ZN(new_n14589_));
  XOR2_X1    g14332(.A1(new_n14589_), .A2(\a[53] ), .Z(new_n14590_));
  INV_X1     g14333(.I(new_n14351_), .ZN(new_n14591_));
  NAND2_X1   g14334(.A1(new_n14352_), .A2(new_n14306_), .ZN(new_n14592_));
  NAND2_X1   g14335(.A1(new_n14592_), .A2(new_n14591_), .ZN(new_n14593_));
  OAI22_X1   g14336(.A1(new_n1518_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1393_), .ZN(new_n14594_));
  NAND2_X1   g14337(.A1(new_n8628_), .A2(\b[20] ), .ZN(new_n14595_));
  AOI21_X1   g14338(.A1(new_n14595_), .A2(new_n14594_), .B(new_n7354_), .ZN(new_n14596_));
  NAND2_X1   g14339(.A1(new_n1517_), .A2(new_n14596_), .ZN(new_n14597_));
  XOR2_X1    g14340(.A1(new_n14597_), .A2(\a[59] ), .Z(new_n14598_));
  NOR2_X1    g14341(.A1(new_n14331_), .A2(new_n14314_), .ZN(new_n14599_));
  NOR2_X1    g14342(.A1(new_n14599_), .A2(new_n14330_), .ZN(new_n14600_));
  OAI22_X1   g14343(.A1(new_n1222_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1124_), .ZN(new_n14601_));
  NAND2_X1   g14344(.A1(new_n9644_), .A2(\b[17] ), .ZN(new_n14602_));
  AOI21_X1   g14345(.A1(new_n14602_), .A2(new_n14601_), .B(new_n8321_), .ZN(new_n14603_));
  NAND2_X1   g14346(.A1(new_n1225_), .A2(new_n14603_), .ZN(new_n14604_));
  XOR2_X1    g14347(.A1(new_n14604_), .A2(\a[62] ), .Z(new_n14605_));
  NAND2_X1   g14348(.A1(new_n14323_), .A2(new_n13758_), .ZN(new_n14606_));
  NAND2_X1   g14349(.A1(new_n14606_), .A2(new_n14322_), .ZN(new_n14607_));
  NOR3_X1    g14350(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n904_), .ZN(new_n14608_));
  NOR2_X1    g14351(.A1(new_n9364_), .A2(new_n904_), .ZN(new_n14609_));
  NOR3_X1    g14352(.A1(new_n14609_), .A2(new_n992_), .A3(new_n8985_), .ZN(new_n14610_));
  NOR2_X1    g14353(.A1(new_n14610_), .A2(new_n14608_), .ZN(new_n14611_));
  INV_X1     g14354(.I(new_n14611_), .ZN(new_n14612_));
  XOR2_X1    g14355(.A1(new_n14607_), .A2(new_n14612_), .Z(new_n14613_));
  NOR2_X1    g14356(.A1(new_n14607_), .A2(new_n14611_), .ZN(new_n14614_));
  NAND2_X1   g14357(.A1(new_n14607_), .A2(new_n14611_), .ZN(new_n14615_));
  INV_X1     g14358(.I(new_n14615_), .ZN(new_n14616_));
  OAI21_X1   g14359(.A1(new_n14614_), .A2(new_n14616_), .B(new_n14605_), .ZN(new_n14617_));
  OAI21_X1   g14360(.A1(new_n14605_), .A2(new_n14613_), .B(new_n14617_), .ZN(new_n14618_));
  NAND2_X1   g14361(.A1(new_n14618_), .A2(new_n14600_), .ZN(new_n14619_));
  NOR2_X1    g14362(.A1(new_n14618_), .A2(new_n14600_), .ZN(new_n14620_));
  INV_X1     g14363(.I(new_n14620_), .ZN(new_n14621_));
  AOI21_X1   g14364(.A1(new_n14621_), .A2(new_n14619_), .B(new_n14598_), .ZN(new_n14622_));
  INV_X1     g14365(.I(new_n14598_), .ZN(new_n14623_));
  XNOR2_X1   g14366(.A1(new_n14618_), .A2(new_n14600_), .ZN(new_n14624_));
  NOR2_X1    g14367(.A1(new_n14624_), .A2(new_n14623_), .ZN(new_n14625_));
  NOR2_X1    g14368(.A1(new_n14625_), .A2(new_n14622_), .ZN(new_n14626_));
  NOR2_X1    g14369(.A1(new_n14343_), .A2(new_n14341_), .ZN(new_n14627_));
  NOR2_X1    g14370(.A1(new_n14627_), .A2(new_n14342_), .ZN(new_n14628_));
  OAI22_X1   g14371(.A1(new_n6721_), .A2(new_n1709_), .B1(new_n6723_), .B2(new_n1825_), .ZN(new_n14629_));
  NAND2_X1   g14372(.A1(new_n7617_), .A2(\b[23] ), .ZN(new_n14630_));
  AOI21_X1   g14373(.A1(new_n14630_), .A2(new_n14629_), .B(new_n6731_), .ZN(new_n14631_));
  NAND2_X1   g14374(.A1(new_n1828_), .A2(new_n14631_), .ZN(new_n14632_));
  XOR2_X1    g14375(.A1(new_n14632_), .A2(\a[56] ), .Z(new_n14633_));
  NOR2_X1    g14376(.A1(new_n14628_), .A2(new_n14633_), .ZN(new_n14634_));
  INV_X1     g14377(.I(new_n14634_), .ZN(new_n14635_));
  NAND2_X1   g14378(.A1(new_n14628_), .A2(new_n14633_), .ZN(new_n14636_));
  AOI21_X1   g14379(.A1(new_n14635_), .A2(new_n14636_), .B(new_n14626_), .ZN(new_n14637_));
  XNOR2_X1   g14380(.A1(new_n14628_), .A2(new_n14633_), .ZN(new_n14638_));
  NOR3_X1    g14381(.A1(new_n14638_), .A2(new_n14622_), .A3(new_n14625_), .ZN(new_n14639_));
  NOR2_X1    g14382(.A1(new_n14639_), .A2(new_n14637_), .ZN(new_n14640_));
  XOR2_X1    g14383(.A1(new_n14640_), .A2(new_n14593_), .Z(new_n14641_));
  INV_X1     g14384(.I(new_n14593_), .ZN(new_n14642_));
  NOR2_X1    g14385(.A1(new_n14640_), .A2(new_n14642_), .ZN(new_n14643_));
  NOR3_X1    g14386(.A1(new_n14639_), .A2(new_n14593_), .A3(new_n14637_), .ZN(new_n14644_));
  OAI21_X1   g14387(.A1(new_n14643_), .A2(new_n14644_), .B(new_n14590_), .ZN(new_n14645_));
  OAI21_X1   g14388(.A1(new_n14641_), .A2(new_n14590_), .B(new_n14645_), .ZN(new_n14646_));
  NOR2_X1    g14389(.A1(new_n14365_), .A2(new_n14304_), .ZN(new_n14647_));
  NOR2_X1    g14390(.A1(new_n14647_), .A2(new_n14364_), .ZN(new_n14648_));
  OAI22_X1   g14391(.A1(new_n5228_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n5225_), .ZN(new_n14649_));
  NAND2_X1   g14392(.A1(new_n5387_), .A2(\b[29] ), .ZN(new_n14650_));
  AOI21_X1   g14393(.A1(new_n14649_), .A2(new_n14650_), .B(new_n5231_), .ZN(new_n14651_));
  NAND2_X1   g14394(.A1(new_n2546_), .A2(new_n14651_), .ZN(new_n14652_));
  XOR2_X1    g14395(.A1(new_n14652_), .A2(\a[50] ), .Z(new_n14653_));
  XOR2_X1    g14396(.A1(new_n14648_), .A2(new_n14653_), .Z(new_n14654_));
  AND2_X2    g14397(.A1(new_n14654_), .A2(new_n14646_), .Z(new_n14655_));
  NOR2_X1    g14398(.A1(new_n14648_), .A2(new_n14653_), .ZN(new_n14656_));
  INV_X1     g14399(.I(new_n14656_), .ZN(new_n14657_));
  NAND2_X1   g14400(.A1(new_n14648_), .A2(new_n14653_), .ZN(new_n14658_));
  AOI21_X1   g14401(.A1(new_n14657_), .A2(new_n14658_), .B(new_n14646_), .ZN(new_n14659_));
  NOR2_X1    g14402(.A1(new_n14655_), .A2(new_n14659_), .ZN(new_n14660_));
  NOR2_X1    g14403(.A1(new_n14367_), .A2(new_n14377_), .ZN(new_n14661_));
  NOR2_X1    g14404(.A1(new_n14661_), .A2(new_n14374_), .ZN(new_n14662_));
  INV_X1     g14405(.I(new_n14662_), .ZN(new_n14663_));
  XOR2_X1    g14406(.A1(new_n14660_), .A2(new_n14663_), .Z(new_n14664_));
  NOR2_X1    g14407(.A1(new_n14664_), .A2(new_n14585_), .ZN(new_n14665_));
  INV_X1     g14408(.I(new_n14585_), .ZN(new_n14666_));
  OAI21_X1   g14409(.A1(new_n14655_), .A2(new_n14659_), .B(new_n14663_), .ZN(new_n14667_));
  NAND2_X1   g14410(.A1(new_n14660_), .A2(new_n14662_), .ZN(new_n14668_));
  AOI21_X1   g14411(.A1(new_n14668_), .A2(new_n14667_), .B(new_n14666_), .ZN(new_n14669_));
  NOR2_X1    g14412(.A1(new_n14665_), .A2(new_n14669_), .ZN(new_n14670_));
  XOR2_X1    g14413(.A1(new_n14670_), .A2(new_n14580_), .Z(new_n14671_));
  NAND2_X1   g14414(.A1(new_n14671_), .A2(new_n14578_), .ZN(new_n14672_));
  OR2_X2     g14415(.A1(new_n14670_), .A2(new_n14580_), .Z(new_n14673_));
  NAND2_X1   g14416(.A1(new_n14670_), .A2(new_n14580_), .ZN(new_n14674_));
  NAND2_X1   g14417(.A1(new_n14673_), .A2(new_n14674_), .ZN(new_n14675_));
  NAND2_X1   g14418(.A1(new_n14675_), .A2(new_n14577_), .ZN(new_n14676_));
  NAND2_X1   g14419(.A1(new_n14676_), .A2(new_n14672_), .ZN(new_n14677_));
  XOR2_X1    g14420(.A1(new_n14677_), .A2(new_n14572_), .Z(new_n14678_));
  NAND2_X1   g14421(.A1(new_n14678_), .A2(new_n14570_), .ZN(new_n14679_));
  AND2_X2    g14422(.A1(new_n14677_), .A2(new_n14572_), .Z(new_n14680_));
  NOR2_X1    g14423(.A1(new_n14677_), .A2(new_n14572_), .ZN(new_n14681_));
  OAI21_X1   g14424(.A1(new_n14680_), .A2(new_n14681_), .B(new_n14569_), .ZN(new_n14682_));
  NAND2_X1   g14425(.A1(new_n14679_), .A2(new_n14682_), .ZN(new_n14683_));
  OAI22_X1   g14426(.A1(new_n3298_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n3293_), .ZN(new_n14684_));
  NAND2_X1   g14427(.A1(new_n4227_), .A2(\b[41] ), .ZN(new_n14685_));
  AOI21_X1   g14428(.A1(new_n14684_), .A2(new_n14685_), .B(new_n3301_), .ZN(new_n14686_));
  NAND2_X1   g14429(.A1(new_n4320_), .A2(new_n14686_), .ZN(new_n14687_));
  XOR2_X1    g14430(.A1(new_n14687_), .A2(\a[38] ), .Z(new_n14688_));
  NOR2_X1    g14431(.A1(new_n14683_), .A2(new_n14688_), .ZN(new_n14689_));
  INV_X1     g14432(.I(new_n14689_), .ZN(new_n14690_));
  NAND2_X1   g14433(.A1(new_n14683_), .A2(new_n14688_), .ZN(new_n14691_));
  AOI21_X1   g14434(.A1(new_n14690_), .A2(new_n14691_), .B(new_n14564_), .ZN(new_n14692_));
  INV_X1     g14435(.I(new_n14564_), .ZN(new_n14693_));
  INV_X1     g14436(.I(new_n14688_), .ZN(new_n14694_));
  XOR2_X1    g14437(.A1(new_n14683_), .A2(new_n14694_), .Z(new_n14695_));
  NOR2_X1    g14438(.A1(new_n14695_), .A2(new_n14693_), .ZN(new_n14696_));
  NOR2_X1    g14439(.A1(new_n14696_), .A2(new_n14692_), .ZN(new_n14697_));
  NAND2_X1   g14440(.A1(new_n14427_), .A2(new_n14424_), .ZN(new_n14698_));
  AOI21_X1   g14441(.A1(new_n14426_), .A2(new_n14698_), .B(new_n14697_), .ZN(new_n14699_));
  NAND2_X1   g14442(.A1(new_n14698_), .A2(new_n14426_), .ZN(new_n14700_));
  NOR3_X1    g14443(.A1(new_n14696_), .A2(new_n14692_), .A3(new_n14700_), .ZN(new_n14701_));
  OAI21_X1   g14444(.A1(new_n14699_), .A2(new_n14701_), .B(new_n14562_), .ZN(new_n14702_));
  XOR2_X1    g14445(.A1(new_n14697_), .A2(new_n14700_), .Z(new_n14703_));
  OAI21_X1   g14446(.A1(new_n14562_), .A2(new_n14703_), .B(new_n14702_), .ZN(new_n14704_));
  XOR2_X1    g14447(.A1(new_n14704_), .A2(new_n14556_), .Z(new_n14705_));
  NAND2_X1   g14448(.A1(new_n14704_), .A2(new_n14556_), .ZN(new_n14706_));
  OR2_X2     g14449(.A1(new_n14704_), .A2(new_n14556_), .Z(new_n14707_));
  AOI21_X1   g14450(.A1(new_n14707_), .A2(new_n14706_), .B(new_n14554_), .ZN(new_n14708_));
  AOI21_X1   g14451(.A1(new_n14554_), .A2(new_n14705_), .B(new_n14708_), .ZN(new_n14709_));
  INV_X1     g14452(.I(new_n14709_), .ZN(new_n14710_));
  NAND2_X1   g14453(.A1(new_n5954_), .A2(new_n2086_), .ZN(new_n14711_));
  AOI22_X1   g14454(.A1(\b[52] ), .A2(new_n2083_), .B1(new_n2670_), .B2(\b[51] ), .ZN(new_n14712_));
  AOI21_X1   g14455(.A1(\b[50] ), .A2(new_n2864_), .B(new_n14712_), .ZN(new_n14713_));
  NAND2_X1   g14456(.A1(new_n14711_), .A2(new_n14713_), .ZN(new_n14714_));
  NOR2_X1    g14457(.A1(new_n14451_), .A2(new_n14442_), .ZN(new_n14715_));
  NOR2_X1    g14458(.A1(new_n14715_), .A2(new_n14450_), .ZN(new_n14716_));
  XOR2_X1    g14459(.A1(new_n14716_), .A2(new_n14714_), .Z(new_n14717_));
  NAND2_X1   g14460(.A1(new_n14717_), .A2(new_n2074_), .ZN(new_n14718_));
  NOR2_X1    g14461(.A1(new_n14717_), .A2(new_n2074_), .ZN(new_n14719_));
  INV_X1     g14462(.I(new_n14719_), .ZN(new_n14720_));
  AOI21_X1   g14463(.A1(new_n14720_), .A2(new_n14718_), .B(new_n14710_), .ZN(new_n14721_));
  INV_X1     g14464(.I(new_n14718_), .ZN(new_n14722_));
  NOR3_X1    g14465(.A1(new_n14722_), .A2(new_n14719_), .A3(new_n14709_), .ZN(new_n14723_));
  OAI21_X1   g14466(.A1(new_n14721_), .A2(new_n14723_), .B(new_n14548_), .ZN(new_n14724_));
  OAI21_X1   g14467(.A1(new_n14722_), .A2(new_n14719_), .B(new_n14709_), .ZN(new_n14725_));
  NAND3_X1   g14468(.A1(new_n14710_), .A2(new_n14720_), .A3(new_n14718_), .ZN(new_n14726_));
  NAND3_X1   g14469(.A1(new_n14726_), .A2(new_n14725_), .A3(new_n14547_), .ZN(new_n14727_));
  AOI21_X1   g14470(.A1(new_n14724_), .A2(new_n14727_), .B(new_n14546_), .ZN(new_n14728_));
  INV_X1     g14471(.I(new_n14546_), .ZN(new_n14729_));
  OAI21_X1   g14472(.A1(new_n14721_), .A2(new_n14723_), .B(new_n14547_), .ZN(new_n14730_));
  NAND3_X1   g14473(.A1(new_n14726_), .A2(new_n14725_), .A3(new_n14548_), .ZN(new_n14731_));
  AOI21_X1   g14474(.A1(new_n14730_), .A2(new_n14731_), .B(new_n14729_), .ZN(new_n14732_));
  NOR2_X1    g14475(.A1(new_n14728_), .A2(new_n14732_), .ZN(new_n14733_));
  NOR2_X1    g14476(.A1(new_n14470_), .A2(new_n14272_), .ZN(new_n14734_));
  NOR2_X1    g14477(.A1(new_n14734_), .A2(new_n14469_), .ZN(new_n14735_));
  OAI22_X1   g14478(.A1(new_n1444_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n1439_), .ZN(new_n14736_));
  OAI21_X1   g14479(.A1(new_n6995_), .A2(new_n1548_), .B(new_n14736_), .ZN(new_n14737_));
  AOI21_X1   g14480(.A1(new_n7559_), .A2(new_n1446_), .B(new_n14737_), .ZN(new_n14738_));
  INV_X1     g14481(.I(new_n14738_), .ZN(new_n14739_));
  NAND2_X1   g14482(.A1(new_n14735_), .A2(new_n14739_), .ZN(new_n14740_));
  INV_X1     g14483(.I(new_n14735_), .ZN(new_n14741_));
  NAND2_X1   g14484(.A1(new_n14741_), .A2(new_n14738_), .ZN(new_n14742_));
  AOI21_X1   g14485(.A1(new_n14742_), .A2(new_n14740_), .B(\a[23] ), .ZN(new_n14743_));
  NAND3_X1   g14486(.A1(new_n14742_), .A2(new_n14740_), .A3(\a[23] ), .ZN(new_n14744_));
  INV_X1     g14487(.I(new_n14744_), .ZN(new_n14745_));
  OAI21_X1   g14488(.A1(new_n14745_), .A2(new_n14743_), .B(new_n14733_), .ZN(new_n14746_));
  OR2_X2     g14489(.A1(new_n14728_), .A2(new_n14732_), .Z(new_n14747_));
  INV_X1     g14490(.I(new_n14743_), .ZN(new_n14748_));
  NAND3_X1   g14491(.A1(new_n14748_), .A2(new_n14747_), .A3(new_n14744_), .ZN(new_n14749_));
  OAI22_X1   g14492(.A1(new_n1168_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n1163_), .ZN(new_n14750_));
  NAND2_X1   g14493(.A1(new_n1774_), .A2(\b[59] ), .ZN(new_n14751_));
  AOI21_X1   g14494(.A1(new_n14750_), .A2(new_n14751_), .B(new_n1171_), .ZN(new_n14752_));
  NAND2_X1   g14495(.A1(new_n8550_), .A2(new_n14752_), .ZN(new_n14753_));
  XOR2_X1    g14496(.A1(new_n14753_), .A2(\a[20] ), .Z(new_n14754_));
  INV_X1     g14497(.I(new_n14754_), .ZN(new_n14755_));
  NAND3_X1   g14498(.A1(new_n14749_), .A2(new_n14746_), .A3(new_n14755_), .ZN(new_n14756_));
  AOI21_X1   g14499(.A1(new_n14748_), .A2(new_n14744_), .B(new_n14747_), .ZN(new_n14757_));
  NOR3_X1    g14500(.A1(new_n14745_), .A2(new_n14743_), .A3(new_n14733_), .ZN(new_n14758_));
  OAI21_X1   g14501(.A1(new_n14757_), .A2(new_n14758_), .B(new_n14754_), .ZN(new_n14759_));
  AOI21_X1   g14502(.A1(new_n14759_), .A2(new_n14756_), .B(new_n14541_), .ZN(new_n14760_));
  INV_X1     g14503(.I(new_n14541_), .ZN(new_n14761_));
  OAI21_X1   g14504(.A1(new_n14757_), .A2(new_n14758_), .B(new_n14755_), .ZN(new_n14762_));
  NAND3_X1   g14505(.A1(new_n14749_), .A2(new_n14746_), .A3(new_n14754_), .ZN(new_n14763_));
  AOI21_X1   g14506(.A1(new_n14762_), .A2(new_n14763_), .B(new_n14761_), .ZN(new_n14764_));
  NOR2_X1    g14507(.A1(new_n1020_), .A2(new_n8932_), .ZN(new_n14765_));
  NOR2_X1    g14508(.A1(new_n935_), .A2(new_n8956_), .ZN(new_n14766_));
  NOR4_X1    g14509(.A1(new_n9323_), .A2(new_n943_), .A3(new_n14765_), .A4(new_n14766_), .ZN(new_n14767_));
  XOR2_X1    g14510(.A1(new_n14767_), .A2(new_n930_), .Z(new_n14768_));
  NOR3_X1    g14511(.A1(new_n14760_), .A2(new_n14764_), .A3(new_n14768_), .ZN(new_n14769_));
  OAI21_X1   g14512(.A1(new_n14760_), .A2(new_n14764_), .B(new_n14768_), .ZN(new_n14770_));
  INV_X1     g14513(.I(new_n14770_), .ZN(new_n14771_));
  OAI21_X1   g14514(.A1(new_n14771_), .A2(new_n14769_), .B(new_n14540_), .ZN(new_n14772_));
  INV_X1     g14515(.I(new_n14768_), .ZN(new_n14773_));
  OAI21_X1   g14516(.A1(new_n14760_), .A2(new_n14764_), .B(new_n14773_), .ZN(new_n14774_));
  INV_X1     g14517(.I(new_n14774_), .ZN(new_n14775_));
  NOR3_X1    g14518(.A1(new_n14760_), .A2(new_n14764_), .A3(new_n14773_), .ZN(new_n14776_));
  OAI21_X1   g14519(.A1(new_n14775_), .A2(new_n14776_), .B(new_n14539_), .ZN(new_n14777_));
  NAND2_X1   g14520(.A1(new_n14772_), .A2(new_n14777_), .ZN(new_n14778_));
  XOR2_X1    g14521(.A1(new_n14524_), .A2(new_n14257_), .Z(new_n14779_));
  NAND3_X1   g14522(.A1(new_n14779_), .A2(new_n13981_), .A3(new_n14528_), .ZN(new_n14780_));
  NOR3_X1    g14523(.A1(new_n14257_), .A2(new_n14519_), .A3(new_n14523_), .ZN(new_n14781_));
  AOI21_X1   g14524(.A1(new_n14531_), .A2(new_n14780_), .B(new_n14781_), .ZN(new_n14782_));
  XOR2_X1    g14525(.A1(new_n14782_), .A2(new_n14778_), .Z(new_n14783_));
  XOR2_X1    g14526(.A1(new_n14783_), .A2(new_n14538_), .Z(\f[79] ));
  NAND2_X1   g14527(.A1(new_n14531_), .A2(new_n14780_), .ZN(new_n14785_));
  NOR2_X1    g14528(.A1(new_n14778_), .A2(new_n14538_), .ZN(new_n14786_));
  INV_X1     g14529(.I(new_n14769_), .ZN(new_n14787_));
  AOI21_X1   g14530(.A1(new_n14787_), .A2(new_n14770_), .B(new_n14539_), .ZN(new_n14788_));
  INV_X1     g14531(.I(new_n14776_), .ZN(new_n14789_));
  AOI21_X1   g14532(.A1(new_n14789_), .A2(new_n14774_), .B(new_n14540_), .ZN(new_n14790_));
  OAI21_X1   g14533(.A1(new_n14788_), .A2(new_n14790_), .B(new_n14538_), .ZN(new_n14791_));
  NAND3_X1   g14534(.A1(new_n14772_), .A2(new_n14777_), .A3(new_n14537_), .ZN(new_n14792_));
  AOI21_X1   g14535(.A1(new_n14791_), .A2(new_n14792_), .B(new_n14781_), .ZN(new_n14793_));
  AOI21_X1   g14536(.A1(new_n14785_), .A2(new_n14793_), .B(new_n14786_), .ZN(new_n14794_));
  AOI21_X1   g14537(.A1(new_n14540_), .A2(new_n14770_), .B(new_n14769_), .ZN(new_n14795_));
  INV_X1     g14538(.I(new_n14795_), .ZN(new_n14796_));
  OAI22_X1   g14539(.A1(new_n1444_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n1439_), .ZN(new_n14797_));
  NAND2_X1   g14540(.A1(new_n2098_), .A2(\b[57] ), .ZN(new_n14798_));
  AOI21_X1   g14541(.A1(new_n14797_), .A2(new_n14798_), .B(new_n1447_), .ZN(new_n14799_));
  NAND2_X1   g14542(.A1(new_n7895_), .A2(new_n14799_), .ZN(new_n14800_));
  XOR2_X1    g14543(.A1(new_n14800_), .A2(\a[23] ), .Z(new_n14801_));
  INV_X1     g14544(.I(new_n14801_), .ZN(new_n14802_));
  OAI22_X1   g14545(.A1(new_n2084_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n2079_), .ZN(new_n14803_));
  NAND2_X1   g14546(.A1(new_n2864_), .A2(\b[51] ), .ZN(new_n14804_));
  AOI21_X1   g14547(.A1(new_n14803_), .A2(new_n14804_), .B(new_n2087_), .ZN(new_n14805_));
  NAND2_X1   g14548(.A1(new_n6219_), .A2(new_n14805_), .ZN(new_n14806_));
  XOR2_X1    g14549(.A1(new_n14806_), .A2(\a[29] ), .Z(new_n14807_));
  OAI22_X1   g14550(.A1(new_n2452_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n2447_), .ZN(new_n14808_));
  NAND2_X1   g14551(.A1(new_n3312_), .A2(\b[48] ), .ZN(new_n14809_));
  AOI21_X1   g14552(.A1(new_n14808_), .A2(new_n14809_), .B(new_n2455_), .ZN(new_n14810_));
  NAND2_X1   g14553(.A1(new_n5537_), .A2(new_n14810_), .ZN(new_n14811_));
  XOR2_X1    g14554(.A1(new_n14811_), .A2(\a[32] ), .Z(new_n14812_));
  NOR2_X1    g14555(.A1(new_n14701_), .A2(new_n14561_), .ZN(new_n14813_));
  NOR2_X1    g14556(.A1(new_n14699_), .A2(new_n14813_), .ZN(new_n14814_));
  INV_X1     g14557(.I(new_n14814_), .ZN(new_n14815_));
  OAI22_X1   g14558(.A1(new_n3298_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n3293_), .ZN(new_n14816_));
  NAND2_X1   g14559(.A1(new_n4227_), .A2(\b[42] ), .ZN(new_n14817_));
  AOI21_X1   g14560(.A1(new_n14816_), .A2(new_n14817_), .B(new_n3301_), .ZN(new_n14818_));
  NAND2_X1   g14561(.A1(new_n4500_), .A2(new_n14818_), .ZN(new_n14819_));
  XOR2_X1    g14562(.A1(new_n14819_), .A2(\a[38] ), .Z(new_n14820_));
  INV_X1     g14563(.I(new_n14681_), .ZN(new_n14821_));
  OAI21_X1   g14564(.A1(new_n14569_), .A2(new_n14680_), .B(new_n14821_), .ZN(new_n14822_));
  OAI22_X1   g14565(.A1(new_n3736_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n3731_), .ZN(new_n14823_));
  NAND2_X1   g14566(.A1(new_n4730_), .A2(\b[39] ), .ZN(new_n14824_));
  AOI21_X1   g14567(.A1(new_n14823_), .A2(new_n14824_), .B(new_n3739_), .ZN(new_n14825_));
  NAND2_X1   g14568(.A1(new_n3996_), .A2(new_n14825_), .ZN(new_n14826_));
  XOR2_X1    g14569(.A1(new_n14826_), .A2(\a[41] ), .Z(new_n14827_));
  OAI22_X1   g14570(.A1(new_n4208_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n4203_), .ZN(new_n14828_));
  NAND2_X1   g14571(.A1(new_n5244_), .A2(\b[36] ), .ZN(new_n14829_));
  AOI21_X1   g14572(.A1(new_n14828_), .A2(new_n14829_), .B(new_n4211_), .ZN(new_n14830_));
  NAND2_X1   g14573(.A1(new_n3565_), .A2(new_n14830_), .ZN(new_n14831_));
  XOR2_X1    g14574(.A1(new_n14831_), .A2(\a[44] ), .Z(new_n14832_));
  INV_X1     g14575(.I(new_n14832_), .ZN(new_n14833_));
  OAI22_X1   g14576(.A1(new_n5228_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n5225_), .ZN(new_n14834_));
  NAND2_X1   g14577(.A1(new_n5387_), .A2(\b[30] ), .ZN(new_n14835_));
  AOI21_X1   g14578(.A1(new_n14834_), .A2(new_n14835_), .B(new_n5231_), .ZN(new_n14836_));
  NAND2_X1   g14579(.A1(new_n2659_), .A2(new_n14836_), .ZN(new_n14837_));
  XOR2_X1    g14580(.A1(new_n14837_), .A2(\a[50] ), .Z(new_n14838_));
  OAI22_X1   g14581(.A1(new_n6721_), .A2(new_n1825_), .B1(new_n6723_), .B2(new_n1927_), .ZN(new_n14839_));
  NAND2_X1   g14582(.A1(new_n7617_), .A2(\b[24] ), .ZN(new_n14840_));
  AOI21_X1   g14583(.A1(new_n14840_), .A2(new_n14839_), .B(new_n6731_), .ZN(new_n14841_));
  NAND2_X1   g14584(.A1(new_n1926_), .A2(new_n14841_), .ZN(new_n14842_));
  XOR2_X1    g14585(.A1(new_n14842_), .A2(\a[56] ), .Z(new_n14843_));
  AOI21_X1   g14586(.A1(new_n14623_), .A2(new_n14619_), .B(new_n14620_), .ZN(new_n14844_));
  OAI22_X1   g14587(.A1(new_n1305_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1222_), .ZN(new_n14845_));
  NAND2_X1   g14588(.A1(new_n9644_), .A2(\b[18] ), .ZN(new_n14846_));
  AOI21_X1   g14589(.A1(new_n14846_), .A2(new_n14845_), .B(new_n8321_), .ZN(new_n14847_));
  NAND2_X1   g14590(.A1(new_n1304_), .A2(new_n14847_), .ZN(new_n14848_));
  XOR2_X1    g14591(.A1(new_n14848_), .A2(\a[62] ), .Z(new_n14849_));
  NOR3_X1    g14592(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n992_), .ZN(new_n14850_));
  NOR2_X1    g14593(.A1(new_n9364_), .A2(new_n992_), .ZN(new_n14851_));
  NOR3_X1    g14594(.A1(new_n14851_), .A2(new_n1044_), .A3(new_n8985_), .ZN(new_n14852_));
  NOR2_X1    g14595(.A1(new_n14852_), .A2(new_n14850_), .ZN(new_n14853_));
  NOR2_X1    g14596(.A1(new_n14612_), .A2(new_n14853_), .ZN(new_n14854_));
  INV_X1     g14597(.I(new_n14853_), .ZN(new_n14855_));
  NOR2_X1    g14598(.A1(new_n14855_), .A2(new_n14611_), .ZN(new_n14856_));
  NOR2_X1    g14599(.A1(new_n14854_), .A2(new_n14856_), .ZN(new_n14857_));
  NOR2_X1    g14600(.A1(new_n14849_), .A2(new_n14857_), .ZN(new_n14858_));
  XOR2_X1    g14601(.A1(new_n14611_), .A2(new_n14853_), .Z(new_n14859_));
  INV_X1     g14602(.I(new_n14859_), .ZN(new_n14860_));
  AOI21_X1   g14603(.A1(new_n14849_), .A2(new_n14860_), .B(new_n14858_), .ZN(new_n14861_));
  OAI22_X1   g14604(.A1(new_n1601_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1518_), .ZN(new_n14862_));
  NAND2_X1   g14605(.A1(new_n8628_), .A2(\b[21] ), .ZN(new_n14863_));
  AOI21_X1   g14606(.A1(new_n14863_), .A2(new_n14862_), .B(new_n7354_), .ZN(new_n14864_));
  NAND2_X1   g14607(.A1(new_n1604_), .A2(new_n14864_), .ZN(new_n14865_));
  XOR2_X1    g14608(.A1(new_n14865_), .A2(\a[59] ), .Z(new_n14866_));
  OAI21_X1   g14609(.A1(new_n14605_), .A2(new_n14614_), .B(new_n14615_), .ZN(new_n14867_));
  XOR2_X1    g14610(.A1(new_n14866_), .A2(new_n14867_), .Z(new_n14868_));
  NOR2_X1    g14611(.A1(new_n14868_), .A2(new_n14861_), .ZN(new_n14869_));
  INV_X1     g14612(.I(new_n14861_), .ZN(new_n14870_));
  INV_X1     g14613(.I(new_n14867_), .ZN(new_n14871_));
  OR2_X2     g14614(.A1(new_n14866_), .A2(new_n14871_), .Z(new_n14872_));
  NAND2_X1   g14615(.A1(new_n14866_), .A2(new_n14871_), .ZN(new_n14873_));
  AOI21_X1   g14616(.A1(new_n14872_), .A2(new_n14873_), .B(new_n14870_), .ZN(new_n14874_));
  NOR2_X1    g14617(.A1(new_n14869_), .A2(new_n14874_), .ZN(new_n14875_));
  XOR2_X1    g14618(.A1(new_n14875_), .A2(new_n14844_), .Z(new_n14876_));
  NOR2_X1    g14619(.A1(new_n14876_), .A2(new_n14843_), .ZN(new_n14877_));
  INV_X1     g14620(.I(new_n14843_), .ZN(new_n14878_));
  OAI21_X1   g14621(.A1(new_n14869_), .A2(new_n14874_), .B(new_n14844_), .ZN(new_n14879_));
  INV_X1     g14622(.I(new_n14844_), .ZN(new_n14880_));
  NAND2_X1   g14623(.A1(new_n14875_), .A2(new_n14880_), .ZN(new_n14881_));
  AOI21_X1   g14624(.A1(new_n14881_), .A2(new_n14879_), .B(new_n14878_), .ZN(new_n14882_));
  NOR2_X1    g14625(.A1(new_n14877_), .A2(new_n14882_), .ZN(new_n14883_));
  INV_X1     g14626(.I(new_n14883_), .ZN(new_n14884_));
  OAI22_X1   g14627(.A1(new_n5786_), .A2(new_n2272_), .B1(new_n2175_), .B2(new_n5792_), .ZN(new_n14885_));
  NAND2_X1   g14628(.A1(new_n6745_), .A2(\b[27] ), .ZN(new_n14886_));
  AOI21_X1   g14629(.A1(new_n14886_), .A2(new_n14885_), .B(new_n5796_), .ZN(new_n14887_));
  NAND2_X1   g14630(.A1(new_n2276_), .A2(new_n14887_), .ZN(new_n14888_));
  XOR2_X1    g14631(.A1(new_n14888_), .A2(\a[53] ), .Z(new_n14889_));
  AOI21_X1   g14632(.A1(new_n14628_), .A2(new_n14633_), .B(new_n14626_), .ZN(new_n14890_));
  NOR2_X1    g14633(.A1(new_n14890_), .A2(new_n14634_), .ZN(new_n14891_));
  XOR2_X1    g14634(.A1(new_n14891_), .A2(new_n14889_), .Z(new_n14892_));
  NAND2_X1   g14635(.A1(new_n14884_), .A2(new_n14892_), .ZN(new_n14893_));
  INV_X1     g14636(.I(new_n14889_), .ZN(new_n14894_));
  INV_X1     g14637(.I(new_n14891_), .ZN(new_n14895_));
  NAND2_X1   g14638(.A1(new_n14895_), .A2(new_n14894_), .ZN(new_n14896_));
  INV_X1     g14639(.I(new_n14896_), .ZN(new_n14897_));
  NAND2_X1   g14640(.A1(new_n14891_), .A2(new_n14889_), .ZN(new_n14898_));
  INV_X1     g14641(.I(new_n14898_), .ZN(new_n14899_));
  OAI21_X1   g14642(.A1(new_n14897_), .A2(new_n14899_), .B(new_n14883_), .ZN(new_n14900_));
  NAND2_X1   g14643(.A1(new_n14893_), .A2(new_n14900_), .ZN(new_n14901_));
  INV_X1     g14644(.I(new_n14901_), .ZN(new_n14902_));
  NOR2_X1    g14645(.A1(new_n14644_), .A2(new_n14590_), .ZN(new_n14903_));
  NOR2_X1    g14646(.A1(new_n14903_), .A2(new_n14643_), .ZN(new_n14904_));
  NOR2_X1    g14647(.A1(new_n14902_), .A2(new_n14904_), .ZN(new_n14905_));
  INV_X1     g14648(.I(new_n14905_), .ZN(new_n14906_));
  NAND2_X1   g14649(.A1(new_n14902_), .A2(new_n14904_), .ZN(new_n14907_));
  AOI21_X1   g14650(.A1(new_n14906_), .A2(new_n14907_), .B(new_n14838_), .ZN(new_n14908_));
  INV_X1     g14651(.I(new_n14838_), .ZN(new_n14909_));
  XOR2_X1    g14652(.A1(new_n14901_), .A2(new_n14904_), .Z(new_n14910_));
  NOR2_X1    g14653(.A1(new_n14910_), .A2(new_n14909_), .ZN(new_n14911_));
  NOR2_X1    g14654(.A1(new_n14908_), .A2(new_n14911_), .ZN(new_n14912_));
  INV_X1     g14655(.I(new_n14912_), .ZN(new_n14913_));
  OAI22_X1   g14656(.A1(new_n4711_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n4706_), .ZN(new_n14914_));
  NAND2_X1   g14657(.A1(new_n5814_), .A2(\b[33] ), .ZN(new_n14915_));
  AOI21_X1   g14658(.A1(new_n14914_), .A2(new_n14915_), .B(new_n4714_), .ZN(new_n14916_));
  NAND2_X1   g14659(.A1(new_n3101_), .A2(new_n14916_), .ZN(new_n14917_));
  XOR2_X1    g14660(.A1(new_n14917_), .A2(\a[47] ), .Z(new_n14918_));
  AOI21_X1   g14661(.A1(new_n14648_), .A2(new_n14653_), .B(new_n14646_), .ZN(new_n14919_));
  NOR2_X1    g14662(.A1(new_n14919_), .A2(new_n14656_), .ZN(new_n14920_));
  NOR2_X1    g14663(.A1(new_n14920_), .A2(new_n14918_), .ZN(new_n14921_));
  NAND2_X1   g14664(.A1(new_n14920_), .A2(new_n14918_), .ZN(new_n14922_));
  INV_X1     g14665(.I(new_n14922_), .ZN(new_n14923_));
  OAI21_X1   g14666(.A1(new_n14923_), .A2(new_n14921_), .B(new_n14913_), .ZN(new_n14924_));
  XOR2_X1    g14667(.A1(new_n14920_), .A2(new_n14918_), .Z(new_n14925_));
  NAND2_X1   g14668(.A1(new_n14925_), .A2(new_n14912_), .ZN(new_n14926_));
  NAND2_X1   g14669(.A1(new_n14668_), .A2(new_n14666_), .ZN(new_n14927_));
  AOI22_X1   g14670(.A1(new_n14927_), .A2(new_n14667_), .B1(new_n14926_), .B2(new_n14924_), .ZN(new_n14928_));
  NAND2_X1   g14671(.A1(new_n14926_), .A2(new_n14924_), .ZN(new_n14929_));
  NAND2_X1   g14672(.A1(new_n14927_), .A2(new_n14667_), .ZN(new_n14930_));
  NOR2_X1    g14673(.A1(new_n14930_), .A2(new_n14929_), .ZN(new_n14931_));
  OAI21_X1   g14674(.A1(new_n14931_), .A2(new_n14928_), .B(new_n14833_), .ZN(new_n14932_));
  XNOR2_X1   g14675(.A1(new_n14930_), .A2(new_n14929_), .ZN(new_n14933_));
  OAI21_X1   g14676(.A1(new_n14933_), .A2(new_n14833_), .B(new_n14932_), .ZN(new_n14934_));
  NAND2_X1   g14677(.A1(new_n14673_), .A2(new_n14578_), .ZN(new_n14935_));
  NAND2_X1   g14678(.A1(new_n14935_), .A2(new_n14674_), .ZN(new_n14936_));
  XNOR2_X1   g14679(.A1(new_n14936_), .A2(new_n14934_), .ZN(new_n14937_));
  NOR2_X1    g14680(.A1(new_n14937_), .A2(new_n14827_), .ZN(new_n14938_));
  INV_X1     g14681(.I(new_n14827_), .ZN(new_n14939_));
  NAND2_X1   g14682(.A1(new_n14936_), .A2(new_n14934_), .ZN(new_n14940_));
  OR2_X2     g14683(.A1(new_n14936_), .A2(new_n14934_), .Z(new_n14941_));
  AOI21_X1   g14684(.A1(new_n14941_), .A2(new_n14940_), .B(new_n14939_), .ZN(new_n14942_));
  NOR2_X1    g14685(.A1(new_n14938_), .A2(new_n14942_), .ZN(new_n14943_));
  XNOR2_X1   g14686(.A1(new_n14943_), .A2(new_n14822_), .ZN(new_n14944_));
  NOR2_X1    g14687(.A1(new_n14944_), .A2(new_n14820_), .ZN(new_n14945_));
  INV_X1     g14688(.I(new_n14822_), .ZN(new_n14946_));
  OR2_X2     g14689(.A1(new_n14938_), .A2(new_n14942_), .Z(new_n14947_));
  NAND2_X1   g14690(.A1(new_n14947_), .A2(new_n14946_), .ZN(new_n14948_));
  NAND2_X1   g14691(.A1(new_n14943_), .A2(new_n14822_), .ZN(new_n14949_));
  NAND2_X1   g14692(.A1(new_n14948_), .A2(new_n14949_), .ZN(new_n14950_));
  AOI21_X1   g14693(.A1(new_n14820_), .A2(new_n14950_), .B(new_n14945_), .ZN(new_n14951_));
  OAI22_X1   g14694(.A1(new_n2846_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n2841_), .ZN(new_n14952_));
  NAND2_X1   g14695(.A1(new_n3755_), .A2(\b[45] ), .ZN(new_n14953_));
  AOI21_X1   g14696(.A1(new_n14952_), .A2(new_n14953_), .B(new_n2849_), .ZN(new_n14954_));
  NAND2_X1   g14697(.A1(new_n5004_), .A2(new_n14954_), .ZN(new_n14955_));
  XOR2_X1    g14698(.A1(new_n14955_), .A2(\a[35] ), .Z(new_n14956_));
  AOI21_X1   g14699(.A1(new_n14693_), .A2(new_n14691_), .B(new_n14689_), .ZN(new_n14957_));
  XNOR2_X1   g14700(.A1(new_n14957_), .A2(new_n14956_), .ZN(new_n14958_));
  NOR2_X1    g14701(.A1(new_n14958_), .A2(new_n14951_), .ZN(new_n14959_));
  NOR2_X1    g14702(.A1(new_n14957_), .A2(new_n14956_), .ZN(new_n14960_));
  INV_X1     g14703(.I(new_n14960_), .ZN(new_n14961_));
  NAND2_X1   g14704(.A1(new_n14957_), .A2(new_n14956_), .ZN(new_n14962_));
  NAND2_X1   g14705(.A1(new_n14961_), .A2(new_n14962_), .ZN(new_n14963_));
  AND2_X2    g14706(.A1(new_n14963_), .A2(new_n14951_), .Z(new_n14964_));
  NOR2_X1    g14707(.A1(new_n14964_), .A2(new_n14959_), .ZN(new_n14965_));
  XOR2_X1    g14708(.A1(new_n14965_), .A2(new_n14815_), .Z(new_n14966_));
  NOR2_X1    g14709(.A1(new_n14966_), .A2(new_n14812_), .ZN(new_n14967_));
  INV_X1     g14710(.I(new_n14812_), .ZN(new_n14968_));
  OAI21_X1   g14711(.A1(new_n14959_), .A2(new_n14964_), .B(new_n14815_), .ZN(new_n14969_));
  NAND2_X1   g14712(.A1(new_n14965_), .A2(new_n14814_), .ZN(new_n14970_));
  AOI21_X1   g14713(.A1(new_n14969_), .A2(new_n14970_), .B(new_n14968_), .ZN(new_n14971_));
  NOR2_X1    g14714(.A1(new_n14967_), .A2(new_n14971_), .ZN(new_n14972_));
  NAND2_X1   g14715(.A1(new_n14707_), .A2(new_n14554_), .ZN(new_n14973_));
  NAND2_X1   g14716(.A1(new_n14973_), .A2(new_n14706_), .ZN(new_n14974_));
  NAND2_X1   g14717(.A1(new_n14972_), .A2(new_n14974_), .ZN(new_n14975_));
  OR2_X2     g14718(.A1(new_n14972_), .A2(new_n14974_), .Z(new_n14976_));
  AOI21_X1   g14719(.A1(new_n14976_), .A2(new_n14975_), .B(new_n14807_), .ZN(new_n14977_));
  INV_X1     g14720(.I(new_n14807_), .ZN(new_n14978_));
  XNOR2_X1   g14721(.A1(new_n14972_), .A2(new_n14974_), .ZN(new_n14979_));
  NOR2_X1    g14722(.A1(new_n14979_), .A2(new_n14978_), .ZN(new_n14980_));
  NOR2_X1    g14723(.A1(new_n14980_), .A2(new_n14977_), .ZN(new_n14981_));
  INV_X1     g14724(.I(new_n14981_), .ZN(new_n14982_));
  OAI22_X1   g14725(.A1(new_n1760_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n1755_), .ZN(new_n14983_));
  OAI21_X1   g14726(.A1(new_n6238_), .A2(new_n1857_), .B(new_n14983_), .ZN(new_n14984_));
  AOI21_X1   g14727(.A1(new_n6994_), .A2(new_n1762_), .B(new_n14984_), .ZN(new_n14985_));
  XOR2_X1    g14728(.A1(new_n14714_), .A2(\a[29] ), .Z(new_n14986_));
  INV_X1     g14729(.I(new_n14986_), .ZN(new_n14987_));
  XOR2_X1    g14730(.A1(new_n14716_), .A2(new_n14987_), .Z(new_n14988_));
  AOI21_X1   g14731(.A1(new_n14710_), .A2(new_n14987_), .B(new_n14988_), .ZN(new_n14989_));
  XOR2_X1    g14732(.A1(new_n14989_), .A2(new_n14985_), .Z(new_n14990_));
  NAND2_X1   g14733(.A1(new_n14990_), .A2(new_n1750_), .ZN(new_n14991_));
  XNOR2_X1   g14734(.A1(new_n14989_), .A2(new_n14985_), .ZN(new_n14992_));
  NAND2_X1   g14735(.A1(new_n14992_), .A2(\a[26] ), .ZN(new_n14993_));
  AOI21_X1   g14736(.A1(new_n14993_), .A2(new_n14991_), .B(new_n14982_), .ZN(new_n14994_));
  NAND3_X1   g14737(.A1(new_n14993_), .A2(new_n14991_), .A3(new_n14982_), .ZN(new_n14995_));
  INV_X1     g14738(.I(new_n14995_), .ZN(new_n14996_));
  NAND2_X1   g14739(.A1(new_n14731_), .A2(new_n14729_), .ZN(new_n14997_));
  NAND2_X1   g14740(.A1(new_n14997_), .A2(new_n14730_), .ZN(new_n14998_));
  INV_X1     g14741(.I(new_n14998_), .ZN(new_n14999_));
  NOR3_X1    g14742(.A1(new_n14996_), .A2(new_n14994_), .A3(new_n14999_), .ZN(new_n15000_));
  INV_X1     g14743(.I(new_n14994_), .ZN(new_n15001_));
  AOI21_X1   g14744(.A1(new_n15001_), .A2(new_n14995_), .B(new_n14998_), .ZN(new_n15002_));
  OAI21_X1   g14745(.A1(new_n15002_), .A2(new_n15000_), .B(new_n14802_), .ZN(new_n15003_));
  AOI21_X1   g14746(.A1(new_n15001_), .A2(new_n14995_), .B(new_n14999_), .ZN(new_n15004_));
  NOR3_X1    g14747(.A1(new_n14996_), .A2(new_n14994_), .A3(new_n14998_), .ZN(new_n15005_));
  OAI21_X1   g14748(.A1(new_n15004_), .A2(new_n15005_), .B(new_n14801_), .ZN(new_n15006_));
  NAND2_X1   g14749(.A1(new_n15003_), .A2(new_n15006_), .ZN(new_n15007_));
  OAI22_X1   g14750(.A1(new_n1168_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n1163_), .ZN(new_n15008_));
  OAI21_X1   g14751(.A1(new_n7930_), .A2(new_n1255_), .B(new_n15008_), .ZN(new_n15009_));
  AOI21_X1   g14752(.A1(new_n8935_), .A2(new_n1170_), .B(new_n15009_), .ZN(new_n15010_));
  XOR2_X1    g14753(.A1(new_n14738_), .A2(\a[23] ), .Z(new_n15011_));
  NAND2_X1   g14754(.A1(new_n14747_), .A2(new_n15011_), .ZN(new_n15012_));
  INV_X1     g14755(.I(new_n15011_), .ZN(new_n15013_));
  NAND2_X1   g14756(.A1(new_n14733_), .A2(new_n15013_), .ZN(new_n15014_));
  INV_X1     g14757(.I(new_n15014_), .ZN(new_n15015_));
  NOR2_X1    g14758(.A1(new_n14733_), .A2(new_n15013_), .ZN(new_n15016_));
  OAI21_X1   g14759(.A1(new_n15015_), .A2(new_n15016_), .B(new_n14735_), .ZN(new_n15017_));
  AOI21_X1   g14760(.A1(new_n15017_), .A2(new_n15012_), .B(new_n15010_), .ZN(new_n15018_));
  INV_X1     g14761(.I(new_n15010_), .ZN(new_n15019_));
  INV_X1     g14762(.I(new_n15016_), .ZN(new_n15020_));
  AOI22_X1   g14763(.A1(new_n15020_), .A2(new_n15014_), .B1(new_n14741_), .B2(new_n15013_), .ZN(new_n15021_));
  NOR2_X1    g14764(.A1(new_n15021_), .A2(new_n15019_), .ZN(new_n15022_));
  OAI21_X1   g14765(.A1(new_n15022_), .A2(new_n15018_), .B(new_n1158_), .ZN(new_n15023_));
  NAND2_X1   g14766(.A1(new_n15021_), .A2(new_n15019_), .ZN(new_n15024_));
  NAND3_X1   g14767(.A1(new_n15017_), .A2(new_n15010_), .A3(new_n15012_), .ZN(new_n15025_));
  NAND3_X1   g14768(.A1(new_n15024_), .A2(new_n15025_), .A3(\a[20] ), .ZN(new_n15026_));
  AOI21_X1   g14769(.A1(new_n15023_), .A2(new_n15026_), .B(new_n15007_), .ZN(new_n15027_));
  NAND3_X1   g14770(.A1(new_n15001_), .A2(new_n14995_), .A3(new_n14998_), .ZN(new_n15028_));
  OAI21_X1   g14771(.A1(new_n14996_), .A2(new_n14994_), .B(new_n14999_), .ZN(new_n15029_));
  AOI21_X1   g14772(.A1(new_n15028_), .A2(new_n15029_), .B(new_n14801_), .ZN(new_n15030_));
  OAI21_X1   g14773(.A1(new_n14996_), .A2(new_n14994_), .B(new_n14998_), .ZN(new_n15031_));
  NAND3_X1   g14774(.A1(new_n15001_), .A2(new_n14995_), .A3(new_n14999_), .ZN(new_n15032_));
  AOI21_X1   g14775(.A1(new_n15032_), .A2(new_n15031_), .B(new_n14802_), .ZN(new_n15033_));
  NOR2_X1    g14776(.A1(new_n15030_), .A2(new_n15033_), .ZN(new_n15034_));
  AOI21_X1   g14777(.A1(new_n15024_), .A2(new_n15025_), .B(\a[20] ), .ZN(new_n15035_));
  NOR3_X1    g14778(.A1(new_n15022_), .A2(new_n15018_), .A3(new_n1158_), .ZN(new_n15036_));
  NOR3_X1    g14779(.A1(new_n15035_), .A2(new_n15036_), .A3(new_n15034_), .ZN(new_n15037_));
  NOR2_X1    g14780(.A1(new_n15037_), .A2(new_n15027_), .ZN(new_n15038_));
  NAND2_X1   g14781(.A1(new_n14763_), .A2(new_n14761_), .ZN(new_n15039_));
  AOI22_X1   g14782(.A1(new_n10814_), .A2(new_n942_), .B1(\b[63] ), .B2(new_n1458_), .ZN(new_n15040_));
  INV_X1     g14783(.I(new_n15040_), .ZN(new_n15041_));
  NAND3_X1   g14784(.A1(new_n15039_), .A2(new_n14762_), .A3(new_n15041_), .ZN(new_n15042_));
  AOI21_X1   g14785(.A1(new_n15039_), .A2(new_n14762_), .B(new_n15041_), .ZN(new_n15043_));
  INV_X1     g14786(.I(new_n15043_), .ZN(new_n15044_));
  AOI21_X1   g14787(.A1(new_n15044_), .A2(new_n15042_), .B(\a[17] ), .ZN(new_n15045_));
  NAND3_X1   g14788(.A1(new_n15044_), .A2(new_n15042_), .A3(\a[17] ), .ZN(new_n15046_));
  INV_X1     g14789(.I(new_n15046_), .ZN(new_n15047_));
  OAI21_X1   g14790(.A1(new_n15045_), .A2(new_n15047_), .B(new_n15038_), .ZN(new_n15048_));
  OAI21_X1   g14791(.A1(new_n15036_), .A2(new_n15035_), .B(new_n15034_), .ZN(new_n15049_));
  NAND3_X1   g14792(.A1(new_n15007_), .A2(new_n15023_), .A3(new_n15026_), .ZN(new_n15050_));
  NAND2_X1   g14793(.A1(new_n15049_), .A2(new_n15050_), .ZN(new_n15051_));
  INV_X1     g14794(.I(new_n15045_), .ZN(new_n15052_));
  NAND3_X1   g14795(.A1(new_n15052_), .A2(new_n15051_), .A3(new_n15046_), .ZN(new_n15053_));
  AOI21_X1   g14796(.A1(new_n15048_), .A2(new_n15053_), .B(new_n14796_), .ZN(new_n15054_));
  AOI21_X1   g14797(.A1(new_n15052_), .A2(new_n15046_), .B(new_n15051_), .ZN(new_n15055_));
  NOR3_X1    g14798(.A1(new_n15038_), .A2(new_n15047_), .A3(new_n15045_), .ZN(new_n15056_));
  NOR3_X1    g14799(.A1(new_n15055_), .A2(new_n15056_), .A3(new_n14795_), .ZN(new_n15057_));
  NOR2_X1    g14800(.A1(new_n15054_), .A2(new_n15057_), .ZN(new_n15058_));
  XOR2_X1    g14801(.A1(new_n14794_), .A2(new_n15058_), .Z(\f[80] ));
  XOR2_X1    g14802(.A1(new_n15040_), .A2(\a[17] ), .Z(new_n15060_));
  NAND2_X1   g14803(.A1(new_n15039_), .A2(new_n14762_), .ZN(new_n15061_));
  NOR2_X1    g14804(.A1(new_n15061_), .A2(new_n15060_), .ZN(new_n15062_));
  INV_X1     g14805(.I(new_n15060_), .ZN(new_n15063_));
  AOI21_X1   g14806(.A1(new_n15039_), .A2(new_n14762_), .B(new_n15063_), .ZN(new_n15064_));
  OAI22_X1   g14807(.A1(new_n15038_), .A2(new_n15060_), .B1(new_n15062_), .B2(new_n15064_), .ZN(new_n15065_));
  INV_X1     g14808(.I(new_n15021_), .ZN(new_n15066_));
  NOR2_X1    g14809(.A1(new_n15034_), .A2(new_n15066_), .ZN(new_n15067_));
  NAND2_X1   g14810(.A1(new_n15034_), .A2(new_n15066_), .ZN(new_n15068_));
  XOR2_X1    g14811(.A1(new_n15010_), .A2(new_n1158_), .Z(new_n15069_));
  INV_X1     g14812(.I(new_n15069_), .ZN(new_n15070_));
  AOI21_X1   g14813(.A1(new_n15068_), .A2(new_n15070_), .B(new_n15067_), .ZN(new_n15071_));
  INV_X1     g14814(.I(new_n15071_), .ZN(new_n15072_));
  OAI22_X1   g14815(.A1(new_n1168_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n1163_), .ZN(new_n15073_));
  NAND2_X1   g14816(.A1(new_n1774_), .A2(\b[61] ), .ZN(new_n15074_));
  AOI21_X1   g14817(.A1(new_n15073_), .A2(new_n15074_), .B(new_n1171_), .ZN(new_n15075_));
  NAND2_X1   g14818(.A1(new_n8963_), .A2(new_n15075_), .ZN(new_n15076_));
  XOR2_X1    g14819(.A1(new_n15076_), .A2(\a[20] ), .Z(new_n15077_));
  OAI22_X1   g14820(.A1(new_n1444_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n1439_), .ZN(new_n15078_));
  NAND2_X1   g14821(.A1(new_n2098_), .A2(\b[58] ), .ZN(new_n15079_));
  AOI21_X1   g14822(.A1(new_n15078_), .A2(new_n15079_), .B(new_n1447_), .ZN(new_n15080_));
  NAND2_X1   g14823(.A1(new_n7929_), .A2(new_n15080_), .ZN(new_n15081_));
  XOR2_X1    g14824(.A1(new_n15081_), .A2(\a[23] ), .Z(new_n15082_));
  INV_X1     g14825(.I(new_n15082_), .ZN(new_n15083_));
  AOI21_X1   g14826(.A1(new_n14802_), .A2(new_n15029_), .B(new_n15000_), .ZN(new_n15084_));
  INV_X1     g14827(.I(new_n14989_), .ZN(new_n15085_));
  NOR2_X1    g14828(.A1(new_n14981_), .A2(new_n15085_), .ZN(new_n15086_));
  NAND2_X1   g14829(.A1(new_n14981_), .A2(new_n15085_), .ZN(new_n15087_));
  XOR2_X1    g14830(.A1(new_n14985_), .A2(new_n1750_), .Z(new_n15088_));
  INV_X1     g14831(.I(new_n15088_), .ZN(new_n15089_));
  AOI21_X1   g14832(.A1(new_n15087_), .A2(new_n15089_), .B(new_n15086_), .ZN(new_n15090_));
  OAI22_X1   g14833(.A1(new_n2084_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n2079_), .ZN(new_n15091_));
  NAND2_X1   g14834(.A1(new_n2864_), .A2(\b[52] ), .ZN(new_n15092_));
  AOI21_X1   g14835(.A1(new_n15091_), .A2(new_n15092_), .B(new_n2087_), .ZN(new_n15093_));
  NAND2_X1   g14836(.A1(new_n6237_), .A2(new_n15093_), .ZN(new_n15094_));
  XOR2_X1    g14837(.A1(new_n15094_), .A2(\a[29] ), .Z(new_n15095_));
  INV_X1     g14838(.I(new_n15095_), .ZN(new_n15096_));
  NAND2_X1   g14839(.A1(new_n14976_), .A2(new_n14978_), .ZN(new_n15097_));
  NAND2_X1   g14840(.A1(new_n15097_), .A2(new_n14975_), .ZN(new_n15098_));
  NOR2_X1    g14841(.A1(new_n14965_), .A2(new_n14814_), .ZN(new_n15099_));
  AOI21_X1   g14842(.A1(new_n14968_), .A2(new_n14970_), .B(new_n15099_), .ZN(new_n15100_));
  INV_X1     g14843(.I(new_n14948_), .ZN(new_n15101_));
  OAI21_X1   g14844(.A1(new_n15101_), .A2(new_n14820_), .B(new_n14949_), .ZN(new_n15102_));
  NAND2_X1   g14845(.A1(new_n14941_), .A2(new_n14939_), .ZN(new_n15103_));
  NOR2_X1    g14846(.A1(new_n14931_), .A2(new_n14832_), .ZN(new_n15104_));
  AOI21_X1   g14847(.A1(new_n14913_), .A2(new_n14922_), .B(new_n14921_), .ZN(new_n15105_));
  AOI21_X1   g14848(.A1(new_n14909_), .A2(new_n14907_), .B(new_n14905_), .ZN(new_n15106_));
  NAND2_X1   g14849(.A1(new_n14879_), .A2(new_n14878_), .ZN(new_n15107_));
  NAND2_X1   g14850(.A1(new_n15107_), .A2(new_n14881_), .ZN(new_n15108_));
  INV_X1     g14851(.I(new_n15108_), .ZN(new_n15109_));
  NAND2_X1   g14852(.A1(new_n14873_), .A2(new_n14870_), .ZN(new_n15110_));
  AND2_X2    g14853(.A1(new_n15110_), .A2(new_n14872_), .Z(new_n15111_));
  NOR2_X1    g14854(.A1(new_n14849_), .A2(new_n14854_), .ZN(new_n15112_));
  NOR2_X1    g14855(.A1(new_n15112_), .A2(new_n14856_), .ZN(new_n15113_));
  OAI22_X1   g14856(.A1(new_n1393_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1305_), .ZN(new_n15114_));
  NAND2_X1   g14857(.A1(new_n9644_), .A2(\b[19] ), .ZN(new_n15115_));
  AOI21_X1   g14858(.A1(new_n15115_), .A2(new_n15114_), .B(new_n8321_), .ZN(new_n15116_));
  NAND2_X1   g14859(.A1(new_n1396_), .A2(new_n15116_), .ZN(new_n15117_));
  XOR2_X1    g14860(.A1(new_n15117_), .A2(new_n8309_), .Z(new_n15118_));
  NOR2_X1    g14861(.A1(new_n8985_), .A2(new_n1124_), .ZN(new_n15119_));
  NOR2_X1    g14862(.A1(new_n9364_), .A2(new_n1044_), .ZN(new_n15120_));
  XNOR2_X1   g14863(.A1(new_n15119_), .A2(new_n15120_), .ZN(new_n15121_));
  XOR2_X1    g14864(.A1(new_n15121_), .A2(\a[17] ), .Z(new_n15122_));
  NOR2_X1    g14865(.A1(new_n15122_), .A2(new_n14853_), .ZN(new_n15123_));
  NOR2_X1    g14866(.A1(new_n15121_), .A2(new_n930_), .ZN(new_n15124_));
  INV_X1     g14867(.I(new_n15124_), .ZN(new_n15125_));
  NAND2_X1   g14868(.A1(new_n15121_), .A2(new_n930_), .ZN(new_n15126_));
  AOI21_X1   g14869(.A1(new_n15125_), .A2(new_n15126_), .B(new_n14855_), .ZN(new_n15127_));
  NOR2_X1    g14870(.A1(new_n15123_), .A2(new_n15127_), .ZN(new_n15128_));
  NOR2_X1    g14871(.A1(new_n15118_), .A2(new_n15128_), .ZN(new_n15129_));
  INV_X1     g14872(.I(new_n15129_), .ZN(new_n15130_));
  NAND2_X1   g14873(.A1(new_n15118_), .A2(new_n15128_), .ZN(new_n15131_));
  AOI21_X1   g14874(.A1(new_n15130_), .A2(new_n15131_), .B(new_n15113_), .ZN(new_n15132_));
  INV_X1     g14875(.I(new_n15132_), .ZN(new_n15133_));
  XOR2_X1    g14876(.A1(new_n15118_), .A2(new_n15128_), .Z(new_n15134_));
  NAND2_X1   g14877(.A1(new_n15134_), .A2(new_n15113_), .ZN(new_n15135_));
  NAND2_X1   g14878(.A1(new_n15133_), .A2(new_n15135_), .ZN(new_n15136_));
  OAI22_X1   g14879(.A1(new_n1709_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1601_), .ZN(new_n15137_));
  NAND2_X1   g14880(.A1(new_n8628_), .A2(\b[22] ), .ZN(new_n15138_));
  AOI21_X1   g14881(.A1(new_n15138_), .A2(new_n15137_), .B(new_n7354_), .ZN(new_n15139_));
  NAND2_X1   g14882(.A1(new_n1708_), .A2(new_n15139_), .ZN(new_n15140_));
  XOR2_X1    g14883(.A1(new_n15140_), .A2(\a[59] ), .Z(new_n15141_));
  INV_X1     g14884(.I(new_n15141_), .ZN(new_n15142_));
  XOR2_X1    g14885(.A1(new_n15136_), .A2(new_n15142_), .Z(new_n15143_));
  INV_X1     g14886(.I(new_n15143_), .ZN(new_n15144_));
  AOI21_X1   g14887(.A1(new_n15133_), .A2(new_n15135_), .B(new_n15141_), .ZN(new_n15145_));
  NOR2_X1    g14888(.A1(new_n15136_), .A2(new_n15142_), .ZN(new_n15146_));
  OAI21_X1   g14889(.A1(new_n15146_), .A2(new_n15145_), .B(new_n15111_), .ZN(new_n15147_));
  OAI21_X1   g14890(.A1(new_n15144_), .A2(new_n15111_), .B(new_n15147_), .ZN(new_n15148_));
  OAI22_X1   g14891(.A1(new_n6721_), .A2(new_n1927_), .B1(new_n6723_), .B2(new_n2039_), .ZN(new_n15149_));
  NAND2_X1   g14892(.A1(new_n7617_), .A2(\b[25] ), .ZN(new_n15150_));
  AOI21_X1   g14893(.A1(new_n15150_), .A2(new_n15149_), .B(new_n6731_), .ZN(new_n15151_));
  NAND2_X1   g14894(.A1(new_n2042_), .A2(new_n15151_), .ZN(new_n15152_));
  XOR2_X1    g14895(.A1(new_n15152_), .A2(\a[56] ), .Z(new_n15153_));
  XNOR2_X1   g14896(.A1(new_n15148_), .A2(new_n15153_), .ZN(new_n15154_));
  NOR2_X1    g14897(.A1(new_n15148_), .A2(new_n15153_), .ZN(new_n15155_));
  NAND2_X1   g14898(.A1(new_n15148_), .A2(new_n15153_), .ZN(new_n15156_));
  INV_X1     g14899(.I(new_n15156_), .ZN(new_n15157_));
  OAI21_X1   g14900(.A1(new_n15157_), .A2(new_n15155_), .B(new_n15109_), .ZN(new_n15158_));
  OAI21_X1   g14901(.A1(new_n15109_), .A2(new_n15154_), .B(new_n15158_), .ZN(new_n15159_));
  OAI22_X1   g14902(.A1(new_n5786_), .A2(new_n2405_), .B1(new_n2272_), .B2(new_n5792_), .ZN(new_n15160_));
  NAND2_X1   g14903(.A1(new_n6745_), .A2(\b[28] ), .ZN(new_n15161_));
  AOI21_X1   g14904(.A1(new_n15161_), .A2(new_n15160_), .B(new_n5796_), .ZN(new_n15162_));
  NAND2_X1   g14905(.A1(new_n2404_), .A2(new_n15162_), .ZN(new_n15163_));
  XOR2_X1    g14906(.A1(new_n15163_), .A2(\a[53] ), .Z(new_n15164_));
  AOI21_X1   g14907(.A1(new_n14883_), .A2(new_n14898_), .B(new_n14897_), .ZN(new_n15165_));
  NOR2_X1    g14908(.A1(new_n15165_), .A2(new_n15164_), .ZN(new_n15166_));
  AND2_X2    g14909(.A1(new_n15165_), .A2(new_n15164_), .Z(new_n15167_));
  OAI21_X1   g14910(.A1(new_n15167_), .A2(new_n15166_), .B(new_n15159_), .ZN(new_n15168_));
  XNOR2_X1   g14911(.A1(new_n15165_), .A2(new_n15164_), .ZN(new_n15169_));
  OAI21_X1   g14912(.A1(new_n15169_), .A2(new_n15159_), .B(new_n15168_), .ZN(new_n15170_));
  OAI22_X1   g14913(.A1(new_n5228_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n5225_), .ZN(new_n15171_));
  NAND2_X1   g14914(.A1(new_n5387_), .A2(\b[31] ), .ZN(new_n15172_));
  AOI21_X1   g14915(.A1(new_n15171_), .A2(new_n15172_), .B(new_n5231_), .ZN(new_n15173_));
  NAND2_X1   g14916(.A1(new_n2797_), .A2(new_n15173_), .ZN(new_n15174_));
  XOR2_X1    g14917(.A1(new_n15174_), .A2(\a[50] ), .Z(new_n15175_));
  NOR2_X1    g14918(.A1(new_n15170_), .A2(new_n15175_), .ZN(new_n15176_));
  NAND2_X1   g14919(.A1(new_n15170_), .A2(new_n15175_), .ZN(new_n15177_));
  INV_X1     g14920(.I(new_n15177_), .ZN(new_n15178_));
  NOR2_X1    g14921(.A1(new_n15178_), .A2(new_n15176_), .ZN(new_n15179_));
  XOR2_X1    g14922(.A1(new_n15170_), .A2(new_n15175_), .Z(new_n15180_));
  NAND2_X1   g14923(.A1(new_n15180_), .A2(new_n15106_), .ZN(new_n15181_));
  OAI21_X1   g14924(.A1(new_n15106_), .A2(new_n15179_), .B(new_n15181_), .ZN(new_n15182_));
  OAI22_X1   g14925(.A1(new_n4711_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n4706_), .ZN(new_n15183_));
  NAND2_X1   g14926(.A1(new_n5814_), .A2(\b[34] ), .ZN(new_n15184_));
  AOI21_X1   g14927(.A1(new_n15183_), .A2(new_n15184_), .B(new_n4714_), .ZN(new_n15185_));
  NAND2_X1   g14928(.A1(new_n3246_), .A2(new_n15185_), .ZN(new_n15186_));
  XOR2_X1    g14929(.A1(new_n15186_), .A2(\a[47] ), .Z(new_n15187_));
  XOR2_X1    g14930(.A1(new_n15182_), .A2(new_n15187_), .Z(new_n15188_));
  NOR2_X1    g14931(.A1(new_n15188_), .A2(new_n15105_), .ZN(new_n15189_));
  INV_X1     g14932(.I(new_n15105_), .ZN(new_n15190_));
  INV_X1     g14933(.I(new_n15187_), .ZN(new_n15191_));
  NAND2_X1   g14934(.A1(new_n15182_), .A2(new_n15191_), .ZN(new_n15192_));
  NOR2_X1    g14935(.A1(new_n15182_), .A2(new_n15191_), .ZN(new_n15193_));
  INV_X1     g14936(.I(new_n15193_), .ZN(new_n15194_));
  AOI21_X1   g14937(.A1(new_n15194_), .A2(new_n15192_), .B(new_n15190_), .ZN(new_n15195_));
  OAI22_X1   g14938(.A1(new_n4208_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n4203_), .ZN(new_n15196_));
  NAND2_X1   g14939(.A1(new_n5244_), .A2(\b[37] ), .ZN(new_n15197_));
  AOI21_X1   g14940(.A1(new_n15196_), .A2(new_n15197_), .B(new_n4211_), .ZN(new_n15198_));
  NAND2_X1   g14941(.A1(new_n3700_), .A2(new_n15198_), .ZN(new_n15199_));
  XOR2_X1    g14942(.A1(new_n15199_), .A2(\a[44] ), .Z(new_n15200_));
  NOR3_X1    g14943(.A1(new_n15189_), .A2(new_n15195_), .A3(new_n15200_), .ZN(new_n15201_));
  NOR2_X1    g14944(.A1(new_n15189_), .A2(new_n15195_), .ZN(new_n15202_));
  INV_X1     g14945(.I(new_n15200_), .ZN(new_n15203_));
  NOR2_X1    g14946(.A1(new_n15202_), .A2(new_n15203_), .ZN(new_n15204_));
  OAI22_X1   g14947(.A1(new_n15201_), .A2(new_n15204_), .B1(new_n14928_), .B2(new_n15104_), .ZN(new_n15205_));
  NOR2_X1    g14948(.A1(new_n15104_), .A2(new_n14928_), .ZN(new_n15206_));
  XOR2_X1    g14949(.A1(new_n15202_), .A2(new_n15203_), .Z(new_n15207_));
  NAND2_X1   g14950(.A1(new_n15207_), .A2(new_n15206_), .ZN(new_n15208_));
  NAND2_X1   g14951(.A1(new_n15208_), .A2(new_n15205_), .ZN(new_n15209_));
  OAI22_X1   g14952(.A1(new_n3736_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n3731_), .ZN(new_n15210_));
  NAND2_X1   g14953(.A1(new_n4730_), .A2(\b[40] ), .ZN(new_n15211_));
  AOI21_X1   g14954(.A1(new_n15210_), .A2(new_n15211_), .B(new_n3739_), .ZN(new_n15212_));
  NAND2_X1   g14955(.A1(new_n4017_), .A2(new_n15212_), .ZN(new_n15213_));
  XOR2_X1    g14956(.A1(new_n15213_), .A2(\a[41] ), .Z(new_n15214_));
  XOR2_X1    g14957(.A1(new_n15209_), .A2(new_n15214_), .Z(new_n15215_));
  AOI21_X1   g14958(.A1(new_n14940_), .A2(new_n15103_), .B(new_n15215_), .ZN(new_n15216_));
  NAND2_X1   g14959(.A1(new_n15103_), .A2(new_n14940_), .ZN(new_n15217_));
  INV_X1     g14960(.I(new_n15209_), .ZN(new_n15218_));
  NOR2_X1    g14961(.A1(new_n15218_), .A2(new_n15214_), .ZN(new_n15219_));
  INV_X1     g14962(.I(new_n15214_), .ZN(new_n15220_));
  NOR2_X1    g14963(.A1(new_n15209_), .A2(new_n15220_), .ZN(new_n15221_));
  NOR2_X1    g14964(.A1(new_n15219_), .A2(new_n15221_), .ZN(new_n15222_));
  NOR2_X1    g14965(.A1(new_n15222_), .A2(new_n15217_), .ZN(new_n15223_));
  NOR2_X1    g14966(.A1(new_n15216_), .A2(new_n15223_), .ZN(new_n15224_));
  OAI22_X1   g14967(.A1(new_n3298_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n3293_), .ZN(new_n15225_));
  NAND2_X1   g14968(.A1(new_n4227_), .A2(\b[43] ), .ZN(new_n15226_));
  AOI21_X1   g14969(.A1(new_n15225_), .A2(new_n15226_), .B(new_n3301_), .ZN(new_n15227_));
  NAND2_X1   g14970(.A1(new_n4513_), .A2(new_n15227_), .ZN(new_n15228_));
  XOR2_X1    g14971(.A1(new_n15228_), .A2(\a[38] ), .Z(new_n15229_));
  INV_X1     g14972(.I(new_n15229_), .ZN(new_n15230_));
  XOR2_X1    g14973(.A1(new_n15224_), .A2(new_n15230_), .Z(new_n15231_));
  AND2_X2    g14974(.A1(new_n15231_), .A2(new_n15102_), .Z(new_n15232_));
  NAND2_X1   g14975(.A1(new_n15224_), .A2(new_n15230_), .ZN(new_n15233_));
  OAI21_X1   g14976(.A1(new_n15216_), .A2(new_n15223_), .B(new_n15229_), .ZN(new_n15234_));
  AOI21_X1   g14977(.A1(new_n15233_), .A2(new_n15234_), .B(new_n15102_), .ZN(new_n15235_));
  NOR2_X1    g14978(.A1(new_n15232_), .A2(new_n15235_), .ZN(new_n15236_));
  OAI22_X1   g14979(.A1(new_n2846_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n2841_), .ZN(new_n15237_));
  NAND2_X1   g14980(.A1(new_n3755_), .A2(\b[46] ), .ZN(new_n15238_));
  AOI21_X1   g14981(.A1(new_n15237_), .A2(new_n15238_), .B(new_n2849_), .ZN(new_n15239_));
  NAND2_X1   g14982(.A1(new_n5177_), .A2(new_n15239_), .ZN(new_n15240_));
  XOR2_X1    g14983(.A1(new_n15240_), .A2(\a[35] ), .Z(new_n15241_));
  AND2_X2    g14984(.A1(new_n14951_), .A2(new_n14962_), .Z(new_n15242_));
  NOR2_X1    g14985(.A1(new_n15242_), .A2(new_n14960_), .ZN(new_n15243_));
  NOR2_X1    g14986(.A1(new_n15243_), .A2(new_n15241_), .ZN(new_n15244_));
  INV_X1     g14987(.I(new_n15244_), .ZN(new_n15245_));
  NAND2_X1   g14988(.A1(new_n15243_), .A2(new_n15241_), .ZN(new_n15246_));
  AOI21_X1   g14989(.A1(new_n15245_), .A2(new_n15246_), .B(new_n15236_), .ZN(new_n15247_));
  INV_X1     g14990(.I(new_n15236_), .ZN(new_n15248_));
  XNOR2_X1   g14991(.A1(new_n15243_), .A2(new_n15241_), .ZN(new_n15249_));
  NOR2_X1    g14992(.A1(new_n15249_), .A2(new_n15248_), .ZN(new_n15250_));
  OAI22_X1   g14993(.A1(new_n2452_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n2447_), .ZN(new_n15251_));
  NAND2_X1   g14994(.A1(new_n3312_), .A2(\b[49] ), .ZN(new_n15252_));
  AOI21_X1   g14995(.A1(new_n15251_), .A2(new_n15252_), .B(new_n2455_), .ZN(new_n15253_));
  NAND2_X1   g14996(.A1(new_n5741_), .A2(new_n15253_), .ZN(new_n15254_));
  XOR2_X1    g14997(.A1(new_n15254_), .A2(\a[32] ), .Z(new_n15255_));
  NOR3_X1    g14998(.A1(new_n15250_), .A2(new_n15247_), .A3(new_n15255_), .ZN(new_n15256_));
  NOR2_X1    g14999(.A1(new_n15250_), .A2(new_n15247_), .ZN(new_n15257_));
  INV_X1     g15000(.I(new_n15255_), .ZN(new_n15258_));
  NOR2_X1    g15001(.A1(new_n15257_), .A2(new_n15258_), .ZN(new_n15259_));
  NOR2_X1    g15002(.A1(new_n15259_), .A2(new_n15256_), .ZN(new_n15260_));
  XOR2_X1    g15003(.A1(new_n15257_), .A2(new_n15258_), .Z(new_n15261_));
  NAND2_X1   g15004(.A1(new_n15261_), .A2(new_n15100_), .ZN(new_n15262_));
  OAI21_X1   g15005(.A1(new_n15100_), .A2(new_n15260_), .B(new_n15262_), .ZN(new_n15263_));
  AND2_X2    g15006(.A1(new_n15263_), .A2(new_n15098_), .Z(new_n15264_));
  NOR2_X1    g15007(.A1(new_n15263_), .A2(new_n15098_), .ZN(new_n15265_));
  OAI21_X1   g15008(.A1(new_n15264_), .A2(new_n15265_), .B(new_n15096_), .ZN(new_n15266_));
  XOR2_X1    g15009(.A1(new_n15263_), .A2(new_n15098_), .Z(new_n15267_));
  NAND2_X1   g15010(.A1(new_n15267_), .A2(new_n15095_), .ZN(new_n15268_));
  OAI22_X1   g15011(.A1(new_n1760_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n1755_), .ZN(new_n15269_));
  NAND2_X1   g15012(.A1(new_n2470_), .A2(\b[55] ), .ZN(new_n15270_));
  AOI21_X1   g15013(.A1(new_n15269_), .A2(new_n15270_), .B(new_n1763_), .ZN(new_n15271_));
  NAND2_X1   g15014(.A1(new_n7308_), .A2(new_n15271_), .ZN(new_n15272_));
  XOR2_X1    g15015(.A1(new_n15272_), .A2(\a[26] ), .Z(new_n15273_));
  AOI21_X1   g15016(.A1(new_n15268_), .A2(new_n15266_), .B(new_n15273_), .ZN(new_n15274_));
  INV_X1     g15017(.I(new_n15274_), .ZN(new_n15275_));
  NAND3_X1   g15018(.A1(new_n15268_), .A2(new_n15266_), .A3(new_n15273_), .ZN(new_n15276_));
  AOI21_X1   g15019(.A1(new_n15275_), .A2(new_n15276_), .B(new_n15090_), .ZN(new_n15277_));
  INV_X1     g15020(.I(new_n15090_), .ZN(new_n15278_));
  INV_X1     g15021(.I(new_n15273_), .ZN(new_n15279_));
  NAND3_X1   g15022(.A1(new_n15268_), .A2(new_n15266_), .A3(new_n15279_), .ZN(new_n15280_));
  INV_X1     g15023(.I(new_n15266_), .ZN(new_n15281_));
  XNOR2_X1   g15024(.A1(new_n15263_), .A2(new_n15098_), .ZN(new_n15282_));
  NOR2_X1    g15025(.A1(new_n15282_), .A2(new_n15096_), .ZN(new_n15283_));
  OAI21_X1   g15026(.A1(new_n15281_), .A2(new_n15283_), .B(new_n15273_), .ZN(new_n15284_));
  AOI21_X1   g15027(.A1(new_n15284_), .A2(new_n15280_), .B(new_n15278_), .ZN(new_n15285_));
  NOR2_X1    g15028(.A1(new_n15277_), .A2(new_n15285_), .ZN(new_n15286_));
  NOR2_X1    g15029(.A1(new_n15286_), .A2(new_n15084_), .ZN(new_n15287_));
  INV_X1     g15030(.I(new_n15084_), .ZN(new_n15288_));
  INV_X1     g15031(.I(new_n15276_), .ZN(new_n15289_));
  OAI21_X1   g15032(.A1(new_n15289_), .A2(new_n15274_), .B(new_n15278_), .ZN(new_n15290_));
  INV_X1     g15033(.I(new_n15280_), .ZN(new_n15291_));
  AOI21_X1   g15034(.A1(new_n15268_), .A2(new_n15266_), .B(new_n15279_), .ZN(new_n15292_));
  OAI21_X1   g15035(.A1(new_n15291_), .A2(new_n15292_), .B(new_n15090_), .ZN(new_n15293_));
  NAND2_X1   g15036(.A1(new_n15290_), .A2(new_n15293_), .ZN(new_n15294_));
  NOR2_X1    g15037(.A1(new_n15294_), .A2(new_n15288_), .ZN(new_n15295_));
  OAI21_X1   g15038(.A1(new_n15295_), .A2(new_n15287_), .B(new_n15083_), .ZN(new_n15296_));
  NOR2_X1    g15039(.A1(new_n15286_), .A2(new_n15288_), .ZN(new_n15297_));
  NOR2_X1    g15040(.A1(new_n15294_), .A2(new_n15084_), .ZN(new_n15298_));
  OAI21_X1   g15041(.A1(new_n15298_), .A2(new_n15297_), .B(new_n15082_), .ZN(new_n15299_));
  AOI21_X1   g15042(.A1(new_n15299_), .A2(new_n15296_), .B(new_n15077_), .ZN(new_n15300_));
  INV_X1     g15043(.I(new_n15077_), .ZN(new_n15301_));
  NAND2_X1   g15044(.A1(new_n15294_), .A2(new_n15288_), .ZN(new_n15302_));
  NAND2_X1   g15045(.A1(new_n15286_), .A2(new_n15084_), .ZN(new_n15303_));
  AOI21_X1   g15046(.A1(new_n15302_), .A2(new_n15303_), .B(new_n15082_), .ZN(new_n15304_));
  NAND2_X1   g15047(.A1(new_n15294_), .A2(new_n15084_), .ZN(new_n15305_));
  NAND2_X1   g15048(.A1(new_n15286_), .A2(new_n15288_), .ZN(new_n15306_));
  AOI21_X1   g15049(.A1(new_n15305_), .A2(new_n15306_), .B(new_n15083_), .ZN(new_n15307_));
  NOR3_X1    g15050(.A1(new_n15304_), .A2(new_n15307_), .A3(new_n15301_), .ZN(new_n15308_));
  OAI21_X1   g15051(.A1(new_n15300_), .A2(new_n15308_), .B(new_n15072_), .ZN(new_n15309_));
  AOI21_X1   g15052(.A1(new_n15299_), .A2(new_n15296_), .B(new_n15301_), .ZN(new_n15310_));
  NOR3_X1    g15053(.A1(new_n15304_), .A2(new_n15307_), .A3(new_n15077_), .ZN(new_n15311_));
  OAI21_X1   g15054(.A1(new_n15310_), .A2(new_n15311_), .B(new_n15071_), .ZN(new_n15312_));
  AOI21_X1   g15055(.A1(new_n15309_), .A2(new_n15312_), .B(new_n15065_), .ZN(new_n15313_));
  INV_X1     g15056(.I(new_n15065_), .ZN(new_n15314_));
  NAND2_X1   g15057(.A1(new_n15309_), .A2(new_n15312_), .ZN(new_n15315_));
  NOR2_X1    g15058(.A1(new_n15315_), .A2(new_n15314_), .ZN(new_n15316_));
  NOR2_X1    g15059(.A1(new_n15316_), .A2(new_n15313_), .ZN(new_n15317_));
  INV_X1     g15060(.I(new_n15054_), .ZN(new_n15318_));
  INV_X1     g15061(.I(new_n14786_), .ZN(new_n15319_));
  AOI21_X1   g15062(.A1(new_n14245_), .A2(new_n14246_), .B(new_n14244_), .ZN(new_n15320_));
  NOR3_X1    g15063(.A1(new_n14242_), .A2(new_n14239_), .A3(new_n13984_), .ZN(new_n15321_));
  NOR2_X1    g15064(.A1(new_n15321_), .A2(new_n15320_), .ZN(new_n15322_));
  AOI21_X1   g15065(.A1(new_n13977_), .A2(new_n13978_), .B(new_n13976_), .ZN(new_n15323_));
  NOR3_X1    g15066(.A1(new_n15323_), .A2(new_n14526_), .A3(new_n13983_), .ZN(new_n15324_));
  AOI21_X1   g15067(.A1(new_n13975_), .A2(new_n14527_), .B(new_n14528_), .ZN(new_n15325_));
  OAI21_X1   g15068(.A1(new_n15325_), .A2(new_n15324_), .B(new_n15322_), .ZN(new_n15326_));
  NOR3_X1    g15069(.A1(new_n14533_), .A2(new_n14525_), .A3(new_n13983_), .ZN(new_n15327_));
  OAI21_X1   g15070(.A1(new_n15326_), .A2(new_n15327_), .B(new_n14793_), .ZN(new_n15328_));
  NAND3_X1   g15071(.A1(new_n15328_), .A2(new_n15319_), .A3(new_n15058_), .ZN(new_n15329_));
  NAND2_X1   g15072(.A1(new_n15329_), .A2(new_n15318_), .ZN(new_n15330_));
  XOR2_X1    g15073(.A1(new_n15330_), .A2(new_n15317_), .Z(\f[81] ));
  NAND3_X1   g15074(.A1(new_n15299_), .A2(new_n15296_), .A3(new_n15077_), .ZN(new_n15332_));
  AOI21_X1   g15075(.A1(new_n15072_), .A2(new_n15332_), .B(new_n15300_), .ZN(new_n15333_));
  NOR2_X1    g15076(.A1(new_n1255_), .A2(new_n8932_), .ZN(new_n15334_));
  NOR2_X1    g15077(.A1(new_n1163_), .A2(new_n8956_), .ZN(new_n15335_));
  NOR4_X1    g15078(.A1(new_n9323_), .A2(new_n1171_), .A3(new_n15334_), .A4(new_n15335_), .ZN(new_n15336_));
  XOR2_X1    g15079(.A1(new_n15336_), .A2(new_n1158_), .Z(new_n15337_));
  INV_X1     g15080(.I(new_n15337_), .ZN(new_n15338_));
  OAI22_X1   g15081(.A1(new_n1444_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n1439_), .ZN(new_n15339_));
  NAND2_X1   g15082(.A1(new_n2098_), .A2(\b[59] ), .ZN(new_n15340_));
  AOI21_X1   g15083(.A1(new_n15339_), .A2(new_n15340_), .B(new_n1447_), .ZN(new_n15341_));
  NAND2_X1   g15084(.A1(new_n8550_), .A2(new_n15341_), .ZN(new_n15342_));
  XOR2_X1    g15085(.A1(new_n15342_), .A2(\a[23] ), .Z(new_n15343_));
  AOI21_X1   g15086(.A1(new_n15278_), .A2(new_n15276_), .B(new_n15274_), .ZN(new_n15344_));
  INV_X1     g15087(.I(new_n15344_), .ZN(new_n15345_));
  OAI22_X1   g15088(.A1(new_n1760_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n1755_), .ZN(new_n15346_));
  NAND2_X1   g15089(.A1(new_n2470_), .A2(\b[56] ), .ZN(new_n15347_));
  AOI21_X1   g15090(.A1(new_n15346_), .A2(new_n15347_), .B(new_n1763_), .ZN(new_n15348_));
  NAND2_X1   g15091(.A1(new_n7559_), .A2(new_n15348_), .ZN(new_n15349_));
  XOR2_X1    g15092(.A1(new_n15349_), .A2(\a[26] ), .Z(new_n15350_));
  NOR2_X1    g15093(.A1(new_n15265_), .A2(new_n15095_), .ZN(new_n15351_));
  NOR2_X1    g15094(.A1(new_n15351_), .A2(new_n15264_), .ZN(new_n15352_));
  OAI22_X1   g15095(.A1(new_n2084_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n2079_), .ZN(new_n15353_));
  NAND2_X1   g15096(.A1(new_n2864_), .A2(\b[53] ), .ZN(new_n15354_));
  AOI21_X1   g15097(.A1(new_n15353_), .A2(new_n15354_), .B(new_n2087_), .ZN(new_n15355_));
  NAND2_X1   g15098(.A1(new_n6471_), .A2(new_n15355_), .ZN(new_n15356_));
  XOR2_X1    g15099(.A1(new_n15356_), .A2(\a[29] ), .Z(new_n15357_));
  NOR2_X1    g15100(.A1(new_n15259_), .A2(new_n15100_), .ZN(new_n15358_));
  NOR2_X1    g15101(.A1(new_n15358_), .A2(new_n15256_), .ZN(new_n15359_));
  OAI22_X1   g15102(.A1(new_n2452_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n2447_), .ZN(new_n15360_));
  NAND2_X1   g15103(.A1(new_n3312_), .A2(\b[50] ), .ZN(new_n15361_));
  AOI21_X1   g15104(.A1(new_n15360_), .A2(new_n15361_), .B(new_n2455_), .ZN(new_n15362_));
  NAND2_X1   g15105(.A1(new_n5954_), .A2(new_n15362_), .ZN(new_n15363_));
  XOR2_X1    g15106(.A1(new_n15363_), .A2(\a[32] ), .Z(new_n15364_));
  AOI21_X1   g15107(.A1(new_n15241_), .A2(new_n15243_), .B(new_n15248_), .ZN(new_n15365_));
  NOR2_X1    g15108(.A1(new_n15365_), .A2(new_n15244_), .ZN(new_n15366_));
  OAI22_X1   g15109(.A1(new_n3298_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n3293_), .ZN(new_n15367_));
  NAND2_X1   g15110(.A1(new_n4227_), .A2(\b[44] ), .ZN(new_n15368_));
  AOI21_X1   g15111(.A1(new_n15367_), .A2(new_n15368_), .B(new_n3301_), .ZN(new_n15369_));
  NAND2_X1   g15112(.A1(new_n4833_), .A2(new_n15369_), .ZN(new_n15370_));
  XOR2_X1    g15113(.A1(new_n15370_), .A2(\a[38] ), .Z(new_n15371_));
  NOR2_X1    g15114(.A1(new_n15204_), .A2(new_n15206_), .ZN(new_n15372_));
  NOR2_X1    g15115(.A1(new_n15372_), .A2(new_n15201_), .ZN(new_n15373_));
  OAI22_X1   g15116(.A1(new_n4208_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n4203_), .ZN(new_n15374_));
  NAND2_X1   g15117(.A1(new_n5244_), .A2(\b[38] ), .ZN(new_n15375_));
  AOI21_X1   g15118(.A1(new_n15374_), .A2(new_n15375_), .B(new_n4211_), .ZN(new_n15376_));
  NAND2_X1   g15119(.A1(new_n3844_), .A2(new_n15376_), .ZN(new_n15377_));
  XOR2_X1    g15120(.A1(new_n15377_), .A2(\a[44] ), .Z(new_n15378_));
  OAI21_X1   g15121(.A1(new_n15105_), .A2(new_n15193_), .B(new_n15192_), .ZN(new_n15379_));
  OAI22_X1   g15122(.A1(new_n5228_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n5225_), .ZN(new_n15380_));
  NAND2_X1   g15123(.A1(new_n5387_), .A2(\b[32] ), .ZN(new_n15381_));
  AOI21_X1   g15124(.A1(new_n15380_), .A2(new_n15381_), .B(new_n5231_), .ZN(new_n15382_));
  NAND2_X1   g15125(.A1(new_n2963_), .A2(new_n15382_), .ZN(new_n15383_));
  XOR2_X1    g15126(.A1(new_n15383_), .A2(\a[50] ), .Z(new_n15384_));
  OAI22_X1   g15127(.A1(new_n6721_), .A2(new_n2039_), .B1(new_n6723_), .B2(new_n2175_), .ZN(new_n15385_));
  NAND2_X1   g15128(.A1(new_n7617_), .A2(\b[26] ), .ZN(new_n15386_));
  AOI21_X1   g15129(.A1(new_n15386_), .A2(new_n15385_), .B(new_n6731_), .ZN(new_n15387_));
  NAND2_X1   g15130(.A1(new_n2174_), .A2(new_n15387_), .ZN(new_n15388_));
  XOR2_X1    g15131(.A1(new_n15388_), .A2(\a[56] ), .Z(new_n15389_));
  NOR2_X1    g15132(.A1(new_n15146_), .A2(new_n15111_), .ZN(new_n15390_));
  NOR2_X1    g15133(.A1(new_n15390_), .A2(new_n15145_), .ZN(new_n15391_));
  OAI22_X1   g15134(.A1(new_n1518_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1393_), .ZN(new_n15392_));
  NAND2_X1   g15135(.A1(new_n9644_), .A2(\b[20] ), .ZN(new_n15393_));
  AOI21_X1   g15136(.A1(new_n15393_), .A2(new_n15392_), .B(new_n8321_), .ZN(new_n15394_));
  NAND2_X1   g15137(.A1(new_n1517_), .A2(new_n15394_), .ZN(new_n15395_));
  XOR2_X1    g15138(.A1(new_n15395_), .A2(new_n8309_), .Z(new_n15396_));
  NAND2_X1   g15139(.A1(new_n15126_), .A2(new_n14855_), .ZN(new_n15397_));
  NAND2_X1   g15140(.A1(new_n15397_), .A2(new_n15125_), .ZN(new_n15398_));
  NOR3_X1    g15141(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n1124_), .ZN(new_n15399_));
  NOR2_X1    g15142(.A1(new_n9364_), .A2(new_n1124_), .ZN(new_n15400_));
  NOR3_X1    g15143(.A1(new_n15400_), .A2(new_n1222_), .A3(new_n8985_), .ZN(new_n15401_));
  NOR2_X1    g15144(.A1(new_n15401_), .A2(new_n15399_), .ZN(new_n15402_));
  INV_X1     g15145(.I(new_n15402_), .ZN(new_n15403_));
  XOR2_X1    g15146(.A1(new_n15398_), .A2(new_n15403_), .Z(new_n15404_));
  INV_X1     g15147(.I(new_n15404_), .ZN(new_n15405_));
  NOR2_X1    g15148(.A1(new_n15398_), .A2(new_n15402_), .ZN(new_n15406_));
  INV_X1     g15149(.I(new_n15406_), .ZN(new_n15407_));
  NAND2_X1   g15150(.A1(new_n15398_), .A2(new_n15402_), .ZN(new_n15408_));
  AOI21_X1   g15151(.A1(new_n15407_), .A2(new_n15408_), .B(new_n15396_), .ZN(new_n15409_));
  AOI21_X1   g15152(.A1(new_n15396_), .A2(new_n15405_), .B(new_n15409_), .ZN(new_n15410_));
  OAI21_X1   g15153(.A1(new_n15113_), .A2(new_n15129_), .B(new_n15131_), .ZN(new_n15411_));
  OAI22_X1   g15154(.A1(new_n1825_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1709_), .ZN(new_n15412_));
  NAND2_X1   g15155(.A1(new_n8628_), .A2(\b[23] ), .ZN(new_n15413_));
  AOI21_X1   g15156(.A1(new_n15413_), .A2(new_n15412_), .B(new_n7354_), .ZN(new_n15414_));
  NAND2_X1   g15157(.A1(new_n1828_), .A2(new_n15414_), .ZN(new_n15415_));
  XOR2_X1    g15158(.A1(new_n15415_), .A2(new_n7343_), .Z(new_n15416_));
  XNOR2_X1   g15159(.A1(new_n15416_), .A2(new_n15411_), .ZN(new_n15417_));
  NOR2_X1    g15160(.A1(new_n15417_), .A2(new_n15410_), .ZN(new_n15418_));
  INV_X1     g15161(.I(new_n15411_), .ZN(new_n15419_));
  INV_X1     g15162(.I(new_n15416_), .ZN(new_n15420_));
  NOR2_X1    g15163(.A1(new_n15420_), .A2(new_n15419_), .ZN(new_n15421_));
  INV_X1     g15164(.I(new_n15421_), .ZN(new_n15422_));
  NOR2_X1    g15165(.A1(new_n15416_), .A2(new_n15411_), .ZN(new_n15423_));
  INV_X1     g15166(.I(new_n15423_), .ZN(new_n15424_));
  NAND2_X1   g15167(.A1(new_n15422_), .A2(new_n15424_), .ZN(new_n15425_));
  AOI21_X1   g15168(.A1(new_n15410_), .A2(new_n15425_), .B(new_n15418_), .ZN(new_n15426_));
  XNOR2_X1   g15169(.A1(new_n15426_), .A2(new_n15391_), .ZN(new_n15427_));
  NOR2_X1    g15170(.A1(new_n15427_), .A2(new_n15389_), .ZN(new_n15428_));
  INV_X1     g15171(.I(new_n15389_), .ZN(new_n15429_));
  NOR2_X1    g15172(.A1(new_n15426_), .A2(new_n15391_), .ZN(new_n15430_));
  INV_X1     g15173(.I(new_n15430_), .ZN(new_n15431_));
  NAND2_X1   g15174(.A1(new_n15426_), .A2(new_n15391_), .ZN(new_n15432_));
  AOI21_X1   g15175(.A1(new_n15431_), .A2(new_n15432_), .B(new_n15429_), .ZN(new_n15433_));
  NOR2_X1    g15176(.A1(new_n15428_), .A2(new_n15433_), .ZN(new_n15434_));
  AOI21_X1   g15177(.A1(new_n15108_), .A2(new_n15156_), .B(new_n15155_), .ZN(new_n15435_));
  OAI22_X1   g15178(.A1(new_n5786_), .A2(new_n2543_), .B1(new_n2405_), .B2(new_n5792_), .ZN(new_n15436_));
  NAND2_X1   g15179(.A1(new_n6745_), .A2(\b[29] ), .ZN(new_n15437_));
  AOI21_X1   g15180(.A1(new_n15437_), .A2(new_n15436_), .B(new_n5796_), .ZN(new_n15438_));
  NAND2_X1   g15181(.A1(new_n2546_), .A2(new_n15438_), .ZN(new_n15439_));
  XOR2_X1    g15182(.A1(new_n15439_), .A2(\a[53] ), .Z(new_n15440_));
  XNOR2_X1   g15183(.A1(new_n15435_), .A2(new_n15440_), .ZN(new_n15441_));
  NOR2_X1    g15184(.A1(new_n15441_), .A2(new_n15434_), .ZN(new_n15442_));
  NOR2_X1    g15185(.A1(new_n15435_), .A2(new_n15440_), .ZN(new_n15443_));
  INV_X1     g15186(.I(new_n15443_), .ZN(new_n15444_));
  NAND2_X1   g15187(.A1(new_n15435_), .A2(new_n15440_), .ZN(new_n15445_));
  NAND2_X1   g15188(.A1(new_n15444_), .A2(new_n15445_), .ZN(new_n15446_));
  AOI21_X1   g15189(.A1(new_n15434_), .A2(new_n15446_), .B(new_n15442_), .ZN(new_n15447_));
  NOR2_X1    g15190(.A1(new_n15167_), .A2(new_n15159_), .ZN(new_n15448_));
  NOR2_X1    g15191(.A1(new_n15448_), .A2(new_n15166_), .ZN(new_n15449_));
  NOR2_X1    g15192(.A1(new_n15447_), .A2(new_n15449_), .ZN(new_n15450_));
  INV_X1     g15193(.I(new_n15450_), .ZN(new_n15451_));
  NAND2_X1   g15194(.A1(new_n15447_), .A2(new_n15449_), .ZN(new_n15452_));
  AOI21_X1   g15195(.A1(new_n15451_), .A2(new_n15452_), .B(new_n15384_), .ZN(new_n15453_));
  INV_X1     g15196(.I(new_n15384_), .ZN(new_n15454_));
  XNOR2_X1   g15197(.A1(new_n15447_), .A2(new_n15449_), .ZN(new_n15455_));
  NOR2_X1    g15198(.A1(new_n15455_), .A2(new_n15454_), .ZN(new_n15456_));
  NOR2_X1    g15199(.A1(new_n15456_), .A2(new_n15453_), .ZN(new_n15457_));
  NOR2_X1    g15200(.A1(new_n15178_), .A2(new_n15106_), .ZN(new_n15458_));
  NOR2_X1    g15201(.A1(new_n15458_), .A2(new_n15176_), .ZN(new_n15459_));
  OAI22_X1   g15202(.A1(new_n4711_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n4706_), .ZN(new_n15460_));
  NAND2_X1   g15203(.A1(new_n5814_), .A2(\b[35] ), .ZN(new_n15461_));
  AOI21_X1   g15204(.A1(new_n15460_), .A2(new_n15461_), .B(new_n4714_), .ZN(new_n15462_));
  NAND2_X1   g15205(.A1(new_n3411_), .A2(new_n15462_), .ZN(new_n15463_));
  XOR2_X1    g15206(.A1(new_n15463_), .A2(\a[47] ), .Z(new_n15464_));
  XNOR2_X1   g15207(.A1(new_n15459_), .A2(new_n15464_), .ZN(new_n15465_));
  NOR2_X1    g15208(.A1(new_n15465_), .A2(new_n15457_), .ZN(new_n15466_));
  INV_X1     g15209(.I(new_n15457_), .ZN(new_n15467_));
  NOR2_X1    g15210(.A1(new_n15459_), .A2(new_n15464_), .ZN(new_n15468_));
  INV_X1     g15211(.I(new_n15468_), .ZN(new_n15469_));
  NAND2_X1   g15212(.A1(new_n15459_), .A2(new_n15464_), .ZN(new_n15470_));
  AOI21_X1   g15213(.A1(new_n15469_), .A2(new_n15470_), .B(new_n15467_), .ZN(new_n15471_));
  NOR2_X1    g15214(.A1(new_n15466_), .A2(new_n15471_), .ZN(new_n15472_));
  XNOR2_X1   g15215(.A1(new_n15472_), .A2(new_n15379_), .ZN(new_n15473_));
  NOR2_X1    g15216(.A1(new_n15472_), .A2(new_n15379_), .ZN(new_n15474_));
  NAND2_X1   g15217(.A1(new_n15472_), .A2(new_n15379_), .ZN(new_n15475_));
  INV_X1     g15218(.I(new_n15475_), .ZN(new_n15476_));
  OAI21_X1   g15219(.A1(new_n15476_), .A2(new_n15474_), .B(new_n15378_), .ZN(new_n15477_));
  OAI21_X1   g15220(.A1(new_n15378_), .A2(new_n15473_), .B(new_n15477_), .ZN(new_n15478_));
  OAI22_X1   g15221(.A1(new_n3736_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n3731_), .ZN(new_n15479_));
  NAND2_X1   g15222(.A1(new_n4730_), .A2(\b[41] ), .ZN(new_n15480_));
  AOI21_X1   g15223(.A1(new_n15479_), .A2(new_n15480_), .B(new_n3739_), .ZN(new_n15481_));
  NAND2_X1   g15224(.A1(new_n4320_), .A2(new_n15481_), .ZN(new_n15482_));
  XOR2_X1    g15225(.A1(new_n15482_), .A2(\a[41] ), .Z(new_n15483_));
  NOR2_X1    g15226(.A1(new_n15478_), .A2(new_n15483_), .ZN(new_n15484_));
  INV_X1     g15227(.I(new_n15484_), .ZN(new_n15485_));
  NAND2_X1   g15228(.A1(new_n15478_), .A2(new_n15483_), .ZN(new_n15486_));
  AOI21_X1   g15229(.A1(new_n15485_), .A2(new_n15486_), .B(new_n15373_), .ZN(new_n15487_));
  INV_X1     g15230(.I(new_n15373_), .ZN(new_n15488_));
  XNOR2_X1   g15231(.A1(new_n15478_), .A2(new_n15483_), .ZN(new_n15489_));
  NOR2_X1    g15232(.A1(new_n15489_), .A2(new_n15488_), .ZN(new_n15490_));
  NOR2_X1    g15233(.A1(new_n15490_), .A2(new_n15487_), .ZN(new_n15491_));
  INV_X1     g15234(.I(new_n15221_), .ZN(new_n15492_));
  AOI21_X1   g15235(.A1(new_n15217_), .A2(new_n15492_), .B(new_n15219_), .ZN(new_n15493_));
  NOR2_X1    g15236(.A1(new_n15491_), .A2(new_n15493_), .ZN(new_n15494_));
  NAND2_X1   g15237(.A1(new_n15491_), .A2(new_n15493_), .ZN(new_n15495_));
  INV_X1     g15238(.I(new_n15495_), .ZN(new_n15496_));
  NOR2_X1    g15239(.A1(new_n15496_), .A2(new_n15494_), .ZN(new_n15497_));
  XOR2_X1    g15240(.A1(new_n15491_), .A2(new_n15493_), .Z(new_n15498_));
  NAND2_X1   g15241(.A1(new_n15498_), .A2(new_n15371_), .ZN(new_n15499_));
  OAI21_X1   g15242(.A1(new_n15371_), .A2(new_n15497_), .B(new_n15499_), .ZN(new_n15500_));
  NAND2_X1   g15243(.A1(new_n15102_), .A2(new_n15234_), .ZN(new_n15501_));
  NAND2_X1   g15244(.A1(new_n15501_), .A2(new_n15233_), .ZN(new_n15502_));
  OAI22_X1   g15245(.A1(new_n2846_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n2841_), .ZN(new_n15503_));
  NAND2_X1   g15246(.A1(new_n3755_), .A2(\b[47] ), .ZN(new_n15504_));
  AOI21_X1   g15247(.A1(new_n15503_), .A2(new_n15504_), .B(new_n2849_), .ZN(new_n15505_));
  NAND2_X1   g15248(.A1(new_n5196_), .A2(new_n15505_), .ZN(new_n15506_));
  XOR2_X1    g15249(.A1(new_n15506_), .A2(\a[35] ), .Z(new_n15507_));
  INV_X1     g15250(.I(new_n15507_), .ZN(new_n15508_));
  NAND2_X1   g15251(.A1(new_n15502_), .A2(new_n15508_), .ZN(new_n15509_));
  INV_X1     g15252(.I(new_n15509_), .ZN(new_n15510_));
  NOR2_X1    g15253(.A1(new_n15502_), .A2(new_n15508_), .ZN(new_n15511_));
  OAI21_X1   g15254(.A1(new_n15510_), .A2(new_n15511_), .B(new_n15500_), .ZN(new_n15512_));
  XOR2_X1    g15255(.A1(new_n15502_), .A2(new_n15507_), .Z(new_n15513_));
  OAI21_X1   g15256(.A1(new_n15500_), .A2(new_n15513_), .B(new_n15512_), .ZN(new_n15514_));
  XOR2_X1    g15257(.A1(new_n15366_), .A2(new_n15514_), .Z(new_n15515_));
  INV_X1     g15258(.I(new_n15514_), .ZN(new_n15516_));
  NOR2_X1    g15259(.A1(new_n15366_), .A2(new_n15516_), .ZN(new_n15517_));
  NOR3_X1    g15260(.A1(new_n15365_), .A2(new_n15244_), .A3(new_n15514_), .ZN(new_n15518_));
  OAI21_X1   g15261(.A1(new_n15517_), .A2(new_n15518_), .B(new_n15364_), .ZN(new_n15519_));
  OAI21_X1   g15262(.A1(new_n15515_), .A2(new_n15364_), .B(new_n15519_), .ZN(new_n15520_));
  NAND2_X1   g15263(.A1(new_n15359_), .A2(new_n15520_), .ZN(new_n15521_));
  OR2_X2     g15264(.A1(new_n15359_), .A2(new_n15520_), .Z(new_n15522_));
  AOI21_X1   g15265(.A1(new_n15522_), .A2(new_n15521_), .B(new_n15357_), .ZN(new_n15523_));
  INV_X1     g15266(.I(new_n15357_), .ZN(new_n15524_));
  XNOR2_X1   g15267(.A1(new_n15359_), .A2(new_n15520_), .ZN(new_n15525_));
  NOR2_X1    g15268(.A1(new_n15525_), .A2(new_n15524_), .ZN(new_n15526_));
  NOR2_X1    g15269(.A1(new_n15526_), .A2(new_n15523_), .ZN(new_n15527_));
  XNOR2_X1   g15270(.A1(new_n15352_), .A2(new_n15527_), .ZN(new_n15528_));
  NOR2_X1    g15271(.A1(new_n15528_), .A2(new_n15350_), .ZN(new_n15529_));
  INV_X1     g15272(.I(new_n15350_), .ZN(new_n15530_));
  OAI22_X1   g15273(.A1(new_n15351_), .A2(new_n15264_), .B1(new_n15526_), .B2(new_n15523_), .ZN(new_n15531_));
  NAND2_X1   g15274(.A1(new_n15352_), .A2(new_n15527_), .ZN(new_n15532_));
  AOI21_X1   g15275(.A1(new_n15532_), .A2(new_n15531_), .B(new_n15530_), .ZN(new_n15533_));
  NOR2_X1    g15276(.A1(new_n15529_), .A2(new_n15533_), .ZN(new_n15534_));
  NOR2_X1    g15277(.A1(new_n15534_), .A2(new_n15345_), .ZN(new_n15535_));
  INV_X1     g15278(.I(new_n15535_), .ZN(new_n15536_));
  NAND2_X1   g15279(.A1(new_n15534_), .A2(new_n15345_), .ZN(new_n15537_));
  AOI21_X1   g15280(.A1(new_n15536_), .A2(new_n15537_), .B(new_n15343_), .ZN(new_n15538_));
  INV_X1     g15281(.I(new_n15343_), .ZN(new_n15539_));
  NOR2_X1    g15282(.A1(new_n15534_), .A2(new_n15344_), .ZN(new_n15540_));
  INV_X1     g15283(.I(new_n15540_), .ZN(new_n15541_));
  NAND2_X1   g15284(.A1(new_n15534_), .A2(new_n15344_), .ZN(new_n15542_));
  AOI21_X1   g15285(.A1(new_n15541_), .A2(new_n15542_), .B(new_n15539_), .ZN(new_n15543_));
  OR2_X2     g15286(.A1(new_n15538_), .A2(new_n15543_), .Z(new_n15544_));
  AOI21_X1   g15287(.A1(new_n15083_), .A2(new_n15303_), .B(new_n15287_), .ZN(new_n15545_));
  NOR2_X1    g15288(.A1(new_n15544_), .A2(new_n15545_), .ZN(new_n15546_));
  NOR2_X1    g15289(.A1(new_n15538_), .A2(new_n15543_), .ZN(new_n15547_));
  INV_X1     g15290(.I(new_n15545_), .ZN(new_n15548_));
  NOR2_X1    g15291(.A1(new_n15547_), .A2(new_n15548_), .ZN(new_n15549_));
  OAI21_X1   g15292(.A1(new_n15546_), .A2(new_n15549_), .B(new_n15338_), .ZN(new_n15550_));
  NOR2_X1    g15293(.A1(new_n15547_), .A2(new_n15545_), .ZN(new_n15551_));
  NAND2_X1   g15294(.A1(new_n15547_), .A2(new_n15545_), .ZN(new_n15552_));
  INV_X1     g15295(.I(new_n15552_), .ZN(new_n15553_));
  OAI21_X1   g15296(.A1(new_n15553_), .A2(new_n15551_), .B(new_n15337_), .ZN(new_n15554_));
  NAND2_X1   g15297(.A1(new_n15554_), .A2(new_n15550_), .ZN(new_n15555_));
  NOR2_X1    g15298(.A1(new_n15316_), .A2(new_n15313_), .ZN(new_n15556_));
  AOI21_X1   g15299(.A1(new_n15330_), .A2(new_n15556_), .B(new_n15555_), .ZN(new_n15557_));
  AOI21_X1   g15300(.A1(new_n14794_), .A2(new_n15058_), .B(new_n15054_), .ZN(new_n15558_));
  OR2_X2     g15301(.A1(new_n15546_), .A2(new_n15549_), .Z(new_n15559_));
  INV_X1     g15302(.I(new_n15551_), .ZN(new_n15560_));
  AOI21_X1   g15303(.A1(new_n15560_), .A2(new_n15552_), .B(new_n15338_), .ZN(new_n15561_));
  AOI21_X1   g15304(.A1(new_n15559_), .A2(new_n15338_), .B(new_n15561_), .ZN(new_n15562_));
  XOR2_X1    g15305(.A1(new_n15315_), .A2(new_n15065_), .Z(new_n15563_));
  NOR3_X1    g15306(.A1(new_n15558_), .A2(new_n15562_), .A3(new_n15563_), .ZN(new_n15564_));
  OAI21_X1   g15307(.A1(new_n15564_), .A2(new_n15557_), .B(new_n15333_), .ZN(new_n15565_));
  INV_X1     g15308(.I(new_n15333_), .ZN(new_n15566_));
  OAI21_X1   g15309(.A1(new_n15558_), .A2(new_n15563_), .B(new_n15562_), .ZN(new_n15567_));
  NAND3_X1   g15310(.A1(new_n15330_), .A2(new_n15555_), .A3(new_n15556_), .ZN(new_n15568_));
  NAND3_X1   g15311(.A1(new_n15567_), .A2(new_n15568_), .A3(new_n15566_), .ZN(new_n15569_));
  NAND2_X1   g15312(.A1(new_n15565_), .A2(new_n15569_), .ZN(\f[82] ));
  NAND2_X1   g15313(.A1(new_n15330_), .A2(new_n15556_), .ZN(new_n15571_));
  AOI22_X1   g15314(.A1(new_n15567_), .A2(new_n15568_), .B1(new_n15571_), .B2(new_n15566_), .ZN(new_n15572_));
  AOI21_X1   g15315(.A1(new_n15338_), .A2(new_n15552_), .B(new_n15551_), .ZN(new_n15573_));
  INV_X1     g15316(.I(new_n15573_), .ZN(new_n15574_));
  INV_X1     g15317(.I(new_n15537_), .ZN(new_n15575_));
  AOI21_X1   g15318(.A1(new_n15539_), .A2(new_n15536_), .B(new_n15575_), .ZN(new_n15576_));
  INV_X1     g15319(.I(new_n15576_), .ZN(new_n15577_));
  OAI22_X1   g15320(.A1(new_n9595_), .A2(new_n1171_), .B1(new_n8956_), .B2(new_n1255_), .ZN(new_n15578_));
  OAI22_X1   g15321(.A1(new_n1760_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n1755_), .ZN(new_n15579_));
  NAND2_X1   g15322(.A1(new_n2470_), .A2(\b[57] ), .ZN(new_n15580_));
  AOI21_X1   g15323(.A1(new_n15579_), .A2(new_n15580_), .B(new_n1763_), .ZN(new_n15581_));
  NAND2_X1   g15324(.A1(new_n7895_), .A2(new_n15581_), .ZN(new_n15582_));
  XOR2_X1    g15325(.A1(new_n15582_), .A2(\a[26] ), .Z(new_n15583_));
  OAI22_X1   g15326(.A1(new_n2084_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n2079_), .ZN(new_n15584_));
  NAND2_X1   g15327(.A1(new_n2864_), .A2(\b[54] ), .ZN(new_n15585_));
  AOI21_X1   g15328(.A1(new_n15584_), .A2(new_n15585_), .B(new_n2087_), .ZN(new_n15586_));
  NAND2_X1   g15329(.A1(new_n6994_), .A2(new_n15586_), .ZN(new_n15587_));
  XOR2_X1    g15330(.A1(new_n15587_), .A2(\a[29] ), .Z(new_n15588_));
  NOR2_X1    g15331(.A1(new_n15518_), .A2(new_n15364_), .ZN(new_n15589_));
  NOR2_X1    g15332(.A1(new_n15589_), .A2(new_n15517_), .ZN(new_n15590_));
  OAI22_X1   g15333(.A1(new_n2452_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n2447_), .ZN(new_n15591_));
  NAND2_X1   g15334(.A1(new_n3312_), .A2(\b[51] ), .ZN(new_n15592_));
  AOI21_X1   g15335(.A1(new_n15591_), .A2(new_n15592_), .B(new_n2455_), .ZN(new_n15593_));
  NAND2_X1   g15336(.A1(new_n6219_), .A2(new_n15593_), .ZN(new_n15594_));
  XOR2_X1    g15337(.A1(new_n15594_), .A2(\a[32] ), .Z(new_n15595_));
  OAI22_X1   g15338(.A1(new_n2846_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n2841_), .ZN(new_n15596_));
  NAND2_X1   g15339(.A1(new_n3755_), .A2(\b[48] ), .ZN(new_n15597_));
  AOI21_X1   g15340(.A1(new_n15596_), .A2(new_n15597_), .B(new_n2849_), .ZN(new_n15598_));
  NAND2_X1   g15341(.A1(new_n5537_), .A2(new_n15598_), .ZN(new_n15599_));
  XOR2_X1    g15342(.A1(new_n15599_), .A2(\a[35] ), .Z(new_n15600_));
  OAI22_X1   g15343(.A1(new_n3736_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n3731_), .ZN(new_n15601_));
  NAND2_X1   g15344(.A1(new_n4730_), .A2(\b[42] ), .ZN(new_n15602_));
  AOI21_X1   g15345(.A1(new_n15601_), .A2(new_n15602_), .B(new_n3739_), .ZN(new_n15603_));
  NAND2_X1   g15346(.A1(new_n4500_), .A2(new_n15603_), .ZN(new_n15604_));
  XOR2_X1    g15347(.A1(new_n15604_), .A2(\a[41] ), .Z(new_n15605_));
  OAI21_X1   g15348(.A1(new_n15378_), .A2(new_n15474_), .B(new_n15475_), .ZN(new_n15606_));
  OAI22_X1   g15349(.A1(new_n4208_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n4203_), .ZN(new_n15607_));
  NAND2_X1   g15350(.A1(new_n5244_), .A2(\b[39] ), .ZN(new_n15608_));
  AOI21_X1   g15351(.A1(new_n15607_), .A2(new_n15608_), .B(new_n4211_), .ZN(new_n15609_));
  NAND2_X1   g15352(.A1(new_n3996_), .A2(new_n15609_), .ZN(new_n15610_));
  XOR2_X1    g15353(.A1(new_n15610_), .A2(\a[44] ), .Z(new_n15611_));
  OAI22_X1   g15354(.A1(new_n4711_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n4706_), .ZN(new_n15612_));
  NAND2_X1   g15355(.A1(new_n5814_), .A2(\b[36] ), .ZN(new_n15613_));
  AOI21_X1   g15356(.A1(new_n15612_), .A2(new_n15613_), .B(new_n4714_), .ZN(new_n15614_));
  NAND2_X1   g15357(.A1(new_n3565_), .A2(new_n15614_), .ZN(new_n15615_));
  XOR2_X1    g15358(.A1(new_n15615_), .A2(\a[47] ), .Z(new_n15616_));
  AOI21_X1   g15359(.A1(new_n15454_), .A2(new_n15452_), .B(new_n15450_), .ZN(new_n15617_));
  INV_X1     g15360(.I(new_n15617_), .ZN(new_n15618_));
  OAI22_X1   g15361(.A1(new_n5228_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n5225_), .ZN(new_n15619_));
  NAND2_X1   g15362(.A1(new_n5387_), .A2(\b[33] ), .ZN(new_n15620_));
  AOI21_X1   g15363(.A1(new_n15619_), .A2(new_n15620_), .B(new_n5231_), .ZN(new_n15621_));
  NAND2_X1   g15364(.A1(new_n3101_), .A2(new_n15621_), .ZN(new_n15622_));
  XOR2_X1    g15365(.A1(new_n15622_), .A2(\a[50] ), .Z(new_n15623_));
  OAI22_X1   g15366(.A1(new_n5786_), .A2(new_n2660_), .B1(new_n2543_), .B2(new_n5792_), .ZN(new_n15624_));
  NAND2_X1   g15367(.A1(new_n6745_), .A2(\b[30] ), .ZN(new_n15625_));
  AOI21_X1   g15368(.A1(new_n15625_), .A2(new_n15624_), .B(new_n5796_), .ZN(new_n15626_));
  NAND2_X1   g15369(.A1(new_n2659_), .A2(new_n15626_), .ZN(new_n15627_));
  XOR2_X1    g15370(.A1(new_n15627_), .A2(\a[53] ), .Z(new_n15628_));
  OAI22_X1   g15371(.A1(new_n1927_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1825_), .ZN(new_n15629_));
  NAND2_X1   g15372(.A1(new_n8628_), .A2(\b[24] ), .ZN(new_n15630_));
  AOI21_X1   g15373(.A1(new_n15630_), .A2(new_n15629_), .B(new_n7354_), .ZN(new_n15631_));
  NAND2_X1   g15374(.A1(new_n1926_), .A2(new_n15631_), .ZN(new_n15632_));
  XOR2_X1    g15375(.A1(new_n15632_), .A2(\a[59] ), .Z(new_n15633_));
  INV_X1     g15376(.I(new_n15408_), .ZN(new_n15634_));
  AOI21_X1   g15377(.A1(new_n15396_), .A2(new_n15407_), .B(new_n15634_), .ZN(new_n15635_));
  OAI22_X1   g15378(.A1(new_n1601_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1518_), .ZN(new_n15636_));
  NAND2_X1   g15379(.A1(new_n9644_), .A2(\b[21] ), .ZN(new_n15637_));
  AOI21_X1   g15380(.A1(new_n15637_), .A2(new_n15636_), .B(new_n8321_), .ZN(new_n15638_));
  NAND2_X1   g15381(.A1(new_n1604_), .A2(new_n15638_), .ZN(new_n15639_));
  XOR2_X1    g15382(.A1(new_n15639_), .A2(\a[62] ), .Z(new_n15640_));
  NOR3_X1    g15383(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n1222_), .ZN(new_n15641_));
  NOR2_X1    g15384(.A1(new_n9364_), .A2(new_n1222_), .ZN(new_n15642_));
  NOR3_X1    g15385(.A1(new_n15642_), .A2(new_n1305_), .A3(new_n8985_), .ZN(new_n15643_));
  NOR2_X1    g15386(.A1(new_n15643_), .A2(new_n15641_), .ZN(new_n15644_));
  XOR2_X1    g15387(.A1(new_n15402_), .A2(new_n15644_), .Z(new_n15645_));
  NOR2_X1    g15388(.A1(new_n15640_), .A2(new_n15645_), .ZN(new_n15646_));
  INV_X1     g15389(.I(new_n15640_), .ZN(new_n15647_));
  NOR2_X1    g15390(.A1(new_n15403_), .A2(new_n15644_), .ZN(new_n15648_));
  INV_X1     g15391(.I(new_n15644_), .ZN(new_n15649_));
  NOR2_X1    g15392(.A1(new_n15649_), .A2(new_n15402_), .ZN(new_n15650_));
  NOR2_X1    g15393(.A1(new_n15648_), .A2(new_n15650_), .ZN(new_n15651_));
  NOR2_X1    g15394(.A1(new_n15647_), .A2(new_n15651_), .ZN(new_n15652_));
  NOR2_X1    g15395(.A1(new_n15652_), .A2(new_n15646_), .ZN(new_n15653_));
  XOR2_X1    g15396(.A1(new_n15653_), .A2(new_n15635_), .Z(new_n15654_));
  INV_X1     g15397(.I(new_n15635_), .ZN(new_n15655_));
  NOR2_X1    g15398(.A1(new_n15653_), .A2(new_n15655_), .ZN(new_n15656_));
  NAND2_X1   g15399(.A1(new_n15653_), .A2(new_n15655_), .ZN(new_n15657_));
  INV_X1     g15400(.I(new_n15657_), .ZN(new_n15658_));
  OAI21_X1   g15401(.A1(new_n15658_), .A2(new_n15656_), .B(new_n15633_), .ZN(new_n15659_));
  OAI21_X1   g15402(.A1(new_n15633_), .A2(new_n15654_), .B(new_n15659_), .ZN(new_n15660_));
  INV_X1     g15403(.I(new_n15660_), .ZN(new_n15661_));
  OAI22_X1   g15404(.A1(new_n6721_), .A2(new_n2175_), .B1(new_n6723_), .B2(new_n2272_), .ZN(new_n15662_));
  NAND2_X1   g15405(.A1(new_n7617_), .A2(\b[27] ), .ZN(new_n15663_));
  AOI21_X1   g15406(.A1(new_n15663_), .A2(new_n15662_), .B(new_n6731_), .ZN(new_n15664_));
  NAND2_X1   g15407(.A1(new_n2276_), .A2(new_n15664_), .ZN(new_n15665_));
  XOR2_X1    g15408(.A1(new_n15665_), .A2(\a[56] ), .Z(new_n15666_));
  AOI21_X1   g15409(.A1(new_n15410_), .A2(new_n15424_), .B(new_n15421_), .ZN(new_n15667_));
  XNOR2_X1   g15410(.A1(new_n15666_), .A2(new_n15667_), .ZN(new_n15668_));
  NOR2_X1    g15411(.A1(new_n15668_), .A2(new_n15661_), .ZN(new_n15669_));
  NOR2_X1    g15412(.A1(new_n15666_), .A2(new_n15667_), .ZN(new_n15670_));
  INV_X1     g15413(.I(new_n15670_), .ZN(new_n15671_));
  NAND2_X1   g15414(.A1(new_n15666_), .A2(new_n15667_), .ZN(new_n15672_));
  AOI21_X1   g15415(.A1(new_n15671_), .A2(new_n15672_), .B(new_n15660_), .ZN(new_n15673_));
  NAND2_X1   g15416(.A1(new_n15432_), .A2(new_n15429_), .ZN(new_n15674_));
  NAND2_X1   g15417(.A1(new_n15674_), .A2(new_n15431_), .ZN(new_n15675_));
  OAI21_X1   g15418(.A1(new_n15669_), .A2(new_n15673_), .B(new_n15675_), .ZN(new_n15676_));
  NOR2_X1    g15419(.A1(new_n15669_), .A2(new_n15673_), .ZN(new_n15677_));
  NAND3_X1   g15420(.A1(new_n15677_), .A2(new_n15431_), .A3(new_n15674_), .ZN(new_n15678_));
  AOI21_X1   g15421(.A1(new_n15678_), .A2(new_n15676_), .B(new_n15628_), .ZN(new_n15679_));
  INV_X1     g15422(.I(new_n15628_), .ZN(new_n15680_));
  XOR2_X1    g15423(.A1(new_n15677_), .A2(new_n15675_), .Z(new_n15681_));
  NOR2_X1    g15424(.A1(new_n15681_), .A2(new_n15680_), .ZN(new_n15682_));
  NOR2_X1    g15425(.A1(new_n15682_), .A2(new_n15679_), .ZN(new_n15683_));
  AOI21_X1   g15426(.A1(new_n15434_), .A2(new_n15445_), .B(new_n15443_), .ZN(new_n15684_));
  INV_X1     g15427(.I(new_n15684_), .ZN(new_n15685_));
  XOR2_X1    g15428(.A1(new_n15683_), .A2(new_n15685_), .Z(new_n15686_));
  NOR2_X1    g15429(.A1(new_n15683_), .A2(new_n15684_), .ZN(new_n15687_));
  NOR3_X1    g15430(.A1(new_n15682_), .A2(new_n15679_), .A3(new_n15685_), .ZN(new_n15688_));
  OAI21_X1   g15431(.A1(new_n15687_), .A2(new_n15688_), .B(new_n15623_), .ZN(new_n15689_));
  OAI21_X1   g15432(.A1(new_n15686_), .A2(new_n15623_), .B(new_n15689_), .ZN(new_n15690_));
  XOR2_X1    g15433(.A1(new_n15690_), .A2(new_n15618_), .Z(new_n15691_));
  AND2_X2    g15434(.A1(new_n15690_), .A2(new_n15617_), .Z(new_n15692_));
  NOR2_X1    g15435(.A1(new_n15690_), .A2(new_n15617_), .ZN(new_n15693_));
  OAI21_X1   g15436(.A1(new_n15692_), .A2(new_n15693_), .B(new_n15616_), .ZN(new_n15694_));
  OAI21_X1   g15437(.A1(new_n15616_), .A2(new_n15691_), .B(new_n15694_), .ZN(new_n15695_));
  AOI21_X1   g15438(.A1(new_n15467_), .A2(new_n15470_), .B(new_n15468_), .ZN(new_n15696_));
  XNOR2_X1   g15439(.A1(new_n15695_), .A2(new_n15696_), .ZN(new_n15697_));
  NOR2_X1    g15440(.A1(new_n15697_), .A2(new_n15611_), .ZN(new_n15698_));
  INV_X1     g15441(.I(new_n15611_), .ZN(new_n15699_));
  NOR2_X1    g15442(.A1(new_n15695_), .A2(new_n15696_), .ZN(new_n15700_));
  INV_X1     g15443(.I(new_n15700_), .ZN(new_n15701_));
  NAND2_X1   g15444(.A1(new_n15695_), .A2(new_n15696_), .ZN(new_n15702_));
  AOI21_X1   g15445(.A1(new_n15701_), .A2(new_n15702_), .B(new_n15699_), .ZN(new_n15703_));
  NOR2_X1    g15446(.A1(new_n15698_), .A2(new_n15703_), .ZN(new_n15704_));
  XNOR2_X1   g15447(.A1(new_n15704_), .A2(new_n15606_), .ZN(new_n15705_));
  NOR2_X1    g15448(.A1(new_n15705_), .A2(new_n15605_), .ZN(new_n15706_));
  INV_X1     g15449(.I(new_n15605_), .ZN(new_n15707_));
  NOR2_X1    g15450(.A1(new_n15704_), .A2(new_n15606_), .ZN(new_n15708_));
  INV_X1     g15451(.I(new_n15708_), .ZN(new_n15709_));
  NAND2_X1   g15452(.A1(new_n15704_), .A2(new_n15606_), .ZN(new_n15710_));
  AOI21_X1   g15453(.A1(new_n15709_), .A2(new_n15710_), .B(new_n15707_), .ZN(new_n15711_));
  NOR2_X1    g15454(.A1(new_n15706_), .A2(new_n15711_), .ZN(new_n15712_));
  OAI22_X1   g15455(.A1(new_n3298_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n3293_), .ZN(new_n15713_));
  NAND2_X1   g15456(.A1(new_n4227_), .A2(\b[45] ), .ZN(new_n15714_));
  AOI21_X1   g15457(.A1(new_n15713_), .A2(new_n15714_), .B(new_n3301_), .ZN(new_n15715_));
  NAND2_X1   g15458(.A1(new_n5004_), .A2(new_n15715_), .ZN(new_n15716_));
  XOR2_X1    g15459(.A1(new_n15716_), .A2(\a[38] ), .Z(new_n15717_));
  NAND2_X1   g15460(.A1(new_n15486_), .A2(new_n15488_), .ZN(new_n15718_));
  NAND2_X1   g15461(.A1(new_n15718_), .A2(new_n15485_), .ZN(new_n15719_));
  XOR2_X1    g15462(.A1(new_n15719_), .A2(new_n15717_), .Z(new_n15720_));
  NOR2_X1    g15463(.A1(new_n15720_), .A2(new_n15712_), .ZN(new_n15721_));
  INV_X1     g15464(.I(new_n15719_), .ZN(new_n15722_));
  NOR2_X1    g15465(.A1(new_n15722_), .A2(new_n15717_), .ZN(new_n15723_));
  INV_X1     g15466(.I(new_n15723_), .ZN(new_n15724_));
  NAND2_X1   g15467(.A1(new_n15722_), .A2(new_n15717_), .ZN(new_n15725_));
  NAND2_X1   g15468(.A1(new_n15724_), .A2(new_n15725_), .ZN(new_n15726_));
  AOI21_X1   g15469(.A1(new_n15712_), .A2(new_n15726_), .B(new_n15721_), .ZN(new_n15727_));
  NOR2_X1    g15470(.A1(new_n15496_), .A2(new_n15371_), .ZN(new_n15728_));
  NOR2_X1    g15471(.A1(new_n15728_), .A2(new_n15494_), .ZN(new_n15729_));
  XNOR2_X1   g15472(.A1(new_n15729_), .A2(new_n15727_), .ZN(new_n15730_));
  NOR2_X1    g15473(.A1(new_n15729_), .A2(new_n15727_), .ZN(new_n15731_));
  NAND2_X1   g15474(.A1(new_n15729_), .A2(new_n15727_), .ZN(new_n15732_));
  INV_X1     g15475(.I(new_n15732_), .ZN(new_n15733_));
  OAI21_X1   g15476(.A1(new_n15733_), .A2(new_n15731_), .B(new_n15600_), .ZN(new_n15734_));
  OAI21_X1   g15477(.A1(new_n15600_), .A2(new_n15730_), .B(new_n15734_), .ZN(new_n15735_));
  INV_X1     g15478(.I(new_n15511_), .ZN(new_n15736_));
  AOI21_X1   g15479(.A1(new_n15500_), .A2(new_n15736_), .B(new_n15510_), .ZN(new_n15737_));
  NOR2_X1    g15480(.A1(new_n15735_), .A2(new_n15737_), .ZN(new_n15738_));
  INV_X1     g15481(.I(new_n15738_), .ZN(new_n15739_));
  NAND2_X1   g15482(.A1(new_n15735_), .A2(new_n15737_), .ZN(new_n15740_));
  AOI21_X1   g15483(.A1(new_n15739_), .A2(new_n15740_), .B(new_n15595_), .ZN(new_n15741_));
  INV_X1     g15484(.I(new_n15595_), .ZN(new_n15742_));
  XNOR2_X1   g15485(.A1(new_n15735_), .A2(new_n15737_), .ZN(new_n15743_));
  NOR2_X1    g15486(.A1(new_n15743_), .A2(new_n15742_), .ZN(new_n15744_));
  NOR2_X1    g15487(.A1(new_n15744_), .A2(new_n15741_), .ZN(new_n15745_));
  NOR2_X1    g15488(.A1(new_n15745_), .A2(new_n15590_), .ZN(new_n15746_));
  INV_X1     g15489(.I(new_n15746_), .ZN(new_n15747_));
  NAND2_X1   g15490(.A1(new_n15745_), .A2(new_n15590_), .ZN(new_n15748_));
  AOI21_X1   g15491(.A1(new_n15747_), .A2(new_n15748_), .B(new_n15588_), .ZN(new_n15749_));
  INV_X1     g15492(.I(new_n15588_), .ZN(new_n15750_));
  XNOR2_X1   g15493(.A1(new_n15745_), .A2(new_n15590_), .ZN(new_n15751_));
  NOR2_X1    g15494(.A1(new_n15751_), .A2(new_n15750_), .ZN(new_n15752_));
  NOR2_X1    g15495(.A1(new_n15752_), .A2(new_n15749_), .ZN(new_n15753_));
  NOR2_X1    g15496(.A1(new_n15359_), .A2(new_n15520_), .ZN(new_n15754_));
  AOI21_X1   g15497(.A1(new_n15524_), .A2(new_n15521_), .B(new_n15754_), .ZN(new_n15755_));
  NOR2_X1    g15498(.A1(new_n15753_), .A2(new_n15755_), .ZN(new_n15756_));
  INV_X1     g15499(.I(new_n15756_), .ZN(new_n15757_));
  NAND2_X1   g15500(.A1(new_n15753_), .A2(new_n15755_), .ZN(new_n15758_));
  AOI21_X1   g15501(.A1(new_n15757_), .A2(new_n15758_), .B(new_n15583_), .ZN(new_n15759_));
  INV_X1     g15502(.I(new_n15583_), .ZN(new_n15760_));
  XNOR2_X1   g15503(.A1(new_n15753_), .A2(new_n15755_), .ZN(new_n15761_));
  NOR2_X1    g15504(.A1(new_n15761_), .A2(new_n15760_), .ZN(new_n15762_));
  NOR2_X1    g15505(.A1(new_n15762_), .A2(new_n15759_), .ZN(new_n15763_));
  INV_X1     g15506(.I(new_n8935_), .ZN(new_n15764_));
  AOI22_X1   g15507(.A1(\b[62] ), .A2(new_n1443_), .B1(new_n1947_), .B2(\b[61] ), .ZN(new_n15765_));
  AOI21_X1   g15508(.A1(\b[60] ), .A2(new_n2098_), .B(new_n15765_), .ZN(new_n15766_));
  OAI21_X1   g15509(.A1(new_n15764_), .A2(new_n1447_), .B(new_n15766_), .ZN(new_n15767_));
  NAND2_X1   g15510(.A1(new_n15532_), .A2(new_n15530_), .ZN(new_n15768_));
  NAND2_X1   g15511(.A1(new_n15768_), .A2(new_n15531_), .ZN(new_n15769_));
  XOR2_X1    g15512(.A1(new_n15769_), .A2(new_n15767_), .Z(new_n15770_));
  XOR2_X1    g15513(.A1(new_n15770_), .A2(\a[23] ), .Z(new_n15771_));
  XOR2_X1    g15514(.A1(new_n15771_), .A2(new_n15763_), .Z(new_n15772_));
  XOR2_X1    g15515(.A1(new_n15772_), .A2(new_n15578_), .Z(new_n15773_));
  NAND2_X1   g15516(.A1(new_n15773_), .A2(new_n1158_), .ZN(new_n15774_));
  XNOR2_X1   g15517(.A1(new_n15772_), .A2(new_n15578_), .ZN(new_n15775_));
  NAND2_X1   g15518(.A1(new_n15775_), .A2(\a[20] ), .ZN(new_n15776_));
  AOI21_X1   g15519(.A1(new_n15776_), .A2(new_n15774_), .B(new_n15577_), .ZN(new_n15777_));
  AND3_X2    g15520(.A1(new_n15776_), .A2(new_n15577_), .A3(new_n15774_), .Z(new_n15778_));
  NOR2_X1    g15521(.A1(new_n15778_), .A2(new_n15777_), .ZN(new_n15779_));
  XOR2_X1    g15522(.A1(new_n15779_), .A2(new_n15574_), .Z(new_n15780_));
  NAND2_X1   g15523(.A1(new_n15780_), .A2(new_n15572_), .ZN(new_n15781_));
  XOR2_X1    g15524(.A1(new_n15779_), .A2(new_n15574_), .Z(new_n15782_));
  OAI21_X1   g15525(.A1(new_n15572_), .A2(new_n15782_), .B(new_n15781_), .ZN(\f[83] ));
  INV_X1     g15526(.I(new_n15769_), .ZN(new_n15784_));
  NOR2_X1    g15527(.A1(new_n15784_), .A2(new_n15763_), .ZN(new_n15785_));
  NAND2_X1   g15528(.A1(new_n15784_), .A2(new_n15763_), .ZN(new_n15786_));
  XOR2_X1    g15529(.A1(new_n15767_), .A2(\a[23] ), .Z(new_n15787_));
  INV_X1     g15530(.I(new_n15787_), .ZN(new_n15788_));
  AOI21_X1   g15531(.A1(new_n15786_), .A2(new_n15788_), .B(new_n15785_), .ZN(new_n15789_));
  INV_X1     g15532(.I(new_n15789_), .ZN(new_n15790_));
  OAI22_X1   g15533(.A1(new_n1444_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n1439_), .ZN(new_n15791_));
  NAND2_X1   g15534(.A1(new_n2098_), .A2(\b[61] ), .ZN(new_n15792_));
  AOI21_X1   g15535(.A1(new_n15791_), .A2(new_n15792_), .B(new_n1447_), .ZN(new_n15793_));
  NAND2_X1   g15536(.A1(new_n8963_), .A2(new_n15793_), .ZN(new_n15794_));
  XOR2_X1    g15537(.A1(new_n15794_), .A2(\a[23] ), .Z(new_n15795_));
  INV_X1     g15538(.I(new_n15795_), .ZN(new_n15796_));
  OAI22_X1   g15539(.A1(new_n1760_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n1755_), .ZN(new_n15797_));
  NAND2_X1   g15540(.A1(new_n2470_), .A2(\b[58] ), .ZN(new_n15798_));
  AOI21_X1   g15541(.A1(new_n15797_), .A2(new_n15798_), .B(new_n1763_), .ZN(new_n15799_));
  NAND2_X1   g15542(.A1(new_n7929_), .A2(new_n15799_), .ZN(new_n15800_));
  XOR2_X1    g15543(.A1(new_n15800_), .A2(\a[26] ), .Z(new_n15801_));
  INV_X1     g15544(.I(new_n15801_), .ZN(new_n15802_));
  NAND2_X1   g15545(.A1(new_n15758_), .A2(new_n15760_), .ZN(new_n15803_));
  NAND2_X1   g15546(.A1(new_n15803_), .A2(new_n15757_), .ZN(new_n15804_));
  AOI21_X1   g15547(.A1(new_n15750_), .A2(new_n15748_), .B(new_n15746_), .ZN(new_n15805_));
  INV_X1     g15548(.I(new_n15805_), .ZN(new_n15806_));
  OAI22_X1   g15549(.A1(new_n2084_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n2079_), .ZN(new_n15807_));
  NAND2_X1   g15550(.A1(new_n2864_), .A2(\b[55] ), .ZN(new_n15808_));
  AOI21_X1   g15551(.A1(new_n15807_), .A2(new_n15808_), .B(new_n2087_), .ZN(new_n15809_));
  NAND2_X1   g15552(.A1(new_n7308_), .A2(new_n15809_), .ZN(new_n15810_));
  XOR2_X1    g15553(.A1(new_n15810_), .A2(\a[29] ), .Z(new_n15811_));
  OAI22_X1   g15554(.A1(new_n2452_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n2447_), .ZN(new_n15812_));
  NAND2_X1   g15555(.A1(new_n3312_), .A2(\b[52] ), .ZN(new_n15813_));
  AOI21_X1   g15556(.A1(new_n15812_), .A2(new_n15813_), .B(new_n2455_), .ZN(new_n15814_));
  NAND2_X1   g15557(.A1(new_n6237_), .A2(new_n15814_), .ZN(new_n15815_));
  XOR2_X1    g15558(.A1(new_n15815_), .A2(\a[32] ), .Z(new_n15816_));
  INV_X1     g15559(.I(new_n15816_), .ZN(new_n15817_));
  NAND2_X1   g15560(.A1(new_n15740_), .A2(new_n15742_), .ZN(new_n15818_));
  NAND2_X1   g15561(.A1(new_n15818_), .A2(new_n15739_), .ZN(new_n15819_));
  NOR2_X1    g15562(.A1(new_n15733_), .A2(new_n15600_), .ZN(new_n15820_));
  NOR2_X1    g15563(.A1(new_n15820_), .A2(new_n15731_), .ZN(new_n15821_));
  INV_X1     g15564(.I(new_n15821_), .ZN(new_n15822_));
  OAI21_X1   g15565(.A1(new_n15605_), .A2(new_n15708_), .B(new_n15710_), .ZN(new_n15823_));
  INV_X1     g15566(.I(new_n15823_), .ZN(new_n15824_));
  NOR2_X1    g15567(.A1(new_n15692_), .A2(new_n15616_), .ZN(new_n15825_));
  NOR2_X1    g15568(.A1(new_n15825_), .A2(new_n15693_), .ZN(new_n15826_));
  INV_X1     g15569(.I(new_n15826_), .ZN(new_n15827_));
  NOR2_X1    g15570(.A1(new_n15688_), .A2(new_n15623_), .ZN(new_n15828_));
  NOR2_X1    g15571(.A1(new_n15828_), .A2(new_n15687_), .ZN(new_n15829_));
  NAND2_X1   g15572(.A1(new_n15678_), .A2(new_n15680_), .ZN(new_n15830_));
  AND2_X2    g15573(.A1(new_n15830_), .A2(new_n15676_), .Z(new_n15831_));
  OAI21_X1   g15574(.A1(new_n15633_), .A2(new_n15656_), .B(new_n15657_), .ZN(new_n15832_));
  INV_X1     g15575(.I(new_n15832_), .ZN(new_n15833_));
  OAI22_X1   g15576(.A1(new_n1709_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1601_), .ZN(new_n15834_));
  NAND2_X1   g15577(.A1(new_n9644_), .A2(\b[22] ), .ZN(new_n15835_));
  AOI21_X1   g15578(.A1(new_n15835_), .A2(new_n15834_), .B(new_n8321_), .ZN(new_n15836_));
  NAND2_X1   g15579(.A1(new_n1708_), .A2(new_n15836_), .ZN(new_n15837_));
  XOR2_X1    g15580(.A1(new_n15837_), .A2(\a[62] ), .Z(new_n15838_));
  NOR2_X1    g15581(.A1(new_n15640_), .A2(new_n15648_), .ZN(new_n15839_));
  NOR2_X1    g15582(.A1(new_n15839_), .A2(new_n15650_), .ZN(new_n15840_));
  NOR2_X1    g15583(.A1(new_n8985_), .A2(new_n1393_), .ZN(new_n15841_));
  NOR2_X1    g15584(.A1(new_n9364_), .A2(new_n1305_), .ZN(new_n15842_));
  XNOR2_X1   g15585(.A1(new_n15841_), .A2(new_n15842_), .ZN(new_n15843_));
  XOR2_X1    g15586(.A1(new_n15843_), .A2(\a[20] ), .Z(new_n15844_));
  NOR2_X1    g15587(.A1(new_n15844_), .A2(new_n15644_), .ZN(new_n15845_));
  NOR2_X1    g15588(.A1(new_n15843_), .A2(new_n1158_), .ZN(new_n15846_));
  INV_X1     g15589(.I(new_n15846_), .ZN(new_n15847_));
  NAND2_X1   g15590(.A1(new_n15843_), .A2(new_n1158_), .ZN(new_n15848_));
  AOI21_X1   g15591(.A1(new_n15847_), .A2(new_n15848_), .B(new_n15649_), .ZN(new_n15849_));
  NOR2_X1    g15592(.A1(new_n15845_), .A2(new_n15849_), .ZN(new_n15850_));
  INV_X1     g15593(.I(new_n15850_), .ZN(new_n15851_));
  NAND2_X1   g15594(.A1(new_n15840_), .A2(new_n15851_), .ZN(new_n15852_));
  NOR2_X1    g15595(.A1(new_n15840_), .A2(new_n15851_), .ZN(new_n15853_));
  INV_X1     g15596(.I(new_n15853_), .ZN(new_n15854_));
  AOI21_X1   g15597(.A1(new_n15854_), .A2(new_n15852_), .B(new_n15838_), .ZN(new_n15855_));
  INV_X1     g15598(.I(new_n15838_), .ZN(new_n15856_));
  XOR2_X1    g15599(.A1(new_n15840_), .A2(new_n15850_), .Z(new_n15857_));
  NOR2_X1    g15600(.A1(new_n15857_), .A2(new_n15856_), .ZN(new_n15858_));
  NOR2_X1    g15601(.A1(new_n15858_), .A2(new_n15855_), .ZN(new_n15859_));
  OAI22_X1   g15602(.A1(new_n2039_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n1927_), .ZN(new_n15860_));
  NAND2_X1   g15603(.A1(new_n8628_), .A2(\b[25] ), .ZN(new_n15861_));
  AOI21_X1   g15604(.A1(new_n15861_), .A2(new_n15860_), .B(new_n7354_), .ZN(new_n15862_));
  NAND2_X1   g15605(.A1(new_n2042_), .A2(new_n15862_), .ZN(new_n15863_));
  XOR2_X1    g15606(.A1(new_n15863_), .A2(\a[59] ), .Z(new_n15864_));
  XNOR2_X1   g15607(.A1(new_n15859_), .A2(new_n15864_), .ZN(new_n15865_));
  NOR2_X1    g15608(.A1(new_n15865_), .A2(new_n15833_), .ZN(new_n15866_));
  NOR2_X1    g15609(.A1(new_n15859_), .A2(new_n15864_), .ZN(new_n15867_));
  INV_X1     g15610(.I(new_n15867_), .ZN(new_n15868_));
  NAND2_X1   g15611(.A1(new_n15859_), .A2(new_n15864_), .ZN(new_n15869_));
  AOI21_X1   g15612(.A1(new_n15868_), .A2(new_n15869_), .B(new_n15832_), .ZN(new_n15870_));
  NOR2_X1    g15613(.A1(new_n15866_), .A2(new_n15870_), .ZN(new_n15871_));
  OAI22_X1   g15614(.A1(new_n6721_), .A2(new_n2272_), .B1(new_n6723_), .B2(new_n2405_), .ZN(new_n15872_));
  NAND2_X1   g15615(.A1(new_n7617_), .A2(\b[28] ), .ZN(new_n15873_));
  AOI21_X1   g15616(.A1(new_n15873_), .A2(new_n15872_), .B(new_n6731_), .ZN(new_n15874_));
  NAND2_X1   g15617(.A1(new_n2404_), .A2(new_n15874_), .ZN(new_n15875_));
  XOR2_X1    g15618(.A1(new_n15875_), .A2(\a[56] ), .Z(new_n15876_));
  AOI21_X1   g15619(.A1(new_n15661_), .A2(new_n15672_), .B(new_n15670_), .ZN(new_n15877_));
  NOR2_X1    g15620(.A1(new_n15877_), .A2(new_n15876_), .ZN(new_n15878_));
  NAND2_X1   g15621(.A1(new_n15877_), .A2(new_n15876_), .ZN(new_n15879_));
  INV_X1     g15622(.I(new_n15879_), .ZN(new_n15880_));
  NOR2_X1    g15623(.A1(new_n15880_), .A2(new_n15878_), .ZN(new_n15881_));
  XOR2_X1    g15624(.A1(new_n15877_), .A2(new_n15876_), .Z(new_n15882_));
  NAND2_X1   g15625(.A1(new_n15882_), .A2(new_n15871_), .ZN(new_n15883_));
  OAI21_X1   g15626(.A1(new_n15871_), .A2(new_n15881_), .B(new_n15883_), .ZN(new_n15884_));
  OAI22_X1   g15627(.A1(new_n5786_), .A2(new_n2794_), .B1(new_n2660_), .B2(new_n5792_), .ZN(new_n15885_));
  NAND2_X1   g15628(.A1(new_n6745_), .A2(\b[31] ), .ZN(new_n15886_));
  AOI21_X1   g15629(.A1(new_n15886_), .A2(new_n15885_), .B(new_n5796_), .ZN(new_n15887_));
  NAND2_X1   g15630(.A1(new_n2797_), .A2(new_n15887_), .ZN(new_n15888_));
  XOR2_X1    g15631(.A1(new_n15888_), .A2(\a[53] ), .Z(new_n15889_));
  NOR2_X1    g15632(.A1(new_n15884_), .A2(new_n15889_), .ZN(new_n15890_));
  INV_X1     g15633(.I(new_n15890_), .ZN(new_n15891_));
  NAND2_X1   g15634(.A1(new_n15884_), .A2(new_n15889_), .ZN(new_n15892_));
  AOI21_X1   g15635(.A1(new_n15891_), .A2(new_n15892_), .B(new_n15831_), .ZN(new_n15893_));
  INV_X1     g15636(.I(new_n15831_), .ZN(new_n15894_));
  XNOR2_X1   g15637(.A1(new_n15884_), .A2(new_n15889_), .ZN(new_n15895_));
  NOR2_X1    g15638(.A1(new_n15895_), .A2(new_n15894_), .ZN(new_n15896_));
  NOR2_X1    g15639(.A1(new_n15896_), .A2(new_n15893_), .ZN(new_n15897_));
  OAI22_X1   g15640(.A1(new_n5228_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n5225_), .ZN(new_n15898_));
  NAND2_X1   g15641(.A1(new_n5387_), .A2(\b[34] ), .ZN(new_n15899_));
  AOI21_X1   g15642(.A1(new_n15898_), .A2(new_n15899_), .B(new_n5231_), .ZN(new_n15900_));
  NAND2_X1   g15643(.A1(new_n3246_), .A2(new_n15900_), .ZN(new_n15901_));
  XOR2_X1    g15644(.A1(new_n15901_), .A2(\a[50] ), .Z(new_n15902_));
  XNOR2_X1   g15645(.A1(new_n15897_), .A2(new_n15902_), .ZN(new_n15903_));
  NOR2_X1    g15646(.A1(new_n15903_), .A2(new_n15829_), .ZN(new_n15904_));
  INV_X1     g15647(.I(new_n15829_), .ZN(new_n15905_));
  NOR2_X1    g15648(.A1(new_n15897_), .A2(new_n15902_), .ZN(new_n15906_));
  INV_X1     g15649(.I(new_n15906_), .ZN(new_n15907_));
  NAND2_X1   g15650(.A1(new_n15897_), .A2(new_n15902_), .ZN(new_n15908_));
  AOI21_X1   g15651(.A1(new_n15907_), .A2(new_n15908_), .B(new_n15905_), .ZN(new_n15909_));
  NOR2_X1    g15652(.A1(new_n15904_), .A2(new_n15909_), .ZN(new_n15910_));
  OAI22_X1   g15653(.A1(new_n4711_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n4706_), .ZN(new_n15911_));
  NAND2_X1   g15654(.A1(new_n5814_), .A2(\b[37] ), .ZN(new_n15912_));
  AOI21_X1   g15655(.A1(new_n15911_), .A2(new_n15912_), .B(new_n4714_), .ZN(new_n15913_));
  NAND2_X1   g15656(.A1(new_n3700_), .A2(new_n15913_), .ZN(new_n15914_));
  XOR2_X1    g15657(.A1(new_n15914_), .A2(\a[47] ), .Z(new_n15915_));
  INV_X1     g15658(.I(new_n15915_), .ZN(new_n15916_));
  XOR2_X1    g15659(.A1(new_n15910_), .A2(new_n15916_), .Z(new_n15917_));
  NAND2_X1   g15660(.A1(new_n15910_), .A2(new_n15916_), .ZN(new_n15918_));
  NOR2_X1    g15661(.A1(new_n15910_), .A2(new_n15916_), .ZN(new_n15919_));
  INV_X1     g15662(.I(new_n15919_), .ZN(new_n15920_));
  AOI21_X1   g15663(.A1(new_n15920_), .A2(new_n15918_), .B(new_n15827_), .ZN(new_n15921_));
  AOI21_X1   g15664(.A1(new_n15827_), .A2(new_n15917_), .B(new_n15921_), .ZN(new_n15922_));
  OAI22_X1   g15665(.A1(new_n4208_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n4203_), .ZN(new_n15923_));
  NAND2_X1   g15666(.A1(new_n5244_), .A2(\b[40] ), .ZN(new_n15924_));
  AOI21_X1   g15667(.A1(new_n15923_), .A2(new_n15924_), .B(new_n4211_), .ZN(new_n15925_));
  NAND2_X1   g15668(.A1(new_n4017_), .A2(new_n15925_), .ZN(new_n15926_));
  XOR2_X1    g15669(.A1(new_n15926_), .A2(\a[44] ), .Z(new_n15927_));
  NAND2_X1   g15670(.A1(new_n15702_), .A2(new_n15699_), .ZN(new_n15928_));
  NAND2_X1   g15671(.A1(new_n15928_), .A2(new_n15701_), .ZN(new_n15929_));
  INV_X1     g15672(.I(new_n15929_), .ZN(new_n15930_));
  NOR2_X1    g15673(.A1(new_n15930_), .A2(new_n15927_), .ZN(new_n15931_));
  INV_X1     g15674(.I(new_n15927_), .ZN(new_n15932_));
  NOR2_X1    g15675(.A1(new_n15929_), .A2(new_n15932_), .ZN(new_n15933_));
  NOR2_X1    g15676(.A1(new_n15931_), .A2(new_n15933_), .ZN(new_n15934_));
  XOR2_X1    g15677(.A1(new_n15929_), .A2(new_n15932_), .Z(new_n15935_));
  NAND2_X1   g15678(.A1(new_n15935_), .A2(new_n15922_), .ZN(new_n15936_));
  OAI21_X1   g15679(.A1(new_n15922_), .A2(new_n15934_), .B(new_n15936_), .ZN(new_n15937_));
  OAI22_X1   g15680(.A1(new_n3736_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n3731_), .ZN(new_n15938_));
  NAND2_X1   g15681(.A1(new_n4730_), .A2(\b[43] ), .ZN(new_n15939_));
  AOI21_X1   g15682(.A1(new_n15938_), .A2(new_n15939_), .B(new_n3739_), .ZN(new_n15940_));
  NAND2_X1   g15683(.A1(new_n4513_), .A2(new_n15940_), .ZN(new_n15941_));
  XOR2_X1    g15684(.A1(new_n15941_), .A2(\a[41] ), .Z(new_n15942_));
  XNOR2_X1   g15685(.A1(new_n15937_), .A2(new_n15942_), .ZN(new_n15943_));
  NOR2_X1    g15686(.A1(new_n15943_), .A2(new_n15824_), .ZN(new_n15944_));
  NOR2_X1    g15687(.A1(new_n15937_), .A2(new_n15942_), .ZN(new_n15945_));
  INV_X1     g15688(.I(new_n15945_), .ZN(new_n15946_));
  NAND2_X1   g15689(.A1(new_n15937_), .A2(new_n15942_), .ZN(new_n15947_));
  AOI21_X1   g15690(.A1(new_n15946_), .A2(new_n15947_), .B(new_n15823_), .ZN(new_n15948_));
  NOR2_X1    g15691(.A1(new_n15944_), .A2(new_n15948_), .ZN(new_n15949_));
  INV_X1     g15692(.I(new_n15949_), .ZN(new_n15950_));
  OAI22_X1   g15693(.A1(new_n3298_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n3293_), .ZN(new_n15951_));
  NAND2_X1   g15694(.A1(new_n4227_), .A2(\b[46] ), .ZN(new_n15952_));
  AOI21_X1   g15695(.A1(new_n15951_), .A2(new_n15952_), .B(new_n3301_), .ZN(new_n15953_));
  NAND2_X1   g15696(.A1(new_n5177_), .A2(new_n15953_), .ZN(new_n15954_));
  XOR2_X1    g15697(.A1(new_n15954_), .A2(\a[38] ), .Z(new_n15955_));
  NAND2_X1   g15698(.A1(new_n15725_), .A2(new_n15712_), .ZN(new_n15956_));
  NAND2_X1   g15699(.A1(new_n15956_), .A2(new_n15724_), .ZN(new_n15957_));
  INV_X1     g15700(.I(new_n15957_), .ZN(new_n15958_));
  NOR2_X1    g15701(.A1(new_n15958_), .A2(new_n15955_), .ZN(new_n15959_));
  INV_X1     g15702(.I(new_n15955_), .ZN(new_n15960_));
  NOR2_X1    g15703(.A1(new_n15957_), .A2(new_n15960_), .ZN(new_n15961_));
  OAI21_X1   g15704(.A1(new_n15961_), .A2(new_n15959_), .B(new_n15950_), .ZN(new_n15962_));
  XOR2_X1    g15705(.A1(new_n15957_), .A2(new_n15955_), .Z(new_n15963_));
  OAI21_X1   g15706(.A1(new_n15950_), .A2(new_n15963_), .B(new_n15962_), .ZN(new_n15964_));
  OAI22_X1   g15707(.A1(new_n2846_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n2841_), .ZN(new_n15965_));
  NAND2_X1   g15708(.A1(new_n3755_), .A2(\b[49] ), .ZN(new_n15966_));
  AOI21_X1   g15709(.A1(new_n15965_), .A2(new_n15966_), .B(new_n2849_), .ZN(new_n15967_));
  NAND2_X1   g15710(.A1(new_n5741_), .A2(new_n15967_), .ZN(new_n15968_));
  XOR2_X1    g15711(.A1(new_n15968_), .A2(\a[35] ), .Z(new_n15969_));
  NOR2_X1    g15712(.A1(new_n15964_), .A2(new_n15969_), .ZN(new_n15970_));
  NAND2_X1   g15713(.A1(new_n15964_), .A2(new_n15969_), .ZN(new_n15971_));
  INV_X1     g15714(.I(new_n15971_), .ZN(new_n15972_));
  OAI21_X1   g15715(.A1(new_n15972_), .A2(new_n15970_), .B(new_n15822_), .ZN(new_n15973_));
  XNOR2_X1   g15716(.A1(new_n15964_), .A2(new_n15969_), .ZN(new_n15974_));
  OAI21_X1   g15717(.A1(new_n15822_), .A2(new_n15974_), .B(new_n15973_), .ZN(new_n15975_));
  XOR2_X1    g15718(.A1(new_n15975_), .A2(new_n15819_), .Z(new_n15976_));
  NAND2_X1   g15719(.A1(new_n15976_), .A2(new_n15817_), .ZN(new_n15977_));
  AND2_X2    g15720(.A1(new_n15975_), .A2(new_n15819_), .Z(new_n15978_));
  NOR2_X1    g15721(.A1(new_n15975_), .A2(new_n15819_), .ZN(new_n15979_));
  OAI21_X1   g15722(.A1(new_n15978_), .A2(new_n15979_), .B(new_n15816_), .ZN(new_n15980_));
  NAND2_X1   g15723(.A1(new_n15977_), .A2(new_n15980_), .ZN(new_n15981_));
  AND2_X2    g15724(.A1(new_n15981_), .A2(new_n15811_), .Z(new_n15982_));
  NOR2_X1    g15725(.A1(new_n15981_), .A2(new_n15811_), .ZN(new_n15983_));
  OAI21_X1   g15726(.A1(new_n15982_), .A2(new_n15983_), .B(new_n15806_), .ZN(new_n15984_));
  XOR2_X1    g15727(.A1(new_n15981_), .A2(new_n15811_), .Z(new_n15985_));
  NAND2_X1   g15728(.A1(new_n15985_), .A2(new_n15805_), .ZN(new_n15986_));
  NAND2_X1   g15729(.A1(new_n15986_), .A2(new_n15984_), .ZN(new_n15987_));
  XOR2_X1    g15730(.A1(new_n15804_), .A2(new_n15987_), .Z(new_n15988_));
  NAND2_X1   g15731(.A1(new_n15988_), .A2(new_n15802_), .ZN(new_n15989_));
  AOI22_X1   g15732(.A1(new_n15803_), .A2(new_n15757_), .B1(new_n15986_), .B2(new_n15984_), .ZN(new_n15990_));
  NOR2_X1    g15733(.A1(new_n15804_), .A2(new_n15987_), .ZN(new_n15991_));
  OAI21_X1   g15734(.A1(new_n15991_), .A2(new_n15990_), .B(new_n15801_), .ZN(new_n15992_));
  AOI21_X1   g15735(.A1(new_n15989_), .A2(new_n15992_), .B(new_n15796_), .ZN(new_n15993_));
  NAND2_X1   g15736(.A1(new_n15989_), .A2(new_n15992_), .ZN(new_n15994_));
  NOR2_X1    g15737(.A1(new_n15994_), .A2(new_n15795_), .ZN(new_n15995_));
  OAI21_X1   g15738(.A1(new_n15995_), .A2(new_n15993_), .B(new_n15790_), .ZN(new_n15996_));
  XOR2_X1    g15739(.A1(new_n15994_), .A2(new_n15796_), .Z(new_n15997_));
  OAI21_X1   g15740(.A1(new_n15997_), .A2(new_n15790_), .B(new_n15996_), .ZN(new_n15998_));
  NAND2_X1   g15741(.A1(new_n15772_), .A2(new_n15577_), .ZN(new_n15999_));
  XOR2_X1    g15742(.A1(new_n15578_), .A2(\a[20] ), .Z(new_n16000_));
  OAI21_X1   g15743(.A1(new_n15772_), .A2(new_n15577_), .B(new_n16000_), .ZN(new_n16001_));
  NAND2_X1   g15744(.A1(new_n16001_), .A2(new_n15999_), .ZN(new_n16002_));
  XNOR2_X1   g15745(.A1(new_n16002_), .A2(new_n15998_), .ZN(new_n16003_));
  AOI21_X1   g15746(.A1(new_n15567_), .A2(new_n15568_), .B(new_n15566_), .ZN(new_n16004_));
  NAND3_X1   g15747(.A1(new_n15330_), .A2(new_n15555_), .A3(new_n15556_), .ZN(new_n16005_));
  INV_X1     g15748(.I(new_n16005_), .ZN(new_n16006_));
  NOR3_X1    g15749(.A1(new_n16004_), .A2(new_n16006_), .A3(new_n15573_), .ZN(new_n16007_));
  AOI21_X1   g15750(.A1(new_n15565_), .A2(new_n16005_), .B(new_n15574_), .ZN(new_n16008_));
  OAI21_X1   g15751(.A1(new_n16008_), .A2(new_n16007_), .B(new_n15779_), .ZN(new_n16009_));
  XNOR2_X1   g15752(.A1(new_n16009_), .A2(new_n16003_), .ZN(new_n16010_));
  NAND2_X1   g15753(.A1(new_n15572_), .A2(new_n15574_), .ZN(new_n16011_));
  XOR2_X1    g15754(.A1(new_n16010_), .A2(new_n16011_), .Z(\f[84] ));
  NOR2_X1    g15755(.A1(new_n1548_), .A2(new_n8932_), .ZN(new_n16013_));
  NOR2_X1    g15756(.A1(new_n1439_), .A2(new_n8956_), .ZN(new_n16014_));
  NOR4_X1    g15757(.A1(new_n9323_), .A2(new_n1447_), .A3(new_n16013_), .A4(new_n16014_), .ZN(new_n16015_));
  XOR2_X1    g15758(.A1(new_n16015_), .A2(new_n1434_), .Z(new_n16016_));
  NOR2_X1    g15759(.A1(new_n15991_), .A2(new_n15801_), .ZN(new_n16017_));
  OAI22_X1   g15760(.A1(new_n1760_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n1755_), .ZN(new_n16018_));
  NAND2_X1   g15761(.A1(new_n2470_), .A2(\b[59] ), .ZN(new_n16019_));
  AOI21_X1   g15762(.A1(new_n16018_), .A2(new_n16019_), .B(new_n1763_), .ZN(new_n16020_));
  NAND2_X1   g15763(.A1(new_n8550_), .A2(new_n16020_), .ZN(new_n16021_));
  XOR2_X1    g15764(.A1(new_n16021_), .A2(\a[26] ), .Z(new_n16022_));
  NOR2_X1    g15765(.A1(new_n15982_), .A2(new_n15805_), .ZN(new_n16023_));
  NOR2_X1    g15766(.A1(new_n16023_), .A2(new_n15983_), .ZN(new_n16024_));
  OAI22_X1   g15767(.A1(new_n2084_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n2079_), .ZN(new_n16025_));
  NAND2_X1   g15768(.A1(new_n2864_), .A2(\b[56] ), .ZN(new_n16026_));
  AOI21_X1   g15769(.A1(new_n16025_), .A2(new_n16026_), .B(new_n2087_), .ZN(new_n16027_));
  NAND2_X1   g15770(.A1(new_n7559_), .A2(new_n16027_), .ZN(new_n16028_));
  XOR2_X1    g15771(.A1(new_n16028_), .A2(\a[29] ), .Z(new_n16029_));
  NOR2_X1    g15772(.A1(new_n15979_), .A2(new_n15816_), .ZN(new_n16030_));
  NOR2_X1    g15773(.A1(new_n16030_), .A2(new_n15978_), .ZN(new_n16031_));
  AOI21_X1   g15774(.A1(new_n15822_), .A2(new_n15971_), .B(new_n15970_), .ZN(new_n16032_));
  OAI22_X1   g15775(.A1(new_n2452_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n2447_), .ZN(new_n16033_));
  NAND2_X1   g15776(.A1(new_n3312_), .A2(\b[53] ), .ZN(new_n16034_));
  AOI21_X1   g15777(.A1(new_n16033_), .A2(new_n16034_), .B(new_n2455_), .ZN(new_n16035_));
  NAND2_X1   g15778(.A1(new_n6471_), .A2(new_n16035_), .ZN(new_n16036_));
  XOR2_X1    g15779(.A1(new_n16036_), .A2(\a[32] ), .Z(new_n16037_));
  INV_X1     g15780(.I(new_n16037_), .ZN(new_n16038_));
  OAI22_X1   g15781(.A1(new_n2846_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n2841_), .ZN(new_n16039_));
  NAND2_X1   g15782(.A1(new_n3755_), .A2(\b[50] ), .ZN(new_n16040_));
  AOI21_X1   g15783(.A1(new_n16039_), .A2(new_n16040_), .B(new_n2849_), .ZN(new_n16041_));
  NAND2_X1   g15784(.A1(new_n5954_), .A2(new_n16041_), .ZN(new_n16042_));
  XOR2_X1    g15785(.A1(new_n16042_), .A2(\a[35] ), .Z(new_n16043_));
  OAI22_X1   g15786(.A1(new_n3736_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n3731_), .ZN(new_n16044_));
  NAND2_X1   g15787(.A1(new_n4730_), .A2(\b[44] ), .ZN(new_n16045_));
  AOI21_X1   g15788(.A1(new_n16044_), .A2(new_n16045_), .B(new_n3739_), .ZN(new_n16046_));
  NAND2_X1   g15789(.A1(new_n4833_), .A2(new_n16046_), .ZN(new_n16047_));
  XOR2_X1    g15790(.A1(new_n16047_), .A2(\a[41] ), .Z(new_n16048_));
  OAI21_X1   g15791(.A1(new_n15826_), .A2(new_n15919_), .B(new_n15918_), .ZN(new_n16049_));
  INV_X1     g15792(.I(new_n16049_), .ZN(new_n16050_));
  OAI22_X1   g15793(.A1(new_n4711_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n4706_), .ZN(new_n16051_));
  NAND2_X1   g15794(.A1(new_n5814_), .A2(\b[38] ), .ZN(new_n16052_));
  AOI21_X1   g15795(.A1(new_n16051_), .A2(new_n16052_), .B(new_n4714_), .ZN(new_n16053_));
  NAND2_X1   g15796(.A1(new_n3844_), .A2(new_n16053_), .ZN(new_n16054_));
  XOR2_X1    g15797(.A1(new_n16054_), .A2(\a[47] ), .Z(new_n16055_));
  NAND2_X1   g15798(.A1(new_n15908_), .A2(new_n15905_), .ZN(new_n16056_));
  NAND2_X1   g15799(.A1(new_n16056_), .A2(new_n15907_), .ZN(new_n16057_));
  OAI22_X1   g15800(.A1(new_n5786_), .A2(new_n2964_), .B1(new_n2794_), .B2(new_n5792_), .ZN(new_n16058_));
  NAND2_X1   g15801(.A1(new_n6745_), .A2(\b[32] ), .ZN(new_n16059_));
  AOI21_X1   g15802(.A1(new_n16059_), .A2(new_n16058_), .B(new_n5796_), .ZN(new_n16060_));
  NAND2_X1   g15803(.A1(new_n2963_), .A2(new_n16060_), .ZN(new_n16061_));
  XOR2_X1    g15804(.A1(new_n16061_), .A2(\a[53] ), .Z(new_n16062_));
  AOI21_X1   g15805(.A1(new_n15832_), .A2(new_n15869_), .B(new_n15867_), .ZN(new_n16063_));
  INV_X1     g15806(.I(new_n16063_), .ZN(new_n16064_));
  OAI22_X1   g15807(.A1(new_n2175_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2039_), .ZN(new_n16065_));
  NAND2_X1   g15808(.A1(new_n8628_), .A2(\b[26] ), .ZN(new_n16066_));
  AOI21_X1   g15809(.A1(new_n16066_), .A2(new_n16065_), .B(new_n7354_), .ZN(new_n16067_));
  NAND2_X1   g15810(.A1(new_n2174_), .A2(new_n16067_), .ZN(new_n16068_));
  XOR2_X1    g15811(.A1(new_n16068_), .A2(\a[59] ), .Z(new_n16069_));
  NAND2_X1   g15812(.A1(new_n15852_), .A2(new_n15856_), .ZN(new_n16070_));
  NAND2_X1   g15813(.A1(new_n16070_), .A2(new_n15854_), .ZN(new_n16071_));
  OAI22_X1   g15814(.A1(new_n1825_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1709_), .ZN(new_n16072_));
  NAND2_X1   g15815(.A1(new_n9644_), .A2(\b[23] ), .ZN(new_n16073_));
  AOI21_X1   g15816(.A1(new_n16073_), .A2(new_n16072_), .B(new_n8321_), .ZN(new_n16074_));
  NAND2_X1   g15817(.A1(new_n1828_), .A2(new_n16074_), .ZN(new_n16075_));
  XOR2_X1    g15818(.A1(new_n16075_), .A2(\a[62] ), .Z(new_n16076_));
  NAND2_X1   g15819(.A1(new_n15848_), .A2(new_n15649_), .ZN(new_n16077_));
  NAND2_X1   g15820(.A1(new_n16077_), .A2(new_n15847_), .ZN(new_n16078_));
  NOR3_X1    g15821(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n1393_), .ZN(new_n16079_));
  NOR2_X1    g15822(.A1(new_n9364_), .A2(new_n1393_), .ZN(new_n16080_));
  NOR3_X1    g15823(.A1(new_n16080_), .A2(new_n1518_), .A3(new_n8985_), .ZN(new_n16081_));
  NOR2_X1    g15824(.A1(new_n16081_), .A2(new_n16079_), .ZN(new_n16082_));
  INV_X1     g15825(.I(new_n16082_), .ZN(new_n16083_));
  XOR2_X1    g15826(.A1(new_n16078_), .A2(new_n16083_), .Z(new_n16084_));
  OR2_X2     g15827(.A1(new_n16076_), .A2(new_n16084_), .Z(new_n16085_));
  NOR2_X1    g15828(.A1(new_n16078_), .A2(new_n16082_), .ZN(new_n16086_));
  NAND2_X1   g15829(.A1(new_n16078_), .A2(new_n16082_), .ZN(new_n16087_));
  INV_X1     g15830(.I(new_n16087_), .ZN(new_n16088_));
  OAI21_X1   g15831(.A1(new_n16086_), .A2(new_n16088_), .B(new_n16076_), .ZN(new_n16089_));
  NAND2_X1   g15832(.A1(new_n16085_), .A2(new_n16089_), .ZN(new_n16090_));
  XOR2_X1    g15833(.A1(new_n16071_), .A2(new_n16090_), .Z(new_n16091_));
  NOR2_X1    g15834(.A1(new_n16091_), .A2(new_n16069_), .ZN(new_n16092_));
  INV_X1     g15835(.I(new_n16069_), .ZN(new_n16093_));
  INV_X1     g15836(.I(new_n16090_), .ZN(new_n16094_));
  NOR2_X1    g15837(.A1(new_n16094_), .A2(new_n16071_), .ZN(new_n16095_));
  INV_X1     g15838(.I(new_n16095_), .ZN(new_n16096_));
  NAND2_X1   g15839(.A1(new_n16094_), .A2(new_n16071_), .ZN(new_n16097_));
  AOI21_X1   g15840(.A1(new_n16096_), .A2(new_n16097_), .B(new_n16093_), .ZN(new_n16098_));
  OAI22_X1   g15841(.A1(new_n6721_), .A2(new_n2405_), .B1(new_n6723_), .B2(new_n2543_), .ZN(new_n16099_));
  NAND2_X1   g15842(.A1(new_n7617_), .A2(\b[29] ), .ZN(new_n16100_));
  AOI21_X1   g15843(.A1(new_n16100_), .A2(new_n16099_), .B(new_n6731_), .ZN(new_n16101_));
  NAND2_X1   g15844(.A1(new_n2546_), .A2(new_n16101_), .ZN(new_n16102_));
  XOR2_X1    g15845(.A1(new_n16102_), .A2(\a[56] ), .Z(new_n16103_));
  NOR3_X1    g15846(.A1(new_n16098_), .A2(new_n16092_), .A3(new_n16103_), .ZN(new_n16104_));
  NOR2_X1    g15847(.A1(new_n16098_), .A2(new_n16092_), .ZN(new_n16105_));
  INV_X1     g15848(.I(new_n16103_), .ZN(new_n16106_));
  NOR2_X1    g15849(.A1(new_n16105_), .A2(new_n16106_), .ZN(new_n16107_));
  OAI21_X1   g15850(.A1(new_n16107_), .A2(new_n16104_), .B(new_n16064_), .ZN(new_n16108_));
  XOR2_X1    g15851(.A1(new_n16105_), .A2(new_n16103_), .Z(new_n16109_));
  OAI21_X1   g15852(.A1(new_n16109_), .A2(new_n16064_), .B(new_n16108_), .ZN(new_n16110_));
  INV_X1     g15853(.I(new_n16110_), .ZN(new_n16111_));
  AOI21_X1   g15854(.A1(new_n15871_), .A2(new_n15879_), .B(new_n15878_), .ZN(new_n16112_));
  NOR2_X1    g15855(.A1(new_n16111_), .A2(new_n16112_), .ZN(new_n16113_));
  INV_X1     g15856(.I(new_n16113_), .ZN(new_n16114_));
  NAND2_X1   g15857(.A1(new_n16111_), .A2(new_n16112_), .ZN(new_n16115_));
  AOI21_X1   g15858(.A1(new_n16114_), .A2(new_n16115_), .B(new_n16062_), .ZN(new_n16116_));
  INV_X1     g15859(.I(new_n16062_), .ZN(new_n16117_));
  XOR2_X1    g15860(.A1(new_n16110_), .A2(new_n16112_), .Z(new_n16118_));
  NOR2_X1    g15861(.A1(new_n16118_), .A2(new_n16117_), .ZN(new_n16119_));
  NAND2_X1   g15862(.A1(new_n15894_), .A2(new_n15892_), .ZN(new_n16120_));
  NAND2_X1   g15863(.A1(new_n16120_), .A2(new_n15891_), .ZN(new_n16121_));
  OAI22_X1   g15864(.A1(new_n5228_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n5225_), .ZN(new_n16122_));
  NAND2_X1   g15865(.A1(new_n5387_), .A2(\b[35] ), .ZN(new_n16123_));
  AOI21_X1   g15866(.A1(new_n16122_), .A2(new_n16123_), .B(new_n5231_), .ZN(new_n16124_));
  NAND2_X1   g15867(.A1(new_n3411_), .A2(new_n16124_), .ZN(new_n16125_));
  XOR2_X1    g15868(.A1(new_n16125_), .A2(\a[50] ), .Z(new_n16126_));
  INV_X1     g15869(.I(new_n16126_), .ZN(new_n16127_));
  XOR2_X1    g15870(.A1(new_n16121_), .A2(new_n16127_), .Z(new_n16128_));
  OAI21_X1   g15871(.A1(new_n16116_), .A2(new_n16119_), .B(new_n16128_), .ZN(new_n16129_));
  NOR2_X1    g15872(.A1(new_n16116_), .A2(new_n16119_), .ZN(new_n16130_));
  AOI21_X1   g15873(.A1(new_n16120_), .A2(new_n15891_), .B(new_n16126_), .ZN(new_n16131_));
  NOR2_X1    g15874(.A1(new_n16121_), .A2(new_n16127_), .ZN(new_n16132_));
  OAI21_X1   g15875(.A1(new_n16132_), .A2(new_n16131_), .B(new_n16130_), .ZN(new_n16133_));
  NAND2_X1   g15876(.A1(new_n16129_), .A2(new_n16133_), .ZN(new_n16134_));
  XOR2_X1    g15877(.A1(new_n16134_), .A2(new_n16057_), .Z(new_n16135_));
  AOI21_X1   g15878(.A1(new_n16129_), .A2(new_n16133_), .B(new_n16057_), .ZN(new_n16136_));
  AOI21_X1   g15879(.A1(new_n15907_), .A2(new_n16056_), .B(new_n16134_), .ZN(new_n16137_));
  OAI21_X1   g15880(.A1(new_n16137_), .A2(new_n16136_), .B(new_n16055_), .ZN(new_n16138_));
  OAI21_X1   g15881(.A1(new_n16055_), .A2(new_n16135_), .B(new_n16138_), .ZN(new_n16139_));
  OAI22_X1   g15882(.A1(new_n4208_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n4203_), .ZN(new_n16140_));
  NAND2_X1   g15883(.A1(new_n5244_), .A2(\b[41] ), .ZN(new_n16141_));
  AOI21_X1   g15884(.A1(new_n16140_), .A2(new_n16141_), .B(new_n4211_), .ZN(new_n16142_));
  NAND2_X1   g15885(.A1(new_n4320_), .A2(new_n16142_), .ZN(new_n16143_));
  XOR2_X1    g15886(.A1(new_n16143_), .A2(\a[44] ), .Z(new_n16144_));
  NOR2_X1    g15887(.A1(new_n16139_), .A2(new_n16144_), .ZN(new_n16145_));
  INV_X1     g15888(.I(new_n16145_), .ZN(new_n16146_));
  NAND2_X1   g15889(.A1(new_n16139_), .A2(new_n16144_), .ZN(new_n16147_));
  AOI21_X1   g15890(.A1(new_n16146_), .A2(new_n16147_), .B(new_n16050_), .ZN(new_n16148_));
  XNOR2_X1   g15891(.A1(new_n16139_), .A2(new_n16144_), .ZN(new_n16149_));
  NOR2_X1    g15892(.A1(new_n16149_), .A2(new_n16049_), .ZN(new_n16150_));
  NOR2_X1    g15893(.A1(new_n16150_), .A2(new_n16148_), .ZN(new_n16151_));
  INV_X1     g15894(.I(new_n16151_), .ZN(new_n16152_));
  OAI21_X1   g15895(.A1(new_n15932_), .A2(new_n15929_), .B(new_n15922_), .ZN(new_n16153_));
  OAI21_X1   g15896(.A1(new_n15927_), .A2(new_n15930_), .B(new_n16153_), .ZN(new_n16154_));
  NAND2_X1   g15897(.A1(new_n16152_), .A2(new_n16154_), .ZN(new_n16155_));
  NOR2_X1    g15898(.A1(new_n16152_), .A2(new_n16154_), .ZN(new_n16156_));
  INV_X1     g15899(.I(new_n16156_), .ZN(new_n16157_));
  AOI21_X1   g15900(.A1(new_n16157_), .A2(new_n16155_), .B(new_n16048_), .ZN(new_n16158_));
  XNOR2_X1   g15901(.A1(new_n16151_), .A2(new_n16154_), .ZN(new_n16159_));
  AOI21_X1   g15902(.A1(new_n16048_), .A2(new_n16159_), .B(new_n16158_), .ZN(new_n16160_));
  AOI21_X1   g15903(.A1(new_n15937_), .A2(new_n15942_), .B(new_n15824_), .ZN(new_n16161_));
  NOR2_X1    g15904(.A1(new_n16161_), .A2(new_n15945_), .ZN(new_n16162_));
  OAI22_X1   g15905(.A1(new_n3298_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n3293_), .ZN(new_n16163_));
  NAND2_X1   g15906(.A1(new_n4227_), .A2(\b[47] ), .ZN(new_n16164_));
  AOI21_X1   g15907(.A1(new_n16163_), .A2(new_n16164_), .B(new_n3301_), .ZN(new_n16165_));
  NAND2_X1   g15908(.A1(new_n5196_), .A2(new_n16165_), .ZN(new_n16166_));
  XOR2_X1    g15909(.A1(new_n16166_), .A2(\a[38] ), .Z(new_n16167_));
  NOR2_X1    g15910(.A1(new_n16162_), .A2(new_n16167_), .ZN(new_n16168_));
  INV_X1     g15911(.I(new_n16162_), .ZN(new_n16169_));
  INV_X1     g15912(.I(new_n16167_), .ZN(new_n16170_));
  NOR2_X1    g15913(.A1(new_n16169_), .A2(new_n16170_), .ZN(new_n16171_));
  NOR2_X1    g15914(.A1(new_n16171_), .A2(new_n16168_), .ZN(new_n16172_));
  XOR2_X1    g15915(.A1(new_n16162_), .A2(new_n16167_), .Z(new_n16173_));
  NAND2_X1   g15916(.A1(new_n16160_), .A2(new_n16173_), .ZN(new_n16174_));
  OAI21_X1   g15917(.A1(new_n16160_), .A2(new_n16172_), .B(new_n16174_), .ZN(new_n16175_));
  NOR2_X1    g15918(.A1(new_n15950_), .A2(new_n15961_), .ZN(new_n16176_));
  NOR2_X1    g15919(.A1(new_n16176_), .A2(new_n15959_), .ZN(new_n16177_));
  INV_X1     g15920(.I(new_n16177_), .ZN(new_n16178_));
  NAND2_X1   g15921(.A1(new_n16178_), .A2(new_n16175_), .ZN(new_n16179_));
  INV_X1     g15922(.I(new_n16175_), .ZN(new_n16180_));
  NAND2_X1   g15923(.A1(new_n16180_), .A2(new_n16177_), .ZN(new_n16181_));
  AOI21_X1   g15924(.A1(new_n16181_), .A2(new_n16179_), .B(new_n16043_), .ZN(new_n16182_));
  INV_X1     g15925(.I(new_n16043_), .ZN(new_n16183_));
  XOR2_X1    g15926(.A1(new_n16175_), .A2(new_n16177_), .Z(new_n16184_));
  NOR2_X1    g15927(.A1(new_n16184_), .A2(new_n16183_), .ZN(new_n16185_));
  NOR2_X1    g15928(.A1(new_n16185_), .A2(new_n16182_), .ZN(new_n16186_));
  XOR2_X1    g15929(.A1(new_n16186_), .A2(new_n16038_), .Z(new_n16187_));
  NOR2_X1    g15930(.A1(new_n16186_), .A2(new_n16037_), .ZN(new_n16188_));
  NOR3_X1    g15931(.A1(new_n16185_), .A2(new_n16038_), .A3(new_n16182_), .ZN(new_n16189_));
  OAI21_X1   g15932(.A1(new_n16188_), .A2(new_n16189_), .B(new_n16032_), .ZN(new_n16190_));
  OAI21_X1   g15933(.A1(new_n16187_), .A2(new_n16032_), .B(new_n16190_), .ZN(new_n16191_));
  NAND2_X1   g15934(.A1(new_n16031_), .A2(new_n16191_), .ZN(new_n16192_));
  NOR2_X1    g15935(.A1(new_n16031_), .A2(new_n16191_), .ZN(new_n16193_));
  INV_X1     g15936(.I(new_n16193_), .ZN(new_n16194_));
  AOI21_X1   g15937(.A1(new_n16194_), .A2(new_n16192_), .B(new_n16029_), .ZN(new_n16195_));
  INV_X1     g15938(.I(new_n16029_), .ZN(new_n16196_));
  XNOR2_X1   g15939(.A1(new_n16031_), .A2(new_n16191_), .ZN(new_n16197_));
  NOR2_X1    g15940(.A1(new_n16197_), .A2(new_n16196_), .ZN(new_n16198_));
  NOR2_X1    g15941(.A1(new_n16198_), .A2(new_n16195_), .ZN(new_n16199_));
  XNOR2_X1   g15942(.A1(new_n16024_), .A2(new_n16199_), .ZN(new_n16200_));
  NOR2_X1    g15943(.A1(new_n16200_), .A2(new_n16022_), .ZN(new_n16201_));
  INV_X1     g15944(.I(new_n16022_), .ZN(new_n16202_));
  NOR2_X1    g15945(.A1(new_n16024_), .A2(new_n16199_), .ZN(new_n16203_));
  INV_X1     g15946(.I(new_n16203_), .ZN(new_n16204_));
  NAND2_X1   g15947(.A1(new_n16024_), .A2(new_n16199_), .ZN(new_n16205_));
  AOI21_X1   g15948(.A1(new_n16204_), .A2(new_n16205_), .B(new_n16202_), .ZN(new_n16206_));
  NOR2_X1    g15949(.A1(new_n16201_), .A2(new_n16206_), .ZN(new_n16207_));
  NOR3_X1    g15950(.A1(new_n16207_), .A2(new_n15990_), .A3(new_n16017_), .ZN(new_n16208_));
  NOR2_X1    g15951(.A1(new_n16017_), .A2(new_n15990_), .ZN(new_n16209_));
  INV_X1     g15952(.I(new_n16207_), .ZN(new_n16210_));
  NOR2_X1    g15953(.A1(new_n16210_), .A2(new_n16209_), .ZN(new_n16211_));
  NOR2_X1    g15954(.A1(new_n16211_), .A2(new_n16208_), .ZN(new_n16212_));
  NOR2_X1    g15955(.A1(new_n16212_), .A2(new_n16016_), .ZN(new_n16213_));
  INV_X1     g15956(.I(new_n16016_), .ZN(new_n16214_));
  XOR2_X1    g15957(.A1(new_n16207_), .A2(new_n16209_), .Z(new_n16215_));
  NOR2_X1    g15958(.A1(new_n16215_), .A2(new_n16214_), .ZN(new_n16216_));
  NOR2_X1    g15959(.A1(new_n16213_), .A2(new_n16216_), .ZN(new_n16217_));
  NOR2_X1    g15960(.A1(new_n15993_), .A2(new_n15789_), .ZN(new_n16218_));
  NOR2_X1    g15961(.A1(new_n16218_), .A2(new_n15995_), .ZN(new_n16219_));
  NAND3_X1   g15962(.A1(new_n15565_), .A2(new_n16005_), .A3(new_n15574_), .ZN(new_n16220_));
  NAND2_X1   g15963(.A1(new_n15572_), .A2(new_n15573_), .ZN(new_n16221_));
  NAND2_X1   g15964(.A1(new_n16221_), .A2(new_n16220_), .ZN(new_n16222_));
  NAND3_X1   g15965(.A1(new_n15572_), .A2(new_n15574_), .A3(new_n16003_), .ZN(new_n16223_));
  NAND3_X1   g15966(.A1(new_n16222_), .A2(new_n15779_), .A3(new_n16223_), .ZN(new_n16224_));
  OR2_X2     g15967(.A1(new_n16002_), .A2(new_n15998_), .Z(new_n16225_));
  NAND2_X1   g15968(.A1(new_n16224_), .A2(new_n16225_), .ZN(new_n16226_));
  XOR2_X1    g15969(.A1(new_n16226_), .A2(new_n16219_), .Z(new_n16227_));
  XOR2_X1    g15970(.A1(new_n16227_), .A2(new_n16217_), .Z(\f[85] ));
  XOR2_X1    g15971(.A1(new_n16217_), .A2(new_n16219_), .Z(new_n16229_));
  NAND2_X1   g15972(.A1(new_n16229_), .A2(new_n16219_), .ZN(new_n16230_));
  INV_X1     g15973(.I(new_n16230_), .ZN(new_n16231_));
  AND2_X2    g15974(.A1(new_n16225_), .A2(new_n16229_), .Z(new_n16232_));
  AOI21_X1   g15975(.A1(new_n16224_), .A2(new_n16232_), .B(new_n16231_), .ZN(new_n16233_));
  NOR2_X1    g15976(.A1(new_n16208_), .A2(new_n16016_), .ZN(new_n16234_));
  NOR2_X1    g15977(.A1(new_n16234_), .A2(new_n16211_), .ZN(new_n16235_));
  AOI21_X1   g15978(.A1(new_n16202_), .A2(new_n16205_), .B(new_n16203_), .ZN(new_n16236_));
  OAI22_X1   g15979(.A1(new_n9595_), .A2(new_n1447_), .B1(new_n8956_), .B2(new_n1548_), .ZN(new_n16237_));
  OAI22_X1   g15980(.A1(new_n2084_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n2079_), .ZN(new_n16238_));
  NAND2_X1   g15981(.A1(new_n2864_), .A2(\b[57] ), .ZN(new_n16239_));
  AOI21_X1   g15982(.A1(new_n16238_), .A2(new_n16239_), .B(new_n2087_), .ZN(new_n16240_));
  NAND2_X1   g15983(.A1(new_n7895_), .A2(new_n16240_), .ZN(new_n16241_));
  XOR2_X1    g15984(.A1(new_n16241_), .A2(\a[29] ), .Z(new_n16242_));
  INV_X1     g15985(.I(new_n16242_), .ZN(new_n16243_));
  OAI22_X1   g15986(.A1(new_n2452_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n2447_), .ZN(new_n16244_));
  NAND2_X1   g15987(.A1(new_n3312_), .A2(\b[54] ), .ZN(new_n16245_));
  AOI21_X1   g15988(.A1(new_n16244_), .A2(new_n16245_), .B(new_n2455_), .ZN(new_n16246_));
  NAND2_X1   g15989(.A1(new_n6994_), .A2(new_n16246_), .ZN(new_n16247_));
  XOR2_X1    g15990(.A1(new_n16247_), .A2(\a[32] ), .Z(new_n16248_));
  NOR2_X1    g15991(.A1(new_n16180_), .A2(new_n16177_), .ZN(new_n16249_));
  AOI21_X1   g15992(.A1(new_n16183_), .A2(new_n16181_), .B(new_n16249_), .ZN(new_n16250_));
  OAI22_X1   g15993(.A1(new_n2846_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n2841_), .ZN(new_n16251_));
  NAND2_X1   g15994(.A1(new_n3755_), .A2(\b[51] ), .ZN(new_n16252_));
  AOI21_X1   g15995(.A1(new_n16251_), .A2(new_n16252_), .B(new_n2849_), .ZN(new_n16253_));
  NAND2_X1   g15996(.A1(new_n6219_), .A2(new_n16253_), .ZN(new_n16254_));
  XOR2_X1    g15997(.A1(new_n16254_), .A2(\a[35] ), .Z(new_n16255_));
  OAI22_X1   g15998(.A1(new_n3298_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n3293_), .ZN(new_n16256_));
  NAND2_X1   g15999(.A1(new_n4227_), .A2(\b[48] ), .ZN(new_n16257_));
  AOI21_X1   g16000(.A1(new_n16256_), .A2(new_n16257_), .B(new_n3301_), .ZN(new_n16258_));
  NAND2_X1   g16001(.A1(new_n5537_), .A2(new_n16258_), .ZN(new_n16259_));
  XOR2_X1    g16002(.A1(new_n16259_), .A2(\a[38] ), .Z(new_n16260_));
  OAI22_X1   g16003(.A1(new_n4208_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n4203_), .ZN(new_n16261_));
  NAND2_X1   g16004(.A1(new_n5244_), .A2(\b[42] ), .ZN(new_n16262_));
  AOI21_X1   g16005(.A1(new_n16261_), .A2(new_n16262_), .B(new_n4211_), .ZN(new_n16263_));
  NAND2_X1   g16006(.A1(new_n4500_), .A2(new_n16263_), .ZN(new_n16264_));
  XOR2_X1    g16007(.A1(new_n16264_), .A2(\a[44] ), .Z(new_n16265_));
  NOR2_X1    g16008(.A1(new_n16136_), .A2(new_n16055_), .ZN(new_n16266_));
  NOR2_X1    g16009(.A1(new_n16266_), .A2(new_n16137_), .ZN(new_n16267_));
  OAI22_X1   g16010(.A1(new_n5228_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n5225_), .ZN(new_n16268_));
  NAND2_X1   g16011(.A1(new_n5387_), .A2(\b[36] ), .ZN(new_n16269_));
  AOI21_X1   g16012(.A1(new_n16268_), .A2(new_n16269_), .B(new_n5231_), .ZN(new_n16270_));
  NAND2_X1   g16013(.A1(new_n3565_), .A2(new_n16270_), .ZN(new_n16271_));
  XOR2_X1    g16014(.A1(new_n16271_), .A2(\a[50] ), .Z(new_n16272_));
  INV_X1     g16015(.I(new_n16272_), .ZN(new_n16273_));
  AOI21_X1   g16016(.A1(new_n16117_), .A2(new_n16115_), .B(new_n16113_), .ZN(new_n16274_));
  INV_X1     g16017(.I(new_n16274_), .ZN(new_n16275_));
  OAI22_X1   g16018(.A1(new_n5786_), .A2(new_n3097_), .B1(new_n2964_), .B2(new_n5792_), .ZN(new_n16276_));
  NAND2_X1   g16019(.A1(new_n6745_), .A2(\b[33] ), .ZN(new_n16277_));
  AOI21_X1   g16020(.A1(new_n16277_), .A2(new_n16276_), .B(new_n5796_), .ZN(new_n16278_));
  NAND2_X1   g16021(.A1(new_n3101_), .A2(new_n16278_), .ZN(new_n16279_));
  XOR2_X1    g16022(.A1(new_n16279_), .A2(\a[53] ), .Z(new_n16280_));
  OAI22_X1   g16023(.A1(new_n6721_), .A2(new_n2543_), .B1(new_n6723_), .B2(new_n2660_), .ZN(new_n16281_));
  NAND2_X1   g16024(.A1(new_n7617_), .A2(\b[30] ), .ZN(new_n16282_));
  AOI21_X1   g16025(.A1(new_n16282_), .A2(new_n16281_), .B(new_n6731_), .ZN(new_n16283_));
  NAND2_X1   g16026(.A1(new_n2659_), .A2(new_n16283_), .ZN(new_n16284_));
  XOR2_X1    g16027(.A1(new_n16284_), .A2(\a[56] ), .Z(new_n16285_));
  OAI22_X1   g16028(.A1(new_n1927_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1825_), .ZN(new_n16286_));
  NAND2_X1   g16029(.A1(new_n9644_), .A2(\b[24] ), .ZN(new_n16287_));
  AOI21_X1   g16030(.A1(new_n16287_), .A2(new_n16286_), .B(new_n8321_), .ZN(new_n16288_));
  NAND2_X1   g16031(.A1(new_n1926_), .A2(new_n16288_), .ZN(new_n16289_));
  XOR2_X1    g16032(.A1(new_n16289_), .A2(\a[62] ), .Z(new_n16290_));
  NOR3_X1    g16033(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n1518_), .ZN(new_n16291_));
  NOR2_X1    g16034(.A1(new_n9364_), .A2(new_n1518_), .ZN(new_n16292_));
  NOR3_X1    g16035(.A1(new_n16292_), .A2(new_n1601_), .A3(new_n8985_), .ZN(new_n16293_));
  NOR2_X1    g16036(.A1(new_n16293_), .A2(new_n16291_), .ZN(new_n16294_));
  XOR2_X1    g16037(.A1(new_n16082_), .A2(new_n16294_), .Z(new_n16295_));
  NOR2_X1    g16038(.A1(new_n16290_), .A2(new_n16295_), .ZN(new_n16296_));
  NOR2_X1    g16039(.A1(new_n16083_), .A2(new_n16294_), .ZN(new_n16297_));
  INV_X1     g16040(.I(new_n16294_), .ZN(new_n16298_));
  NOR2_X1    g16041(.A1(new_n16298_), .A2(new_n16082_), .ZN(new_n16299_));
  NOR2_X1    g16042(.A1(new_n16297_), .A2(new_n16299_), .ZN(new_n16300_));
  INV_X1     g16043(.I(new_n16300_), .ZN(new_n16301_));
  AOI21_X1   g16044(.A1(new_n16290_), .A2(new_n16301_), .B(new_n16296_), .ZN(new_n16302_));
  OAI22_X1   g16045(.A1(new_n2272_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2175_), .ZN(new_n16303_));
  NAND2_X1   g16046(.A1(new_n8628_), .A2(\b[27] ), .ZN(new_n16304_));
  AOI21_X1   g16047(.A1(new_n16304_), .A2(new_n16303_), .B(new_n7354_), .ZN(new_n16305_));
  NAND2_X1   g16048(.A1(new_n2276_), .A2(new_n16305_), .ZN(new_n16306_));
  XOR2_X1    g16049(.A1(new_n16306_), .A2(\a[59] ), .Z(new_n16307_));
  OAI21_X1   g16050(.A1(new_n16076_), .A2(new_n16086_), .B(new_n16087_), .ZN(new_n16308_));
  XOR2_X1    g16051(.A1(new_n16307_), .A2(new_n16308_), .Z(new_n16309_));
  NOR2_X1    g16052(.A1(new_n16309_), .A2(new_n16302_), .ZN(new_n16310_));
  INV_X1     g16053(.I(new_n16308_), .ZN(new_n16311_));
  NOR2_X1    g16054(.A1(new_n16307_), .A2(new_n16311_), .ZN(new_n16312_));
  INV_X1     g16055(.I(new_n16312_), .ZN(new_n16313_));
  NAND2_X1   g16056(.A1(new_n16307_), .A2(new_n16311_), .ZN(new_n16314_));
  NAND2_X1   g16057(.A1(new_n16313_), .A2(new_n16314_), .ZN(new_n16315_));
  AOI21_X1   g16058(.A1(new_n16302_), .A2(new_n16315_), .B(new_n16310_), .ZN(new_n16316_));
  OAI21_X1   g16059(.A1(new_n16069_), .A2(new_n16095_), .B(new_n16097_), .ZN(new_n16317_));
  XOR2_X1    g16060(.A1(new_n16316_), .A2(new_n16317_), .Z(new_n16318_));
  NOR2_X1    g16061(.A1(new_n16318_), .A2(new_n16285_), .ZN(new_n16319_));
  INV_X1     g16062(.I(new_n16285_), .ZN(new_n16320_));
  INV_X1     g16063(.I(new_n16317_), .ZN(new_n16321_));
  NOR2_X1    g16064(.A1(new_n16316_), .A2(new_n16321_), .ZN(new_n16322_));
  INV_X1     g16065(.I(new_n16322_), .ZN(new_n16323_));
  NAND2_X1   g16066(.A1(new_n16316_), .A2(new_n16321_), .ZN(new_n16324_));
  AOI21_X1   g16067(.A1(new_n16323_), .A2(new_n16324_), .B(new_n16320_), .ZN(new_n16325_));
  NOR2_X1    g16068(.A1(new_n16319_), .A2(new_n16325_), .ZN(new_n16326_));
  NOR2_X1    g16069(.A1(new_n16107_), .A2(new_n16063_), .ZN(new_n16327_));
  NOR2_X1    g16070(.A1(new_n16327_), .A2(new_n16104_), .ZN(new_n16328_));
  XOR2_X1    g16071(.A1(new_n16326_), .A2(new_n16328_), .Z(new_n16329_));
  NOR2_X1    g16072(.A1(new_n16329_), .A2(new_n16280_), .ZN(new_n16330_));
  INV_X1     g16073(.I(new_n16280_), .ZN(new_n16331_));
  INV_X1     g16074(.I(new_n16326_), .ZN(new_n16332_));
  NOR2_X1    g16075(.A1(new_n16332_), .A2(new_n16328_), .ZN(new_n16333_));
  INV_X1     g16076(.I(new_n16333_), .ZN(new_n16334_));
  NAND2_X1   g16077(.A1(new_n16332_), .A2(new_n16328_), .ZN(new_n16335_));
  AOI21_X1   g16078(.A1(new_n16334_), .A2(new_n16335_), .B(new_n16331_), .ZN(new_n16336_));
  NOR2_X1    g16079(.A1(new_n16336_), .A2(new_n16330_), .ZN(new_n16337_));
  NOR2_X1    g16080(.A1(new_n16337_), .A2(new_n16275_), .ZN(new_n16338_));
  NOR3_X1    g16081(.A1(new_n16336_), .A2(new_n16330_), .A3(new_n16274_), .ZN(new_n16339_));
  OAI21_X1   g16082(.A1(new_n16338_), .A2(new_n16339_), .B(new_n16273_), .ZN(new_n16340_));
  XOR2_X1    g16083(.A1(new_n16337_), .A2(new_n16275_), .Z(new_n16341_));
  NAND2_X1   g16084(.A1(new_n16341_), .A2(new_n16272_), .ZN(new_n16342_));
  NAND2_X1   g16085(.A1(new_n16342_), .A2(new_n16340_), .ZN(new_n16343_));
  OAI22_X1   g16086(.A1(new_n4711_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n4706_), .ZN(new_n16344_));
  NAND2_X1   g16087(.A1(new_n5814_), .A2(\b[39] ), .ZN(new_n16345_));
  AOI21_X1   g16088(.A1(new_n16344_), .A2(new_n16345_), .B(new_n4714_), .ZN(new_n16346_));
  NAND2_X1   g16089(.A1(new_n3996_), .A2(new_n16346_), .ZN(new_n16347_));
  XOR2_X1    g16090(.A1(new_n16347_), .A2(\a[47] ), .Z(new_n16348_));
  NOR2_X1    g16091(.A1(new_n16132_), .A2(new_n16130_), .ZN(new_n16349_));
  NOR2_X1    g16092(.A1(new_n16349_), .A2(new_n16131_), .ZN(new_n16350_));
  NOR2_X1    g16093(.A1(new_n16350_), .A2(new_n16348_), .ZN(new_n16351_));
  INV_X1     g16094(.I(new_n16351_), .ZN(new_n16352_));
  NAND2_X1   g16095(.A1(new_n16350_), .A2(new_n16348_), .ZN(new_n16353_));
  NAND2_X1   g16096(.A1(new_n16352_), .A2(new_n16353_), .ZN(new_n16354_));
  XNOR2_X1   g16097(.A1(new_n16350_), .A2(new_n16348_), .ZN(new_n16355_));
  NOR2_X1    g16098(.A1(new_n16343_), .A2(new_n16355_), .ZN(new_n16356_));
  AOI21_X1   g16099(.A1(new_n16343_), .A2(new_n16354_), .B(new_n16356_), .ZN(new_n16357_));
  XNOR2_X1   g16100(.A1(new_n16357_), .A2(new_n16267_), .ZN(new_n16358_));
  NOR2_X1    g16101(.A1(new_n16358_), .A2(new_n16265_), .ZN(new_n16359_));
  INV_X1     g16102(.I(new_n16265_), .ZN(new_n16360_));
  NOR2_X1    g16103(.A1(new_n16357_), .A2(new_n16267_), .ZN(new_n16361_));
  INV_X1     g16104(.I(new_n16361_), .ZN(new_n16362_));
  NAND2_X1   g16105(.A1(new_n16357_), .A2(new_n16267_), .ZN(new_n16363_));
  AOI21_X1   g16106(.A1(new_n16362_), .A2(new_n16363_), .B(new_n16360_), .ZN(new_n16364_));
  NOR2_X1    g16107(.A1(new_n16359_), .A2(new_n16364_), .ZN(new_n16365_));
  INV_X1     g16108(.I(new_n16365_), .ZN(new_n16366_));
  OAI22_X1   g16109(.A1(new_n3736_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n3731_), .ZN(new_n16367_));
  NAND2_X1   g16110(.A1(new_n4730_), .A2(\b[45] ), .ZN(new_n16368_));
  AOI21_X1   g16111(.A1(new_n16367_), .A2(new_n16368_), .B(new_n3739_), .ZN(new_n16369_));
  NAND2_X1   g16112(.A1(new_n5004_), .A2(new_n16369_), .ZN(new_n16370_));
  XOR2_X1    g16113(.A1(new_n16370_), .A2(\a[41] ), .Z(new_n16371_));
  INV_X1     g16114(.I(new_n16371_), .ZN(new_n16372_));
  NAND2_X1   g16115(.A1(new_n16147_), .A2(new_n16049_), .ZN(new_n16373_));
  NAND2_X1   g16116(.A1(new_n16373_), .A2(new_n16146_), .ZN(new_n16374_));
  XOR2_X1    g16117(.A1(new_n16374_), .A2(new_n16372_), .Z(new_n16375_));
  NAND2_X1   g16118(.A1(new_n16366_), .A2(new_n16375_), .ZN(new_n16376_));
  AOI21_X1   g16119(.A1(new_n16373_), .A2(new_n16146_), .B(new_n16371_), .ZN(new_n16377_));
  NOR2_X1    g16120(.A1(new_n16374_), .A2(new_n16372_), .ZN(new_n16378_));
  OAI21_X1   g16121(.A1(new_n16377_), .A2(new_n16378_), .B(new_n16365_), .ZN(new_n16379_));
  NAND2_X1   g16122(.A1(new_n16376_), .A2(new_n16379_), .ZN(new_n16380_));
  OAI21_X1   g16123(.A1(new_n16048_), .A2(new_n16156_), .B(new_n16155_), .ZN(new_n16381_));
  XNOR2_X1   g16124(.A1(new_n16380_), .A2(new_n16381_), .ZN(new_n16382_));
  NOR2_X1    g16125(.A1(new_n16382_), .A2(new_n16260_), .ZN(new_n16383_));
  INV_X1     g16126(.I(new_n16260_), .ZN(new_n16384_));
  INV_X1     g16127(.I(new_n16380_), .ZN(new_n16385_));
  INV_X1     g16128(.I(new_n16381_), .ZN(new_n16386_));
  NOR2_X1    g16129(.A1(new_n16385_), .A2(new_n16386_), .ZN(new_n16387_));
  NOR2_X1    g16130(.A1(new_n16380_), .A2(new_n16381_), .ZN(new_n16388_));
  NOR2_X1    g16131(.A1(new_n16387_), .A2(new_n16388_), .ZN(new_n16389_));
  NOR2_X1    g16132(.A1(new_n16389_), .A2(new_n16384_), .ZN(new_n16390_));
  NOR2_X1    g16133(.A1(new_n16390_), .A2(new_n16383_), .ZN(new_n16391_));
  INV_X1     g16134(.I(new_n16391_), .ZN(new_n16392_));
  INV_X1     g16135(.I(new_n16168_), .ZN(new_n16393_));
  OAI21_X1   g16136(.A1(new_n16160_), .A2(new_n16171_), .B(new_n16393_), .ZN(new_n16394_));
  INV_X1     g16137(.I(new_n16394_), .ZN(new_n16395_));
  NOR2_X1    g16138(.A1(new_n16392_), .A2(new_n16395_), .ZN(new_n16396_));
  NOR2_X1    g16139(.A1(new_n16391_), .A2(new_n16394_), .ZN(new_n16397_));
  NOR2_X1    g16140(.A1(new_n16396_), .A2(new_n16397_), .ZN(new_n16398_));
  NOR2_X1    g16141(.A1(new_n16398_), .A2(new_n16255_), .ZN(new_n16399_));
  INV_X1     g16142(.I(new_n16255_), .ZN(new_n16400_));
  XOR2_X1    g16143(.A1(new_n16391_), .A2(new_n16395_), .Z(new_n16401_));
  NOR2_X1    g16144(.A1(new_n16401_), .A2(new_n16400_), .ZN(new_n16402_));
  NOR2_X1    g16145(.A1(new_n16399_), .A2(new_n16402_), .ZN(new_n16403_));
  NOR2_X1    g16146(.A1(new_n16403_), .A2(new_n16250_), .ZN(new_n16404_));
  INV_X1     g16147(.I(new_n16404_), .ZN(new_n16405_));
  NAND2_X1   g16148(.A1(new_n16403_), .A2(new_n16250_), .ZN(new_n16406_));
  AOI21_X1   g16149(.A1(new_n16405_), .A2(new_n16406_), .B(new_n16248_), .ZN(new_n16407_));
  INV_X1     g16150(.I(new_n16248_), .ZN(new_n16408_));
  XNOR2_X1   g16151(.A1(new_n16403_), .A2(new_n16250_), .ZN(new_n16409_));
  NOR2_X1    g16152(.A1(new_n16409_), .A2(new_n16408_), .ZN(new_n16410_));
  NOR2_X1    g16153(.A1(new_n16410_), .A2(new_n16407_), .ZN(new_n16411_));
  NOR2_X1    g16154(.A1(new_n16189_), .A2(new_n16032_), .ZN(new_n16412_));
  NOR2_X1    g16155(.A1(new_n16412_), .A2(new_n16188_), .ZN(new_n16413_));
  NOR2_X1    g16156(.A1(new_n16411_), .A2(new_n16413_), .ZN(new_n16414_));
  NAND2_X1   g16157(.A1(new_n16411_), .A2(new_n16413_), .ZN(new_n16415_));
  INV_X1     g16158(.I(new_n16415_), .ZN(new_n16416_));
  OAI21_X1   g16159(.A1(new_n16416_), .A2(new_n16414_), .B(new_n16243_), .ZN(new_n16417_));
  XNOR2_X1   g16160(.A1(new_n16411_), .A2(new_n16413_), .ZN(new_n16418_));
  OAI21_X1   g16161(.A1(new_n16243_), .A2(new_n16418_), .B(new_n16417_), .ZN(new_n16419_));
  AOI22_X1   g16162(.A1(\b[62] ), .A2(new_n1759_), .B1(new_n2289_), .B2(\b[61] ), .ZN(new_n16420_));
  AOI21_X1   g16163(.A1(\b[60] ), .A2(new_n2470_), .B(new_n16420_), .ZN(new_n16421_));
  OAI21_X1   g16164(.A1(new_n15764_), .A2(new_n1763_), .B(new_n16421_), .ZN(new_n16422_));
  NAND2_X1   g16165(.A1(new_n16192_), .A2(new_n16196_), .ZN(new_n16423_));
  NAND2_X1   g16166(.A1(new_n16423_), .A2(new_n16194_), .ZN(new_n16424_));
  XOR2_X1    g16167(.A1(new_n16424_), .A2(new_n16422_), .Z(new_n16425_));
  XOR2_X1    g16168(.A1(new_n16425_), .A2(\a[26] ), .Z(new_n16426_));
  XOR2_X1    g16169(.A1(new_n16426_), .A2(new_n16419_), .Z(new_n16427_));
  XOR2_X1    g16170(.A1(new_n16427_), .A2(new_n16237_), .Z(new_n16428_));
  XOR2_X1    g16171(.A1(new_n16428_), .A2(new_n1434_), .Z(new_n16429_));
  XOR2_X1    g16172(.A1(new_n16429_), .A2(new_n16236_), .Z(new_n16430_));
  NOR2_X1    g16173(.A1(new_n16430_), .A2(new_n16235_), .ZN(new_n16431_));
  NAND2_X1   g16174(.A1(new_n16430_), .A2(new_n16235_), .ZN(new_n16432_));
  INV_X1     g16175(.I(new_n16432_), .ZN(new_n16433_));
  NOR2_X1    g16176(.A1(new_n16433_), .A2(new_n16431_), .ZN(new_n16434_));
  XOR2_X1    g16177(.A1(new_n16233_), .A2(new_n16434_), .Z(\f[86] ));
  NOR2_X1    g16178(.A1(new_n16427_), .A2(new_n16236_), .ZN(new_n16436_));
  XOR2_X1    g16179(.A1(new_n16237_), .A2(new_n1434_), .Z(new_n16437_));
  AOI21_X1   g16180(.A1(new_n16427_), .A2(new_n16236_), .B(new_n16437_), .ZN(new_n16438_));
  NOR2_X1    g16181(.A1(new_n16438_), .A2(new_n16436_), .ZN(new_n16439_));
  NAND2_X1   g16182(.A1(new_n16419_), .A2(new_n16424_), .ZN(new_n16440_));
  XOR2_X1    g16183(.A1(new_n16422_), .A2(new_n1750_), .Z(new_n16441_));
  OAI21_X1   g16184(.A1(new_n16419_), .A2(new_n16424_), .B(new_n16441_), .ZN(new_n16442_));
  NAND2_X1   g16185(.A1(new_n16442_), .A2(new_n16440_), .ZN(new_n16443_));
  OAI22_X1   g16186(.A1(new_n1760_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n1755_), .ZN(new_n16444_));
  NAND2_X1   g16187(.A1(new_n2470_), .A2(\b[61] ), .ZN(new_n16445_));
  AOI21_X1   g16188(.A1(new_n16444_), .A2(new_n16445_), .B(new_n1763_), .ZN(new_n16446_));
  NAND2_X1   g16189(.A1(new_n8963_), .A2(new_n16446_), .ZN(new_n16447_));
  XOR2_X1    g16190(.A1(new_n16447_), .A2(\a[26] ), .Z(new_n16448_));
  AOI21_X1   g16191(.A1(new_n16243_), .A2(new_n16415_), .B(new_n16414_), .ZN(new_n16449_));
  OAI22_X1   g16192(.A1(new_n2084_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n2079_), .ZN(new_n16450_));
  NAND2_X1   g16193(.A1(new_n2864_), .A2(\b[58] ), .ZN(new_n16451_));
  AOI21_X1   g16194(.A1(new_n16450_), .A2(new_n16451_), .B(new_n2087_), .ZN(new_n16452_));
  NAND2_X1   g16195(.A1(new_n7929_), .A2(new_n16452_), .ZN(new_n16453_));
  XOR2_X1    g16196(.A1(new_n16453_), .A2(\a[29] ), .Z(new_n16454_));
  INV_X1     g16197(.I(new_n16454_), .ZN(new_n16455_));
  AOI21_X1   g16198(.A1(new_n16408_), .A2(new_n16406_), .B(new_n16404_), .ZN(new_n16456_));
  OAI22_X1   g16199(.A1(new_n2452_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n2447_), .ZN(new_n16457_));
  NAND2_X1   g16200(.A1(new_n3312_), .A2(\b[55] ), .ZN(new_n16458_));
  AOI21_X1   g16201(.A1(new_n16457_), .A2(new_n16458_), .B(new_n2455_), .ZN(new_n16459_));
  NAND2_X1   g16202(.A1(new_n7308_), .A2(new_n16459_), .ZN(new_n16460_));
  XOR2_X1    g16203(.A1(new_n16460_), .A2(\a[32] ), .Z(new_n16461_));
  INV_X1     g16204(.I(new_n16397_), .ZN(new_n16462_));
  AOI21_X1   g16205(.A1(new_n16400_), .A2(new_n16462_), .B(new_n16396_), .ZN(new_n16463_));
  INV_X1     g16206(.I(new_n16388_), .ZN(new_n16464_));
  AOI21_X1   g16207(.A1(new_n16384_), .A2(new_n16464_), .B(new_n16387_), .ZN(new_n16465_));
  AOI21_X1   g16208(.A1(new_n16360_), .A2(new_n16363_), .B(new_n16361_), .ZN(new_n16466_));
  AOI21_X1   g16209(.A1(new_n16343_), .A2(new_n16353_), .B(new_n16351_), .ZN(new_n16467_));
  NOR2_X1    g16210(.A1(new_n16338_), .A2(new_n16272_), .ZN(new_n16468_));
  NOR2_X1    g16211(.A1(new_n16468_), .A2(new_n16339_), .ZN(new_n16469_));
  AOI21_X1   g16212(.A1(new_n16320_), .A2(new_n16324_), .B(new_n16322_), .ZN(new_n16470_));
  AOI21_X1   g16213(.A1(new_n16302_), .A2(new_n16314_), .B(new_n16312_), .ZN(new_n16471_));
  NOR2_X1    g16214(.A1(new_n16290_), .A2(new_n16297_), .ZN(new_n16472_));
  NOR2_X1    g16215(.A1(new_n16472_), .A2(new_n16299_), .ZN(new_n16473_));
  OAI22_X1   g16216(.A1(new_n2039_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n1927_), .ZN(new_n16474_));
  NAND2_X1   g16217(.A1(new_n9644_), .A2(\b[25] ), .ZN(new_n16475_));
  AOI21_X1   g16218(.A1(new_n16475_), .A2(new_n16474_), .B(new_n8321_), .ZN(new_n16476_));
  NAND2_X1   g16219(.A1(new_n2042_), .A2(new_n16476_), .ZN(new_n16477_));
  XOR2_X1    g16220(.A1(new_n16477_), .A2(\a[62] ), .Z(new_n16478_));
  INV_X1     g16221(.I(new_n16478_), .ZN(new_n16479_));
  NOR2_X1    g16222(.A1(new_n8985_), .A2(new_n1709_), .ZN(new_n16480_));
  NOR2_X1    g16223(.A1(new_n9364_), .A2(new_n1601_), .ZN(new_n16481_));
  XNOR2_X1   g16224(.A1(new_n16480_), .A2(new_n16481_), .ZN(new_n16482_));
  XOR2_X1    g16225(.A1(new_n16482_), .A2(\a[23] ), .Z(new_n16483_));
  NOR2_X1    g16226(.A1(new_n16483_), .A2(new_n16294_), .ZN(new_n16484_));
  NOR2_X1    g16227(.A1(new_n16482_), .A2(new_n1434_), .ZN(new_n16485_));
  INV_X1     g16228(.I(new_n16485_), .ZN(new_n16486_));
  NAND2_X1   g16229(.A1(new_n16482_), .A2(new_n1434_), .ZN(new_n16487_));
  AOI21_X1   g16230(.A1(new_n16486_), .A2(new_n16487_), .B(new_n16298_), .ZN(new_n16488_));
  NOR2_X1    g16231(.A1(new_n16484_), .A2(new_n16488_), .ZN(new_n16489_));
  NOR2_X1    g16232(.A1(new_n16479_), .A2(new_n16489_), .ZN(new_n16490_));
  INV_X1     g16233(.I(new_n16490_), .ZN(new_n16491_));
  NAND2_X1   g16234(.A1(new_n16479_), .A2(new_n16489_), .ZN(new_n16492_));
  AOI21_X1   g16235(.A1(new_n16491_), .A2(new_n16492_), .B(new_n16473_), .ZN(new_n16493_));
  XOR2_X1    g16236(.A1(new_n16478_), .A2(new_n16489_), .Z(new_n16494_));
  INV_X1     g16237(.I(new_n16494_), .ZN(new_n16495_));
  AOI21_X1   g16238(.A1(new_n16473_), .A2(new_n16495_), .B(new_n16493_), .ZN(new_n16496_));
  OAI22_X1   g16239(.A1(new_n2405_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2272_), .ZN(new_n16497_));
  NAND2_X1   g16240(.A1(new_n8628_), .A2(\b[28] ), .ZN(new_n16498_));
  AOI21_X1   g16241(.A1(new_n16498_), .A2(new_n16497_), .B(new_n7354_), .ZN(new_n16499_));
  NAND2_X1   g16242(.A1(new_n2404_), .A2(new_n16499_), .ZN(new_n16500_));
  XOR2_X1    g16243(.A1(new_n16500_), .A2(\a[59] ), .Z(new_n16501_));
  XNOR2_X1   g16244(.A1(new_n16496_), .A2(new_n16501_), .ZN(new_n16502_));
  NOR2_X1    g16245(.A1(new_n16502_), .A2(new_n16471_), .ZN(new_n16503_));
  INV_X1     g16246(.I(new_n16471_), .ZN(new_n16504_));
  NOR2_X1    g16247(.A1(new_n16496_), .A2(new_n16501_), .ZN(new_n16505_));
  INV_X1     g16248(.I(new_n16505_), .ZN(new_n16506_));
  NAND2_X1   g16249(.A1(new_n16496_), .A2(new_n16501_), .ZN(new_n16507_));
  AOI21_X1   g16250(.A1(new_n16506_), .A2(new_n16507_), .B(new_n16504_), .ZN(new_n16508_));
  NOR2_X1    g16251(.A1(new_n16503_), .A2(new_n16508_), .ZN(new_n16509_));
  OAI22_X1   g16252(.A1(new_n6721_), .A2(new_n2660_), .B1(new_n6723_), .B2(new_n2794_), .ZN(new_n16510_));
  NAND2_X1   g16253(.A1(new_n7617_), .A2(\b[31] ), .ZN(new_n16511_));
  AOI21_X1   g16254(.A1(new_n16511_), .A2(new_n16510_), .B(new_n6731_), .ZN(new_n16512_));
  NAND2_X1   g16255(.A1(new_n2797_), .A2(new_n16512_), .ZN(new_n16513_));
  XOR2_X1    g16256(.A1(new_n16513_), .A2(\a[56] ), .Z(new_n16514_));
  XOR2_X1    g16257(.A1(new_n16509_), .A2(new_n16514_), .Z(new_n16515_));
  NOR2_X1    g16258(.A1(new_n16515_), .A2(new_n16470_), .ZN(new_n16516_));
  INV_X1     g16259(.I(new_n16470_), .ZN(new_n16517_));
  INV_X1     g16260(.I(new_n16509_), .ZN(new_n16518_));
  NOR2_X1    g16261(.A1(new_n16518_), .A2(new_n16514_), .ZN(new_n16519_));
  INV_X1     g16262(.I(new_n16519_), .ZN(new_n16520_));
  NAND2_X1   g16263(.A1(new_n16518_), .A2(new_n16514_), .ZN(new_n16521_));
  AOI21_X1   g16264(.A1(new_n16520_), .A2(new_n16521_), .B(new_n16517_), .ZN(new_n16522_));
  NOR2_X1    g16265(.A1(new_n16522_), .A2(new_n16516_), .ZN(new_n16523_));
  OAI22_X1   g16266(.A1(new_n5786_), .A2(new_n3247_), .B1(new_n3097_), .B2(new_n5792_), .ZN(new_n16524_));
  NAND2_X1   g16267(.A1(new_n6745_), .A2(\b[34] ), .ZN(new_n16525_));
  AOI21_X1   g16268(.A1(new_n16525_), .A2(new_n16524_), .B(new_n5796_), .ZN(new_n16526_));
  NAND2_X1   g16269(.A1(new_n3246_), .A2(new_n16526_), .ZN(new_n16527_));
  XOR2_X1    g16270(.A1(new_n16527_), .A2(\a[53] ), .Z(new_n16528_));
  NAND2_X1   g16271(.A1(new_n16335_), .A2(new_n16331_), .ZN(new_n16529_));
  NAND2_X1   g16272(.A1(new_n16529_), .A2(new_n16334_), .ZN(new_n16530_));
  INV_X1     g16273(.I(new_n16530_), .ZN(new_n16531_));
  NOR2_X1    g16274(.A1(new_n16531_), .A2(new_n16528_), .ZN(new_n16532_));
  INV_X1     g16275(.I(new_n16528_), .ZN(new_n16533_));
  NOR2_X1    g16276(.A1(new_n16530_), .A2(new_n16533_), .ZN(new_n16534_));
  NOR2_X1    g16277(.A1(new_n16532_), .A2(new_n16534_), .ZN(new_n16535_));
  NOR2_X1    g16278(.A1(new_n16535_), .A2(new_n16523_), .ZN(new_n16536_));
  XOR2_X1    g16279(.A1(new_n16530_), .A2(new_n16528_), .Z(new_n16537_));
  NOR3_X1    g16280(.A1(new_n16537_), .A2(new_n16516_), .A3(new_n16522_), .ZN(new_n16538_));
  NOR2_X1    g16281(.A1(new_n16536_), .A2(new_n16538_), .ZN(new_n16539_));
  OAI22_X1   g16282(.A1(new_n5228_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n5225_), .ZN(new_n16540_));
  NAND2_X1   g16283(.A1(new_n5387_), .A2(\b[37] ), .ZN(new_n16541_));
  AOI21_X1   g16284(.A1(new_n16540_), .A2(new_n16541_), .B(new_n5231_), .ZN(new_n16542_));
  NAND2_X1   g16285(.A1(new_n3700_), .A2(new_n16542_), .ZN(new_n16543_));
  XOR2_X1    g16286(.A1(new_n16543_), .A2(\a[50] ), .Z(new_n16544_));
  XOR2_X1    g16287(.A1(new_n16539_), .A2(new_n16544_), .Z(new_n16545_));
  NOR3_X1    g16288(.A1(new_n16536_), .A2(new_n16538_), .A3(new_n16544_), .ZN(new_n16546_));
  INV_X1     g16289(.I(new_n16544_), .ZN(new_n16547_));
  NOR2_X1    g16290(.A1(new_n16539_), .A2(new_n16547_), .ZN(new_n16548_));
  OAI21_X1   g16291(.A1(new_n16548_), .A2(new_n16546_), .B(new_n16469_), .ZN(new_n16549_));
  OAI21_X1   g16292(.A1(new_n16545_), .A2(new_n16469_), .B(new_n16549_), .ZN(new_n16550_));
  OAI22_X1   g16293(.A1(new_n4711_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n4706_), .ZN(new_n16551_));
  NAND2_X1   g16294(.A1(new_n5814_), .A2(\b[40] ), .ZN(new_n16552_));
  AOI21_X1   g16295(.A1(new_n16551_), .A2(new_n16552_), .B(new_n4714_), .ZN(new_n16553_));
  NAND2_X1   g16296(.A1(new_n4017_), .A2(new_n16553_), .ZN(new_n16554_));
  XOR2_X1    g16297(.A1(new_n16554_), .A2(\a[47] ), .Z(new_n16555_));
  NOR2_X1    g16298(.A1(new_n16550_), .A2(new_n16555_), .ZN(new_n16556_));
  INV_X1     g16299(.I(new_n16556_), .ZN(new_n16557_));
  NAND2_X1   g16300(.A1(new_n16550_), .A2(new_n16555_), .ZN(new_n16558_));
  AOI21_X1   g16301(.A1(new_n16557_), .A2(new_n16558_), .B(new_n16467_), .ZN(new_n16559_));
  INV_X1     g16302(.I(new_n16467_), .ZN(new_n16560_));
  XNOR2_X1   g16303(.A1(new_n16550_), .A2(new_n16555_), .ZN(new_n16561_));
  NOR2_X1    g16304(.A1(new_n16561_), .A2(new_n16560_), .ZN(new_n16562_));
  NOR2_X1    g16305(.A1(new_n16562_), .A2(new_n16559_), .ZN(new_n16563_));
  OAI22_X1   g16306(.A1(new_n4208_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n4203_), .ZN(new_n16564_));
  NAND2_X1   g16307(.A1(new_n5244_), .A2(\b[43] ), .ZN(new_n16565_));
  AOI21_X1   g16308(.A1(new_n16564_), .A2(new_n16565_), .B(new_n4211_), .ZN(new_n16566_));
  NAND2_X1   g16309(.A1(new_n4513_), .A2(new_n16566_), .ZN(new_n16567_));
  XOR2_X1    g16310(.A1(new_n16567_), .A2(\a[44] ), .Z(new_n16568_));
  XNOR2_X1   g16311(.A1(new_n16563_), .A2(new_n16568_), .ZN(new_n16569_));
  NOR2_X1    g16312(.A1(new_n16569_), .A2(new_n16466_), .ZN(new_n16570_));
  INV_X1     g16313(.I(new_n16466_), .ZN(new_n16571_));
  NOR2_X1    g16314(.A1(new_n16563_), .A2(new_n16568_), .ZN(new_n16572_));
  INV_X1     g16315(.I(new_n16572_), .ZN(new_n16573_));
  NAND2_X1   g16316(.A1(new_n16563_), .A2(new_n16568_), .ZN(new_n16574_));
  AOI21_X1   g16317(.A1(new_n16573_), .A2(new_n16574_), .B(new_n16571_), .ZN(new_n16575_));
  NOR2_X1    g16318(.A1(new_n16570_), .A2(new_n16575_), .ZN(new_n16576_));
  INV_X1     g16319(.I(new_n16576_), .ZN(new_n16577_));
  OAI22_X1   g16320(.A1(new_n3736_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n3731_), .ZN(new_n16578_));
  NAND2_X1   g16321(.A1(new_n4730_), .A2(\b[46] ), .ZN(new_n16579_));
  AOI21_X1   g16322(.A1(new_n16578_), .A2(new_n16579_), .B(new_n3739_), .ZN(new_n16580_));
  NAND2_X1   g16323(.A1(new_n5177_), .A2(new_n16580_), .ZN(new_n16581_));
  XOR2_X1    g16324(.A1(new_n16581_), .A2(\a[41] ), .Z(new_n16582_));
  NOR2_X1    g16325(.A1(new_n16366_), .A2(new_n16378_), .ZN(new_n16583_));
  NOR2_X1    g16326(.A1(new_n16583_), .A2(new_n16377_), .ZN(new_n16584_));
  NOR2_X1    g16327(.A1(new_n16584_), .A2(new_n16582_), .ZN(new_n16585_));
  INV_X1     g16328(.I(new_n16582_), .ZN(new_n16586_));
  NOR3_X1    g16329(.A1(new_n16583_), .A2(new_n16377_), .A3(new_n16586_), .ZN(new_n16587_));
  OAI21_X1   g16330(.A1(new_n16585_), .A2(new_n16587_), .B(new_n16577_), .ZN(new_n16588_));
  XOR2_X1    g16331(.A1(new_n16584_), .A2(new_n16586_), .Z(new_n16589_));
  OAI21_X1   g16332(.A1(new_n16577_), .A2(new_n16589_), .B(new_n16588_), .ZN(new_n16590_));
  OAI22_X1   g16333(.A1(new_n3298_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n3293_), .ZN(new_n16591_));
  NAND2_X1   g16334(.A1(new_n4227_), .A2(\b[49] ), .ZN(new_n16592_));
  AOI21_X1   g16335(.A1(new_n16591_), .A2(new_n16592_), .B(new_n3301_), .ZN(new_n16593_));
  NAND2_X1   g16336(.A1(new_n5741_), .A2(new_n16593_), .ZN(new_n16594_));
  XOR2_X1    g16337(.A1(new_n16594_), .A2(\a[38] ), .Z(new_n16595_));
  NOR2_X1    g16338(.A1(new_n16590_), .A2(new_n16595_), .ZN(new_n16596_));
  INV_X1     g16339(.I(new_n16596_), .ZN(new_n16597_));
  NAND2_X1   g16340(.A1(new_n16590_), .A2(new_n16595_), .ZN(new_n16598_));
  AOI21_X1   g16341(.A1(new_n16597_), .A2(new_n16598_), .B(new_n16465_), .ZN(new_n16599_));
  INV_X1     g16342(.I(new_n16465_), .ZN(new_n16600_));
  XNOR2_X1   g16343(.A1(new_n16590_), .A2(new_n16595_), .ZN(new_n16601_));
  NOR2_X1    g16344(.A1(new_n16601_), .A2(new_n16600_), .ZN(new_n16602_));
  NOR2_X1    g16345(.A1(new_n16602_), .A2(new_n16599_), .ZN(new_n16603_));
  OAI22_X1   g16346(.A1(new_n2846_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n2841_), .ZN(new_n16604_));
  NAND2_X1   g16347(.A1(new_n3755_), .A2(\b[52] ), .ZN(new_n16605_));
  AOI21_X1   g16348(.A1(new_n16604_), .A2(new_n16605_), .B(new_n2849_), .ZN(new_n16606_));
  NAND2_X1   g16349(.A1(new_n6237_), .A2(new_n16606_), .ZN(new_n16607_));
  XOR2_X1    g16350(.A1(new_n16607_), .A2(\a[35] ), .Z(new_n16608_));
  XNOR2_X1   g16351(.A1(new_n16603_), .A2(new_n16608_), .ZN(new_n16609_));
  NOR2_X1    g16352(.A1(new_n16609_), .A2(new_n16463_), .ZN(new_n16610_));
  INV_X1     g16353(.I(new_n16463_), .ZN(new_n16611_));
  NOR2_X1    g16354(.A1(new_n16603_), .A2(new_n16608_), .ZN(new_n16612_));
  INV_X1     g16355(.I(new_n16612_), .ZN(new_n16613_));
  NAND2_X1   g16356(.A1(new_n16603_), .A2(new_n16608_), .ZN(new_n16614_));
  AOI21_X1   g16357(.A1(new_n16613_), .A2(new_n16614_), .B(new_n16611_), .ZN(new_n16615_));
  NOR2_X1    g16358(.A1(new_n16610_), .A2(new_n16615_), .ZN(new_n16616_));
  XOR2_X1    g16359(.A1(new_n16616_), .A2(new_n16461_), .Z(new_n16617_));
  NOR2_X1    g16360(.A1(new_n16617_), .A2(new_n16456_), .ZN(new_n16618_));
  INV_X1     g16361(.I(new_n16456_), .ZN(new_n16619_));
  INV_X1     g16362(.I(new_n16461_), .ZN(new_n16620_));
  NOR2_X1    g16363(.A1(new_n16616_), .A2(new_n16620_), .ZN(new_n16621_));
  INV_X1     g16364(.I(new_n16621_), .ZN(new_n16622_));
  NAND2_X1   g16365(.A1(new_n16616_), .A2(new_n16620_), .ZN(new_n16623_));
  AOI21_X1   g16366(.A1(new_n16622_), .A2(new_n16623_), .B(new_n16619_), .ZN(new_n16624_));
  NOR2_X1    g16367(.A1(new_n16618_), .A2(new_n16624_), .ZN(new_n16625_));
  NOR2_X1    g16368(.A1(new_n16625_), .A2(new_n16455_), .ZN(new_n16626_));
  INV_X1     g16369(.I(new_n16625_), .ZN(new_n16627_));
  NOR2_X1    g16370(.A1(new_n16627_), .A2(new_n16454_), .ZN(new_n16628_));
  NOR2_X1    g16371(.A1(new_n16628_), .A2(new_n16626_), .ZN(new_n16629_));
  NOR2_X1    g16372(.A1(new_n16629_), .A2(new_n16449_), .ZN(new_n16630_));
  INV_X1     g16373(.I(new_n16449_), .ZN(new_n16631_));
  XOR2_X1    g16374(.A1(new_n16625_), .A2(new_n16454_), .Z(new_n16632_));
  NOR2_X1    g16375(.A1(new_n16632_), .A2(new_n16631_), .ZN(new_n16633_));
  NOR2_X1    g16376(.A1(new_n16630_), .A2(new_n16633_), .ZN(new_n16634_));
  NOR2_X1    g16377(.A1(new_n16634_), .A2(new_n16448_), .ZN(new_n16635_));
  INV_X1     g16378(.I(new_n16635_), .ZN(new_n16636_));
  NAND2_X1   g16379(.A1(new_n16634_), .A2(new_n16448_), .ZN(new_n16637_));
  NAND2_X1   g16380(.A1(new_n16636_), .A2(new_n16637_), .ZN(new_n16638_));
  XNOR2_X1   g16381(.A1(new_n16634_), .A2(new_n16448_), .ZN(new_n16639_));
  NOR2_X1    g16382(.A1(new_n16639_), .A2(new_n16443_), .ZN(new_n16640_));
  AOI21_X1   g16383(.A1(new_n16443_), .A2(new_n16638_), .B(new_n16640_), .ZN(new_n16641_));
  NOR2_X1    g16384(.A1(new_n16641_), .A2(new_n16439_), .ZN(new_n16642_));
  NAND2_X1   g16385(.A1(new_n16641_), .A2(new_n16439_), .ZN(new_n16643_));
  INV_X1     g16386(.I(new_n16643_), .ZN(new_n16644_));
  NOR2_X1    g16387(.A1(new_n16644_), .A2(new_n16642_), .ZN(new_n16645_));
  INV_X1     g16388(.I(new_n16223_), .ZN(new_n16646_));
  OAI21_X1   g16389(.A1(new_n16009_), .A2(new_n16646_), .B(new_n16232_), .ZN(new_n16647_));
  NAND3_X1   g16390(.A1(new_n16647_), .A2(new_n16230_), .A3(new_n16434_), .ZN(new_n16648_));
  NAND2_X1   g16391(.A1(new_n16648_), .A2(new_n16432_), .ZN(new_n16649_));
  XOR2_X1    g16392(.A1(new_n16649_), .A2(new_n16645_), .Z(\f[87] ));
  AOI21_X1   g16393(.A1(new_n16443_), .A2(new_n16637_), .B(new_n16635_), .ZN(new_n16651_));
  NOR2_X1    g16394(.A1(new_n1857_), .A2(new_n8932_), .ZN(new_n16652_));
  NOR2_X1    g16395(.A1(new_n1755_), .A2(new_n8956_), .ZN(new_n16653_));
  NOR4_X1    g16396(.A1(new_n9323_), .A2(new_n1763_), .A3(new_n16652_), .A4(new_n16653_), .ZN(new_n16654_));
  XOR2_X1    g16397(.A1(new_n16654_), .A2(new_n1750_), .Z(new_n16655_));
  OAI22_X1   g16398(.A1(new_n2084_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n2079_), .ZN(new_n16656_));
  NAND2_X1   g16399(.A1(new_n2864_), .A2(\b[59] ), .ZN(new_n16657_));
  AOI21_X1   g16400(.A1(new_n16656_), .A2(new_n16657_), .B(new_n2087_), .ZN(new_n16658_));
  NAND2_X1   g16401(.A1(new_n8550_), .A2(new_n16658_), .ZN(new_n16659_));
  XOR2_X1    g16402(.A1(new_n16659_), .A2(\a[29] ), .Z(new_n16660_));
  INV_X1     g16403(.I(new_n16660_), .ZN(new_n16661_));
  OAI21_X1   g16404(.A1(new_n16456_), .A2(new_n16621_), .B(new_n16623_), .ZN(new_n16662_));
  OAI22_X1   g16405(.A1(new_n2452_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n2447_), .ZN(new_n16663_));
  NAND2_X1   g16406(.A1(new_n3312_), .A2(\b[56] ), .ZN(new_n16664_));
  AOI21_X1   g16407(.A1(new_n16663_), .A2(new_n16664_), .B(new_n2455_), .ZN(new_n16665_));
  NAND2_X1   g16408(.A1(new_n7559_), .A2(new_n16665_), .ZN(new_n16666_));
  XOR2_X1    g16409(.A1(new_n16666_), .A2(\a[32] ), .Z(new_n16667_));
  AOI21_X1   g16410(.A1(new_n16611_), .A2(new_n16614_), .B(new_n16612_), .ZN(new_n16668_));
  AOI21_X1   g16411(.A1(new_n16600_), .A2(new_n16598_), .B(new_n16596_), .ZN(new_n16669_));
  OAI22_X1   g16412(.A1(new_n3298_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n3293_), .ZN(new_n16670_));
  NAND2_X1   g16413(.A1(new_n4227_), .A2(\b[50] ), .ZN(new_n16671_));
  AOI21_X1   g16414(.A1(new_n16670_), .A2(new_n16671_), .B(new_n3301_), .ZN(new_n16672_));
  NAND2_X1   g16415(.A1(new_n5954_), .A2(new_n16672_), .ZN(new_n16673_));
  XOR2_X1    g16416(.A1(new_n16673_), .A2(\a[38] ), .Z(new_n16674_));
  OAI22_X1   g16417(.A1(new_n4208_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n4203_), .ZN(new_n16675_));
  NAND2_X1   g16418(.A1(new_n5244_), .A2(\b[44] ), .ZN(new_n16676_));
  AOI21_X1   g16419(.A1(new_n16675_), .A2(new_n16676_), .B(new_n4211_), .ZN(new_n16677_));
  NAND2_X1   g16420(.A1(new_n4833_), .A2(new_n16677_), .ZN(new_n16678_));
  XOR2_X1    g16421(.A1(new_n16678_), .A2(\a[44] ), .Z(new_n16679_));
  NOR2_X1    g16422(.A1(new_n16548_), .A2(new_n16469_), .ZN(new_n16680_));
  NOR2_X1    g16423(.A1(new_n16680_), .A2(new_n16546_), .ZN(new_n16681_));
  OAI22_X1   g16424(.A1(new_n5228_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n5225_), .ZN(new_n16682_));
  NAND2_X1   g16425(.A1(new_n5387_), .A2(\b[38] ), .ZN(new_n16683_));
  AOI21_X1   g16426(.A1(new_n16682_), .A2(new_n16683_), .B(new_n5231_), .ZN(new_n16684_));
  NAND2_X1   g16427(.A1(new_n3844_), .A2(new_n16684_), .ZN(new_n16685_));
  XOR2_X1    g16428(.A1(new_n16685_), .A2(\a[50] ), .Z(new_n16686_));
  INV_X1     g16429(.I(new_n16534_), .ZN(new_n16687_));
  AOI21_X1   g16430(.A1(new_n16523_), .A2(new_n16687_), .B(new_n16532_), .ZN(new_n16688_));
  OAI22_X1   g16431(.A1(new_n6721_), .A2(new_n2794_), .B1(new_n6723_), .B2(new_n2964_), .ZN(new_n16689_));
  NAND2_X1   g16432(.A1(new_n7617_), .A2(\b[32] ), .ZN(new_n16690_));
  AOI21_X1   g16433(.A1(new_n16690_), .A2(new_n16689_), .B(new_n6731_), .ZN(new_n16691_));
  NAND2_X1   g16434(.A1(new_n2963_), .A2(new_n16691_), .ZN(new_n16692_));
  XOR2_X1    g16435(.A1(new_n16692_), .A2(\a[56] ), .Z(new_n16693_));
  INV_X1     g16436(.I(new_n16693_), .ZN(new_n16694_));
  OAI21_X1   g16437(.A1(new_n16473_), .A2(new_n16490_), .B(new_n16492_), .ZN(new_n16695_));
  INV_X1     g16438(.I(new_n16695_), .ZN(new_n16696_));
  OAI22_X1   g16439(.A1(new_n2175_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2039_), .ZN(new_n16697_));
  NAND2_X1   g16440(.A1(new_n9644_), .A2(\b[26] ), .ZN(new_n16698_));
  AOI21_X1   g16441(.A1(new_n16698_), .A2(new_n16697_), .B(new_n8321_), .ZN(new_n16699_));
  NAND2_X1   g16442(.A1(new_n2174_), .A2(new_n16699_), .ZN(new_n16700_));
  XOR2_X1    g16443(.A1(new_n16700_), .A2(new_n8309_), .Z(new_n16701_));
  NAND2_X1   g16444(.A1(new_n16487_), .A2(new_n16298_), .ZN(new_n16702_));
  NAND2_X1   g16445(.A1(new_n16702_), .A2(new_n16486_), .ZN(new_n16703_));
  NOR3_X1    g16446(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n1709_), .ZN(new_n16704_));
  NOR2_X1    g16447(.A1(new_n9364_), .A2(new_n1709_), .ZN(new_n16705_));
  NOR3_X1    g16448(.A1(new_n16705_), .A2(new_n1825_), .A3(new_n8985_), .ZN(new_n16706_));
  NOR2_X1    g16449(.A1(new_n16706_), .A2(new_n16704_), .ZN(new_n16707_));
  INV_X1     g16450(.I(new_n16707_), .ZN(new_n16708_));
  XOR2_X1    g16451(.A1(new_n16703_), .A2(new_n16708_), .Z(new_n16709_));
  INV_X1     g16452(.I(new_n16709_), .ZN(new_n16710_));
  NOR2_X1    g16453(.A1(new_n16703_), .A2(new_n16707_), .ZN(new_n16711_));
  INV_X1     g16454(.I(new_n16711_), .ZN(new_n16712_));
  NAND2_X1   g16455(.A1(new_n16703_), .A2(new_n16707_), .ZN(new_n16713_));
  AOI21_X1   g16456(.A1(new_n16712_), .A2(new_n16713_), .B(new_n16701_), .ZN(new_n16714_));
  AOI21_X1   g16457(.A1(new_n16701_), .A2(new_n16710_), .B(new_n16714_), .ZN(new_n16715_));
  INV_X1     g16458(.I(new_n16715_), .ZN(new_n16716_));
  OAI22_X1   g16459(.A1(new_n2543_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2405_), .ZN(new_n16717_));
  NAND2_X1   g16460(.A1(new_n8628_), .A2(\b[29] ), .ZN(new_n16718_));
  AOI21_X1   g16461(.A1(new_n16718_), .A2(new_n16717_), .B(new_n7354_), .ZN(new_n16719_));
  NAND2_X1   g16462(.A1(new_n2546_), .A2(new_n16719_), .ZN(new_n16720_));
  XOR2_X1    g16463(.A1(new_n16720_), .A2(\a[59] ), .Z(new_n16721_));
  NOR2_X1    g16464(.A1(new_n16721_), .A2(new_n16716_), .ZN(new_n16722_));
  AND2_X2    g16465(.A1(new_n16721_), .A2(new_n16716_), .Z(new_n16723_));
  NOR2_X1    g16466(.A1(new_n16723_), .A2(new_n16722_), .ZN(new_n16724_));
  NOR2_X1    g16467(.A1(new_n16724_), .A2(new_n16696_), .ZN(new_n16725_));
  XOR2_X1    g16468(.A1(new_n16721_), .A2(new_n16715_), .Z(new_n16726_));
  NOR2_X1    g16469(.A1(new_n16726_), .A2(new_n16695_), .ZN(new_n16727_));
  NOR2_X1    g16470(.A1(new_n16725_), .A2(new_n16727_), .ZN(new_n16728_));
  NAND2_X1   g16471(.A1(new_n16507_), .A2(new_n16504_), .ZN(new_n16729_));
  NAND2_X1   g16472(.A1(new_n16729_), .A2(new_n16506_), .ZN(new_n16730_));
  INV_X1     g16473(.I(new_n16730_), .ZN(new_n16731_));
  NOR2_X1    g16474(.A1(new_n16731_), .A2(new_n16728_), .ZN(new_n16732_));
  INV_X1     g16475(.I(new_n16728_), .ZN(new_n16733_));
  NOR2_X1    g16476(.A1(new_n16733_), .A2(new_n16730_), .ZN(new_n16734_));
  OAI21_X1   g16477(.A1(new_n16734_), .A2(new_n16732_), .B(new_n16694_), .ZN(new_n16735_));
  XNOR2_X1   g16478(.A1(new_n16728_), .A2(new_n16730_), .ZN(new_n16736_));
  NAND2_X1   g16479(.A1(new_n16736_), .A2(new_n16693_), .ZN(new_n16737_));
  NAND2_X1   g16480(.A1(new_n16737_), .A2(new_n16735_), .ZN(new_n16738_));
  NAND2_X1   g16481(.A1(new_n16521_), .A2(new_n16517_), .ZN(new_n16739_));
  NAND2_X1   g16482(.A1(new_n16739_), .A2(new_n16520_), .ZN(new_n16740_));
  OAI22_X1   g16483(.A1(new_n5786_), .A2(new_n3408_), .B1(new_n3247_), .B2(new_n5792_), .ZN(new_n16741_));
  NAND2_X1   g16484(.A1(new_n6745_), .A2(\b[35] ), .ZN(new_n16742_));
  AOI21_X1   g16485(.A1(new_n16742_), .A2(new_n16741_), .B(new_n5796_), .ZN(new_n16743_));
  NAND2_X1   g16486(.A1(new_n3411_), .A2(new_n16743_), .ZN(new_n16744_));
  XOR2_X1    g16487(.A1(new_n16744_), .A2(\a[53] ), .Z(new_n16745_));
  INV_X1     g16488(.I(new_n16745_), .ZN(new_n16746_));
  XOR2_X1    g16489(.A1(new_n16740_), .A2(new_n16746_), .Z(new_n16747_));
  NAND2_X1   g16490(.A1(new_n16747_), .A2(new_n16738_), .ZN(new_n16748_));
  INV_X1     g16491(.I(new_n16738_), .ZN(new_n16749_));
  AOI21_X1   g16492(.A1(new_n16739_), .A2(new_n16520_), .B(new_n16745_), .ZN(new_n16750_));
  NOR2_X1    g16493(.A1(new_n16740_), .A2(new_n16746_), .ZN(new_n16751_));
  OAI21_X1   g16494(.A1(new_n16751_), .A2(new_n16750_), .B(new_n16749_), .ZN(new_n16752_));
  NAND2_X1   g16495(.A1(new_n16748_), .A2(new_n16752_), .ZN(new_n16753_));
  XNOR2_X1   g16496(.A1(new_n16688_), .A2(new_n16753_), .ZN(new_n16754_));
  AND2_X2    g16497(.A1(new_n16688_), .A2(new_n16753_), .Z(new_n16755_));
  NOR2_X1    g16498(.A1(new_n16688_), .A2(new_n16753_), .ZN(new_n16756_));
  OAI21_X1   g16499(.A1(new_n16755_), .A2(new_n16756_), .B(new_n16686_), .ZN(new_n16757_));
  OAI21_X1   g16500(.A1(new_n16686_), .A2(new_n16754_), .B(new_n16757_), .ZN(new_n16758_));
  OAI22_X1   g16501(.A1(new_n4711_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n4706_), .ZN(new_n16759_));
  NAND2_X1   g16502(.A1(new_n5814_), .A2(\b[41] ), .ZN(new_n16760_));
  AOI21_X1   g16503(.A1(new_n16759_), .A2(new_n16760_), .B(new_n4714_), .ZN(new_n16761_));
  NAND2_X1   g16504(.A1(new_n4320_), .A2(new_n16761_), .ZN(new_n16762_));
  XOR2_X1    g16505(.A1(new_n16762_), .A2(\a[47] ), .Z(new_n16763_));
  NOR2_X1    g16506(.A1(new_n16758_), .A2(new_n16763_), .ZN(new_n16764_));
  INV_X1     g16507(.I(new_n16764_), .ZN(new_n16765_));
  NAND2_X1   g16508(.A1(new_n16758_), .A2(new_n16763_), .ZN(new_n16766_));
  AOI21_X1   g16509(.A1(new_n16765_), .A2(new_n16766_), .B(new_n16681_), .ZN(new_n16767_));
  INV_X1     g16510(.I(new_n16681_), .ZN(new_n16768_));
  XNOR2_X1   g16511(.A1(new_n16758_), .A2(new_n16763_), .ZN(new_n16769_));
  NOR2_X1    g16512(.A1(new_n16769_), .A2(new_n16768_), .ZN(new_n16770_));
  NOR2_X1    g16513(.A1(new_n16770_), .A2(new_n16767_), .ZN(new_n16771_));
  AOI21_X1   g16514(.A1(new_n16560_), .A2(new_n16558_), .B(new_n16556_), .ZN(new_n16772_));
  NOR2_X1    g16515(.A1(new_n16771_), .A2(new_n16772_), .ZN(new_n16773_));
  INV_X1     g16516(.I(new_n16773_), .ZN(new_n16774_));
  NAND2_X1   g16517(.A1(new_n16771_), .A2(new_n16772_), .ZN(new_n16775_));
  AOI21_X1   g16518(.A1(new_n16774_), .A2(new_n16775_), .B(new_n16679_), .ZN(new_n16776_));
  INV_X1     g16519(.I(new_n16679_), .ZN(new_n16777_));
  XNOR2_X1   g16520(.A1(new_n16771_), .A2(new_n16772_), .ZN(new_n16778_));
  NOR2_X1    g16521(.A1(new_n16778_), .A2(new_n16777_), .ZN(new_n16779_));
  NOR2_X1    g16522(.A1(new_n16779_), .A2(new_n16776_), .ZN(new_n16780_));
  NAND2_X1   g16523(.A1(new_n16574_), .A2(new_n16571_), .ZN(new_n16781_));
  NAND2_X1   g16524(.A1(new_n16781_), .A2(new_n16573_), .ZN(new_n16782_));
  INV_X1     g16525(.I(new_n16782_), .ZN(new_n16783_));
  OAI22_X1   g16526(.A1(new_n3736_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n3731_), .ZN(new_n16784_));
  NAND2_X1   g16527(.A1(new_n4730_), .A2(\b[47] ), .ZN(new_n16785_));
  AOI21_X1   g16528(.A1(new_n16784_), .A2(new_n16785_), .B(new_n3739_), .ZN(new_n16786_));
  NAND2_X1   g16529(.A1(new_n5196_), .A2(new_n16786_), .ZN(new_n16787_));
  XOR2_X1    g16530(.A1(new_n16787_), .A2(\a[41] ), .Z(new_n16788_));
  NOR2_X1    g16531(.A1(new_n16783_), .A2(new_n16788_), .ZN(new_n16789_));
  INV_X1     g16532(.I(new_n16789_), .ZN(new_n16790_));
  NAND2_X1   g16533(.A1(new_n16783_), .A2(new_n16788_), .ZN(new_n16791_));
  AOI21_X1   g16534(.A1(new_n16790_), .A2(new_n16791_), .B(new_n16780_), .ZN(new_n16792_));
  XNOR2_X1   g16535(.A1(new_n16782_), .A2(new_n16788_), .ZN(new_n16793_));
  AOI21_X1   g16536(.A1(new_n16780_), .A2(new_n16793_), .B(new_n16792_), .ZN(new_n16794_));
  NOR2_X1    g16537(.A1(new_n16577_), .A2(new_n16587_), .ZN(new_n16795_));
  NOR2_X1    g16538(.A1(new_n16795_), .A2(new_n16585_), .ZN(new_n16796_));
  NOR2_X1    g16539(.A1(new_n16794_), .A2(new_n16796_), .ZN(new_n16797_));
  INV_X1     g16540(.I(new_n16797_), .ZN(new_n16798_));
  NAND2_X1   g16541(.A1(new_n16794_), .A2(new_n16796_), .ZN(new_n16799_));
  AOI21_X1   g16542(.A1(new_n16798_), .A2(new_n16799_), .B(new_n16674_), .ZN(new_n16800_));
  INV_X1     g16543(.I(new_n16674_), .ZN(new_n16801_));
  XNOR2_X1   g16544(.A1(new_n16794_), .A2(new_n16796_), .ZN(new_n16802_));
  NOR2_X1    g16545(.A1(new_n16802_), .A2(new_n16801_), .ZN(new_n16803_));
  NOR2_X1    g16546(.A1(new_n16803_), .A2(new_n16800_), .ZN(new_n16804_));
  OAI22_X1   g16547(.A1(new_n2846_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n2841_), .ZN(new_n16805_));
  NAND2_X1   g16548(.A1(new_n3755_), .A2(\b[53] ), .ZN(new_n16806_));
  AOI21_X1   g16549(.A1(new_n16805_), .A2(new_n16806_), .B(new_n2849_), .ZN(new_n16807_));
  NAND2_X1   g16550(.A1(new_n6471_), .A2(new_n16807_), .ZN(new_n16808_));
  XOR2_X1    g16551(.A1(new_n16808_), .A2(\a[35] ), .Z(new_n16809_));
  XNOR2_X1   g16552(.A1(new_n16804_), .A2(new_n16809_), .ZN(new_n16810_));
  NOR2_X1    g16553(.A1(new_n16810_), .A2(new_n16669_), .ZN(new_n16811_));
  INV_X1     g16554(.I(new_n16669_), .ZN(new_n16812_));
  NOR2_X1    g16555(.A1(new_n16804_), .A2(new_n16809_), .ZN(new_n16813_));
  INV_X1     g16556(.I(new_n16813_), .ZN(new_n16814_));
  NAND2_X1   g16557(.A1(new_n16804_), .A2(new_n16809_), .ZN(new_n16815_));
  AOI21_X1   g16558(.A1(new_n16814_), .A2(new_n16815_), .B(new_n16812_), .ZN(new_n16816_));
  NOR2_X1    g16559(.A1(new_n16811_), .A2(new_n16816_), .ZN(new_n16817_));
  XOR2_X1    g16560(.A1(new_n16817_), .A2(new_n16668_), .Z(new_n16818_));
  NOR2_X1    g16561(.A1(new_n16818_), .A2(new_n16667_), .ZN(new_n16819_));
  INV_X1     g16562(.I(new_n16668_), .ZN(new_n16820_));
  NOR2_X1    g16563(.A1(new_n16817_), .A2(new_n16820_), .ZN(new_n16821_));
  INV_X1     g16564(.I(new_n16821_), .ZN(new_n16822_));
  NAND2_X1   g16565(.A1(new_n16817_), .A2(new_n16820_), .ZN(new_n16823_));
  NAND2_X1   g16566(.A1(new_n16822_), .A2(new_n16823_), .ZN(new_n16824_));
  AOI21_X1   g16567(.A1(new_n16667_), .A2(new_n16824_), .B(new_n16819_), .ZN(new_n16825_));
  NOR2_X1    g16568(.A1(new_n16825_), .A2(new_n16662_), .ZN(new_n16826_));
  NAND2_X1   g16569(.A1(new_n16825_), .A2(new_n16662_), .ZN(new_n16827_));
  INV_X1     g16570(.I(new_n16827_), .ZN(new_n16828_));
  OAI21_X1   g16571(.A1(new_n16828_), .A2(new_n16826_), .B(new_n16661_), .ZN(new_n16829_));
  XNOR2_X1   g16572(.A1(new_n16825_), .A2(new_n16662_), .ZN(new_n16830_));
  OAI21_X1   g16573(.A1(new_n16661_), .A2(new_n16830_), .B(new_n16829_), .ZN(new_n16831_));
  NOR2_X1    g16574(.A1(new_n16626_), .A2(new_n16449_), .ZN(new_n16832_));
  NOR2_X1    g16575(.A1(new_n16832_), .A2(new_n16628_), .ZN(new_n16833_));
  XOR2_X1    g16576(.A1(new_n16831_), .A2(new_n16833_), .Z(new_n16834_));
  NOR2_X1    g16577(.A1(new_n16834_), .A2(new_n16655_), .ZN(new_n16835_));
  INV_X1     g16578(.I(new_n16655_), .ZN(new_n16836_));
  INV_X1     g16579(.I(new_n16831_), .ZN(new_n16837_));
  NOR2_X1    g16580(.A1(new_n16837_), .A2(new_n16833_), .ZN(new_n16838_));
  INV_X1     g16581(.I(new_n16838_), .ZN(new_n16839_));
  NAND2_X1   g16582(.A1(new_n16837_), .A2(new_n16833_), .ZN(new_n16840_));
  AOI21_X1   g16583(.A1(new_n16839_), .A2(new_n16840_), .B(new_n16836_), .ZN(new_n16841_));
  NOR2_X1    g16584(.A1(new_n16841_), .A2(new_n16835_), .ZN(new_n16842_));
  INV_X1     g16585(.I(new_n16842_), .ZN(new_n16843_));
  NOR2_X1    g16586(.A1(new_n16644_), .A2(new_n16642_), .ZN(new_n16844_));
  AOI21_X1   g16587(.A1(new_n16649_), .A2(new_n16844_), .B(new_n16843_), .ZN(new_n16845_));
  AOI21_X1   g16588(.A1(new_n16233_), .A2(new_n16434_), .B(new_n16433_), .ZN(new_n16846_));
  INV_X1     g16589(.I(new_n16844_), .ZN(new_n16847_));
  NOR3_X1    g16590(.A1(new_n16846_), .A2(new_n16842_), .A3(new_n16847_), .ZN(new_n16848_));
  OAI21_X1   g16591(.A1(new_n16848_), .A2(new_n16845_), .B(new_n16651_), .ZN(new_n16849_));
  INV_X1     g16592(.I(new_n16651_), .ZN(new_n16850_));
  OAI21_X1   g16593(.A1(new_n16846_), .A2(new_n16847_), .B(new_n16842_), .ZN(new_n16851_));
  NAND3_X1   g16594(.A1(new_n16649_), .A2(new_n16843_), .A3(new_n16844_), .ZN(new_n16852_));
  NAND3_X1   g16595(.A1(new_n16851_), .A2(new_n16852_), .A3(new_n16850_), .ZN(new_n16853_));
  NAND2_X1   g16596(.A1(new_n16849_), .A2(new_n16853_), .ZN(\f[88] ));
  NAND2_X1   g16597(.A1(new_n16649_), .A2(new_n16844_), .ZN(new_n16855_));
  AOI22_X1   g16598(.A1(new_n16851_), .A2(new_n16852_), .B1(new_n16855_), .B2(new_n16850_), .ZN(new_n16856_));
  AOI21_X1   g16599(.A1(new_n16836_), .A2(new_n16840_), .B(new_n16838_), .ZN(new_n16857_));
  INV_X1     g16600(.I(new_n16857_), .ZN(new_n16858_));
  NOR2_X1    g16601(.A1(new_n16826_), .A2(new_n16660_), .ZN(new_n16859_));
  NOR2_X1    g16602(.A1(new_n16859_), .A2(new_n16828_), .ZN(new_n16860_));
  OAI22_X1   g16603(.A1(new_n9595_), .A2(new_n1763_), .B1(new_n8956_), .B2(new_n1857_), .ZN(new_n16861_));
  OAI22_X1   g16604(.A1(new_n2084_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n2079_), .ZN(new_n16862_));
  NAND2_X1   g16605(.A1(new_n2864_), .A2(\b[60] ), .ZN(new_n16863_));
  AOI21_X1   g16606(.A1(new_n16862_), .A2(new_n16863_), .B(new_n2087_), .ZN(new_n16864_));
  NAND2_X1   g16607(.A1(new_n8935_), .A2(new_n16864_), .ZN(new_n16865_));
  XOR2_X1    g16608(.A1(new_n16865_), .A2(\a[29] ), .Z(new_n16866_));
  OAI21_X1   g16609(.A1(new_n16667_), .A2(new_n16821_), .B(new_n16823_), .ZN(new_n16867_));
  OAI22_X1   g16610(.A1(new_n2452_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n2447_), .ZN(new_n16868_));
  NAND2_X1   g16611(.A1(new_n3312_), .A2(\b[57] ), .ZN(new_n16869_));
  AOI21_X1   g16612(.A1(new_n16868_), .A2(new_n16869_), .B(new_n2455_), .ZN(new_n16870_));
  NAND2_X1   g16613(.A1(new_n7895_), .A2(new_n16870_), .ZN(new_n16871_));
  XOR2_X1    g16614(.A1(new_n16871_), .A2(\a[32] ), .Z(new_n16872_));
  OAI22_X1   g16615(.A1(new_n2846_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n2841_), .ZN(new_n16873_));
  NAND2_X1   g16616(.A1(new_n3755_), .A2(\b[54] ), .ZN(new_n16874_));
  AOI21_X1   g16617(.A1(new_n16873_), .A2(new_n16874_), .B(new_n2849_), .ZN(new_n16875_));
  NAND2_X1   g16618(.A1(new_n6994_), .A2(new_n16875_), .ZN(new_n16876_));
  XOR2_X1    g16619(.A1(new_n16876_), .A2(\a[35] ), .Z(new_n16877_));
  AOI21_X1   g16620(.A1(new_n16801_), .A2(new_n16799_), .B(new_n16797_), .ZN(new_n16878_));
  INV_X1     g16621(.I(new_n16878_), .ZN(new_n16879_));
  OAI22_X1   g16622(.A1(new_n3298_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n3293_), .ZN(new_n16880_));
  NAND2_X1   g16623(.A1(new_n4227_), .A2(\b[51] ), .ZN(new_n16881_));
  AOI21_X1   g16624(.A1(new_n16880_), .A2(new_n16881_), .B(new_n3301_), .ZN(new_n16882_));
  NAND2_X1   g16625(.A1(new_n6219_), .A2(new_n16882_), .ZN(new_n16883_));
  XOR2_X1    g16626(.A1(new_n16883_), .A2(\a[38] ), .Z(new_n16884_));
  OAI22_X1   g16627(.A1(new_n3736_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n3731_), .ZN(new_n16885_));
  NAND2_X1   g16628(.A1(new_n4730_), .A2(\b[48] ), .ZN(new_n16886_));
  AOI21_X1   g16629(.A1(new_n16885_), .A2(new_n16886_), .B(new_n3739_), .ZN(new_n16887_));
  NAND2_X1   g16630(.A1(new_n5537_), .A2(new_n16887_), .ZN(new_n16888_));
  XOR2_X1    g16631(.A1(new_n16888_), .A2(\a[41] ), .Z(new_n16889_));
  OAI22_X1   g16632(.A1(new_n4711_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n4706_), .ZN(new_n16890_));
  NAND2_X1   g16633(.A1(new_n5814_), .A2(\b[42] ), .ZN(new_n16891_));
  AOI21_X1   g16634(.A1(new_n16890_), .A2(new_n16891_), .B(new_n4714_), .ZN(new_n16892_));
  NAND2_X1   g16635(.A1(new_n4500_), .A2(new_n16892_), .ZN(new_n16893_));
  XOR2_X1    g16636(.A1(new_n16893_), .A2(\a[47] ), .Z(new_n16894_));
  NOR2_X1    g16637(.A1(new_n16755_), .A2(new_n16686_), .ZN(new_n16895_));
  NOR2_X1    g16638(.A1(new_n16895_), .A2(new_n16756_), .ZN(new_n16896_));
  OAI22_X1   g16639(.A1(new_n5786_), .A2(new_n3566_), .B1(new_n3408_), .B2(new_n5792_), .ZN(new_n16897_));
  NAND2_X1   g16640(.A1(new_n6745_), .A2(\b[36] ), .ZN(new_n16898_));
  AOI21_X1   g16641(.A1(new_n16898_), .A2(new_n16897_), .B(new_n5796_), .ZN(new_n16899_));
  NAND2_X1   g16642(.A1(new_n3565_), .A2(new_n16899_), .ZN(new_n16900_));
  XOR2_X1    g16643(.A1(new_n16900_), .A2(\a[53] ), .Z(new_n16901_));
  INV_X1     g16644(.I(new_n16732_), .ZN(new_n16902_));
  OAI21_X1   g16645(.A1(new_n16693_), .A2(new_n16734_), .B(new_n16902_), .ZN(new_n16903_));
  OAI22_X1   g16646(.A1(new_n6721_), .A2(new_n2964_), .B1(new_n6723_), .B2(new_n3097_), .ZN(new_n16904_));
  NAND2_X1   g16647(.A1(new_n7617_), .A2(\b[33] ), .ZN(new_n16905_));
  AOI21_X1   g16648(.A1(new_n16905_), .A2(new_n16904_), .B(new_n6731_), .ZN(new_n16906_));
  NAND2_X1   g16649(.A1(new_n3101_), .A2(new_n16906_), .ZN(new_n16907_));
  XOR2_X1    g16650(.A1(new_n16907_), .A2(\a[56] ), .Z(new_n16908_));
  OAI22_X1   g16651(.A1(new_n2660_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2543_), .ZN(new_n16909_));
  NAND2_X1   g16652(.A1(new_n8628_), .A2(\b[30] ), .ZN(new_n16910_));
  AOI21_X1   g16653(.A1(new_n16910_), .A2(new_n16909_), .B(new_n7354_), .ZN(new_n16911_));
  NAND2_X1   g16654(.A1(new_n2659_), .A2(new_n16911_), .ZN(new_n16912_));
  XOR2_X1    g16655(.A1(new_n16912_), .A2(\a[59] ), .Z(new_n16913_));
  INV_X1     g16656(.I(new_n16713_), .ZN(new_n16914_));
  AOI21_X1   g16657(.A1(new_n16701_), .A2(new_n16712_), .B(new_n16914_), .ZN(new_n16915_));
  OAI22_X1   g16658(.A1(new_n2272_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2175_), .ZN(new_n16916_));
  NAND2_X1   g16659(.A1(new_n9644_), .A2(\b[27] ), .ZN(new_n16917_));
  AOI21_X1   g16660(.A1(new_n16917_), .A2(new_n16916_), .B(new_n8321_), .ZN(new_n16918_));
  NAND2_X1   g16661(.A1(new_n2276_), .A2(new_n16918_), .ZN(new_n16919_));
  XOR2_X1    g16662(.A1(new_n16919_), .A2(\a[62] ), .Z(new_n16920_));
  NOR3_X1    g16663(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n1825_), .ZN(new_n16921_));
  NOR2_X1    g16664(.A1(new_n9364_), .A2(new_n1825_), .ZN(new_n16922_));
  NOR3_X1    g16665(.A1(new_n16922_), .A2(new_n1927_), .A3(new_n8985_), .ZN(new_n16923_));
  NOR2_X1    g16666(.A1(new_n16923_), .A2(new_n16921_), .ZN(new_n16924_));
  XOR2_X1    g16667(.A1(new_n16707_), .A2(new_n16924_), .Z(new_n16925_));
  NOR2_X1    g16668(.A1(new_n16920_), .A2(new_n16925_), .ZN(new_n16926_));
  INV_X1     g16669(.I(new_n16920_), .ZN(new_n16927_));
  NOR2_X1    g16670(.A1(new_n16708_), .A2(new_n16924_), .ZN(new_n16928_));
  INV_X1     g16671(.I(new_n16924_), .ZN(new_n16929_));
  NOR2_X1    g16672(.A1(new_n16929_), .A2(new_n16707_), .ZN(new_n16930_));
  NOR2_X1    g16673(.A1(new_n16928_), .A2(new_n16930_), .ZN(new_n16931_));
  NOR2_X1    g16674(.A1(new_n16927_), .A2(new_n16931_), .ZN(new_n16932_));
  NOR2_X1    g16675(.A1(new_n16932_), .A2(new_n16926_), .ZN(new_n16933_));
  XOR2_X1    g16676(.A1(new_n16933_), .A2(new_n16915_), .Z(new_n16934_));
  NOR2_X1    g16677(.A1(new_n16934_), .A2(new_n16913_), .ZN(new_n16935_));
  INV_X1     g16678(.I(new_n16913_), .ZN(new_n16936_));
  INV_X1     g16679(.I(new_n16915_), .ZN(new_n16937_));
  NOR2_X1    g16680(.A1(new_n16933_), .A2(new_n16937_), .ZN(new_n16938_));
  INV_X1     g16681(.I(new_n16938_), .ZN(new_n16939_));
  NAND2_X1   g16682(.A1(new_n16933_), .A2(new_n16937_), .ZN(new_n16940_));
  AOI21_X1   g16683(.A1(new_n16939_), .A2(new_n16940_), .B(new_n16936_), .ZN(new_n16941_));
  NOR2_X1    g16684(.A1(new_n16935_), .A2(new_n16941_), .ZN(new_n16942_));
  NOR2_X1    g16685(.A1(new_n16723_), .A2(new_n16696_), .ZN(new_n16943_));
  NOR2_X1    g16686(.A1(new_n16943_), .A2(new_n16722_), .ZN(new_n16944_));
  XOR2_X1    g16687(.A1(new_n16942_), .A2(new_n16944_), .Z(new_n16945_));
  NOR2_X1    g16688(.A1(new_n16945_), .A2(new_n16908_), .ZN(new_n16946_));
  INV_X1     g16689(.I(new_n16908_), .ZN(new_n16947_));
  INV_X1     g16690(.I(new_n16942_), .ZN(new_n16948_));
  NOR2_X1    g16691(.A1(new_n16948_), .A2(new_n16944_), .ZN(new_n16949_));
  INV_X1     g16692(.I(new_n16949_), .ZN(new_n16950_));
  NAND2_X1   g16693(.A1(new_n16948_), .A2(new_n16944_), .ZN(new_n16951_));
  AOI21_X1   g16694(.A1(new_n16950_), .A2(new_n16951_), .B(new_n16947_), .ZN(new_n16952_));
  NOR2_X1    g16695(.A1(new_n16952_), .A2(new_n16946_), .ZN(new_n16953_));
  NOR2_X1    g16696(.A1(new_n16953_), .A2(new_n16903_), .ZN(new_n16954_));
  INV_X1     g16697(.I(new_n16954_), .ZN(new_n16955_));
  NAND2_X1   g16698(.A1(new_n16953_), .A2(new_n16903_), .ZN(new_n16956_));
  AOI21_X1   g16699(.A1(new_n16955_), .A2(new_n16956_), .B(new_n16901_), .ZN(new_n16957_));
  INV_X1     g16700(.I(new_n16901_), .ZN(new_n16958_));
  XNOR2_X1   g16701(.A1(new_n16953_), .A2(new_n16903_), .ZN(new_n16959_));
  NOR2_X1    g16702(.A1(new_n16959_), .A2(new_n16958_), .ZN(new_n16960_));
  OAI22_X1   g16703(.A1(new_n5228_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n5225_), .ZN(new_n16961_));
  NAND2_X1   g16704(.A1(new_n5387_), .A2(\b[39] ), .ZN(new_n16962_));
  AOI21_X1   g16705(.A1(new_n16961_), .A2(new_n16962_), .B(new_n5231_), .ZN(new_n16963_));
  NAND2_X1   g16706(.A1(new_n3996_), .A2(new_n16963_), .ZN(new_n16964_));
  XOR2_X1    g16707(.A1(new_n16964_), .A2(\a[50] ), .Z(new_n16965_));
  NOR2_X1    g16708(.A1(new_n16751_), .A2(new_n16749_), .ZN(new_n16966_));
  NOR2_X1    g16709(.A1(new_n16966_), .A2(new_n16750_), .ZN(new_n16967_));
  NOR2_X1    g16710(.A1(new_n16967_), .A2(new_n16965_), .ZN(new_n16968_));
  AND2_X2    g16711(.A1(new_n16967_), .A2(new_n16965_), .Z(new_n16969_));
  OAI22_X1   g16712(.A1(new_n16969_), .A2(new_n16968_), .B1(new_n16957_), .B2(new_n16960_), .ZN(new_n16970_));
  NOR2_X1    g16713(.A1(new_n16960_), .A2(new_n16957_), .ZN(new_n16971_));
  XOR2_X1    g16714(.A1(new_n16967_), .A2(new_n16965_), .Z(new_n16972_));
  NAND2_X1   g16715(.A1(new_n16972_), .A2(new_n16971_), .ZN(new_n16973_));
  NAND2_X1   g16716(.A1(new_n16973_), .A2(new_n16970_), .ZN(new_n16974_));
  XOR2_X1    g16717(.A1(new_n16896_), .A2(new_n16974_), .Z(new_n16975_));
  INV_X1     g16718(.I(new_n16974_), .ZN(new_n16976_));
  NOR2_X1    g16719(.A1(new_n16896_), .A2(new_n16976_), .ZN(new_n16977_));
  NAND2_X1   g16720(.A1(new_n16896_), .A2(new_n16976_), .ZN(new_n16978_));
  INV_X1     g16721(.I(new_n16978_), .ZN(new_n16979_));
  OAI21_X1   g16722(.A1(new_n16979_), .A2(new_n16977_), .B(new_n16894_), .ZN(new_n16980_));
  OAI21_X1   g16723(.A1(new_n16894_), .A2(new_n16975_), .B(new_n16980_), .ZN(new_n16981_));
  OAI22_X1   g16724(.A1(new_n4208_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n4203_), .ZN(new_n16982_));
  NAND2_X1   g16725(.A1(new_n5244_), .A2(\b[45] ), .ZN(new_n16983_));
  AOI21_X1   g16726(.A1(new_n16982_), .A2(new_n16983_), .B(new_n4211_), .ZN(new_n16984_));
  NAND2_X1   g16727(.A1(new_n5004_), .A2(new_n16984_), .ZN(new_n16985_));
  XOR2_X1    g16728(.A1(new_n16985_), .A2(\a[44] ), .Z(new_n16986_));
  INV_X1     g16729(.I(new_n16986_), .ZN(new_n16987_));
  NAND2_X1   g16730(.A1(new_n16768_), .A2(new_n16766_), .ZN(new_n16988_));
  NAND2_X1   g16731(.A1(new_n16988_), .A2(new_n16765_), .ZN(new_n16989_));
  XOR2_X1    g16732(.A1(new_n16989_), .A2(new_n16987_), .Z(new_n16990_));
  NAND2_X1   g16733(.A1(new_n16990_), .A2(new_n16981_), .ZN(new_n16991_));
  AOI21_X1   g16734(.A1(new_n16988_), .A2(new_n16765_), .B(new_n16986_), .ZN(new_n16992_));
  NOR2_X1    g16735(.A1(new_n16989_), .A2(new_n16987_), .ZN(new_n16993_));
  NOR2_X1    g16736(.A1(new_n16993_), .A2(new_n16992_), .ZN(new_n16994_));
  OAI21_X1   g16737(.A1(new_n16981_), .A2(new_n16994_), .B(new_n16991_), .ZN(new_n16995_));
  NAND2_X1   g16738(.A1(new_n16775_), .A2(new_n16777_), .ZN(new_n16996_));
  NAND2_X1   g16739(.A1(new_n16996_), .A2(new_n16774_), .ZN(new_n16997_));
  XNOR2_X1   g16740(.A1(new_n16995_), .A2(new_n16997_), .ZN(new_n16998_));
  NOR2_X1    g16741(.A1(new_n16998_), .A2(new_n16889_), .ZN(new_n16999_));
  INV_X1     g16742(.I(new_n16889_), .ZN(new_n17000_));
  INV_X1     g16743(.I(new_n16995_), .ZN(new_n17001_));
  INV_X1     g16744(.I(new_n16997_), .ZN(new_n17002_));
  NOR2_X1    g16745(.A1(new_n17001_), .A2(new_n17002_), .ZN(new_n17003_));
  NOR2_X1    g16746(.A1(new_n16995_), .A2(new_n16997_), .ZN(new_n17004_));
  NOR2_X1    g16747(.A1(new_n17003_), .A2(new_n17004_), .ZN(new_n17005_));
  NOR2_X1    g16748(.A1(new_n17005_), .A2(new_n17000_), .ZN(new_n17006_));
  NOR2_X1    g16749(.A1(new_n17006_), .A2(new_n16999_), .ZN(new_n17007_));
  INV_X1     g16750(.I(new_n16780_), .ZN(new_n17008_));
  AOI21_X1   g16751(.A1(new_n17008_), .A2(new_n16791_), .B(new_n16789_), .ZN(new_n17009_));
  XOR2_X1    g16752(.A1(new_n17007_), .A2(new_n17009_), .Z(new_n17010_));
  NOR2_X1    g16753(.A1(new_n17010_), .A2(new_n16884_), .ZN(new_n17011_));
  INV_X1     g16754(.I(new_n16884_), .ZN(new_n17012_));
  INV_X1     g16755(.I(new_n17007_), .ZN(new_n17013_));
  NOR2_X1    g16756(.A1(new_n17013_), .A2(new_n17009_), .ZN(new_n17014_));
  INV_X1     g16757(.I(new_n17014_), .ZN(new_n17015_));
  NAND2_X1   g16758(.A1(new_n17013_), .A2(new_n17009_), .ZN(new_n17016_));
  AOI21_X1   g16759(.A1(new_n17015_), .A2(new_n17016_), .B(new_n17012_), .ZN(new_n17017_));
  NOR2_X1    g16760(.A1(new_n17017_), .A2(new_n17011_), .ZN(new_n17018_));
  NOR2_X1    g16761(.A1(new_n17018_), .A2(new_n16879_), .ZN(new_n17019_));
  INV_X1     g16762(.I(new_n17018_), .ZN(new_n17020_));
  NOR2_X1    g16763(.A1(new_n17020_), .A2(new_n16878_), .ZN(new_n17021_));
  NOR2_X1    g16764(.A1(new_n17021_), .A2(new_n17019_), .ZN(new_n17022_));
  NOR2_X1    g16765(.A1(new_n17022_), .A2(new_n16877_), .ZN(new_n17023_));
  INV_X1     g16766(.I(new_n16877_), .ZN(new_n17024_));
  XOR2_X1    g16767(.A1(new_n17018_), .A2(new_n16878_), .Z(new_n17025_));
  NOR2_X1    g16768(.A1(new_n17025_), .A2(new_n17024_), .ZN(new_n17026_));
  NOR2_X1    g16769(.A1(new_n17023_), .A2(new_n17026_), .ZN(new_n17027_));
  AOI21_X1   g16770(.A1(new_n16812_), .A2(new_n16815_), .B(new_n16813_), .ZN(new_n17028_));
  NOR2_X1    g16771(.A1(new_n17027_), .A2(new_n17028_), .ZN(new_n17029_));
  INV_X1     g16772(.I(new_n17028_), .ZN(new_n17030_));
  NOR3_X1    g16773(.A1(new_n17030_), .A2(new_n17023_), .A3(new_n17026_), .ZN(new_n17031_));
  NOR2_X1    g16774(.A1(new_n17029_), .A2(new_n17031_), .ZN(new_n17032_));
  NOR2_X1    g16775(.A1(new_n17032_), .A2(new_n16872_), .ZN(new_n17033_));
  INV_X1     g16776(.I(new_n16872_), .ZN(new_n17034_));
  XOR2_X1    g16777(.A1(new_n17027_), .A2(new_n17030_), .Z(new_n17035_));
  NOR2_X1    g16778(.A1(new_n17035_), .A2(new_n17034_), .ZN(new_n17036_));
  NOR2_X1    g16779(.A1(new_n17036_), .A2(new_n17033_), .ZN(new_n17037_));
  XOR2_X1    g16780(.A1(new_n17037_), .A2(new_n16867_), .Z(new_n17038_));
  NOR2_X1    g16781(.A1(new_n17038_), .A2(new_n16866_), .ZN(new_n17039_));
  INV_X1     g16782(.I(new_n16866_), .ZN(new_n17040_));
  INV_X1     g16783(.I(new_n16867_), .ZN(new_n17041_));
  NOR2_X1    g16784(.A1(new_n17037_), .A2(new_n17041_), .ZN(new_n17042_));
  INV_X1     g16785(.I(new_n17042_), .ZN(new_n17043_));
  NAND2_X1   g16786(.A1(new_n17037_), .A2(new_n17041_), .ZN(new_n17044_));
  AOI21_X1   g16787(.A1(new_n17043_), .A2(new_n17044_), .B(new_n17040_), .ZN(new_n17045_));
  NOR2_X1    g16788(.A1(new_n17039_), .A2(new_n17045_), .ZN(new_n17046_));
  XOR2_X1    g16789(.A1(new_n17046_), .A2(new_n16861_), .Z(new_n17047_));
  XOR2_X1    g16790(.A1(new_n17047_), .A2(\a[26] ), .Z(new_n17048_));
  XNOR2_X1   g16791(.A1(new_n17048_), .A2(new_n16860_), .ZN(new_n17049_));
  XOR2_X1    g16792(.A1(new_n17049_), .A2(new_n16858_), .Z(new_n17050_));
  NAND2_X1   g16793(.A1(new_n16856_), .A2(new_n17050_), .ZN(new_n17051_));
  XOR2_X1    g16794(.A1(new_n17049_), .A2(new_n16858_), .Z(new_n17052_));
  OAI21_X1   g16795(.A1(new_n16856_), .A2(new_n17052_), .B(new_n17051_), .ZN(\f[89] ));
  XOR2_X1    g16796(.A1(new_n16861_), .A2(new_n1750_), .Z(new_n17054_));
  XNOR2_X1   g16797(.A1(new_n16860_), .A2(new_n17054_), .ZN(new_n17055_));
  INV_X1     g16798(.I(new_n17055_), .ZN(new_n17056_));
  OAI21_X1   g16799(.A1(new_n17046_), .A2(new_n17054_), .B(new_n17056_), .ZN(new_n17057_));
  AOI21_X1   g16800(.A1(new_n17040_), .A2(new_n17044_), .B(new_n17042_), .ZN(new_n17058_));
  OAI22_X1   g16801(.A1(new_n2084_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n2079_), .ZN(new_n17059_));
  NAND2_X1   g16802(.A1(new_n2864_), .A2(\b[61] ), .ZN(new_n17060_));
  AOI21_X1   g16803(.A1(new_n17059_), .A2(new_n17060_), .B(new_n2087_), .ZN(new_n17061_));
  NAND2_X1   g16804(.A1(new_n8963_), .A2(new_n17061_), .ZN(new_n17062_));
  XOR2_X1    g16805(.A1(new_n17062_), .A2(\a[29] ), .Z(new_n17063_));
  NOR2_X1    g16806(.A1(new_n17019_), .A2(new_n16877_), .ZN(new_n17064_));
  NOR2_X1    g16807(.A1(new_n17064_), .A2(new_n17021_), .ZN(new_n17065_));
  INV_X1     g16808(.I(new_n17065_), .ZN(new_n17066_));
  AOI21_X1   g16809(.A1(new_n17012_), .A2(new_n17016_), .B(new_n17014_), .ZN(new_n17067_));
  INV_X1     g16810(.I(new_n17004_), .ZN(new_n17068_));
  AOI21_X1   g16811(.A1(new_n17000_), .A2(new_n17068_), .B(new_n17003_), .ZN(new_n17069_));
  INV_X1     g16812(.I(new_n16894_), .ZN(new_n17070_));
  AOI21_X1   g16813(.A1(new_n17070_), .A2(new_n16978_), .B(new_n16977_), .ZN(new_n17071_));
  INV_X1     g16814(.I(new_n17071_), .ZN(new_n17072_));
  NOR2_X1    g16815(.A1(new_n16971_), .A2(new_n16969_), .ZN(new_n17073_));
  NOR2_X1    g16816(.A1(new_n17073_), .A2(new_n16968_), .ZN(new_n17074_));
  OAI21_X1   g16817(.A1(new_n16901_), .A2(new_n16954_), .B(new_n16956_), .ZN(new_n17075_));
  INV_X1     g16818(.I(new_n17075_), .ZN(new_n17076_));
  OAI21_X1   g16819(.A1(new_n16913_), .A2(new_n16938_), .B(new_n16940_), .ZN(new_n17077_));
  INV_X1     g16820(.I(new_n17077_), .ZN(new_n17078_));
  OAI22_X1   g16821(.A1(new_n2794_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2660_), .ZN(new_n17079_));
  NAND2_X1   g16822(.A1(new_n8628_), .A2(\b[31] ), .ZN(new_n17080_));
  AOI21_X1   g16823(.A1(new_n17080_), .A2(new_n17079_), .B(new_n7354_), .ZN(new_n17081_));
  NAND2_X1   g16824(.A1(new_n2797_), .A2(new_n17081_), .ZN(new_n17082_));
  XOR2_X1    g16825(.A1(new_n17082_), .A2(\a[59] ), .Z(new_n17083_));
  INV_X1     g16826(.I(new_n16928_), .ZN(new_n17084_));
  AOI21_X1   g16827(.A1(new_n16927_), .A2(new_n17084_), .B(new_n16930_), .ZN(new_n17085_));
  INV_X1     g16828(.I(new_n17085_), .ZN(new_n17086_));
  OAI22_X1   g16829(.A1(new_n2405_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2272_), .ZN(new_n17087_));
  NAND2_X1   g16830(.A1(new_n9644_), .A2(\b[28] ), .ZN(new_n17088_));
  AOI21_X1   g16831(.A1(new_n17088_), .A2(new_n17087_), .B(new_n8321_), .ZN(new_n17089_));
  NAND2_X1   g16832(.A1(new_n2404_), .A2(new_n17089_), .ZN(new_n17090_));
  XOR2_X1    g16833(.A1(new_n17090_), .A2(\a[62] ), .Z(new_n17091_));
  INV_X1     g16834(.I(new_n17091_), .ZN(new_n17092_));
  NOR2_X1    g16835(.A1(new_n8985_), .A2(new_n2039_), .ZN(new_n17093_));
  NOR2_X1    g16836(.A1(new_n9364_), .A2(new_n1927_), .ZN(new_n17094_));
  XNOR2_X1   g16837(.A1(new_n17093_), .A2(new_n17094_), .ZN(new_n17095_));
  XOR2_X1    g16838(.A1(new_n17095_), .A2(\a[26] ), .Z(new_n17096_));
  NOR2_X1    g16839(.A1(new_n17096_), .A2(new_n16924_), .ZN(new_n17097_));
  NOR2_X1    g16840(.A1(new_n17095_), .A2(new_n1750_), .ZN(new_n17098_));
  INV_X1     g16841(.I(new_n17098_), .ZN(new_n17099_));
  NAND2_X1   g16842(.A1(new_n17095_), .A2(new_n1750_), .ZN(new_n17100_));
  AOI21_X1   g16843(.A1(new_n17099_), .A2(new_n17100_), .B(new_n16929_), .ZN(new_n17101_));
  NOR2_X1    g16844(.A1(new_n17097_), .A2(new_n17101_), .ZN(new_n17102_));
  NOR2_X1    g16845(.A1(new_n17092_), .A2(new_n17102_), .ZN(new_n17103_));
  INV_X1     g16846(.I(new_n17103_), .ZN(new_n17104_));
  NAND2_X1   g16847(.A1(new_n17092_), .A2(new_n17102_), .ZN(new_n17105_));
  NAND2_X1   g16848(.A1(new_n17104_), .A2(new_n17105_), .ZN(new_n17106_));
  NAND2_X1   g16849(.A1(new_n17086_), .A2(new_n17106_), .ZN(new_n17107_));
  XNOR2_X1   g16850(.A1(new_n17091_), .A2(new_n17102_), .ZN(new_n17108_));
  NAND2_X1   g16851(.A1(new_n17085_), .A2(new_n17108_), .ZN(new_n17109_));
  NAND2_X1   g16852(.A1(new_n17107_), .A2(new_n17109_), .ZN(new_n17110_));
  XOR2_X1    g16853(.A1(new_n17110_), .A2(new_n17083_), .Z(new_n17111_));
  NOR2_X1    g16854(.A1(new_n17111_), .A2(new_n17078_), .ZN(new_n17112_));
  AOI21_X1   g16855(.A1(new_n17107_), .A2(new_n17109_), .B(new_n17083_), .ZN(new_n17113_));
  INV_X1     g16856(.I(new_n17113_), .ZN(new_n17114_));
  INV_X1     g16857(.I(new_n17083_), .ZN(new_n17115_));
  NOR2_X1    g16858(.A1(new_n17110_), .A2(new_n17115_), .ZN(new_n17116_));
  INV_X1     g16859(.I(new_n17116_), .ZN(new_n17117_));
  AOI21_X1   g16860(.A1(new_n17117_), .A2(new_n17114_), .B(new_n17077_), .ZN(new_n17118_));
  NOR2_X1    g16861(.A1(new_n17112_), .A2(new_n17118_), .ZN(new_n17119_));
  OAI22_X1   g16862(.A1(new_n6721_), .A2(new_n3097_), .B1(new_n6723_), .B2(new_n3247_), .ZN(new_n17120_));
  NAND2_X1   g16863(.A1(new_n7617_), .A2(\b[34] ), .ZN(new_n17121_));
  AOI21_X1   g16864(.A1(new_n17121_), .A2(new_n17120_), .B(new_n6731_), .ZN(new_n17122_));
  NAND2_X1   g16865(.A1(new_n3246_), .A2(new_n17122_), .ZN(new_n17123_));
  XOR2_X1    g16866(.A1(new_n17123_), .A2(\a[56] ), .Z(new_n17124_));
  NAND2_X1   g16867(.A1(new_n16951_), .A2(new_n16947_), .ZN(new_n17125_));
  NAND2_X1   g16868(.A1(new_n17125_), .A2(new_n16950_), .ZN(new_n17126_));
  INV_X1     g16869(.I(new_n17126_), .ZN(new_n17127_));
  NOR2_X1    g16870(.A1(new_n17127_), .A2(new_n17124_), .ZN(new_n17128_));
  INV_X1     g16871(.I(new_n17124_), .ZN(new_n17129_));
  NOR2_X1    g16872(.A1(new_n17126_), .A2(new_n17129_), .ZN(new_n17130_));
  NOR2_X1    g16873(.A1(new_n17128_), .A2(new_n17130_), .ZN(new_n17131_));
  NOR2_X1    g16874(.A1(new_n17131_), .A2(new_n17119_), .ZN(new_n17132_));
  XOR2_X1    g16875(.A1(new_n17126_), .A2(new_n17124_), .Z(new_n17133_));
  NOR3_X1    g16876(.A1(new_n17133_), .A2(new_n17112_), .A3(new_n17118_), .ZN(new_n17134_));
  NOR2_X1    g16877(.A1(new_n17132_), .A2(new_n17134_), .ZN(new_n17135_));
  OAI22_X1   g16878(.A1(new_n5786_), .A2(new_n3696_), .B1(new_n3566_), .B2(new_n5792_), .ZN(new_n17136_));
  NAND2_X1   g16879(.A1(new_n6745_), .A2(\b[37] ), .ZN(new_n17137_));
  AOI21_X1   g16880(.A1(new_n17137_), .A2(new_n17136_), .B(new_n5796_), .ZN(new_n17138_));
  NAND2_X1   g16881(.A1(new_n3700_), .A2(new_n17138_), .ZN(new_n17139_));
  XOR2_X1    g16882(.A1(new_n17139_), .A2(\a[53] ), .Z(new_n17140_));
  XOR2_X1    g16883(.A1(new_n17135_), .A2(new_n17140_), .Z(new_n17141_));
  NOR3_X1    g16884(.A1(new_n17132_), .A2(new_n17134_), .A3(new_n17140_), .ZN(new_n17142_));
  INV_X1     g16885(.I(new_n17140_), .ZN(new_n17143_));
  NOR2_X1    g16886(.A1(new_n17135_), .A2(new_n17143_), .ZN(new_n17144_));
  OAI21_X1   g16887(.A1(new_n17144_), .A2(new_n17142_), .B(new_n17076_), .ZN(new_n17145_));
  OAI21_X1   g16888(.A1(new_n17076_), .A2(new_n17141_), .B(new_n17145_), .ZN(new_n17146_));
  OAI22_X1   g16889(.A1(new_n5228_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n5225_), .ZN(new_n17147_));
  NAND2_X1   g16890(.A1(new_n5387_), .A2(\b[40] ), .ZN(new_n17148_));
  AOI21_X1   g16891(.A1(new_n17147_), .A2(new_n17148_), .B(new_n5231_), .ZN(new_n17149_));
  NAND2_X1   g16892(.A1(new_n4017_), .A2(new_n17149_), .ZN(new_n17150_));
  XOR2_X1    g16893(.A1(new_n17150_), .A2(\a[50] ), .Z(new_n17151_));
  NOR2_X1    g16894(.A1(new_n17146_), .A2(new_n17151_), .ZN(new_n17152_));
  INV_X1     g16895(.I(new_n17152_), .ZN(new_n17153_));
  NAND2_X1   g16896(.A1(new_n17146_), .A2(new_n17151_), .ZN(new_n17154_));
  AOI21_X1   g16897(.A1(new_n17153_), .A2(new_n17154_), .B(new_n17074_), .ZN(new_n17155_));
  INV_X1     g16898(.I(new_n17074_), .ZN(new_n17156_));
  XNOR2_X1   g16899(.A1(new_n17146_), .A2(new_n17151_), .ZN(new_n17157_));
  NOR2_X1    g16900(.A1(new_n17157_), .A2(new_n17156_), .ZN(new_n17158_));
  NOR2_X1    g16901(.A1(new_n17158_), .A2(new_n17155_), .ZN(new_n17159_));
  OAI22_X1   g16902(.A1(new_n4711_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n4706_), .ZN(new_n17160_));
  NAND2_X1   g16903(.A1(new_n5814_), .A2(\b[43] ), .ZN(new_n17161_));
  AOI21_X1   g16904(.A1(new_n17160_), .A2(new_n17161_), .B(new_n4714_), .ZN(new_n17162_));
  NAND2_X1   g16905(.A1(new_n4513_), .A2(new_n17162_), .ZN(new_n17163_));
  XOR2_X1    g16906(.A1(new_n17163_), .A2(\a[47] ), .Z(new_n17164_));
  XNOR2_X1   g16907(.A1(new_n17159_), .A2(new_n17164_), .ZN(new_n17165_));
  INV_X1     g16908(.I(new_n17165_), .ZN(new_n17166_));
  NOR2_X1    g16909(.A1(new_n17159_), .A2(new_n17164_), .ZN(new_n17167_));
  NAND2_X1   g16910(.A1(new_n17159_), .A2(new_n17164_), .ZN(new_n17168_));
  INV_X1     g16911(.I(new_n17168_), .ZN(new_n17169_));
  NOR2_X1    g16912(.A1(new_n17169_), .A2(new_n17167_), .ZN(new_n17170_));
  NOR2_X1    g16913(.A1(new_n17170_), .A2(new_n17072_), .ZN(new_n17171_));
  AOI21_X1   g16914(.A1(new_n17072_), .A2(new_n17166_), .B(new_n17171_), .ZN(new_n17172_));
  OAI22_X1   g16915(.A1(new_n4208_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n4203_), .ZN(new_n17173_));
  NAND2_X1   g16916(.A1(new_n5244_), .A2(\b[46] ), .ZN(new_n17174_));
  AOI21_X1   g16917(.A1(new_n17173_), .A2(new_n17174_), .B(new_n4211_), .ZN(new_n17175_));
  NAND2_X1   g16918(.A1(new_n5177_), .A2(new_n17175_), .ZN(new_n17176_));
  XOR2_X1    g16919(.A1(new_n17176_), .A2(\a[44] ), .Z(new_n17177_));
  NOR2_X1    g16920(.A1(new_n16993_), .A2(new_n16981_), .ZN(new_n17178_));
  NOR2_X1    g16921(.A1(new_n17178_), .A2(new_n16992_), .ZN(new_n17179_));
  NOR2_X1    g16922(.A1(new_n17179_), .A2(new_n17177_), .ZN(new_n17180_));
  INV_X1     g16923(.I(new_n17180_), .ZN(new_n17181_));
  NAND2_X1   g16924(.A1(new_n17179_), .A2(new_n17177_), .ZN(new_n17182_));
  AOI21_X1   g16925(.A1(new_n17181_), .A2(new_n17182_), .B(new_n17172_), .ZN(new_n17183_));
  INV_X1     g16926(.I(new_n17172_), .ZN(new_n17184_));
  XNOR2_X1   g16927(.A1(new_n17179_), .A2(new_n17177_), .ZN(new_n17185_));
  NOR2_X1    g16928(.A1(new_n17184_), .A2(new_n17185_), .ZN(new_n17186_));
  NOR2_X1    g16929(.A1(new_n17186_), .A2(new_n17183_), .ZN(new_n17187_));
  INV_X1     g16930(.I(new_n17187_), .ZN(new_n17188_));
  OAI22_X1   g16931(.A1(new_n3736_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n3731_), .ZN(new_n17189_));
  NAND2_X1   g16932(.A1(new_n4730_), .A2(\b[49] ), .ZN(new_n17190_));
  AOI21_X1   g16933(.A1(new_n17189_), .A2(new_n17190_), .B(new_n3739_), .ZN(new_n17191_));
  NAND2_X1   g16934(.A1(new_n5741_), .A2(new_n17191_), .ZN(new_n17192_));
  XOR2_X1    g16935(.A1(new_n17192_), .A2(\a[41] ), .Z(new_n17193_));
  NOR2_X1    g16936(.A1(new_n17188_), .A2(new_n17193_), .ZN(new_n17194_));
  INV_X1     g16937(.I(new_n17193_), .ZN(new_n17195_));
  NOR2_X1    g16938(.A1(new_n17187_), .A2(new_n17195_), .ZN(new_n17196_));
  NOR2_X1    g16939(.A1(new_n17194_), .A2(new_n17196_), .ZN(new_n17197_));
  NOR2_X1    g16940(.A1(new_n17197_), .A2(new_n17069_), .ZN(new_n17198_));
  INV_X1     g16941(.I(new_n17069_), .ZN(new_n17199_));
  XOR2_X1    g16942(.A1(new_n17187_), .A2(new_n17193_), .Z(new_n17200_));
  NOR2_X1    g16943(.A1(new_n17200_), .A2(new_n17199_), .ZN(new_n17201_));
  NOR2_X1    g16944(.A1(new_n17198_), .A2(new_n17201_), .ZN(new_n17202_));
  OAI22_X1   g16945(.A1(new_n3298_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n3293_), .ZN(new_n17203_));
  NAND2_X1   g16946(.A1(new_n4227_), .A2(\b[52] ), .ZN(new_n17204_));
  AOI21_X1   g16947(.A1(new_n17203_), .A2(new_n17204_), .B(new_n3301_), .ZN(new_n17205_));
  NAND2_X1   g16948(.A1(new_n6237_), .A2(new_n17205_), .ZN(new_n17206_));
  XOR2_X1    g16949(.A1(new_n17206_), .A2(\a[38] ), .Z(new_n17207_));
  XNOR2_X1   g16950(.A1(new_n17202_), .A2(new_n17207_), .ZN(new_n17208_));
  NOR2_X1    g16951(.A1(new_n17208_), .A2(new_n17067_), .ZN(new_n17209_));
  INV_X1     g16952(.I(new_n17067_), .ZN(new_n17210_));
  NOR2_X1    g16953(.A1(new_n17202_), .A2(new_n17207_), .ZN(new_n17211_));
  INV_X1     g16954(.I(new_n17211_), .ZN(new_n17212_));
  NAND2_X1   g16955(.A1(new_n17202_), .A2(new_n17207_), .ZN(new_n17213_));
  AOI21_X1   g16956(.A1(new_n17212_), .A2(new_n17213_), .B(new_n17210_), .ZN(new_n17214_));
  NOR2_X1    g16957(.A1(new_n17209_), .A2(new_n17214_), .ZN(new_n17215_));
  OAI22_X1   g16958(.A1(new_n2846_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n2841_), .ZN(new_n17216_));
  NAND2_X1   g16959(.A1(new_n3755_), .A2(\b[55] ), .ZN(new_n17217_));
  AOI21_X1   g16960(.A1(new_n17216_), .A2(new_n17217_), .B(new_n2849_), .ZN(new_n17218_));
  NAND2_X1   g16961(.A1(new_n7308_), .A2(new_n17218_), .ZN(new_n17219_));
  XOR2_X1    g16962(.A1(new_n17219_), .A2(\a[35] ), .Z(new_n17220_));
  XOR2_X1    g16963(.A1(new_n17215_), .A2(new_n17220_), .Z(new_n17221_));
  INV_X1     g16964(.I(new_n17221_), .ZN(new_n17222_));
  INV_X1     g16965(.I(new_n17215_), .ZN(new_n17223_));
  NOR2_X1    g16966(.A1(new_n17223_), .A2(new_n17220_), .ZN(new_n17224_));
  INV_X1     g16967(.I(new_n17224_), .ZN(new_n17225_));
  NAND2_X1   g16968(.A1(new_n17223_), .A2(new_n17220_), .ZN(new_n17226_));
  AOI21_X1   g16969(.A1(new_n17225_), .A2(new_n17226_), .B(new_n17066_), .ZN(new_n17227_));
  AOI21_X1   g16970(.A1(new_n17066_), .A2(new_n17222_), .B(new_n17227_), .ZN(new_n17228_));
  OAI22_X1   g16971(.A1(new_n2452_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n2447_), .ZN(new_n17229_));
  NAND2_X1   g16972(.A1(new_n3312_), .A2(\b[58] ), .ZN(new_n17230_));
  AOI21_X1   g16973(.A1(new_n17229_), .A2(new_n17230_), .B(new_n2455_), .ZN(new_n17231_));
  NAND2_X1   g16974(.A1(new_n7929_), .A2(new_n17231_), .ZN(new_n17232_));
  XOR2_X1    g16975(.A1(new_n17232_), .A2(\a[32] ), .Z(new_n17233_));
  NOR2_X1    g16976(.A1(new_n17031_), .A2(new_n16872_), .ZN(new_n17234_));
  NOR2_X1    g16977(.A1(new_n17234_), .A2(new_n17029_), .ZN(new_n17235_));
  XNOR2_X1   g16978(.A1(new_n17235_), .A2(new_n17233_), .ZN(new_n17236_));
  NOR2_X1    g16979(.A1(new_n17236_), .A2(new_n17228_), .ZN(new_n17237_));
  NOR2_X1    g16980(.A1(new_n17235_), .A2(new_n17233_), .ZN(new_n17238_));
  INV_X1     g16981(.I(new_n17238_), .ZN(new_n17239_));
  NAND2_X1   g16982(.A1(new_n17235_), .A2(new_n17233_), .ZN(new_n17240_));
  NAND2_X1   g16983(.A1(new_n17239_), .A2(new_n17240_), .ZN(new_n17241_));
  AOI21_X1   g16984(.A1(new_n17228_), .A2(new_n17241_), .B(new_n17237_), .ZN(new_n17242_));
  XNOR2_X1   g16985(.A1(new_n17242_), .A2(new_n17063_), .ZN(new_n17243_));
  NOR2_X1    g16986(.A1(new_n17243_), .A2(new_n17058_), .ZN(new_n17244_));
  INV_X1     g16987(.I(new_n17058_), .ZN(new_n17245_));
  NOR2_X1    g16988(.A1(new_n17242_), .A2(new_n17063_), .ZN(new_n17246_));
  INV_X1     g16989(.I(new_n17246_), .ZN(new_n17247_));
  NAND2_X1   g16990(.A1(new_n17242_), .A2(new_n17063_), .ZN(new_n17248_));
  AOI21_X1   g16991(.A1(new_n17247_), .A2(new_n17248_), .B(new_n17245_), .ZN(new_n17249_));
  NOR2_X1    g16992(.A1(new_n17244_), .A2(new_n17249_), .ZN(new_n17250_));
  XOR2_X1    g16993(.A1(new_n17057_), .A2(new_n17250_), .Z(new_n17251_));
  AOI21_X1   g16994(.A1(new_n16851_), .A2(new_n16852_), .B(new_n16850_), .ZN(new_n17252_));
  NAND3_X1   g16995(.A1(new_n16649_), .A2(new_n16843_), .A3(new_n16844_), .ZN(new_n17253_));
  INV_X1     g16996(.I(new_n17253_), .ZN(new_n17254_));
  NOR3_X1    g16997(.A1(new_n17252_), .A2(new_n17254_), .A3(new_n16857_), .ZN(new_n17255_));
  AOI21_X1   g16998(.A1(new_n16849_), .A2(new_n17253_), .B(new_n16858_), .ZN(new_n17256_));
  OAI21_X1   g16999(.A1(new_n17256_), .A2(new_n17255_), .B(new_n17049_), .ZN(new_n17257_));
  XNOR2_X1   g17000(.A1(new_n17257_), .A2(new_n17251_), .ZN(new_n17258_));
  NAND2_X1   g17001(.A1(new_n16856_), .A2(new_n16858_), .ZN(new_n17259_));
  XOR2_X1    g17002(.A1(new_n17258_), .A2(new_n17259_), .Z(\f[90] ));
  NOR2_X1    g17003(.A1(new_n2214_), .A2(new_n8932_), .ZN(new_n17261_));
  NOR2_X1    g17004(.A1(new_n2079_), .A2(new_n8956_), .ZN(new_n17262_));
  NOR4_X1    g17005(.A1(new_n9323_), .A2(new_n2087_), .A3(new_n17261_), .A4(new_n17262_), .ZN(new_n17263_));
  XOR2_X1    g17006(.A1(new_n17263_), .A2(new_n2074_), .Z(new_n17264_));
  NAND2_X1   g17007(.A1(new_n17228_), .A2(new_n17240_), .ZN(new_n17265_));
  NAND2_X1   g17008(.A1(new_n17265_), .A2(new_n17239_), .ZN(new_n17266_));
  OAI22_X1   g17009(.A1(new_n2452_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n2447_), .ZN(new_n17267_));
  NAND2_X1   g17010(.A1(new_n3312_), .A2(\b[59] ), .ZN(new_n17268_));
  AOI21_X1   g17011(.A1(new_n17267_), .A2(new_n17268_), .B(new_n2455_), .ZN(new_n17269_));
  NAND2_X1   g17012(.A1(new_n8550_), .A2(new_n17269_), .ZN(new_n17270_));
  XOR2_X1    g17013(.A1(new_n17270_), .A2(\a[32] ), .Z(new_n17271_));
  AOI21_X1   g17014(.A1(new_n17066_), .A2(new_n17226_), .B(new_n17224_), .ZN(new_n17272_));
  OAI22_X1   g17015(.A1(new_n2846_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n2841_), .ZN(new_n17273_));
  NAND2_X1   g17016(.A1(new_n3755_), .A2(\b[56] ), .ZN(new_n17274_));
  AOI21_X1   g17017(.A1(new_n17273_), .A2(new_n17274_), .B(new_n2849_), .ZN(new_n17275_));
  NAND2_X1   g17018(.A1(new_n7559_), .A2(new_n17275_), .ZN(new_n17276_));
  XOR2_X1    g17019(.A1(new_n17276_), .A2(\a[35] ), .Z(new_n17277_));
  AOI21_X1   g17020(.A1(new_n17210_), .A2(new_n17213_), .B(new_n17211_), .ZN(new_n17278_));
  INV_X1     g17021(.I(new_n17278_), .ZN(new_n17279_));
  INV_X1     g17022(.I(new_n17196_), .ZN(new_n17280_));
  AOI21_X1   g17023(.A1(new_n17199_), .A2(new_n17280_), .B(new_n17194_), .ZN(new_n17281_));
  OAI22_X1   g17024(.A1(new_n3736_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n3731_), .ZN(new_n17282_));
  NAND2_X1   g17025(.A1(new_n4730_), .A2(\b[50] ), .ZN(new_n17283_));
  AOI21_X1   g17026(.A1(new_n17282_), .A2(new_n17283_), .B(new_n3739_), .ZN(new_n17284_));
  NAND2_X1   g17027(.A1(new_n5954_), .A2(new_n17284_), .ZN(new_n17285_));
  XOR2_X1    g17028(.A1(new_n17285_), .A2(\a[41] ), .Z(new_n17286_));
  OAI22_X1   g17029(.A1(new_n4711_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n4706_), .ZN(new_n17287_));
  NAND2_X1   g17030(.A1(new_n5814_), .A2(\b[44] ), .ZN(new_n17288_));
  AOI21_X1   g17031(.A1(new_n17287_), .A2(new_n17288_), .B(new_n4714_), .ZN(new_n17289_));
  NAND2_X1   g17032(.A1(new_n4833_), .A2(new_n17289_), .ZN(new_n17290_));
  XOR2_X1    g17033(.A1(new_n17290_), .A2(\a[47] ), .Z(new_n17291_));
  NOR2_X1    g17034(.A1(new_n17144_), .A2(new_n17076_), .ZN(new_n17292_));
  NOR2_X1    g17035(.A1(new_n17292_), .A2(new_n17142_), .ZN(new_n17293_));
  OAI22_X1   g17036(.A1(new_n5786_), .A2(new_n3845_), .B1(new_n3696_), .B2(new_n5792_), .ZN(new_n17294_));
  NAND2_X1   g17037(.A1(new_n6745_), .A2(\b[38] ), .ZN(new_n17295_));
  AOI21_X1   g17038(.A1(new_n17295_), .A2(new_n17294_), .B(new_n5796_), .ZN(new_n17296_));
  NAND2_X1   g17039(.A1(new_n3844_), .A2(new_n17296_), .ZN(new_n17297_));
  XOR2_X1    g17040(.A1(new_n17297_), .A2(\a[53] ), .Z(new_n17298_));
  INV_X1     g17041(.I(new_n17130_), .ZN(new_n17299_));
  AOI21_X1   g17042(.A1(new_n17119_), .A2(new_n17299_), .B(new_n17128_), .ZN(new_n17300_));
  OAI22_X1   g17043(.A1(new_n2964_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2794_), .ZN(new_n17301_));
  NAND2_X1   g17044(.A1(new_n8628_), .A2(\b[32] ), .ZN(new_n17302_));
  AOI21_X1   g17045(.A1(new_n17302_), .A2(new_n17301_), .B(new_n7354_), .ZN(new_n17303_));
  NAND2_X1   g17046(.A1(new_n2963_), .A2(new_n17303_), .ZN(new_n17304_));
  XOR2_X1    g17047(.A1(new_n17304_), .A2(\a[59] ), .Z(new_n17305_));
  INV_X1     g17048(.I(new_n17305_), .ZN(new_n17306_));
  OAI22_X1   g17049(.A1(new_n2543_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2405_), .ZN(new_n17307_));
  NAND2_X1   g17050(.A1(new_n9644_), .A2(\b[29] ), .ZN(new_n17308_));
  AOI21_X1   g17051(.A1(new_n17308_), .A2(new_n17307_), .B(new_n8321_), .ZN(new_n17309_));
  NAND2_X1   g17052(.A1(new_n2546_), .A2(new_n17309_), .ZN(new_n17310_));
  XOR2_X1    g17053(.A1(new_n17310_), .A2(\a[62] ), .Z(new_n17311_));
  NAND2_X1   g17054(.A1(new_n17100_), .A2(new_n16929_), .ZN(new_n17312_));
  NAND2_X1   g17055(.A1(new_n17312_), .A2(new_n17099_), .ZN(new_n17313_));
  NOR3_X1    g17056(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n2039_), .ZN(new_n17314_));
  NOR2_X1    g17057(.A1(new_n9364_), .A2(new_n2039_), .ZN(new_n17315_));
  NOR3_X1    g17058(.A1(new_n17315_), .A2(new_n2175_), .A3(new_n8985_), .ZN(new_n17316_));
  NOR2_X1    g17059(.A1(new_n17316_), .A2(new_n17314_), .ZN(new_n17317_));
  INV_X1     g17060(.I(new_n17317_), .ZN(new_n17318_));
  XOR2_X1    g17061(.A1(new_n17313_), .A2(new_n17318_), .Z(new_n17319_));
  NOR2_X1    g17062(.A1(new_n17313_), .A2(new_n17317_), .ZN(new_n17320_));
  NAND2_X1   g17063(.A1(new_n17313_), .A2(new_n17317_), .ZN(new_n17321_));
  INV_X1     g17064(.I(new_n17321_), .ZN(new_n17322_));
  OAI21_X1   g17065(.A1(new_n17320_), .A2(new_n17322_), .B(new_n17311_), .ZN(new_n17323_));
  OAI21_X1   g17066(.A1(new_n17311_), .A2(new_n17319_), .B(new_n17323_), .ZN(new_n17324_));
  NAND2_X1   g17067(.A1(new_n17086_), .A2(new_n17104_), .ZN(new_n17325_));
  NAND2_X1   g17068(.A1(new_n17325_), .A2(new_n17105_), .ZN(new_n17326_));
  INV_X1     g17069(.I(new_n17326_), .ZN(new_n17327_));
  NOR2_X1    g17070(.A1(new_n17327_), .A2(new_n17324_), .ZN(new_n17328_));
  INV_X1     g17071(.I(new_n17328_), .ZN(new_n17329_));
  NAND2_X1   g17072(.A1(new_n17327_), .A2(new_n17324_), .ZN(new_n17330_));
  NAND2_X1   g17073(.A1(new_n17329_), .A2(new_n17330_), .ZN(new_n17331_));
  NAND2_X1   g17074(.A1(new_n17331_), .A2(new_n17306_), .ZN(new_n17332_));
  XNOR2_X1   g17075(.A1(new_n17324_), .A2(new_n17326_), .ZN(new_n17333_));
  NAND2_X1   g17076(.A1(new_n17333_), .A2(new_n17305_), .ZN(new_n17334_));
  NAND2_X1   g17077(.A1(new_n17332_), .A2(new_n17334_), .ZN(new_n17335_));
  NAND2_X1   g17078(.A1(new_n17117_), .A2(new_n17077_), .ZN(new_n17336_));
  NAND2_X1   g17079(.A1(new_n17336_), .A2(new_n17114_), .ZN(new_n17337_));
  INV_X1     g17080(.I(new_n17337_), .ZN(new_n17338_));
  OAI22_X1   g17081(.A1(new_n6721_), .A2(new_n3247_), .B1(new_n6723_), .B2(new_n3408_), .ZN(new_n17339_));
  NAND2_X1   g17082(.A1(new_n7617_), .A2(\b[35] ), .ZN(new_n17340_));
  AOI21_X1   g17083(.A1(new_n17340_), .A2(new_n17339_), .B(new_n6731_), .ZN(new_n17341_));
  NAND2_X1   g17084(.A1(new_n3411_), .A2(new_n17341_), .ZN(new_n17342_));
  XOR2_X1    g17085(.A1(new_n17342_), .A2(\a[56] ), .Z(new_n17343_));
  NOR2_X1    g17086(.A1(new_n17338_), .A2(new_n17343_), .ZN(new_n17344_));
  INV_X1     g17087(.I(new_n17343_), .ZN(new_n17345_));
  NOR2_X1    g17088(.A1(new_n17337_), .A2(new_n17345_), .ZN(new_n17346_));
  OAI21_X1   g17089(.A1(new_n17344_), .A2(new_n17346_), .B(new_n17335_), .ZN(new_n17347_));
  XOR2_X1    g17090(.A1(new_n17337_), .A2(new_n17343_), .Z(new_n17348_));
  OAI21_X1   g17091(.A1(new_n17335_), .A2(new_n17348_), .B(new_n17347_), .ZN(new_n17349_));
  XOR2_X1    g17092(.A1(new_n17300_), .A2(new_n17349_), .Z(new_n17350_));
  INV_X1     g17093(.I(new_n17349_), .ZN(new_n17351_));
  NOR2_X1    g17094(.A1(new_n17300_), .A2(new_n17351_), .ZN(new_n17352_));
  INV_X1     g17095(.I(new_n17352_), .ZN(new_n17353_));
  NAND2_X1   g17096(.A1(new_n17300_), .A2(new_n17351_), .ZN(new_n17354_));
  NAND2_X1   g17097(.A1(new_n17353_), .A2(new_n17354_), .ZN(new_n17355_));
  NAND2_X1   g17098(.A1(new_n17355_), .A2(new_n17298_), .ZN(new_n17356_));
  OAI21_X1   g17099(.A1(new_n17298_), .A2(new_n17350_), .B(new_n17356_), .ZN(new_n17357_));
  OAI22_X1   g17100(.A1(new_n5228_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n5225_), .ZN(new_n17358_));
  NAND2_X1   g17101(.A1(new_n5387_), .A2(\b[41] ), .ZN(new_n17359_));
  AOI21_X1   g17102(.A1(new_n17358_), .A2(new_n17359_), .B(new_n5231_), .ZN(new_n17360_));
  NAND2_X1   g17103(.A1(new_n4320_), .A2(new_n17360_), .ZN(new_n17361_));
  XOR2_X1    g17104(.A1(new_n17361_), .A2(\a[50] ), .Z(new_n17362_));
  NOR2_X1    g17105(.A1(new_n17357_), .A2(new_n17362_), .ZN(new_n17363_));
  INV_X1     g17106(.I(new_n17363_), .ZN(new_n17364_));
  NAND2_X1   g17107(.A1(new_n17357_), .A2(new_n17362_), .ZN(new_n17365_));
  AOI21_X1   g17108(.A1(new_n17364_), .A2(new_n17365_), .B(new_n17293_), .ZN(new_n17366_));
  INV_X1     g17109(.I(new_n17293_), .ZN(new_n17367_));
  XNOR2_X1   g17110(.A1(new_n17357_), .A2(new_n17362_), .ZN(new_n17368_));
  NOR2_X1    g17111(.A1(new_n17368_), .A2(new_n17367_), .ZN(new_n17369_));
  NOR2_X1    g17112(.A1(new_n17369_), .A2(new_n17366_), .ZN(new_n17370_));
  AOI21_X1   g17113(.A1(new_n17156_), .A2(new_n17154_), .B(new_n17152_), .ZN(new_n17371_));
  NOR2_X1    g17114(.A1(new_n17370_), .A2(new_n17371_), .ZN(new_n17372_));
  INV_X1     g17115(.I(new_n17372_), .ZN(new_n17373_));
  NAND2_X1   g17116(.A1(new_n17370_), .A2(new_n17371_), .ZN(new_n17374_));
  AOI21_X1   g17117(.A1(new_n17373_), .A2(new_n17374_), .B(new_n17291_), .ZN(new_n17375_));
  INV_X1     g17118(.I(new_n17291_), .ZN(new_n17376_));
  XNOR2_X1   g17119(.A1(new_n17370_), .A2(new_n17371_), .ZN(new_n17377_));
  NOR2_X1    g17120(.A1(new_n17377_), .A2(new_n17376_), .ZN(new_n17378_));
  NOR2_X1    g17121(.A1(new_n17378_), .A2(new_n17375_), .ZN(new_n17379_));
  NOR2_X1    g17122(.A1(new_n17169_), .A2(new_n17071_), .ZN(new_n17380_));
  NOR2_X1    g17123(.A1(new_n17380_), .A2(new_n17167_), .ZN(new_n17381_));
  OAI22_X1   g17124(.A1(new_n4208_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n4203_), .ZN(new_n17382_));
  NAND2_X1   g17125(.A1(new_n5244_), .A2(\b[47] ), .ZN(new_n17383_));
  AOI21_X1   g17126(.A1(new_n17382_), .A2(new_n17383_), .B(new_n4211_), .ZN(new_n17384_));
  NAND2_X1   g17127(.A1(new_n5196_), .A2(new_n17384_), .ZN(new_n17385_));
  XOR2_X1    g17128(.A1(new_n17385_), .A2(\a[44] ), .Z(new_n17386_));
  NOR2_X1    g17129(.A1(new_n17381_), .A2(new_n17386_), .ZN(new_n17387_));
  INV_X1     g17130(.I(new_n17386_), .ZN(new_n17388_));
  NOR3_X1    g17131(.A1(new_n17380_), .A2(new_n17167_), .A3(new_n17388_), .ZN(new_n17389_));
  NOR2_X1    g17132(.A1(new_n17387_), .A2(new_n17389_), .ZN(new_n17390_));
  NOR2_X1    g17133(.A1(new_n17390_), .A2(new_n17379_), .ZN(new_n17391_));
  INV_X1     g17134(.I(new_n17379_), .ZN(new_n17392_));
  XOR2_X1    g17135(.A1(new_n17381_), .A2(new_n17388_), .Z(new_n17393_));
  NOR2_X1    g17136(.A1(new_n17393_), .A2(new_n17392_), .ZN(new_n17394_));
  NOR2_X1    g17137(.A1(new_n17394_), .A2(new_n17391_), .ZN(new_n17395_));
  NAND2_X1   g17138(.A1(new_n17172_), .A2(new_n17182_), .ZN(new_n17396_));
  NAND2_X1   g17139(.A1(new_n17396_), .A2(new_n17181_), .ZN(new_n17397_));
  INV_X1     g17140(.I(new_n17397_), .ZN(new_n17398_));
  NOR2_X1    g17141(.A1(new_n17395_), .A2(new_n17398_), .ZN(new_n17399_));
  NOR3_X1    g17142(.A1(new_n17394_), .A2(new_n17397_), .A3(new_n17391_), .ZN(new_n17400_));
  NOR2_X1    g17143(.A1(new_n17399_), .A2(new_n17400_), .ZN(new_n17401_));
  NOR2_X1    g17144(.A1(new_n17401_), .A2(new_n17286_), .ZN(new_n17402_));
  XOR2_X1    g17145(.A1(new_n17395_), .A2(new_n17398_), .Z(new_n17403_));
  AOI21_X1   g17146(.A1(new_n17286_), .A2(new_n17403_), .B(new_n17402_), .ZN(new_n17404_));
  OAI22_X1   g17147(.A1(new_n3298_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n3293_), .ZN(new_n17405_));
  NAND2_X1   g17148(.A1(new_n4227_), .A2(\b[53] ), .ZN(new_n17406_));
  AOI21_X1   g17149(.A1(new_n17405_), .A2(new_n17406_), .B(new_n3301_), .ZN(new_n17407_));
  NAND2_X1   g17150(.A1(new_n6471_), .A2(new_n17407_), .ZN(new_n17408_));
  XOR2_X1    g17151(.A1(new_n17408_), .A2(\a[38] ), .Z(new_n17409_));
  XNOR2_X1   g17152(.A1(new_n17404_), .A2(new_n17409_), .ZN(new_n17410_));
  NOR2_X1    g17153(.A1(new_n17410_), .A2(new_n17281_), .ZN(new_n17411_));
  INV_X1     g17154(.I(new_n17281_), .ZN(new_n17412_));
  NOR2_X1    g17155(.A1(new_n17404_), .A2(new_n17409_), .ZN(new_n17413_));
  INV_X1     g17156(.I(new_n17413_), .ZN(new_n17414_));
  NAND2_X1   g17157(.A1(new_n17404_), .A2(new_n17409_), .ZN(new_n17415_));
  AOI21_X1   g17158(.A1(new_n17414_), .A2(new_n17415_), .B(new_n17412_), .ZN(new_n17416_));
  NOR2_X1    g17159(.A1(new_n17411_), .A2(new_n17416_), .ZN(new_n17417_));
  NOR2_X1    g17160(.A1(new_n17417_), .A2(new_n17279_), .ZN(new_n17418_));
  INV_X1     g17161(.I(new_n17418_), .ZN(new_n17419_));
  NAND2_X1   g17162(.A1(new_n17417_), .A2(new_n17279_), .ZN(new_n17420_));
  AOI21_X1   g17163(.A1(new_n17419_), .A2(new_n17420_), .B(new_n17277_), .ZN(new_n17421_));
  XOR2_X1    g17164(.A1(new_n17417_), .A2(new_n17278_), .Z(new_n17422_));
  INV_X1     g17165(.I(new_n17422_), .ZN(new_n17423_));
  AOI21_X1   g17166(.A1(new_n17423_), .A2(new_n17277_), .B(new_n17421_), .ZN(new_n17424_));
  XNOR2_X1   g17167(.A1(new_n17424_), .A2(new_n17272_), .ZN(new_n17425_));
  NOR2_X1    g17168(.A1(new_n17425_), .A2(new_n17271_), .ZN(new_n17426_));
  INV_X1     g17169(.I(new_n17271_), .ZN(new_n17427_));
  NOR2_X1    g17170(.A1(new_n17424_), .A2(new_n17272_), .ZN(new_n17428_));
  INV_X1     g17171(.I(new_n17428_), .ZN(new_n17429_));
  NAND2_X1   g17172(.A1(new_n17424_), .A2(new_n17272_), .ZN(new_n17430_));
  AOI21_X1   g17173(.A1(new_n17429_), .A2(new_n17430_), .B(new_n17427_), .ZN(new_n17431_));
  NOR2_X1    g17174(.A1(new_n17426_), .A2(new_n17431_), .ZN(new_n17432_));
  NOR2_X1    g17175(.A1(new_n17432_), .A2(new_n17266_), .ZN(new_n17433_));
  INV_X1     g17176(.I(new_n17266_), .ZN(new_n17434_));
  INV_X1     g17177(.I(new_n17432_), .ZN(new_n17435_));
  NOR2_X1    g17178(.A1(new_n17435_), .A2(new_n17434_), .ZN(new_n17436_));
  NOR2_X1    g17179(.A1(new_n17436_), .A2(new_n17433_), .ZN(new_n17437_));
  NOR2_X1    g17180(.A1(new_n17437_), .A2(new_n17264_), .ZN(new_n17438_));
  INV_X1     g17181(.I(new_n17264_), .ZN(new_n17439_));
  XOR2_X1    g17182(.A1(new_n17432_), .A2(new_n17434_), .Z(new_n17440_));
  NOR2_X1    g17183(.A1(new_n17440_), .A2(new_n17439_), .ZN(new_n17441_));
  NOR2_X1    g17184(.A1(new_n17438_), .A2(new_n17441_), .ZN(new_n17442_));
  AOI21_X1   g17185(.A1(new_n17245_), .A2(new_n17248_), .B(new_n17246_), .ZN(new_n17443_));
  NAND3_X1   g17186(.A1(new_n16849_), .A2(new_n17253_), .A3(new_n16858_), .ZN(new_n17444_));
  NAND2_X1   g17187(.A1(new_n16856_), .A2(new_n16857_), .ZN(new_n17445_));
  NAND2_X1   g17188(.A1(new_n17445_), .A2(new_n17444_), .ZN(new_n17446_));
  NAND3_X1   g17189(.A1(new_n16856_), .A2(new_n16858_), .A3(new_n17251_), .ZN(new_n17447_));
  NAND3_X1   g17190(.A1(new_n17446_), .A2(new_n17049_), .A3(new_n17447_), .ZN(new_n17448_));
  OAI21_X1   g17191(.A1(new_n17244_), .A2(new_n17249_), .B(new_n17057_), .ZN(new_n17449_));
  NAND2_X1   g17192(.A1(new_n17448_), .A2(new_n17449_), .ZN(new_n17450_));
  XOR2_X1    g17193(.A1(new_n17450_), .A2(new_n17443_), .Z(new_n17451_));
  XOR2_X1    g17194(.A1(new_n17451_), .A2(new_n17442_), .Z(\f[91] ));
  XOR2_X1    g17195(.A1(new_n17442_), .A2(new_n17443_), .Z(new_n17453_));
  NAND2_X1   g17196(.A1(new_n17453_), .A2(new_n17443_), .ZN(new_n17454_));
  INV_X1     g17197(.I(new_n17454_), .ZN(new_n17455_));
  NAND2_X1   g17198(.A1(new_n17449_), .A2(new_n17453_), .ZN(new_n17456_));
  INV_X1     g17199(.I(new_n17456_), .ZN(new_n17457_));
  AOI21_X1   g17200(.A1(new_n17448_), .A2(new_n17457_), .B(new_n17455_), .ZN(new_n17458_));
  NOR2_X1    g17201(.A1(new_n17433_), .A2(new_n17264_), .ZN(new_n17459_));
  NOR2_X1    g17202(.A1(new_n17459_), .A2(new_n17436_), .ZN(new_n17460_));
  INV_X1     g17203(.I(new_n17460_), .ZN(new_n17461_));
  NAND2_X1   g17204(.A1(new_n17430_), .A2(new_n17427_), .ZN(new_n17462_));
  NAND2_X1   g17205(.A1(new_n17462_), .A2(new_n17429_), .ZN(new_n17463_));
  OAI22_X1   g17206(.A1(new_n9595_), .A2(new_n2087_), .B1(new_n8956_), .B2(new_n2214_), .ZN(new_n17464_));
  OAI22_X1   g17207(.A1(new_n2452_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n2447_), .ZN(new_n17465_));
  NAND2_X1   g17208(.A1(new_n3312_), .A2(\b[60] ), .ZN(new_n17466_));
  AOI21_X1   g17209(.A1(new_n17465_), .A2(new_n17466_), .B(new_n2455_), .ZN(new_n17467_));
  NAND2_X1   g17210(.A1(new_n8935_), .A2(new_n17467_), .ZN(new_n17468_));
  XOR2_X1    g17211(.A1(new_n17468_), .A2(\a[32] ), .Z(new_n17469_));
  OAI21_X1   g17212(.A1(new_n17277_), .A2(new_n17418_), .B(new_n17420_), .ZN(new_n17470_));
  OAI22_X1   g17213(.A1(new_n3298_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n3293_), .ZN(new_n17471_));
  NAND2_X1   g17214(.A1(new_n4227_), .A2(\b[54] ), .ZN(new_n17472_));
  AOI21_X1   g17215(.A1(new_n17471_), .A2(new_n17472_), .B(new_n3301_), .ZN(new_n17473_));
  NAND2_X1   g17216(.A1(new_n6994_), .A2(new_n17473_), .ZN(new_n17474_));
  XOR2_X1    g17217(.A1(new_n17474_), .A2(\a[38] ), .Z(new_n17475_));
  INV_X1     g17218(.I(new_n17286_), .ZN(new_n17476_));
  INV_X1     g17219(.I(new_n17400_), .ZN(new_n17477_));
  AOI21_X1   g17220(.A1(new_n17477_), .A2(new_n17476_), .B(new_n17399_), .ZN(new_n17478_));
  OAI22_X1   g17221(.A1(new_n3736_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n3731_), .ZN(new_n17479_));
  NAND2_X1   g17222(.A1(new_n4730_), .A2(\b[51] ), .ZN(new_n17480_));
  AOI21_X1   g17223(.A1(new_n17479_), .A2(new_n17480_), .B(new_n3739_), .ZN(new_n17481_));
  NAND2_X1   g17224(.A1(new_n6219_), .A2(new_n17481_), .ZN(new_n17482_));
  XOR2_X1    g17225(.A1(new_n17482_), .A2(\a[41] ), .Z(new_n17483_));
  OAI22_X1   g17226(.A1(new_n4208_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n4203_), .ZN(new_n17484_));
  NAND2_X1   g17227(.A1(new_n5244_), .A2(\b[48] ), .ZN(new_n17485_));
  AOI21_X1   g17228(.A1(new_n17484_), .A2(new_n17485_), .B(new_n4211_), .ZN(new_n17486_));
  NAND2_X1   g17229(.A1(new_n5537_), .A2(new_n17486_), .ZN(new_n17487_));
  XOR2_X1    g17230(.A1(new_n17487_), .A2(\a[44] ), .Z(new_n17488_));
  OAI22_X1   g17231(.A1(new_n5228_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n5225_), .ZN(new_n17489_));
  NAND2_X1   g17232(.A1(new_n5387_), .A2(\b[42] ), .ZN(new_n17490_));
  AOI21_X1   g17233(.A1(new_n17489_), .A2(new_n17490_), .B(new_n5231_), .ZN(new_n17491_));
  NAND2_X1   g17234(.A1(new_n4500_), .A2(new_n17491_), .ZN(new_n17492_));
  XOR2_X1    g17235(.A1(new_n17492_), .A2(\a[50] ), .Z(new_n17493_));
  INV_X1     g17236(.I(new_n17354_), .ZN(new_n17494_));
  OAI21_X1   g17237(.A1(new_n17298_), .A2(new_n17494_), .B(new_n17353_), .ZN(new_n17495_));
  OAI22_X1   g17238(.A1(new_n6721_), .A2(new_n3408_), .B1(new_n6723_), .B2(new_n3566_), .ZN(new_n17496_));
  NAND2_X1   g17239(.A1(new_n7617_), .A2(\b[36] ), .ZN(new_n17497_));
  AOI21_X1   g17240(.A1(new_n17497_), .A2(new_n17496_), .B(new_n6731_), .ZN(new_n17498_));
  NAND2_X1   g17241(.A1(new_n3565_), .A2(new_n17498_), .ZN(new_n17499_));
  XOR2_X1    g17242(.A1(new_n17499_), .A2(\a[56] ), .Z(new_n17500_));
  INV_X1     g17243(.I(new_n17500_), .ZN(new_n17501_));
  AOI21_X1   g17244(.A1(new_n17306_), .A2(new_n17330_), .B(new_n17328_), .ZN(new_n17502_));
  INV_X1     g17245(.I(new_n17502_), .ZN(new_n17503_));
  OAI22_X1   g17246(.A1(new_n3097_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n2964_), .ZN(new_n17504_));
  NAND2_X1   g17247(.A1(new_n8628_), .A2(\b[33] ), .ZN(new_n17505_));
  AOI21_X1   g17248(.A1(new_n17505_), .A2(new_n17504_), .B(new_n7354_), .ZN(new_n17506_));
  NAND2_X1   g17249(.A1(new_n3101_), .A2(new_n17506_), .ZN(new_n17507_));
  XOR2_X1    g17250(.A1(new_n17507_), .A2(\a[59] ), .Z(new_n17508_));
  OAI21_X1   g17251(.A1(new_n17311_), .A2(new_n17320_), .B(new_n17321_), .ZN(new_n17509_));
  NOR3_X1    g17252(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n2175_), .ZN(new_n17510_));
  NOR2_X1    g17253(.A1(new_n9364_), .A2(new_n2175_), .ZN(new_n17511_));
  NOR3_X1    g17254(.A1(new_n17511_), .A2(new_n2272_), .A3(new_n8985_), .ZN(new_n17512_));
  NOR2_X1    g17255(.A1(new_n17512_), .A2(new_n17510_), .ZN(new_n17513_));
  NOR2_X1    g17256(.A1(new_n17318_), .A2(new_n17513_), .ZN(new_n17514_));
  INV_X1     g17257(.I(new_n17514_), .ZN(new_n17515_));
  INV_X1     g17258(.I(new_n17513_), .ZN(new_n17516_));
  NOR2_X1    g17259(.A1(new_n17516_), .A2(new_n17317_), .ZN(new_n17517_));
  INV_X1     g17260(.I(new_n17517_), .ZN(new_n17518_));
  NAND2_X1   g17261(.A1(new_n17515_), .A2(new_n17518_), .ZN(new_n17519_));
  XOR2_X1    g17262(.A1(new_n17317_), .A2(new_n17513_), .Z(new_n17520_));
  NOR2_X1    g17263(.A1(new_n17509_), .A2(new_n17520_), .ZN(new_n17521_));
  AOI21_X1   g17264(.A1(new_n17509_), .A2(new_n17519_), .B(new_n17521_), .ZN(new_n17522_));
  OAI22_X1   g17265(.A1(new_n2660_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2543_), .ZN(new_n17523_));
  NAND2_X1   g17266(.A1(new_n9644_), .A2(\b[30] ), .ZN(new_n17524_));
  AOI21_X1   g17267(.A1(new_n17524_), .A2(new_n17523_), .B(new_n8321_), .ZN(new_n17525_));
  NAND2_X1   g17268(.A1(new_n2659_), .A2(new_n17525_), .ZN(new_n17526_));
  XOR2_X1    g17269(.A1(new_n17526_), .A2(\a[62] ), .Z(new_n17527_));
  XNOR2_X1   g17270(.A1(new_n17522_), .A2(new_n17527_), .ZN(new_n17528_));
  NOR2_X1    g17271(.A1(new_n17528_), .A2(new_n17508_), .ZN(new_n17529_));
  INV_X1     g17272(.I(new_n17508_), .ZN(new_n17530_));
  NOR2_X1    g17273(.A1(new_n17522_), .A2(new_n17527_), .ZN(new_n17531_));
  INV_X1     g17274(.I(new_n17531_), .ZN(new_n17532_));
  NAND2_X1   g17275(.A1(new_n17522_), .A2(new_n17527_), .ZN(new_n17533_));
  AOI21_X1   g17276(.A1(new_n17532_), .A2(new_n17533_), .B(new_n17530_), .ZN(new_n17534_));
  NOR2_X1    g17277(.A1(new_n17529_), .A2(new_n17534_), .ZN(new_n17535_));
  NOR2_X1    g17278(.A1(new_n17535_), .A2(new_n17503_), .ZN(new_n17536_));
  NAND2_X1   g17279(.A1(new_n17535_), .A2(new_n17503_), .ZN(new_n17537_));
  INV_X1     g17280(.I(new_n17537_), .ZN(new_n17538_));
  OAI21_X1   g17281(.A1(new_n17538_), .A2(new_n17536_), .B(new_n17501_), .ZN(new_n17539_));
  XOR2_X1    g17282(.A1(new_n17535_), .A2(new_n17502_), .Z(new_n17540_));
  OAI21_X1   g17283(.A1(new_n17501_), .A2(new_n17540_), .B(new_n17539_), .ZN(new_n17541_));
  INV_X1     g17284(.I(new_n17344_), .ZN(new_n17542_));
  OAI22_X1   g17285(.A1(new_n5786_), .A2(new_n3997_), .B1(new_n3845_), .B2(new_n5792_), .ZN(new_n17543_));
  NAND2_X1   g17286(.A1(new_n6745_), .A2(\b[39] ), .ZN(new_n17544_));
  AOI21_X1   g17287(.A1(new_n17544_), .A2(new_n17543_), .B(new_n5796_), .ZN(new_n17545_));
  NAND2_X1   g17288(.A1(new_n3996_), .A2(new_n17545_), .ZN(new_n17546_));
  XOR2_X1    g17289(.A1(new_n17546_), .A2(\a[53] ), .Z(new_n17547_));
  OAI21_X1   g17290(.A1(new_n17337_), .A2(new_n17345_), .B(new_n17335_), .ZN(new_n17548_));
  AOI21_X1   g17291(.A1(new_n17548_), .A2(new_n17542_), .B(new_n17547_), .ZN(new_n17549_));
  INV_X1     g17292(.I(new_n17547_), .ZN(new_n17550_));
  NAND2_X1   g17293(.A1(new_n17548_), .A2(new_n17542_), .ZN(new_n17551_));
  NOR2_X1    g17294(.A1(new_n17551_), .A2(new_n17550_), .ZN(new_n17552_));
  OAI21_X1   g17295(.A1(new_n17549_), .A2(new_n17552_), .B(new_n17541_), .ZN(new_n17553_));
  XOR2_X1    g17296(.A1(new_n17551_), .A2(new_n17547_), .Z(new_n17554_));
  OAI21_X1   g17297(.A1(new_n17541_), .A2(new_n17554_), .B(new_n17553_), .ZN(new_n17555_));
  XNOR2_X1   g17298(.A1(new_n17555_), .A2(new_n17495_), .ZN(new_n17556_));
  NOR2_X1    g17299(.A1(new_n17556_), .A2(new_n17493_), .ZN(new_n17557_));
  INV_X1     g17300(.I(new_n17493_), .ZN(new_n17558_));
  NAND2_X1   g17301(.A1(new_n17555_), .A2(new_n17495_), .ZN(new_n17559_));
  NOR2_X1    g17302(.A1(new_n17555_), .A2(new_n17495_), .ZN(new_n17560_));
  INV_X1     g17303(.I(new_n17560_), .ZN(new_n17561_));
  AOI21_X1   g17304(.A1(new_n17561_), .A2(new_n17559_), .B(new_n17558_), .ZN(new_n17562_));
  NOR2_X1    g17305(.A1(new_n17557_), .A2(new_n17562_), .ZN(new_n17563_));
  OAI22_X1   g17306(.A1(new_n4711_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n4706_), .ZN(new_n17564_));
  NAND2_X1   g17307(.A1(new_n5814_), .A2(\b[45] ), .ZN(new_n17565_));
  AOI21_X1   g17308(.A1(new_n17564_), .A2(new_n17565_), .B(new_n4714_), .ZN(new_n17566_));
  NAND2_X1   g17309(.A1(new_n5004_), .A2(new_n17566_), .ZN(new_n17567_));
  XOR2_X1    g17310(.A1(new_n17567_), .A2(\a[47] ), .Z(new_n17568_));
  NAND2_X1   g17311(.A1(new_n17365_), .A2(new_n17367_), .ZN(new_n17569_));
  NAND2_X1   g17312(.A1(new_n17569_), .A2(new_n17364_), .ZN(new_n17570_));
  XOR2_X1    g17313(.A1(new_n17570_), .A2(new_n17568_), .Z(new_n17571_));
  NOR2_X1    g17314(.A1(new_n17571_), .A2(new_n17563_), .ZN(new_n17572_));
  INV_X1     g17315(.I(new_n17570_), .ZN(new_n17573_));
  NOR2_X1    g17316(.A1(new_n17573_), .A2(new_n17568_), .ZN(new_n17574_));
  INV_X1     g17317(.I(new_n17574_), .ZN(new_n17575_));
  NAND2_X1   g17318(.A1(new_n17573_), .A2(new_n17568_), .ZN(new_n17576_));
  NAND2_X1   g17319(.A1(new_n17575_), .A2(new_n17576_), .ZN(new_n17577_));
  AOI21_X1   g17320(.A1(new_n17563_), .A2(new_n17577_), .B(new_n17572_), .ZN(new_n17578_));
  NAND2_X1   g17321(.A1(new_n17374_), .A2(new_n17376_), .ZN(new_n17579_));
  NAND2_X1   g17322(.A1(new_n17579_), .A2(new_n17373_), .ZN(new_n17580_));
  XOR2_X1    g17323(.A1(new_n17578_), .A2(new_n17580_), .Z(new_n17581_));
  NOR2_X1    g17324(.A1(new_n17581_), .A2(new_n17488_), .ZN(new_n17582_));
  INV_X1     g17325(.I(new_n17488_), .ZN(new_n17583_));
  INV_X1     g17326(.I(new_n17580_), .ZN(new_n17584_));
  NOR2_X1    g17327(.A1(new_n17584_), .A2(new_n17578_), .ZN(new_n17585_));
  INV_X1     g17328(.I(new_n17585_), .ZN(new_n17586_));
  NAND2_X1   g17329(.A1(new_n17584_), .A2(new_n17578_), .ZN(new_n17587_));
  AOI21_X1   g17330(.A1(new_n17586_), .A2(new_n17587_), .B(new_n17583_), .ZN(new_n17588_));
  NOR2_X1    g17331(.A1(new_n17582_), .A2(new_n17588_), .ZN(new_n17589_));
  NOR2_X1    g17332(.A1(new_n17379_), .A2(new_n17389_), .ZN(new_n17590_));
  NOR2_X1    g17333(.A1(new_n17590_), .A2(new_n17387_), .ZN(new_n17591_));
  XOR2_X1    g17334(.A1(new_n17589_), .A2(new_n17591_), .Z(new_n17592_));
  NOR2_X1    g17335(.A1(new_n17592_), .A2(new_n17483_), .ZN(new_n17593_));
  INV_X1     g17336(.I(new_n17483_), .ZN(new_n17594_));
  INV_X1     g17337(.I(new_n17589_), .ZN(new_n17595_));
  NOR2_X1    g17338(.A1(new_n17595_), .A2(new_n17591_), .ZN(new_n17596_));
  INV_X1     g17339(.I(new_n17596_), .ZN(new_n17597_));
  NAND2_X1   g17340(.A1(new_n17595_), .A2(new_n17591_), .ZN(new_n17598_));
  AOI21_X1   g17341(.A1(new_n17597_), .A2(new_n17598_), .B(new_n17594_), .ZN(new_n17599_));
  NOR2_X1    g17342(.A1(new_n17599_), .A2(new_n17593_), .ZN(new_n17600_));
  XOR2_X1    g17343(.A1(new_n17600_), .A2(new_n17478_), .Z(new_n17601_));
  NOR2_X1    g17344(.A1(new_n17601_), .A2(new_n17475_), .ZN(new_n17602_));
  INV_X1     g17345(.I(new_n17475_), .ZN(new_n17603_));
  INV_X1     g17346(.I(new_n17478_), .ZN(new_n17604_));
  NOR2_X1    g17347(.A1(new_n17600_), .A2(new_n17604_), .ZN(new_n17605_));
  INV_X1     g17348(.I(new_n17605_), .ZN(new_n17606_));
  NAND2_X1   g17349(.A1(new_n17600_), .A2(new_n17604_), .ZN(new_n17607_));
  AOI21_X1   g17350(.A1(new_n17606_), .A2(new_n17607_), .B(new_n17603_), .ZN(new_n17608_));
  NOR2_X1    g17351(.A1(new_n17602_), .A2(new_n17608_), .ZN(new_n17609_));
  OAI22_X1   g17352(.A1(new_n2846_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n2841_), .ZN(new_n17610_));
  NAND2_X1   g17353(.A1(new_n3755_), .A2(\b[57] ), .ZN(new_n17611_));
  AOI21_X1   g17354(.A1(new_n17610_), .A2(new_n17611_), .B(new_n2849_), .ZN(new_n17612_));
  NAND2_X1   g17355(.A1(new_n7895_), .A2(new_n17612_), .ZN(new_n17613_));
  XOR2_X1    g17356(.A1(new_n17613_), .A2(\a[35] ), .Z(new_n17614_));
  NAND2_X1   g17357(.A1(new_n17415_), .A2(new_n17412_), .ZN(new_n17615_));
  NAND2_X1   g17358(.A1(new_n17615_), .A2(new_n17414_), .ZN(new_n17616_));
  XOR2_X1    g17359(.A1(new_n17616_), .A2(new_n17614_), .Z(new_n17617_));
  NOR2_X1    g17360(.A1(new_n17617_), .A2(new_n17609_), .ZN(new_n17618_));
  INV_X1     g17361(.I(new_n17616_), .ZN(new_n17619_));
  NOR2_X1    g17362(.A1(new_n17619_), .A2(new_n17614_), .ZN(new_n17620_));
  INV_X1     g17363(.I(new_n17620_), .ZN(new_n17621_));
  NAND2_X1   g17364(.A1(new_n17619_), .A2(new_n17614_), .ZN(new_n17622_));
  NAND2_X1   g17365(.A1(new_n17621_), .A2(new_n17622_), .ZN(new_n17623_));
  AOI21_X1   g17366(.A1(new_n17609_), .A2(new_n17623_), .B(new_n17618_), .ZN(new_n17624_));
  XOR2_X1    g17367(.A1(new_n17624_), .A2(new_n17470_), .Z(new_n17625_));
  NOR2_X1    g17368(.A1(new_n17625_), .A2(new_n17469_), .ZN(new_n17626_));
  INV_X1     g17369(.I(new_n17469_), .ZN(new_n17627_));
  INV_X1     g17370(.I(new_n17470_), .ZN(new_n17628_));
  NOR2_X1    g17371(.A1(new_n17624_), .A2(new_n17628_), .ZN(new_n17629_));
  INV_X1     g17372(.I(new_n17629_), .ZN(new_n17630_));
  NAND2_X1   g17373(.A1(new_n17624_), .A2(new_n17628_), .ZN(new_n17631_));
  AOI21_X1   g17374(.A1(new_n17630_), .A2(new_n17631_), .B(new_n17627_), .ZN(new_n17632_));
  NOR2_X1    g17375(.A1(new_n17626_), .A2(new_n17632_), .ZN(new_n17633_));
  XOR2_X1    g17376(.A1(new_n17633_), .A2(new_n17464_), .Z(new_n17634_));
  XOR2_X1    g17377(.A1(new_n17634_), .A2(\a[29] ), .Z(new_n17635_));
  XOR2_X1    g17378(.A1(new_n17635_), .A2(new_n17463_), .Z(new_n17636_));
  XOR2_X1    g17379(.A1(new_n17636_), .A2(new_n17461_), .Z(new_n17637_));
  XOR2_X1    g17380(.A1(new_n17458_), .A2(new_n17637_), .Z(\f[92] ));
  XOR2_X1    g17381(.A1(new_n17464_), .A2(new_n2074_), .Z(new_n17639_));
  XOR2_X1    g17382(.A1(new_n17463_), .A2(new_n17639_), .Z(new_n17640_));
  INV_X1     g17383(.I(new_n17640_), .ZN(new_n17641_));
  OAI21_X1   g17384(.A1(new_n17633_), .A2(new_n17639_), .B(new_n17641_), .ZN(new_n17642_));
  AOI21_X1   g17385(.A1(new_n17627_), .A2(new_n17631_), .B(new_n17629_), .ZN(new_n17643_));
  OAI22_X1   g17386(.A1(new_n2452_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n2447_), .ZN(new_n17644_));
  NAND2_X1   g17387(.A1(new_n3312_), .A2(\b[61] ), .ZN(new_n17645_));
  AOI21_X1   g17388(.A1(new_n17644_), .A2(new_n17645_), .B(new_n2455_), .ZN(new_n17646_));
  NAND2_X1   g17389(.A1(new_n8963_), .A2(new_n17646_), .ZN(new_n17647_));
  XOR2_X1    g17390(.A1(new_n17647_), .A2(\a[32] ), .Z(new_n17648_));
  OAI21_X1   g17391(.A1(new_n17475_), .A2(new_n17605_), .B(new_n17607_), .ZN(new_n17649_));
  AOI21_X1   g17392(.A1(new_n17594_), .A2(new_n17598_), .B(new_n17596_), .ZN(new_n17650_));
  AOI21_X1   g17393(.A1(new_n17583_), .A2(new_n17587_), .B(new_n17585_), .ZN(new_n17651_));
  OAI21_X1   g17394(.A1(new_n17493_), .A2(new_n17560_), .B(new_n17559_), .ZN(new_n17652_));
  INV_X1     g17395(.I(new_n17652_), .ZN(new_n17653_));
  INV_X1     g17396(.I(new_n17552_), .ZN(new_n17654_));
  AOI21_X1   g17397(.A1(new_n17541_), .A2(new_n17654_), .B(new_n17549_), .ZN(new_n17655_));
  OAI21_X1   g17398(.A1(new_n17500_), .A2(new_n17536_), .B(new_n17537_), .ZN(new_n17656_));
  INV_X1     g17399(.I(new_n17656_), .ZN(new_n17657_));
  AOI21_X1   g17400(.A1(new_n17530_), .A2(new_n17533_), .B(new_n17531_), .ZN(new_n17658_));
  AOI21_X1   g17401(.A1(new_n17509_), .A2(new_n17515_), .B(new_n17517_), .ZN(new_n17659_));
  OAI22_X1   g17402(.A1(new_n2794_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2660_), .ZN(new_n17660_));
  NAND2_X1   g17403(.A1(new_n9644_), .A2(\b[31] ), .ZN(new_n17661_));
  AOI21_X1   g17404(.A1(new_n17661_), .A2(new_n17660_), .B(new_n8321_), .ZN(new_n17662_));
  NAND2_X1   g17405(.A1(new_n2797_), .A2(new_n17662_), .ZN(new_n17663_));
  XOR2_X1    g17406(.A1(new_n17663_), .A2(\a[62] ), .Z(new_n17664_));
  NOR2_X1    g17407(.A1(new_n8985_), .A2(new_n2405_), .ZN(new_n17665_));
  NOR2_X1    g17408(.A1(new_n9364_), .A2(new_n2272_), .ZN(new_n17666_));
  XNOR2_X1   g17409(.A1(new_n17665_), .A2(new_n17666_), .ZN(new_n17667_));
  NOR2_X1    g17410(.A1(new_n17667_), .A2(new_n2074_), .ZN(new_n17668_));
  INV_X1     g17411(.I(new_n17668_), .ZN(new_n17669_));
  NAND2_X1   g17412(.A1(new_n17667_), .A2(new_n2074_), .ZN(new_n17670_));
  AOI21_X1   g17413(.A1(new_n17669_), .A2(new_n17670_), .B(new_n17513_), .ZN(new_n17671_));
  XOR2_X1    g17414(.A1(new_n17667_), .A2(\a[29] ), .Z(new_n17672_));
  NOR2_X1    g17415(.A1(new_n17672_), .A2(new_n17516_), .ZN(new_n17673_));
  NOR2_X1    g17416(.A1(new_n17673_), .A2(new_n17671_), .ZN(new_n17674_));
  NOR2_X1    g17417(.A1(new_n17664_), .A2(new_n17674_), .ZN(new_n17675_));
  INV_X1     g17418(.I(new_n17664_), .ZN(new_n17676_));
  INV_X1     g17419(.I(new_n17674_), .ZN(new_n17677_));
  NOR2_X1    g17420(.A1(new_n17676_), .A2(new_n17677_), .ZN(new_n17678_));
  NOR2_X1    g17421(.A1(new_n17678_), .A2(new_n17675_), .ZN(new_n17679_));
  NOR2_X1    g17422(.A1(new_n17679_), .A2(new_n17659_), .ZN(new_n17680_));
  XOR2_X1    g17423(.A1(new_n17664_), .A2(new_n17674_), .Z(new_n17681_));
  AOI21_X1   g17424(.A1(new_n17659_), .A2(new_n17681_), .B(new_n17680_), .ZN(new_n17682_));
  OAI22_X1   g17425(.A1(new_n3247_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n3097_), .ZN(new_n17683_));
  NAND2_X1   g17426(.A1(new_n8628_), .A2(\b[34] ), .ZN(new_n17684_));
  AOI21_X1   g17427(.A1(new_n17684_), .A2(new_n17683_), .B(new_n7354_), .ZN(new_n17685_));
  NAND2_X1   g17428(.A1(new_n3246_), .A2(new_n17685_), .ZN(new_n17686_));
  XOR2_X1    g17429(.A1(new_n17686_), .A2(\a[59] ), .Z(new_n17687_));
  XNOR2_X1   g17430(.A1(new_n17682_), .A2(new_n17687_), .ZN(new_n17688_));
  NOR2_X1    g17431(.A1(new_n17688_), .A2(new_n17658_), .ZN(new_n17689_));
  INV_X1     g17432(.I(new_n17658_), .ZN(new_n17690_));
  NOR2_X1    g17433(.A1(new_n17682_), .A2(new_n17687_), .ZN(new_n17691_));
  INV_X1     g17434(.I(new_n17691_), .ZN(new_n17692_));
  NAND2_X1   g17435(.A1(new_n17682_), .A2(new_n17687_), .ZN(new_n17693_));
  AOI21_X1   g17436(.A1(new_n17692_), .A2(new_n17693_), .B(new_n17690_), .ZN(new_n17694_));
  NOR2_X1    g17437(.A1(new_n17689_), .A2(new_n17694_), .ZN(new_n17695_));
  OAI22_X1   g17438(.A1(new_n6721_), .A2(new_n3566_), .B1(new_n6723_), .B2(new_n3696_), .ZN(new_n17696_));
  NAND2_X1   g17439(.A1(new_n7617_), .A2(\b[37] ), .ZN(new_n17697_));
  AOI21_X1   g17440(.A1(new_n17697_), .A2(new_n17696_), .B(new_n6731_), .ZN(new_n17698_));
  NAND2_X1   g17441(.A1(new_n3700_), .A2(new_n17698_), .ZN(new_n17699_));
  XOR2_X1    g17442(.A1(new_n17699_), .A2(\a[56] ), .Z(new_n17700_));
  XOR2_X1    g17443(.A1(new_n17695_), .A2(new_n17700_), .Z(new_n17701_));
  NOR3_X1    g17444(.A1(new_n17689_), .A2(new_n17694_), .A3(new_n17700_), .ZN(new_n17702_));
  INV_X1     g17445(.I(new_n17700_), .ZN(new_n17703_));
  NOR2_X1    g17446(.A1(new_n17695_), .A2(new_n17703_), .ZN(new_n17704_));
  OAI21_X1   g17447(.A1(new_n17704_), .A2(new_n17702_), .B(new_n17657_), .ZN(new_n17705_));
  OAI21_X1   g17448(.A1(new_n17657_), .A2(new_n17701_), .B(new_n17705_), .ZN(new_n17706_));
  OAI22_X1   g17449(.A1(new_n5786_), .A2(new_n4018_), .B1(new_n3997_), .B2(new_n5792_), .ZN(new_n17707_));
  NAND2_X1   g17450(.A1(new_n6745_), .A2(\b[40] ), .ZN(new_n17708_));
  AOI21_X1   g17451(.A1(new_n17708_), .A2(new_n17707_), .B(new_n5796_), .ZN(new_n17709_));
  NAND2_X1   g17452(.A1(new_n4017_), .A2(new_n17709_), .ZN(new_n17710_));
  XOR2_X1    g17453(.A1(new_n17710_), .A2(\a[53] ), .Z(new_n17711_));
  NOR2_X1    g17454(.A1(new_n17706_), .A2(new_n17711_), .ZN(new_n17712_));
  INV_X1     g17455(.I(new_n17712_), .ZN(new_n17713_));
  NAND2_X1   g17456(.A1(new_n17706_), .A2(new_n17711_), .ZN(new_n17714_));
  AOI21_X1   g17457(.A1(new_n17713_), .A2(new_n17714_), .B(new_n17655_), .ZN(new_n17715_));
  INV_X1     g17458(.I(new_n17655_), .ZN(new_n17716_));
  XNOR2_X1   g17459(.A1(new_n17706_), .A2(new_n17711_), .ZN(new_n17717_));
  NOR2_X1    g17460(.A1(new_n17717_), .A2(new_n17716_), .ZN(new_n17718_));
  NOR2_X1    g17461(.A1(new_n17718_), .A2(new_n17715_), .ZN(new_n17719_));
  OAI22_X1   g17462(.A1(new_n5228_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n5225_), .ZN(new_n17720_));
  NAND2_X1   g17463(.A1(new_n5387_), .A2(\b[43] ), .ZN(new_n17721_));
  AOI21_X1   g17464(.A1(new_n17720_), .A2(new_n17721_), .B(new_n5231_), .ZN(new_n17722_));
  NAND2_X1   g17465(.A1(new_n4513_), .A2(new_n17722_), .ZN(new_n17723_));
  XOR2_X1    g17466(.A1(new_n17723_), .A2(\a[50] ), .Z(new_n17724_));
  XNOR2_X1   g17467(.A1(new_n17719_), .A2(new_n17724_), .ZN(new_n17725_));
  NOR2_X1    g17468(.A1(new_n17725_), .A2(new_n17653_), .ZN(new_n17726_));
  NOR2_X1    g17469(.A1(new_n17719_), .A2(new_n17724_), .ZN(new_n17727_));
  INV_X1     g17470(.I(new_n17727_), .ZN(new_n17728_));
  NAND2_X1   g17471(.A1(new_n17719_), .A2(new_n17724_), .ZN(new_n17729_));
  AOI21_X1   g17472(.A1(new_n17728_), .A2(new_n17729_), .B(new_n17652_), .ZN(new_n17730_));
  NOR2_X1    g17473(.A1(new_n17726_), .A2(new_n17730_), .ZN(new_n17731_));
  OAI22_X1   g17474(.A1(new_n4711_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n4706_), .ZN(new_n17732_));
  NAND2_X1   g17475(.A1(new_n5814_), .A2(\b[46] ), .ZN(new_n17733_));
  AOI21_X1   g17476(.A1(new_n17732_), .A2(new_n17733_), .B(new_n4714_), .ZN(new_n17734_));
  NAND2_X1   g17477(.A1(new_n5177_), .A2(new_n17734_), .ZN(new_n17735_));
  XOR2_X1    g17478(.A1(new_n17735_), .A2(\a[47] ), .Z(new_n17736_));
  NAND2_X1   g17479(.A1(new_n17576_), .A2(new_n17563_), .ZN(new_n17737_));
  NAND2_X1   g17480(.A1(new_n17737_), .A2(new_n17575_), .ZN(new_n17738_));
  INV_X1     g17481(.I(new_n17738_), .ZN(new_n17739_));
  NOR2_X1    g17482(.A1(new_n17739_), .A2(new_n17736_), .ZN(new_n17740_));
  INV_X1     g17483(.I(new_n17736_), .ZN(new_n17741_));
  NOR2_X1    g17484(.A1(new_n17738_), .A2(new_n17741_), .ZN(new_n17742_));
  NOR2_X1    g17485(.A1(new_n17740_), .A2(new_n17742_), .ZN(new_n17743_));
  NOR2_X1    g17486(.A1(new_n17743_), .A2(new_n17731_), .ZN(new_n17744_));
  XOR2_X1    g17487(.A1(new_n17738_), .A2(new_n17736_), .Z(new_n17745_));
  NOR3_X1    g17488(.A1(new_n17745_), .A2(new_n17726_), .A3(new_n17730_), .ZN(new_n17746_));
  NOR2_X1    g17489(.A1(new_n17744_), .A2(new_n17746_), .ZN(new_n17747_));
  INV_X1     g17490(.I(new_n17747_), .ZN(new_n17748_));
  OAI22_X1   g17491(.A1(new_n4208_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n4203_), .ZN(new_n17749_));
  NAND2_X1   g17492(.A1(new_n5244_), .A2(\b[49] ), .ZN(new_n17750_));
  AOI21_X1   g17493(.A1(new_n17749_), .A2(new_n17750_), .B(new_n4211_), .ZN(new_n17751_));
  NAND2_X1   g17494(.A1(new_n5741_), .A2(new_n17751_), .ZN(new_n17752_));
  XOR2_X1    g17495(.A1(new_n17752_), .A2(\a[44] ), .Z(new_n17753_));
  NOR2_X1    g17496(.A1(new_n17748_), .A2(new_n17753_), .ZN(new_n17754_));
  INV_X1     g17497(.I(new_n17753_), .ZN(new_n17755_));
  NOR2_X1    g17498(.A1(new_n17747_), .A2(new_n17755_), .ZN(new_n17756_));
  NOR2_X1    g17499(.A1(new_n17754_), .A2(new_n17756_), .ZN(new_n17757_));
  NOR2_X1    g17500(.A1(new_n17757_), .A2(new_n17651_), .ZN(new_n17758_));
  INV_X1     g17501(.I(new_n17651_), .ZN(new_n17759_));
  XOR2_X1    g17502(.A1(new_n17747_), .A2(new_n17753_), .Z(new_n17760_));
  NOR2_X1    g17503(.A1(new_n17760_), .A2(new_n17759_), .ZN(new_n17761_));
  NOR2_X1    g17504(.A1(new_n17758_), .A2(new_n17761_), .ZN(new_n17762_));
  OAI22_X1   g17505(.A1(new_n3736_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n3731_), .ZN(new_n17763_));
  NAND2_X1   g17506(.A1(new_n4730_), .A2(\b[52] ), .ZN(new_n17764_));
  AOI21_X1   g17507(.A1(new_n17763_), .A2(new_n17764_), .B(new_n3739_), .ZN(new_n17765_));
  NAND2_X1   g17508(.A1(new_n6237_), .A2(new_n17765_), .ZN(new_n17766_));
  XOR2_X1    g17509(.A1(new_n17766_), .A2(\a[41] ), .Z(new_n17767_));
  XNOR2_X1   g17510(.A1(new_n17762_), .A2(new_n17767_), .ZN(new_n17768_));
  NOR2_X1    g17511(.A1(new_n17768_), .A2(new_n17650_), .ZN(new_n17769_));
  INV_X1     g17512(.I(new_n17650_), .ZN(new_n17770_));
  NOR2_X1    g17513(.A1(new_n17762_), .A2(new_n17767_), .ZN(new_n17771_));
  INV_X1     g17514(.I(new_n17771_), .ZN(new_n17772_));
  NAND2_X1   g17515(.A1(new_n17762_), .A2(new_n17767_), .ZN(new_n17773_));
  AOI21_X1   g17516(.A1(new_n17772_), .A2(new_n17773_), .B(new_n17770_), .ZN(new_n17774_));
  NOR2_X1    g17517(.A1(new_n17769_), .A2(new_n17774_), .ZN(new_n17775_));
  OAI22_X1   g17518(.A1(new_n3298_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n3293_), .ZN(new_n17776_));
  NAND2_X1   g17519(.A1(new_n4227_), .A2(\b[55] ), .ZN(new_n17777_));
  AOI21_X1   g17520(.A1(new_n17776_), .A2(new_n17777_), .B(new_n3301_), .ZN(new_n17778_));
  NAND2_X1   g17521(.A1(new_n7308_), .A2(new_n17778_), .ZN(new_n17779_));
  XOR2_X1    g17522(.A1(new_n17779_), .A2(\a[38] ), .Z(new_n17780_));
  XOR2_X1    g17523(.A1(new_n17775_), .A2(new_n17780_), .Z(new_n17781_));
  INV_X1     g17524(.I(new_n17781_), .ZN(new_n17782_));
  INV_X1     g17525(.I(new_n17775_), .ZN(new_n17783_));
  NOR2_X1    g17526(.A1(new_n17783_), .A2(new_n17780_), .ZN(new_n17784_));
  INV_X1     g17527(.I(new_n17784_), .ZN(new_n17785_));
  NAND2_X1   g17528(.A1(new_n17783_), .A2(new_n17780_), .ZN(new_n17786_));
  AOI21_X1   g17529(.A1(new_n17785_), .A2(new_n17786_), .B(new_n17649_), .ZN(new_n17787_));
  AOI21_X1   g17530(.A1(new_n17649_), .A2(new_n17782_), .B(new_n17787_), .ZN(new_n17788_));
  OAI22_X1   g17531(.A1(new_n2846_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n2841_), .ZN(new_n17789_));
  NAND2_X1   g17532(.A1(new_n3755_), .A2(\b[58] ), .ZN(new_n17790_));
  AOI21_X1   g17533(.A1(new_n17789_), .A2(new_n17790_), .B(new_n2849_), .ZN(new_n17791_));
  NAND2_X1   g17534(.A1(new_n7929_), .A2(new_n17791_), .ZN(new_n17792_));
  XOR2_X1    g17535(.A1(new_n17792_), .A2(\a[35] ), .Z(new_n17793_));
  NAND2_X1   g17536(.A1(new_n17622_), .A2(new_n17609_), .ZN(new_n17794_));
  NAND2_X1   g17537(.A1(new_n17794_), .A2(new_n17621_), .ZN(new_n17795_));
  INV_X1     g17538(.I(new_n17795_), .ZN(new_n17796_));
  NOR2_X1    g17539(.A1(new_n17796_), .A2(new_n17793_), .ZN(new_n17797_));
  INV_X1     g17540(.I(new_n17793_), .ZN(new_n17798_));
  NOR2_X1    g17541(.A1(new_n17795_), .A2(new_n17798_), .ZN(new_n17799_));
  NOR2_X1    g17542(.A1(new_n17797_), .A2(new_n17799_), .ZN(new_n17800_));
  NOR2_X1    g17543(.A1(new_n17800_), .A2(new_n17788_), .ZN(new_n17801_));
  XOR2_X1    g17544(.A1(new_n17795_), .A2(new_n17793_), .Z(new_n17802_));
  INV_X1     g17545(.I(new_n17802_), .ZN(new_n17803_));
  AOI21_X1   g17546(.A1(new_n17788_), .A2(new_n17803_), .B(new_n17801_), .ZN(new_n17804_));
  XOR2_X1    g17547(.A1(new_n17804_), .A2(new_n17648_), .Z(new_n17805_));
  INV_X1     g17548(.I(new_n17648_), .ZN(new_n17806_));
  NOR2_X1    g17549(.A1(new_n17804_), .A2(new_n17806_), .ZN(new_n17807_));
  NAND2_X1   g17550(.A1(new_n17804_), .A2(new_n17806_), .ZN(new_n17808_));
  INV_X1     g17551(.I(new_n17808_), .ZN(new_n17809_));
  OAI21_X1   g17552(.A1(new_n17809_), .A2(new_n17807_), .B(new_n17643_), .ZN(new_n17810_));
  OAI21_X1   g17553(.A1(new_n17643_), .A2(new_n17805_), .B(new_n17810_), .ZN(new_n17811_));
  XNOR2_X1   g17554(.A1(new_n17642_), .A2(new_n17811_), .ZN(new_n17812_));
  NOR2_X1    g17555(.A1(new_n17636_), .A2(new_n17461_), .ZN(new_n17813_));
  AOI21_X1   g17556(.A1(new_n17458_), .A2(new_n17637_), .B(new_n17813_), .ZN(new_n17814_));
  XNOR2_X1   g17557(.A1(new_n17814_), .A2(new_n17812_), .ZN(\f[93] ));
  NOR2_X1    g17558(.A1(new_n2602_), .A2(new_n8932_), .ZN(new_n17816_));
  NOR2_X1    g17559(.A1(new_n2447_), .A2(new_n8956_), .ZN(new_n17817_));
  NOR4_X1    g17560(.A1(new_n9323_), .A2(new_n2455_), .A3(new_n17816_), .A4(new_n17817_), .ZN(new_n17818_));
  XOR2_X1    g17561(.A1(new_n17818_), .A2(new_n2442_), .Z(new_n17819_));
  INV_X1     g17562(.I(new_n17799_), .ZN(new_n17820_));
  AOI21_X1   g17563(.A1(new_n17788_), .A2(new_n17820_), .B(new_n17797_), .ZN(new_n17821_));
  INV_X1     g17564(.I(new_n17821_), .ZN(new_n17822_));
  OAI22_X1   g17565(.A1(new_n3298_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n3293_), .ZN(new_n17823_));
  NAND2_X1   g17566(.A1(new_n4227_), .A2(\b[56] ), .ZN(new_n17824_));
  AOI21_X1   g17567(.A1(new_n17823_), .A2(new_n17824_), .B(new_n3301_), .ZN(new_n17825_));
  NAND2_X1   g17568(.A1(new_n7559_), .A2(new_n17825_), .ZN(new_n17826_));
  XOR2_X1    g17569(.A1(new_n17826_), .A2(\a[38] ), .Z(new_n17827_));
  AOI21_X1   g17570(.A1(new_n17770_), .A2(new_n17773_), .B(new_n17771_), .ZN(new_n17828_));
  INV_X1     g17571(.I(new_n17828_), .ZN(new_n17829_));
  INV_X1     g17572(.I(new_n17756_), .ZN(new_n17830_));
  AOI21_X1   g17573(.A1(new_n17759_), .A2(new_n17830_), .B(new_n17754_), .ZN(new_n17831_));
  OAI22_X1   g17574(.A1(new_n4208_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n4203_), .ZN(new_n17832_));
  NAND2_X1   g17575(.A1(new_n5244_), .A2(\b[50] ), .ZN(new_n17833_));
  AOI21_X1   g17576(.A1(new_n17832_), .A2(new_n17833_), .B(new_n4211_), .ZN(new_n17834_));
  NAND2_X1   g17577(.A1(new_n5954_), .A2(new_n17834_), .ZN(new_n17835_));
  XOR2_X1    g17578(.A1(new_n17835_), .A2(\a[44] ), .Z(new_n17836_));
  OAI22_X1   g17579(.A1(new_n5228_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n5225_), .ZN(new_n17837_));
  NAND2_X1   g17580(.A1(new_n5387_), .A2(\b[44] ), .ZN(new_n17838_));
  AOI21_X1   g17581(.A1(new_n17837_), .A2(new_n17838_), .B(new_n5231_), .ZN(new_n17839_));
  NAND2_X1   g17582(.A1(new_n4833_), .A2(new_n17839_), .ZN(new_n17840_));
  XOR2_X1    g17583(.A1(new_n17840_), .A2(\a[50] ), .Z(new_n17841_));
  NOR2_X1    g17584(.A1(new_n17704_), .A2(new_n17657_), .ZN(new_n17842_));
  NOR2_X1    g17585(.A1(new_n17842_), .A2(new_n17702_), .ZN(new_n17843_));
  OAI22_X1   g17586(.A1(new_n6721_), .A2(new_n3696_), .B1(new_n6723_), .B2(new_n3845_), .ZN(new_n17844_));
  NAND2_X1   g17587(.A1(new_n7617_), .A2(\b[38] ), .ZN(new_n17845_));
  AOI21_X1   g17588(.A1(new_n17845_), .A2(new_n17844_), .B(new_n6731_), .ZN(new_n17846_));
  NAND2_X1   g17589(.A1(new_n3844_), .A2(new_n17846_), .ZN(new_n17847_));
  XOR2_X1    g17590(.A1(new_n17847_), .A2(\a[56] ), .Z(new_n17848_));
  NAND2_X1   g17591(.A1(new_n17693_), .A2(new_n17690_), .ZN(new_n17849_));
  NAND2_X1   g17592(.A1(new_n17849_), .A2(new_n17692_), .ZN(new_n17850_));
  OAI22_X1   g17593(.A1(new_n3408_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n3247_), .ZN(new_n17851_));
  NAND2_X1   g17594(.A1(new_n8628_), .A2(\b[35] ), .ZN(new_n17852_));
  AOI21_X1   g17595(.A1(new_n17852_), .A2(new_n17851_), .B(new_n7354_), .ZN(new_n17853_));
  NAND2_X1   g17596(.A1(new_n3411_), .A2(new_n17853_), .ZN(new_n17854_));
  XOR2_X1    g17597(.A1(new_n17854_), .A2(\a[59] ), .Z(new_n17855_));
  INV_X1     g17598(.I(new_n17675_), .ZN(new_n17856_));
  OAI21_X1   g17599(.A1(new_n17659_), .A2(new_n17678_), .B(new_n17856_), .ZN(new_n17857_));
  OAI22_X1   g17600(.A1(new_n2964_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2794_), .ZN(new_n17858_));
  NAND2_X1   g17601(.A1(new_n9644_), .A2(\b[32] ), .ZN(new_n17859_));
  AOI21_X1   g17602(.A1(new_n17859_), .A2(new_n17858_), .B(new_n8321_), .ZN(new_n17860_));
  NAND2_X1   g17603(.A1(new_n2963_), .A2(new_n17860_), .ZN(new_n17861_));
  XOR2_X1    g17604(.A1(new_n17861_), .A2(new_n8309_), .Z(new_n17862_));
  NAND2_X1   g17605(.A1(new_n17670_), .A2(new_n17516_), .ZN(new_n17863_));
  NAND2_X1   g17606(.A1(new_n17863_), .A2(new_n17669_), .ZN(new_n17864_));
  NOR3_X1    g17607(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n2405_), .ZN(new_n17865_));
  NOR2_X1    g17608(.A1(new_n9364_), .A2(new_n2405_), .ZN(new_n17866_));
  NOR3_X1    g17609(.A1(new_n17866_), .A2(new_n2543_), .A3(new_n8985_), .ZN(new_n17867_));
  NOR2_X1    g17610(.A1(new_n17867_), .A2(new_n17865_), .ZN(new_n17868_));
  INV_X1     g17611(.I(new_n17868_), .ZN(new_n17869_));
  XOR2_X1    g17612(.A1(new_n17864_), .A2(new_n17869_), .Z(new_n17870_));
  INV_X1     g17613(.I(new_n17870_), .ZN(new_n17871_));
  NOR2_X1    g17614(.A1(new_n17864_), .A2(new_n17868_), .ZN(new_n17872_));
  INV_X1     g17615(.I(new_n17872_), .ZN(new_n17873_));
  NAND2_X1   g17616(.A1(new_n17864_), .A2(new_n17868_), .ZN(new_n17874_));
  AOI21_X1   g17617(.A1(new_n17873_), .A2(new_n17874_), .B(new_n17862_), .ZN(new_n17875_));
  AOI21_X1   g17618(.A1(new_n17862_), .A2(new_n17871_), .B(new_n17875_), .ZN(new_n17876_));
  XNOR2_X1   g17619(.A1(new_n17857_), .A2(new_n17876_), .ZN(new_n17877_));
  NOR2_X1    g17620(.A1(new_n17877_), .A2(new_n17855_), .ZN(new_n17878_));
  NOR2_X1    g17621(.A1(new_n17857_), .A2(new_n17876_), .ZN(new_n17879_));
  INV_X1     g17622(.I(new_n17879_), .ZN(new_n17880_));
  NAND2_X1   g17623(.A1(new_n17857_), .A2(new_n17876_), .ZN(new_n17881_));
  NAND2_X1   g17624(.A1(new_n17880_), .A2(new_n17881_), .ZN(new_n17882_));
  AOI21_X1   g17625(.A1(new_n17855_), .A2(new_n17882_), .B(new_n17878_), .ZN(new_n17883_));
  XNOR2_X1   g17626(.A1(new_n17883_), .A2(new_n17850_), .ZN(new_n17884_));
  NOR2_X1    g17627(.A1(new_n17883_), .A2(new_n17850_), .ZN(new_n17885_));
  NAND2_X1   g17628(.A1(new_n17883_), .A2(new_n17850_), .ZN(new_n17886_));
  INV_X1     g17629(.I(new_n17886_), .ZN(new_n17887_));
  OAI21_X1   g17630(.A1(new_n17887_), .A2(new_n17885_), .B(new_n17848_), .ZN(new_n17888_));
  OAI21_X1   g17631(.A1(new_n17848_), .A2(new_n17884_), .B(new_n17888_), .ZN(new_n17889_));
  OAI22_X1   g17632(.A1(new_n5786_), .A2(new_n4316_), .B1(new_n4018_), .B2(new_n5792_), .ZN(new_n17890_));
  NAND2_X1   g17633(.A1(new_n6745_), .A2(\b[41] ), .ZN(new_n17891_));
  AOI21_X1   g17634(.A1(new_n17891_), .A2(new_n17890_), .B(new_n5796_), .ZN(new_n17892_));
  NAND2_X1   g17635(.A1(new_n4320_), .A2(new_n17892_), .ZN(new_n17893_));
  XOR2_X1    g17636(.A1(new_n17893_), .A2(\a[53] ), .Z(new_n17894_));
  NOR2_X1    g17637(.A1(new_n17889_), .A2(new_n17894_), .ZN(new_n17895_));
  INV_X1     g17638(.I(new_n17895_), .ZN(new_n17896_));
  NAND2_X1   g17639(.A1(new_n17889_), .A2(new_n17894_), .ZN(new_n17897_));
  AOI21_X1   g17640(.A1(new_n17896_), .A2(new_n17897_), .B(new_n17843_), .ZN(new_n17898_));
  INV_X1     g17641(.I(new_n17843_), .ZN(new_n17899_));
  XNOR2_X1   g17642(.A1(new_n17889_), .A2(new_n17894_), .ZN(new_n17900_));
  NOR2_X1    g17643(.A1(new_n17900_), .A2(new_n17899_), .ZN(new_n17901_));
  NOR2_X1    g17644(.A1(new_n17901_), .A2(new_n17898_), .ZN(new_n17902_));
  AOI21_X1   g17645(.A1(new_n17716_), .A2(new_n17714_), .B(new_n17712_), .ZN(new_n17903_));
  NOR2_X1    g17646(.A1(new_n17902_), .A2(new_n17903_), .ZN(new_n17904_));
  INV_X1     g17647(.I(new_n17904_), .ZN(new_n17905_));
  NAND2_X1   g17648(.A1(new_n17902_), .A2(new_n17903_), .ZN(new_n17906_));
  AOI21_X1   g17649(.A1(new_n17905_), .A2(new_n17906_), .B(new_n17841_), .ZN(new_n17907_));
  INV_X1     g17650(.I(new_n17841_), .ZN(new_n17908_));
  XNOR2_X1   g17651(.A1(new_n17902_), .A2(new_n17903_), .ZN(new_n17909_));
  NOR2_X1    g17652(.A1(new_n17909_), .A2(new_n17908_), .ZN(new_n17910_));
  NOR2_X1    g17653(.A1(new_n17910_), .A2(new_n17907_), .ZN(new_n17911_));
  NAND2_X1   g17654(.A1(new_n17729_), .A2(new_n17652_), .ZN(new_n17912_));
  NAND2_X1   g17655(.A1(new_n17912_), .A2(new_n17728_), .ZN(new_n17913_));
  INV_X1     g17656(.I(new_n17913_), .ZN(new_n17914_));
  OAI22_X1   g17657(.A1(new_n4711_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n4706_), .ZN(new_n17915_));
  NAND2_X1   g17658(.A1(new_n5814_), .A2(\b[47] ), .ZN(new_n17916_));
  AOI21_X1   g17659(.A1(new_n17915_), .A2(new_n17916_), .B(new_n4714_), .ZN(new_n17917_));
  NAND2_X1   g17660(.A1(new_n5196_), .A2(new_n17917_), .ZN(new_n17918_));
  XOR2_X1    g17661(.A1(new_n17918_), .A2(\a[47] ), .Z(new_n17919_));
  NOR2_X1    g17662(.A1(new_n17914_), .A2(new_n17919_), .ZN(new_n17920_));
  INV_X1     g17663(.I(new_n17919_), .ZN(new_n17921_));
  NOR2_X1    g17664(.A1(new_n17913_), .A2(new_n17921_), .ZN(new_n17922_));
  NOR2_X1    g17665(.A1(new_n17920_), .A2(new_n17922_), .ZN(new_n17923_));
  NOR2_X1    g17666(.A1(new_n17923_), .A2(new_n17911_), .ZN(new_n17924_));
  INV_X1     g17667(.I(new_n17911_), .ZN(new_n17925_));
  XOR2_X1    g17668(.A1(new_n17913_), .A2(new_n17919_), .Z(new_n17926_));
  NOR2_X1    g17669(.A1(new_n17926_), .A2(new_n17925_), .ZN(new_n17927_));
  NOR2_X1    g17670(.A1(new_n17924_), .A2(new_n17927_), .ZN(new_n17928_));
  INV_X1     g17671(.I(new_n17742_), .ZN(new_n17929_));
  AOI21_X1   g17672(.A1(new_n17731_), .A2(new_n17929_), .B(new_n17740_), .ZN(new_n17930_));
  NOR2_X1    g17673(.A1(new_n17930_), .A2(new_n17928_), .ZN(new_n17931_));
  AND2_X2    g17674(.A1(new_n17930_), .A2(new_n17928_), .Z(new_n17932_));
  NOR2_X1    g17675(.A1(new_n17932_), .A2(new_n17931_), .ZN(new_n17933_));
  NOR2_X1    g17676(.A1(new_n17933_), .A2(new_n17836_), .ZN(new_n17934_));
  INV_X1     g17677(.I(new_n17836_), .ZN(new_n17935_));
  XNOR2_X1   g17678(.A1(new_n17930_), .A2(new_n17928_), .ZN(new_n17936_));
  NOR2_X1    g17679(.A1(new_n17936_), .A2(new_n17935_), .ZN(new_n17937_));
  NOR2_X1    g17680(.A1(new_n17934_), .A2(new_n17937_), .ZN(new_n17938_));
  OAI22_X1   g17681(.A1(new_n3736_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n3731_), .ZN(new_n17939_));
  NAND2_X1   g17682(.A1(new_n4730_), .A2(\b[53] ), .ZN(new_n17940_));
  AOI21_X1   g17683(.A1(new_n17939_), .A2(new_n17940_), .B(new_n3739_), .ZN(new_n17941_));
  NAND2_X1   g17684(.A1(new_n6471_), .A2(new_n17941_), .ZN(new_n17942_));
  XOR2_X1    g17685(.A1(new_n17942_), .A2(\a[41] ), .Z(new_n17943_));
  XNOR2_X1   g17686(.A1(new_n17938_), .A2(new_n17943_), .ZN(new_n17944_));
  NOR2_X1    g17687(.A1(new_n17944_), .A2(new_n17831_), .ZN(new_n17945_));
  INV_X1     g17688(.I(new_n17831_), .ZN(new_n17946_));
  NOR2_X1    g17689(.A1(new_n17938_), .A2(new_n17943_), .ZN(new_n17947_));
  INV_X1     g17690(.I(new_n17947_), .ZN(new_n17948_));
  NAND2_X1   g17691(.A1(new_n17938_), .A2(new_n17943_), .ZN(new_n17949_));
  AOI21_X1   g17692(.A1(new_n17948_), .A2(new_n17949_), .B(new_n17946_), .ZN(new_n17950_));
  NOR2_X1    g17693(.A1(new_n17945_), .A2(new_n17950_), .ZN(new_n17951_));
  NOR2_X1    g17694(.A1(new_n17829_), .A2(new_n17951_), .ZN(new_n17952_));
  INV_X1     g17695(.I(new_n17951_), .ZN(new_n17953_));
  NOR2_X1    g17696(.A1(new_n17953_), .A2(new_n17828_), .ZN(new_n17954_));
  NOR2_X1    g17697(.A1(new_n17954_), .A2(new_n17952_), .ZN(new_n17955_));
  NOR2_X1    g17698(.A1(new_n17955_), .A2(new_n17827_), .ZN(new_n17956_));
  INV_X1     g17699(.I(new_n17827_), .ZN(new_n17957_));
  XOR2_X1    g17700(.A1(new_n17951_), .A2(new_n17828_), .Z(new_n17958_));
  NOR2_X1    g17701(.A1(new_n17958_), .A2(new_n17957_), .ZN(new_n17959_));
  NOR2_X1    g17702(.A1(new_n17956_), .A2(new_n17959_), .ZN(new_n17960_));
  AOI21_X1   g17703(.A1(new_n17649_), .A2(new_n17786_), .B(new_n17784_), .ZN(new_n17961_));
  OAI22_X1   g17704(.A1(new_n2846_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n2841_), .ZN(new_n17962_));
  NAND2_X1   g17705(.A1(new_n3755_), .A2(\b[59] ), .ZN(new_n17963_));
  AOI21_X1   g17706(.A1(new_n17962_), .A2(new_n17963_), .B(new_n2849_), .ZN(new_n17964_));
  NAND2_X1   g17707(.A1(new_n8550_), .A2(new_n17964_), .ZN(new_n17965_));
  XOR2_X1    g17708(.A1(new_n17965_), .A2(\a[35] ), .Z(new_n17966_));
  XNOR2_X1   g17709(.A1(new_n17961_), .A2(new_n17966_), .ZN(new_n17967_));
  NOR2_X1    g17710(.A1(new_n17967_), .A2(new_n17960_), .ZN(new_n17968_));
  INV_X1     g17711(.I(new_n17960_), .ZN(new_n17969_));
  NOR2_X1    g17712(.A1(new_n17961_), .A2(new_n17966_), .ZN(new_n17970_));
  INV_X1     g17713(.I(new_n17970_), .ZN(new_n17971_));
  NAND2_X1   g17714(.A1(new_n17961_), .A2(new_n17966_), .ZN(new_n17972_));
  AOI21_X1   g17715(.A1(new_n17971_), .A2(new_n17972_), .B(new_n17969_), .ZN(new_n17973_));
  NOR2_X1    g17716(.A1(new_n17968_), .A2(new_n17973_), .ZN(new_n17974_));
  NOR2_X1    g17717(.A1(new_n17974_), .A2(new_n17822_), .ZN(new_n17975_));
  INV_X1     g17718(.I(new_n17974_), .ZN(new_n17976_));
  NOR2_X1    g17719(.A1(new_n17976_), .A2(new_n17821_), .ZN(new_n17977_));
  NOR2_X1    g17720(.A1(new_n17977_), .A2(new_n17975_), .ZN(new_n17978_));
  NOR2_X1    g17721(.A1(new_n17978_), .A2(new_n17819_), .ZN(new_n17979_));
  INV_X1     g17722(.I(new_n17819_), .ZN(new_n17980_));
  XOR2_X1    g17723(.A1(new_n17974_), .A2(new_n17821_), .Z(new_n17981_));
  NOR2_X1    g17724(.A1(new_n17981_), .A2(new_n17980_), .ZN(new_n17982_));
  NOR2_X1    g17725(.A1(new_n17979_), .A2(new_n17982_), .ZN(new_n17983_));
  OAI21_X1   g17726(.A1(new_n17643_), .A2(new_n17807_), .B(new_n17808_), .ZN(new_n17984_));
  INV_X1     g17727(.I(new_n17813_), .ZN(new_n17985_));
  INV_X1     g17728(.I(new_n17447_), .ZN(new_n17986_));
  OAI21_X1   g17729(.A1(new_n17257_), .A2(new_n17986_), .B(new_n17457_), .ZN(new_n17987_));
  NAND3_X1   g17730(.A1(new_n17987_), .A2(new_n17454_), .A3(new_n17637_), .ZN(new_n17988_));
  NAND3_X1   g17731(.A1(new_n17988_), .A2(new_n17985_), .A3(new_n17812_), .ZN(new_n17989_));
  NAND2_X1   g17732(.A1(new_n17642_), .A2(new_n17811_), .ZN(new_n17990_));
  NAND2_X1   g17733(.A1(new_n17989_), .A2(new_n17990_), .ZN(new_n17991_));
  XNOR2_X1   g17734(.A1(new_n17991_), .A2(new_n17984_), .ZN(new_n17992_));
  XOR2_X1    g17735(.A1(new_n17992_), .A2(new_n17983_), .Z(\f[94] ));
  NOR2_X1    g17736(.A1(new_n17983_), .A2(new_n17984_), .ZN(new_n17994_));
  INV_X1     g17737(.I(new_n17994_), .ZN(new_n17995_));
  XOR2_X1    g17738(.A1(new_n17983_), .A2(new_n17984_), .Z(new_n17996_));
  AOI21_X1   g17739(.A1(new_n17642_), .A2(new_n17811_), .B(new_n17996_), .ZN(new_n17997_));
  NAND2_X1   g17740(.A1(new_n17989_), .A2(new_n17997_), .ZN(new_n17998_));
  NAND2_X1   g17741(.A1(new_n17998_), .A2(new_n17995_), .ZN(new_n17999_));
  NOR2_X1    g17742(.A1(new_n17975_), .A2(new_n17819_), .ZN(new_n18000_));
  NOR2_X1    g17743(.A1(new_n18000_), .A2(new_n17977_), .ZN(new_n18001_));
  AOI21_X1   g17744(.A1(new_n17969_), .A2(new_n17972_), .B(new_n17970_), .ZN(new_n18002_));
  OAI22_X1   g17745(.A1(new_n9595_), .A2(new_n2455_), .B1(new_n8956_), .B2(new_n2602_), .ZN(new_n18003_));
  OAI22_X1   g17746(.A1(new_n2846_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n2841_), .ZN(new_n18004_));
  NAND2_X1   g17747(.A1(new_n3755_), .A2(\b[60] ), .ZN(new_n18005_));
  AOI21_X1   g17748(.A1(new_n18004_), .A2(new_n18005_), .B(new_n2849_), .ZN(new_n18006_));
  NAND2_X1   g17749(.A1(new_n8935_), .A2(new_n18006_), .ZN(new_n18007_));
  XOR2_X1    g17750(.A1(new_n18007_), .A2(\a[35] ), .Z(new_n18008_));
  OAI22_X1   g17751(.A1(new_n3736_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n3731_), .ZN(new_n18009_));
  NAND2_X1   g17752(.A1(new_n4730_), .A2(\b[54] ), .ZN(new_n18010_));
  AOI21_X1   g17753(.A1(new_n18009_), .A2(new_n18010_), .B(new_n3739_), .ZN(new_n18011_));
  NAND2_X1   g17754(.A1(new_n6994_), .A2(new_n18011_), .ZN(new_n18012_));
  XOR2_X1    g17755(.A1(new_n18012_), .A2(\a[41] ), .Z(new_n18013_));
  INV_X1     g17756(.I(new_n17932_), .ZN(new_n18014_));
  AOI21_X1   g17757(.A1(new_n18014_), .A2(new_n17935_), .B(new_n17931_), .ZN(new_n18015_));
  OAI22_X1   g17758(.A1(new_n4208_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n4203_), .ZN(new_n18016_));
  NAND2_X1   g17759(.A1(new_n5244_), .A2(\b[51] ), .ZN(new_n18017_));
  AOI21_X1   g17760(.A1(new_n18016_), .A2(new_n18017_), .B(new_n4211_), .ZN(new_n18018_));
  NAND2_X1   g17761(.A1(new_n6219_), .A2(new_n18018_), .ZN(new_n18019_));
  XOR2_X1    g17762(.A1(new_n18019_), .A2(\a[44] ), .Z(new_n18020_));
  OAI22_X1   g17763(.A1(new_n4711_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n4706_), .ZN(new_n18021_));
  NAND2_X1   g17764(.A1(new_n5814_), .A2(\b[48] ), .ZN(new_n18022_));
  AOI21_X1   g17765(.A1(new_n18021_), .A2(new_n18022_), .B(new_n4714_), .ZN(new_n18023_));
  NAND2_X1   g17766(.A1(new_n5537_), .A2(new_n18023_), .ZN(new_n18024_));
  XOR2_X1    g17767(.A1(new_n18024_), .A2(\a[47] ), .Z(new_n18025_));
  OAI22_X1   g17768(.A1(new_n5786_), .A2(new_n4501_), .B1(new_n4316_), .B2(new_n5792_), .ZN(new_n18026_));
  NAND2_X1   g17769(.A1(new_n6745_), .A2(\b[42] ), .ZN(new_n18027_));
  AOI21_X1   g17770(.A1(new_n18027_), .A2(new_n18026_), .B(new_n5796_), .ZN(new_n18028_));
  NAND2_X1   g17771(.A1(new_n4500_), .A2(new_n18028_), .ZN(new_n18029_));
  XOR2_X1    g17772(.A1(new_n18029_), .A2(\a[53] ), .Z(new_n18030_));
  OAI21_X1   g17773(.A1(new_n17848_), .A2(new_n17885_), .B(new_n17886_), .ZN(new_n18031_));
  OAI22_X1   g17774(.A1(new_n6721_), .A2(new_n3845_), .B1(new_n6723_), .B2(new_n3997_), .ZN(new_n18032_));
  NAND2_X1   g17775(.A1(new_n7617_), .A2(\b[39] ), .ZN(new_n18033_));
  AOI21_X1   g17776(.A1(new_n18033_), .A2(new_n18032_), .B(new_n6731_), .ZN(new_n18034_));
  NAND2_X1   g17777(.A1(new_n3996_), .A2(new_n18034_), .ZN(new_n18035_));
  XOR2_X1    g17778(.A1(new_n18035_), .A2(\a[56] ), .Z(new_n18036_));
  NAND2_X1   g17779(.A1(new_n17862_), .A2(new_n17873_), .ZN(new_n18037_));
  NAND2_X1   g17780(.A1(new_n18037_), .A2(new_n17874_), .ZN(new_n18038_));
  NOR3_X1    g17781(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n2543_), .ZN(new_n18039_));
  NOR2_X1    g17782(.A1(new_n9364_), .A2(new_n2543_), .ZN(new_n18040_));
  NOR3_X1    g17783(.A1(new_n18040_), .A2(new_n2660_), .A3(new_n8985_), .ZN(new_n18041_));
  NOR2_X1    g17784(.A1(new_n18041_), .A2(new_n18039_), .ZN(new_n18042_));
  NOR2_X1    g17785(.A1(new_n17869_), .A2(new_n18042_), .ZN(new_n18043_));
  INV_X1     g17786(.I(new_n18042_), .ZN(new_n18044_));
  NOR2_X1    g17787(.A1(new_n18044_), .A2(new_n17868_), .ZN(new_n18045_));
  NOR2_X1    g17788(.A1(new_n18043_), .A2(new_n18045_), .ZN(new_n18046_));
  INV_X1     g17789(.I(new_n18046_), .ZN(new_n18047_));
  XOR2_X1    g17790(.A1(new_n17868_), .A2(new_n18042_), .Z(new_n18048_));
  NOR2_X1    g17791(.A1(new_n18038_), .A2(new_n18048_), .ZN(new_n18049_));
  AOI21_X1   g17792(.A1(new_n18038_), .A2(new_n18047_), .B(new_n18049_), .ZN(new_n18050_));
  INV_X1     g17793(.I(new_n18050_), .ZN(new_n18051_));
  OAI22_X1   g17794(.A1(new_n3566_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n3408_), .ZN(new_n18052_));
  NAND2_X1   g17795(.A1(new_n8628_), .A2(\b[36] ), .ZN(new_n18053_));
  AOI21_X1   g17796(.A1(new_n18053_), .A2(new_n18052_), .B(new_n7354_), .ZN(new_n18054_));
  NAND2_X1   g17797(.A1(new_n3565_), .A2(new_n18054_), .ZN(new_n18055_));
  XOR2_X1    g17798(.A1(new_n18055_), .A2(\a[59] ), .Z(new_n18056_));
  OAI22_X1   g17799(.A1(new_n3097_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n2964_), .ZN(new_n18057_));
  NAND2_X1   g17800(.A1(new_n9644_), .A2(\b[33] ), .ZN(new_n18058_));
  AOI21_X1   g17801(.A1(new_n18058_), .A2(new_n18057_), .B(new_n8321_), .ZN(new_n18059_));
  NAND2_X1   g17802(.A1(new_n3101_), .A2(new_n18059_), .ZN(new_n18060_));
  XOR2_X1    g17803(.A1(new_n18060_), .A2(\a[62] ), .Z(new_n18061_));
  NOR2_X1    g17804(.A1(new_n18056_), .A2(new_n18061_), .ZN(new_n18062_));
  AND2_X2    g17805(.A1(new_n18056_), .A2(new_n18061_), .Z(new_n18063_));
  OAI21_X1   g17806(.A1(new_n18063_), .A2(new_n18062_), .B(new_n18051_), .ZN(new_n18064_));
  XOR2_X1    g17807(.A1(new_n18056_), .A2(new_n18061_), .Z(new_n18065_));
  NAND2_X1   g17808(.A1(new_n18065_), .A2(new_n18050_), .ZN(new_n18066_));
  NAND2_X1   g17809(.A1(new_n18066_), .A2(new_n18064_), .ZN(new_n18067_));
  OAI21_X1   g17810(.A1(new_n17855_), .A2(new_n17879_), .B(new_n17881_), .ZN(new_n18068_));
  INV_X1     g17811(.I(new_n18068_), .ZN(new_n18069_));
  XOR2_X1    g17812(.A1(new_n18067_), .A2(new_n18069_), .Z(new_n18070_));
  NOR2_X1    g17813(.A1(new_n18070_), .A2(new_n18036_), .ZN(new_n18071_));
  INV_X1     g17814(.I(new_n18036_), .ZN(new_n18072_));
  INV_X1     g17815(.I(new_n18067_), .ZN(new_n18073_));
  NOR2_X1    g17816(.A1(new_n18073_), .A2(new_n18069_), .ZN(new_n18074_));
  NOR2_X1    g17817(.A1(new_n18067_), .A2(new_n18068_), .ZN(new_n18075_));
  NOR2_X1    g17818(.A1(new_n18074_), .A2(new_n18075_), .ZN(new_n18076_));
  NOR2_X1    g17819(.A1(new_n18076_), .A2(new_n18072_), .ZN(new_n18077_));
  NOR2_X1    g17820(.A1(new_n18077_), .A2(new_n18071_), .ZN(new_n18078_));
  XNOR2_X1   g17821(.A1(new_n18078_), .A2(new_n18031_), .ZN(new_n18079_));
  NOR2_X1    g17822(.A1(new_n18079_), .A2(new_n18030_), .ZN(new_n18080_));
  INV_X1     g17823(.I(new_n18030_), .ZN(new_n18081_));
  NOR2_X1    g17824(.A1(new_n18078_), .A2(new_n18031_), .ZN(new_n18082_));
  INV_X1     g17825(.I(new_n18082_), .ZN(new_n18083_));
  NAND2_X1   g17826(.A1(new_n18078_), .A2(new_n18031_), .ZN(new_n18084_));
  AOI21_X1   g17827(.A1(new_n18083_), .A2(new_n18084_), .B(new_n18081_), .ZN(new_n18085_));
  NOR2_X1    g17828(.A1(new_n18080_), .A2(new_n18085_), .ZN(new_n18086_));
  INV_X1     g17829(.I(new_n18086_), .ZN(new_n18087_));
  OAI22_X1   g17830(.A1(new_n5228_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n5225_), .ZN(new_n18088_));
  NAND2_X1   g17831(.A1(new_n5387_), .A2(\b[45] ), .ZN(new_n18089_));
  AOI21_X1   g17832(.A1(new_n18088_), .A2(new_n18089_), .B(new_n5231_), .ZN(new_n18090_));
  NAND2_X1   g17833(.A1(new_n5004_), .A2(new_n18090_), .ZN(new_n18091_));
  XOR2_X1    g17834(.A1(new_n18091_), .A2(\a[50] ), .Z(new_n18092_));
  NAND2_X1   g17835(.A1(new_n17897_), .A2(new_n17899_), .ZN(new_n18093_));
  NAND2_X1   g17836(.A1(new_n18093_), .A2(new_n17896_), .ZN(new_n18094_));
  XNOR2_X1   g17837(.A1(new_n18094_), .A2(new_n18092_), .ZN(new_n18095_));
  NAND2_X1   g17838(.A1(new_n18095_), .A2(new_n18087_), .ZN(new_n18096_));
  INV_X1     g17839(.I(new_n18094_), .ZN(new_n18097_));
  NOR2_X1    g17840(.A1(new_n18097_), .A2(new_n18092_), .ZN(new_n18098_));
  NAND2_X1   g17841(.A1(new_n18097_), .A2(new_n18092_), .ZN(new_n18099_));
  INV_X1     g17842(.I(new_n18099_), .ZN(new_n18100_));
  OAI21_X1   g17843(.A1(new_n18100_), .A2(new_n18098_), .B(new_n18086_), .ZN(new_n18101_));
  NAND2_X1   g17844(.A1(new_n18101_), .A2(new_n18096_), .ZN(new_n18102_));
  NAND2_X1   g17845(.A1(new_n17906_), .A2(new_n17908_), .ZN(new_n18103_));
  NAND2_X1   g17846(.A1(new_n18103_), .A2(new_n17905_), .ZN(new_n18104_));
  XNOR2_X1   g17847(.A1(new_n18102_), .A2(new_n18104_), .ZN(new_n18105_));
  NOR2_X1    g17848(.A1(new_n18105_), .A2(new_n18025_), .ZN(new_n18106_));
  INV_X1     g17849(.I(new_n18025_), .ZN(new_n18107_));
  INV_X1     g17850(.I(new_n18102_), .ZN(new_n18108_));
  INV_X1     g17851(.I(new_n18104_), .ZN(new_n18109_));
  NOR2_X1    g17852(.A1(new_n18108_), .A2(new_n18109_), .ZN(new_n18110_));
  NOR2_X1    g17853(.A1(new_n18102_), .A2(new_n18104_), .ZN(new_n18111_));
  NOR2_X1    g17854(.A1(new_n18110_), .A2(new_n18111_), .ZN(new_n18112_));
  NOR2_X1    g17855(.A1(new_n18112_), .A2(new_n18107_), .ZN(new_n18113_));
  NOR2_X1    g17856(.A1(new_n18113_), .A2(new_n18106_), .ZN(new_n18114_));
  NOR2_X1    g17857(.A1(new_n17922_), .A2(new_n17911_), .ZN(new_n18115_));
  NOR2_X1    g17858(.A1(new_n18115_), .A2(new_n17920_), .ZN(new_n18116_));
  XOR2_X1    g17859(.A1(new_n18114_), .A2(new_n18116_), .Z(new_n18117_));
  NOR2_X1    g17860(.A1(new_n18117_), .A2(new_n18020_), .ZN(new_n18118_));
  INV_X1     g17861(.I(new_n18020_), .ZN(new_n18119_));
  INV_X1     g17862(.I(new_n18114_), .ZN(new_n18120_));
  NOR2_X1    g17863(.A1(new_n18120_), .A2(new_n18116_), .ZN(new_n18121_));
  INV_X1     g17864(.I(new_n18121_), .ZN(new_n18122_));
  NAND2_X1   g17865(.A1(new_n18120_), .A2(new_n18116_), .ZN(new_n18123_));
  AOI21_X1   g17866(.A1(new_n18122_), .A2(new_n18123_), .B(new_n18119_), .ZN(new_n18124_));
  NOR2_X1    g17867(.A1(new_n18124_), .A2(new_n18118_), .ZN(new_n18125_));
  XOR2_X1    g17868(.A1(new_n18125_), .A2(new_n18015_), .Z(new_n18126_));
  NOR2_X1    g17869(.A1(new_n18126_), .A2(new_n18013_), .ZN(new_n18127_));
  INV_X1     g17870(.I(new_n18013_), .ZN(new_n18128_));
  INV_X1     g17871(.I(new_n18015_), .ZN(new_n18129_));
  NOR2_X1    g17872(.A1(new_n18129_), .A2(new_n18125_), .ZN(new_n18130_));
  INV_X1     g17873(.I(new_n18130_), .ZN(new_n18131_));
  NAND2_X1   g17874(.A1(new_n18129_), .A2(new_n18125_), .ZN(new_n18132_));
  AOI21_X1   g17875(.A1(new_n18131_), .A2(new_n18132_), .B(new_n18128_), .ZN(new_n18133_));
  NOR2_X1    g17876(.A1(new_n18133_), .A2(new_n18127_), .ZN(new_n18134_));
  OAI22_X1   g17877(.A1(new_n3298_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n3293_), .ZN(new_n18135_));
  NAND2_X1   g17878(.A1(new_n4227_), .A2(\b[57] ), .ZN(new_n18136_));
  AOI21_X1   g17879(.A1(new_n18135_), .A2(new_n18136_), .B(new_n3301_), .ZN(new_n18137_));
  NAND2_X1   g17880(.A1(new_n7895_), .A2(new_n18137_), .ZN(new_n18138_));
  XOR2_X1    g17881(.A1(new_n18138_), .A2(\a[38] ), .Z(new_n18139_));
  NAND2_X1   g17882(.A1(new_n17949_), .A2(new_n17946_), .ZN(new_n18140_));
  NAND2_X1   g17883(.A1(new_n18140_), .A2(new_n17948_), .ZN(new_n18141_));
  XOR2_X1    g17884(.A1(new_n18141_), .A2(new_n18139_), .Z(new_n18142_));
  NOR2_X1    g17885(.A1(new_n18142_), .A2(new_n18134_), .ZN(new_n18143_));
  INV_X1     g17886(.I(new_n18134_), .ZN(new_n18144_));
  INV_X1     g17887(.I(new_n18141_), .ZN(new_n18145_));
  NOR2_X1    g17888(.A1(new_n18145_), .A2(new_n18139_), .ZN(new_n18146_));
  INV_X1     g17889(.I(new_n18146_), .ZN(new_n18147_));
  NAND2_X1   g17890(.A1(new_n18145_), .A2(new_n18139_), .ZN(new_n18148_));
  AOI21_X1   g17891(.A1(new_n18147_), .A2(new_n18148_), .B(new_n18144_), .ZN(new_n18149_));
  NOR2_X1    g17892(.A1(new_n18149_), .A2(new_n18143_), .ZN(new_n18150_));
  INV_X1     g17893(.I(new_n17952_), .ZN(new_n18151_));
  AOI21_X1   g17894(.A1(new_n18151_), .A2(new_n17957_), .B(new_n17954_), .ZN(new_n18152_));
  NOR2_X1    g17895(.A1(new_n18152_), .A2(new_n18150_), .ZN(new_n18153_));
  AND2_X2    g17896(.A1(new_n18152_), .A2(new_n18150_), .Z(new_n18154_));
  NOR2_X1    g17897(.A1(new_n18154_), .A2(new_n18153_), .ZN(new_n18155_));
  NOR2_X1    g17898(.A1(new_n18155_), .A2(new_n18008_), .ZN(new_n18156_));
  INV_X1     g17899(.I(new_n18008_), .ZN(new_n18157_));
  XNOR2_X1   g17900(.A1(new_n18152_), .A2(new_n18150_), .ZN(new_n18158_));
  NOR2_X1    g17901(.A1(new_n18158_), .A2(new_n18157_), .ZN(new_n18159_));
  NOR2_X1    g17902(.A1(new_n18156_), .A2(new_n18159_), .ZN(new_n18160_));
  XOR2_X1    g17903(.A1(new_n18160_), .A2(new_n18003_), .Z(new_n18161_));
  XOR2_X1    g17904(.A1(new_n18161_), .A2(new_n2442_), .Z(new_n18162_));
  XOR2_X1    g17905(.A1(new_n18162_), .A2(new_n18002_), .Z(new_n18163_));
  NOR2_X1    g17906(.A1(new_n18163_), .A2(new_n18001_), .ZN(new_n18164_));
  NAND2_X1   g17907(.A1(new_n18163_), .A2(new_n18001_), .ZN(new_n18165_));
  INV_X1     g17908(.I(new_n18165_), .ZN(new_n18166_));
  NOR2_X1    g17909(.A1(new_n18166_), .A2(new_n18164_), .ZN(new_n18167_));
  INV_X1     g17910(.I(new_n18167_), .ZN(new_n18168_));
  XOR2_X1    g17911(.A1(new_n17999_), .A2(new_n18168_), .Z(\f[95] ));
  NAND2_X1   g17912(.A1(new_n18160_), .A2(new_n18002_), .ZN(new_n18170_));
  XOR2_X1    g17913(.A1(new_n18003_), .A2(\a[32] ), .Z(new_n18171_));
  NAND2_X1   g17914(.A1(new_n18170_), .A2(new_n18171_), .ZN(new_n18172_));
  OAI21_X1   g17915(.A1(new_n18002_), .A2(new_n18160_), .B(new_n18172_), .ZN(new_n18173_));
  INV_X1     g17916(.I(new_n18154_), .ZN(new_n18174_));
  AOI21_X1   g17917(.A1(new_n18174_), .A2(new_n18157_), .B(new_n18153_), .ZN(new_n18175_));
  OAI22_X1   g17918(.A1(new_n2846_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n2841_), .ZN(new_n18176_));
  NAND2_X1   g17919(.A1(new_n3755_), .A2(\b[61] ), .ZN(new_n18177_));
  AOI21_X1   g17920(.A1(new_n18176_), .A2(new_n18177_), .B(new_n2849_), .ZN(new_n18178_));
  NAND2_X1   g17921(.A1(new_n8963_), .A2(new_n18178_), .ZN(new_n18179_));
  XOR2_X1    g17922(.A1(new_n18179_), .A2(\a[35] ), .Z(new_n18180_));
  INV_X1     g17923(.I(new_n18180_), .ZN(new_n18181_));
  OAI21_X1   g17924(.A1(new_n18013_), .A2(new_n18130_), .B(new_n18132_), .ZN(new_n18182_));
  AOI21_X1   g17925(.A1(new_n18119_), .A2(new_n18123_), .B(new_n18121_), .ZN(new_n18183_));
  INV_X1     g17926(.I(new_n18111_), .ZN(new_n18184_));
  AOI21_X1   g17927(.A1(new_n18107_), .A2(new_n18184_), .B(new_n18110_), .ZN(new_n18185_));
  OAI21_X1   g17928(.A1(new_n18030_), .A2(new_n18082_), .B(new_n18084_), .ZN(new_n18186_));
  NOR2_X1    g17929(.A1(new_n18063_), .A2(new_n18050_), .ZN(new_n18187_));
  NOR2_X1    g17930(.A1(new_n18187_), .A2(new_n18062_), .ZN(new_n18188_));
  INV_X1     g17931(.I(new_n18043_), .ZN(new_n18189_));
  AOI21_X1   g17932(.A1(new_n18038_), .A2(new_n18189_), .B(new_n18045_), .ZN(new_n18190_));
  OAI22_X1   g17933(.A1(new_n3247_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n3097_), .ZN(new_n18191_));
  NAND2_X1   g17934(.A1(new_n9644_), .A2(\b[34] ), .ZN(new_n18192_));
  AOI21_X1   g17935(.A1(new_n18192_), .A2(new_n18191_), .B(new_n8321_), .ZN(new_n18193_));
  NAND2_X1   g17936(.A1(new_n3246_), .A2(new_n18193_), .ZN(new_n18194_));
  XOR2_X1    g17937(.A1(new_n18194_), .A2(\a[62] ), .Z(new_n18195_));
  NOR2_X1    g17938(.A1(new_n8985_), .A2(new_n2794_), .ZN(new_n18196_));
  NOR2_X1    g17939(.A1(new_n9364_), .A2(new_n2660_), .ZN(new_n18197_));
  XNOR2_X1   g17940(.A1(new_n18196_), .A2(new_n18197_), .ZN(new_n18198_));
  NOR2_X1    g17941(.A1(new_n18198_), .A2(new_n2442_), .ZN(new_n18199_));
  INV_X1     g17942(.I(new_n18199_), .ZN(new_n18200_));
  NAND2_X1   g17943(.A1(new_n18198_), .A2(new_n2442_), .ZN(new_n18201_));
  AOI21_X1   g17944(.A1(new_n18200_), .A2(new_n18201_), .B(new_n18042_), .ZN(new_n18202_));
  XOR2_X1    g17945(.A1(new_n18198_), .A2(\a[32] ), .Z(new_n18203_));
  NOR2_X1    g17946(.A1(new_n18203_), .A2(new_n18044_), .ZN(new_n18204_));
  NOR2_X1    g17947(.A1(new_n18204_), .A2(new_n18202_), .ZN(new_n18205_));
  NOR2_X1    g17948(.A1(new_n18195_), .A2(new_n18205_), .ZN(new_n18206_));
  AND2_X2    g17949(.A1(new_n18195_), .A2(new_n18205_), .Z(new_n18207_));
  NOR2_X1    g17950(.A1(new_n18207_), .A2(new_n18206_), .ZN(new_n18208_));
  XOR2_X1    g17951(.A1(new_n18195_), .A2(new_n18205_), .Z(new_n18209_));
  NAND2_X1   g17952(.A1(new_n18209_), .A2(new_n18190_), .ZN(new_n18210_));
  OAI21_X1   g17953(.A1(new_n18190_), .A2(new_n18208_), .B(new_n18210_), .ZN(new_n18211_));
  OAI22_X1   g17954(.A1(new_n3696_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n3566_), .ZN(new_n18212_));
  NAND2_X1   g17955(.A1(new_n8628_), .A2(\b[37] ), .ZN(new_n18213_));
  AOI21_X1   g17956(.A1(new_n18213_), .A2(new_n18212_), .B(new_n7354_), .ZN(new_n18214_));
  NAND2_X1   g17957(.A1(new_n3700_), .A2(new_n18214_), .ZN(new_n18215_));
  XOR2_X1    g17958(.A1(new_n18215_), .A2(\a[59] ), .Z(new_n18216_));
  XOR2_X1    g17959(.A1(new_n18211_), .A2(new_n18216_), .Z(new_n18217_));
  NOR2_X1    g17960(.A1(new_n18217_), .A2(new_n18188_), .ZN(new_n18218_));
  INV_X1     g17961(.I(new_n18188_), .ZN(new_n18219_));
  INV_X1     g17962(.I(new_n18211_), .ZN(new_n18220_));
  NOR2_X1    g17963(.A1(new_n18220_), .A2(new_n18216_), .ZN(new_n18221_));
  INV_X1     g17964(.I(new_n18221_), .ZN(new_n18222_));
  NAND2_X1   g17965(.A1(new_n18220_), .A2(new_n18216_), .ZN(new_n18223_));
  AOI21_X1   g17966(.A1(new_n18222_), .A2(new_n18223_), .B(new_n18219_), .ZN(new_n18224_));
  NOR2_X1    g17967(.A1(new_n18224_), .A2(new_n18218_), .ZN(new_n18225_));
  OAI22_X1   g17968(.A1(new_n6721_), .A2(new_n3997_), .B1(new_n6723_), .B2(new_n4018_), .ZN(new_n18226_));
  NAND2_X1   g17969(.A1(new_n7617_), .A2(\b[40] ), .ZN(new_n18227_));
  AOI21_X1   g17970(.A1(new_n18227_), .A2(new_n18226_), .B(new_n6731_), .ZN(new_n18228_));
  NAND2_X1   g17971(.A1(new_n4017_), .A2(new_n18228_), .ZN(new_n18229_));
  XOR2_X1    g17972(.A1(new_n18229_), .A2(\a[56] ), .Z(new_n18230_));
  INV_X1     g17973(.I(new_n18075_), .ZN(new_n18231_));
  AOI21_X1   g17974(.A1(new_n18072_), .A2(new_n18231_), .B(new_n18074_), .ZN(new_n18232_));
  NOR2_X1    g17975(.A1(new_n18232_), .A2(new_n18230_), .ZN(new_n18233_));
  AND2_X2    g17976(.A1(new_n18232_), .A2(new_n18230_), .Z(new_n18234_));
  NOR2_X1    g17977(.A1(new_n18234_), .A2(new_n18233_), .ZN(new_n18235_));
  NOR2_X1    g17978(.A1(new_n18235_), .A2(new_n18225_), .ZN(new_n18236_));
  XNOR2_X1   g17979(.A1(new_n18232_), .A2(new_n18230_), .ZN(new_n18237_));
  NOR3_X1    g17980(.A1(new_n18237_), .A2(new_n18218_), .A3(new_n18224_), .ZN(new_n18238_));
  NOR2_X1    g17981(.A1(new_n18238_), .A2(new_n18236_), .ZN(new_n18239_));
  OAI22_X1   g17982(.A1(new_n5786_), .A2(new_n4509_), .B1(new_n4501_), .B2(new_n5792_), .ZN(new_n18240_));
  NAND2_X1   g17983(.A1(new_n6745_), .A2(\b[43] ), .ZN(new_n18241_));
  AOI21_X1   g17984(.A1(new_n18241_), .A2(new_n18240_), .B(new_n5796_), .ZN(new_n18242_));
  NAND2_X1   g17985(.A1(new_n4513_), .A2(new_n18242_), .ZN(new_n18243_));
  XOR2_X1    g17986(.A1(new_n18243_), .A2(\a[53] ), .Z(new_n18244_));
  INV_X1     g17987(.I(new_n18244_), .ZN(new_n18245_));
  XOR2_X1    g17988(.A1(new_n18239_), .A2(new_n18245_), .Z(new_n18246_));
  AND2_X2    g17989(.A1(new_n18246_), .A2(new_n18186_), .Z(new_n18247_));
  NAND2_X1   g17990(.A1(new_n18239_), .A2(new_n18245_), .ZN(new_n18248_));
  OAI21_X1   g17991(.A1(new_n18238_), .A2(new_n18236_), .B(new_n18244_), .ZN(new_n18249_));
  AOI21_X1   g17992(.A1(new_n18248_), .A2(new_n18249_), .B(new_n18186_), .ZN(new_n18250_));
  NOR2_X1    g17993(.A1(new_n18247_), .A2(new_n18250_), .ZN(new_n18251_));
  OAI22_X1   g17994(.A1(new_n5228_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n5225_), .ZN(new_n18252_));
  NAND2_X1   g17995(.A1(new_n5387_), .A2(\b[46] ), .ZN(new_n18253_));
  AOI21_X1   g17996(.A1(new_n18252_), .A2(new_n18253_), .B(new_n5231_), .ZN(new_n18254_));
  NAND2_X1   g17997(.A1(new_n5177_), .A2(new_n18254_), .ZN(new_n18255_));
  XOR2_X1    g17998(.A1(new_n18255_), .A2(\a[50] ), .Z(new_n18256_));
  NOR2_X1    g17999(.A1(new_n18100_), .A2(new_n18087_), .ZN(new_n18257_));
  NOR2_X1    g18000(.A1(new_n18257_), .A2(new_n18098_), .ZN(new_n18258_));
  NOR2_X1    g18001(.A1(new_n18258_), .A2(new_n18256_), .ZN(new_n18259_));
  INV_X1     g18002(.I(new_n18256_), .ZN(new_n18260_));
  NOR3_X1    g18003(.A1(new_n18257_), .A2(new_n18098_), .A3(new_n18260_), .ZN(new_n18261_));
  NOR2_X1    g18004(.A1(new_n18259_), .A2(new_n18261_), .ZN(new_n18262_));
  NOR2_X1    g18005(.A1(new_n18262_), .A2(new_n18251_), .ZN(new_n18263_));
  XOR2_X1    g18006(.A1(new_n18258_), .A2(new_n18260_), .Z(new_n18264_));
  NOR3_X1    g18007(.A1(new_n18264_), .A2(new_n18247_), .A3(new_n18250_), .ZN(new_n18265_));
  NOR2_X1    g18008(.A1(new_n18265_), .A2(new_n18263_), .ZN(new_n18266_));
  INV_X1     g18009(.I(new_n18266_), .ZN(new_n18267_));
  OAI22_X1   g18010(.A1(new_n4711_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n4706_), .ZN(new_n18268_));
  NAND2_X1   g18011(.A1(new_n5814_), .A2(\b[49] ), .ZN(new_n18269_));
  AOI21_X1   g18012(.A1(new_n18268_), .A2(new_n18269_), .B(new_n4714_), .ZN(new_n18270_));
  NAND2_X1   g18013(.A1(new_n5741_), .A2(new_n18270_), .ZN(new_n18271_));
  XOR2_X1    g18014(.A1(new_n18271_), .A2(\a[47] ), .Z(new_n18272_));
  NOR2_X1    g18015(.A1(new_n18267_), .A2(new_n18272_), .ZN(new_n18273_));
  INV_X1     g18016(.I(new_n18272_), .ZN(new_n18274_));
  NOR2_X1    g18017(.A1(new_n18266_), .A2(new_n18274_), .ZN(new_n18275_));
  NOR2_X1    g18018(.A1(new_n18273_), .A2(new_n18275_), .ZN(new_n18276_));
  NOR2_X1    g18019(.A1(new_n18276_), .A2(new_n18185_), .ZN(new_n18277_));
  INV_X1     g18020(.I(new_n18185_), .ZN(new_n18278_));
  XOR2_X1    g18021(.A1(new_n18266_), .A2(new_n18272_), .Z(new_n18279_));
  NOR2_X1    g18022(.A1(new_n18279_), .A2(new_n18278_), .ZN(new_n18280_));
  NOR2_X1    g18023(.A1(new_n18277_), .A2(new_n18280_), .ZN(new_n18281_));
  OAI22_X1   g18024(.A1(new_n4208_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n4203_), .ZN(new_n18282_));
  NAND2_X1   g18025(.A1(new_n5244_), .A2(\b[52] ), .ZN(new_n18283_));
  AOI21_X1   g18026(.A1(new_n18282_), .A2(new_n18283_), .B(new_n4211_), .ZN(new_n18284_));
  NAND2_X1   g18027(.A1(new_n6237_), .A2(new_n18284_), .ZN(new_n18285_));
  XOR2_X1    g18028(.A1(new_n18285_), .A2(\a[44] ), .Z(new_n18286_));
  XNOR2_X1   g18029(.A1(new_n18281_), .A2(new_n18286_), .ZN(new_n18287_));
  NOR2_X1    g18030(.A1(new_n18287_), .A2(new_n18183_), .ZN(new_n18288_));
  INV_X1     g18031(.I(new_n18183_), .ZN(new_n18289_));
  NOR2_X1    g18032(.A1(new_n18281_), .A2(new_n18286_), .ZN(new_n18290_));
  INV_X1     g18033(.I(new_n18290_), .ZN(new_n18291_));
  NAND2_X1   g18034(.A1(new_n18281_), .A2(new_n18286_), .ZN(new_n18292_));
  AOI21_X1   g18035(.A1(new_n18291_), .A2(new_n18292_), .B(new_n18289_), .ZN(new_n18293_));
  NOR2_X1    g18036(.A1(new_n18288_), .A2(new_n18293_), .ZN(new_n18294_));
  OAI22_X1   g18037(.A1(new_n3736_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n3731_), .ZN(new_n18295_));
  NAND2_X1   g18038(.A1(new_n4730_), .A2(\b[55] ), .ZN(new_n18296_));
  AOI21_X1   g18039(.A1(new_n18295_), .A2(new_n18296_), .B(new_n3739_), .ZN(new_n18297_));
  NAND2_X1   g18040(.A1(new_n7308_), .A2(new_n18297_), .ZN(new_n18298_));
  XOR2_X1    g18041(.A1(new_n18298_), .A2(\a[41] ), .Z(new_n18299_));
  XOR2_X1    g18042(.A1(new_n18294_), .A2(new_n18299_), .Z(new_n18300_));
  INV_X1     g18043(.I(new_n18300_), .ZN(new_n18301_));
  INV_X1     g18044(.I(new_n18294_), .ZN(new_n18302_));
  NOR2_X1    g18045(.A1(new_n18302_), .A2(new_n18299_), .ZN(new_n18303_));
  INV_X1     g18046(.I(new_n18303_), .ZN(new_n18304_));
  NAND2_X1   g18047(.A1(new_n18302_), .A2(new_n18299_), .ZN(new_n18305_));
  AOI21_X1   g18048(.A1(new_n18304_), .A2(new_n18305_), .B(new_n18182_), .ZN(new_n18306_));
  AOI21_X1   g18049(.A1(new_n18182_), .A2(new_n18301_), .B(new_n18306_), .ZN(new_n18307_));
  INV_X1     g18050(.I(new_n18307_), .ZN(new_n18308_));
  OAI22_X1   g18051(.A1(new_n3298_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n3293_), .ZN(new_n18309_));
  NAND2_X1   g18052(.A1(new_n4227_), .A2(\b[58] ), .ZN(new_n18310_));
  AOI21_X1   g18053(.A1(new_n18309_), .A2(new_n18310_), .B(new_n3301_), .ZN(new_n18311_));
  NAND2_X1   g18054(.A1(new_n7929_), .A2(new_n18311_), .ZN(new_n18312_));
  XOR2_X1    g18055(.A1(new_n18312_), .A2(\a[38] ), .Z(new_n18313_));
  NAND2_X1   g18056(.A1(new_n18148_), .A2(new_n18134_), .ZN(new_n18314_));
  AOI21_X1   g18057(.A1(new_n18314_), .A2(new_n18147_), .B(new_n18313_), .ZN(new_n18315_));
  INV_X1     g18058(.I(new_n18313_), .ZN(new_n18316_));
  NAND2_X1   g18059(.A1(new_n18314_), .A2(new_n18147_), .ZN(new_n18317_));
  NOR2_X1    g18060(.A1(new_n18317_), .A2(new_n18316_), .ZN(new_n18318_));
  OAI21_X1   g18061(.A1(new_n18315_), .A2(new_n18318_), .B(new_n18308_), .ZN(new_n18319_));
  XOR2_X1    g18062(.A1(new_n18317_), .A2(new_n18313_), .Z(new_n18320_));
  OAI21_X1   g18063(.A1(new_n18308_), .A2(new_n18320_), .B(new_n18319_), .ZN(new_n18321_));
  XOR2_X1    g18064(.A1(new_n18321_), .A2(new_n18181_), .Z(new_n18322_));
  NOR2_X1    g18065(.A1(new_n18322_), .A2(new_n18175_), .ZN(new_n18323_));
  INV_X1     g18066(.I(new_n18175_), .ZN(new_n18324_));
  AND2_X2    g18067(.A1(new_n18321_), .A2(new_n18180_), .Z(new_n18325_));
  NOR2_X1    g18068(.A1(new_n18321_), .A2(new_n18180_), .ZN(new_n18326_));
  NOR2_X1    g18069(.A1(new_n18325_), .A2(new_n18326_), .ZN(new_n18327_));
  NOR2_X1    g18070(.A1(new_n18327_), .A2(new_n18324_), .ZN(new_n18328_));
  NOR2_X1    g18071(.A1(new_n18328_), .A2(new_n18323_), .ZN(new_n18329_));
  XNOR2_X1   g18072(.A1(new_n18329_), .A2(new_n18173_), .ZN(new_n18330_));
  NAND3_X1   g18073(.A1(new_n17998_), .A2(new_n17995_), .A3(new_n18167_), .ZN(new_n18331_));
  NAND3_X1   g18074(.A1(new_n18331_), .A2(new_n18165_), .A3(new_n18330_), .ZN(new_n18332_));
  INV_X1     g18075(.I(new_n18330_), .ZN(new_n18333_));
  INV_X1     g18076(.I(new_n17997_), .ZN(new_n18334_));
  AOI21_X1   g18077(.A1(new_n17814_), .A2(new_n17812_), .B(new_n18334_), .ZN(new_n18335_));
  NOR3_X1    g18078(.A1(new_n18335_), .A2(new_n17994_), .A3(new_n18168_), .ZN(new_n18336_));
  OAI21_X1   g18079(.A1(new_n18336_), .A2(new_n18166_), .B(new_n18333_), .ZN(new_n18337_));
  NAND2_X1   g18080(.A1(new_n18337_), .A2(new_n18332_), .ZN(\f[96] ));
  NOR2_X1    g18081(.A1(new_n3015_), .A2(new_n8932_), .ZN(new_n18339_));
  NOR2_X1    g18082(.A1(new_n2841_), .A2(new_n8956_), .ZN(new_n18340_));
  NOR4_X1    g18083(.A1(new_n9323_), .A2(new_n2849_), .A3(new_n18339_), .A4(new_n18340_), .ZN(new_n18341_));
  XOR2_X1    g18084(.A1(new_n18341_), .A2(new_n2836_), .Z(new_n18342_));
  NOR2_X1    g18085(.A1(new_n18308_), .A2(new_n18318_), .ZN(new_n18343_));
  OAI22_X1   g18086(.A1(new_n3736_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n3731_), .ZN(new_n18344_));
  NAND2_X1   g18087(.A1(new_n4730_), .A2(\b[56] ), .ZN(new_n18345_));
  AOI21_X1   g18088(.A1(new_n18344_), .A2(new_n18345_), .B(new_n3739_), .ZN(new_n18346_));
  NAND2_X1   g18089(.A1(new_n7559_), .A2(new_n18346_), .ZN(new_n18347_));
  XOR2_X1    g18090(.A1(new_n18347_), .A2(\a[41] ), .Z(new_n18348_));
  AOI21_X1   g18091(.A1(new_n18289_), .A2(new_n18292_), .B(new_n18290_), .ZN(new_n18349_));
  INV_X1     g18092(.I(new_n18349_), .ZN(new_n18350_));
  INV_X1     g18093(.I(new_n18275_), .ZN(new_n18351_));
  AOI21_X1   g18094(.A1(new_n18278_), .A2(new_n18351_), .B(new_n18273_), .ZN(new_n18352_));
  OAI22_X1   g18095(.A1(new_n4711_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n4706_), .ZN(new_n18353_));
  NAND2_X1   g18096(.A1(new_n5814_), .A2(\b[50] ), .ZN(new_n18354_));
  AOI21_X1   g18097(.A1(new_n18353_), .A2(new_n18354_), .B(new_n4714_), .ZN(new_n18355_));
  NAND2_X1   g18098(.A1(new_n5954_), .A2(new_n18355_), .ZN(new_n18356_));
  XOR2_X1    g18099(.A1(new_n18356_), .A2(\a[47] ), .Z(new_n18357_));
  OAI22_X1   g18100(.A1(new_n5786_), .A2(new_n4834_), .B1(new_n4509_), .B2(new_n5792_), .ZN(new_n18358_));
  NAND2_X1   g18101(.A1(new_n6745_), .A2(\b[44] ), .ZN(new_n18359_));
  AOI21_X1   g18102(.A1(new_n18359_), .A2(new_n18358_), .B(new_n5796_), .ZN(new_n18360_));
  NAND2_X1   g18103(.A1(new_n4833_), .A2(new_n18360_), .ZN(new_n18361_));
  XOR2_X1    g18104(.A1(new_n18361_), .A2(\a[53] ), .Z(new_n18362_));
  AOI21_X1   g18105(.A1(new_n18219_), .A2(new_n18223_), .B(new_n18221_), .ZN(new_n18363_));
  OAI22_X1   g18106(.A1(new_n3845_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n3696_), .ZN(new_n18364_));
  NAND2_X1   g18107(.A1(new_n8628_), .A2(\b[38] ), .ZN(new_n18365_));
  AOI21_X1   g18108(.A1(new_n18365_), .A2(new_n18364_), .B(new_n7354_), .ZN(new_n18366_));
  NAND2_X1   g18109(.A1(new_n3844_), .A2(new_n18366_), .ZN(new_n18367_));
  XOR2_X1    g18110(.A1(new_n18367_), .A2(\a[59] ), .Z(new_n18368_));
  NOR2_X1    g18111(.A1(new_n18190_), .A2(new_n18207_), .ZN(new_n18369_));
  NOR2_X1    g18112(.A1(new_n18369_), .A2(new_n18206_), .ZN(new_n18370_));
  OAI22_X1   g18113(.A1(new_n3408_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n3247_), .ZN(new_n18371_));
  NAND2_X1   g18114(.A1(new_n9644_), .A2(\b[35] ), .ZN(new_n18372_));
  AOI21_X1   g18115(.A1(new_n18372_), .A2(new_n18371_), .B(new_n8321_), .ZN(new_n18373_));
  NAND2_X1   g18116(.A1(new_n3411_), .A2(new_n18373_), .ZN(new_n18374_));
  XOR2_X1    g18117(.A1(new_n18374_), .A2(\a[62] ), .Z(new_n18375_));
  NAND2_X1   g18118(.A1(new_n18201_), .A2(new_n18044_), .ZN(new_n18376_));
  NAND2_X1   g18119(.A1(new_n18376_), .A2(new_n18200_), .ZN(new_n18377_));
  NOR3_X1    g18120(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n2794_), .ZN(new_n18378_));
  NOR2_X1    g18121(.A1(new_n9364_), .A2(new_n2794_), .ZN(new_n18379_));
  NOR3_X1    g18122(.A1(new_n18379_), .A2(new_n2964_), .A3(new_n8985_), .ZN(new_n18380_));
  NOR2_X1    g18123(.A1(new_n18380_), .A2(new_n18378_), .ZN(new_n18381_));
  INV_X1     g18124(.I(new_n18381_), .ZN(new_n18382_));
  XOR2_X1    g18125(.A1(new_n18377_), .A2(new_n18382_), .Z(new_n18383_));
  NOR2_X1    g18126(.A1(new_n18375_), .A2(new_n18383_), .ZN(new_n18384_));
  NOR2_X1    g18127(.A1(new_n18377_), .A2(new_n18381_), .ZN(new_n18385_));
  INV_X1     g18128(.I(new_n18385_), .ZN(new_n18386_));
  NAND2_X1   g18129(.A1(new_n18377_), .A2(new_n18381_), .ZN(new_n18387_));
  NAND2_X1   g18130(.A1(new_n18386_), .A2(new_n18387_), .ZN(new_n18388_));
  AOI21_X1   g18131(.A1(new_n18375_), .A2(new_n18388_), .B(new_n18384_), .ZN(new_n18389_));
  XOR2_X1    g18132(.A1(new_n18389_), .A2(new_n18370_), .Z(new_n18390_));
  NOR2_X1    g18133(.A1(new_n18390_), .A2(new_n18368_), .ZN(new_n18391_));
  INV_X1     g18134(.I(new_n18368_), .ZN(new_n18392_));
  INV_X1     g18135(.I(new_n18370_), .ZN(new_n18393_));
  NOR2_X1    g18136(.A1(new_n18389_), .A2(new_n18393_), .ZN(new_n18394_));
  INV_X1     g18137(.I(new_n18394_), .ZN(new_n18395_));
  NAND2_X1   g18138(.A1(new_n18389_), .A2(new_n18393_), .ZN(new_n18396_));
  AOI21_X1   g18139(.A1(new_n18395_), .A2(new_n18396_), .B(new_n18392_), .ZN(new_n18397_));
  NOR2_X1    g18140(.A1(new_n18391_), .A2(new_n18397_), .ZN(new_n18398_));
  INV_X1     g18141(.I(new_n18398_), .ZN(new_n18399_));
  OAI22_X1   g18142(.A1(new_n6721_), .A2(new_n4018_), .B1(new_n6723_), .B2(new_n4316_), .ZN(new_n18400_));
  NAND2_X1   g18143(.A1(new_n7617_), .A2(\b[41] ), .ZN(new_n18401_));
  AOI21_X1   g18144(.A1(new_n18401_), .A2(new_n18400_), .B(new_n6731_), .ZN(new_n18402_));
  NAND2_X1   g18145(.A1(new_n4320_), .A2(new_n18402_), .ZN(new_n18403_));
  XOR2_X1    g18146(.A1(new_n18403_), .A2(\a[56] ), .Z(new_n18404_));
  NOR2_X1    g18147(.A1(new_n18399_), .A2(new_n18404_), .ZN(new_n18405_));
  INV_X1     g18148(.I(new_n18404_), .ZN(new_n18406_));
  NOR2_X1    g18149(.A1(new_n18398_), .A2(new_n18406_), .ZN(new_n18407_));
  NOR2_X1    g18150(.A1(new_n18405_), .A2(new_n18407_), .ZN(new_n18408_));
  NOR2_X1    g18151(.A1(new_n18408_), .A2(new_n18363_), .ZN(new_n18409_));
  INV_X1     g18152(.I(new_n18363_), .ZN(new_n18410_));
  XOR2_X1    g18153(.A1(new_n18398_), .A2(new_n18404_), .Z(new_n18411_));
  NOR2_X1    g18154(.A1(new_n18411_), .A2(new_n18410_), .ZN(new_n18412_));
  NOR2_X1    g18155(.A1(new_n18409_), .A2(new_n18412_), .ZN(new_n18413_));
  INV_X1     g18156(.I(new_n18234_), .ZN(new_n18414_));
  AOI21_X1   g18157(.A1(new_n18414_), .A2(new_n18225_), .B(new_n18233_), .ZN(new_n18415_));
  NOR2_X1    g18158(.A1(new_n18413_), .A2(new_n18415_), .ZN(new_n18416_));
  INV_X1     g18159(.I(new_n18416_), .ZN(new_n18417_));
  NAND2_X1   g18160(.A1(new_n18413_), .A2(new_n18415_), .ZN(new_n18418_));
  AOI21_X1   g18161(.A1(new_n18417_), .A2(new_n18418_), .B(new_n18362_), .ZN(new_n18419_));
  INV_X1     g18162(.I(new_n18362_), .ZN(new_n18420_));
  XNOR2_X1   g18163(.A1(new_n18413_), .A2(new_n18415_), .ZN(new_n18421_));
  NOR2_X1    g18164(.A1(new_n18421_), .A2(new_n18420_), .ZN(new_n18422_));
  NOR2_X1    g18165(.A1(new_n18422_), .A2(new_n18419_), .ZN(new_n18423_));
  NAND2_X1   g18166(.A1(new_n18249_), .A2(new_n18186_), .ZN(new_n18424_));
  NAND2_X1   g18167(.A1(new_n18424_), .A2(new_n18248_), .ZN(new_n18425_));
  OAI22_X1   g18168(.A1(new_n5228_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n5225_), .ZN(new_n18426_));
  NAND2_X1   g18169(.A1(new_n5387_), .A2(\b[47] ), .ZN(new_n18427_));
  AOI21_X1   g18170(.A1(new_n18426_), .A2(new_n18427_), .B(new_n5231_), .ZN(new_n18428_));
  NAND2_X1   g18171(.A1(new_n5196_), .A2(new_n18428_), .ZN(new_n18429_));
  XOR2_X1    g18172(.A1(new_n18429_), .A2(\a[50] ), .Z(new_n18430_));
  INV_X1     g18173(.I(new_n18430_), .ZN(new_n18431_));
  NAND2_X1   g18174(.A1(new_n18425_), .A2(new_n18431_), .ZN(new_n18432_));
  NOR2_X1    g18175(.A1(new_n18425_), .A2(new_n18431_), .ZN(new_n18433_));
  INV_X1     g18176(.I(new_n18433_), .ZN(new_n18434_));
  AOI21_X1   g18177(.A1(new_n18434_), .A2(new_n18432_), .B(new_n18423_), .ZN(new_n18435_));
  XOR2_X1    g18178(.A1(new_n18425_), .A2(new_n18430_), .Z(new_n18436_));
  NOR3_X1    g18179(.A1(new_n18436_), .A2(new_n18419_), .A3(new_n18422_), .ZN(new_n18437_));
  NOR2_X1    g18180(.A1(new_n18435_), .A2(new_n18437_), .ZN(new_n18438_));
  INV_X1     g18181(.I(new_n18261_), .ZN(new_n18439_));
  AOI21_X1   g18182(.A1(new_n18439_), .A2(new_n18251_), .B(new_n18259_), .ZN(new_n18440_));
  NOR2_X1    g18183(.A1(new_n18440_), .A2(new_n18438_), .ZN(new_n18441_));
  INV_X1     g18184(.I(new_n18438_), .ZN(new_n18442_));
  INV_X1     g18185(.I(new_n18440_), .ZN(new_n18443_));
  NOR2_X1    g18186(.A1(new_n18443_), .A2(new_n18442_), .ZN(new_n18444_));
  NOR2_X1    g18187(.A1(new_n18444_), .A2(new_n18441_), .ZN(new_n18445_));
  NOR2_X1    g18188(.A1(new_n18445_), .A2(new_n18357_), .ZN(new_n18446_));
  XOR2_X1    g18189(.A1(new_n18440_), .A2(new_n18438_), .Z(new_n18447_));
  AOI21_X1   g18190(.A1(new_n18357_), .A2(new_n18447_), .B(new_n18446_), .ZN(new_n18448_));
  OAI22_X1   g18191(.A1(new_n4208_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n4203_), .ZN(new_n18449_));
  NAND2_X1   g18192(.A1(new_n5244_), .A2(\b[53] ), .ZN(new_n18450_));
  AOI21_X1   g18193(.A1(new_n18449_), .A2(new_n18450_), .B(new_n4211_), .ZN(new_n18451_));
  NAND2_X1   g18194(.A1(new_n6471_), .A2(new_n18451_), .ZN(new_n18452_));
  XOR2_X1    g18195(.A1(new_n18452_), .A2(\a[44] ), .Z(new_n18453_));
  XNOR2_X1   g18196(.A1(new_n18448_), .A2(new_n18453_), .ZN(new_n18454_));
  NOR2_X1    g18197(.A1(new_n18454_), .A2(new_n18352_), .ZN(new_n18455_));
  INV_X1     g18198(.I(new_n18352_), .ZN(new_n18456_));
  NOR2_X1    g18199(.A1(new_n18448_), .A2(new_n18453_), .ZN(new_n18457_));
  INV_X1     g18200(.I(new_n18457_), .ZN(new_n18458_));
  NAND2_X1   g18201(.A1(new_n18448_), .A2(new_n18453_), .ZN(new_n18459_));
  AOI21_X1   g18202(.A1(new_n18458_), .A2(new_n18459_), .B(new_n18456_), .ZN(new_n18460_));
  NOR2_X1    g18203(.A1(new_n18455_), .A2(new_n18460_), .ZN(new_n18461_));
  NOR2_X1    g18204(.A1(new_n18350_), .A2(new_n18461_), .ZN(new_n18462_));
  INV_X1     g18205(.I(new_n18462_), .ZN(new_n18463_));
  NAND2_X1   g18206(.A1(new_n18350_), .A2(new_n18461_), .ZN(new_n18464_));
  AOI21_X1   g18207(.A1(new_n18463_), .A2(new_n18464_), .B(new_n18348_), .ZN(new_n18465_));
  INV_X1     g18208(.I(new_n18348_), .ZN(new_n18466_));
  XOR2_X1    g18209(.A1(new_n18461_), .A2(new_n18349_), .Z(new_n18467_));
  NOR2_X1    g18210(.A1(new_n18467_), .A2(new_n18466_), .ZN(new_n18468_));
  NOR2_X1    g18211(.A1(new_n18468_), .A2(new_n18465_), .ZN(new_n18469_));
  AOI21_X1   g18212(.A1(new_n18182_), .A2(new_n18305_), .B(new_n18303_), .ZN(new_n18470_));
  OAI22_X1   g18213(.A1(new_n3298_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n3293_), .ZN(new_n18471_));
  NAND2_X1   g18214(.A1(new_n4227_), .A2(\b[59] ), .ZN(new_n18472_));
  AOI21_X1   g18215(.A1(new_n18471_), .A2(new_n18472_), .B(new_n3301_), .ZN(new_n18473_));
  NAND2_X1   g18216(.A1(new_n8550_), .A2(new_n18473_), .ZN(new_n18474_));
  XOR2_X1    g18217(.A1(new_n18474_), .A2(\a[38] ), .Z(new_n18475_));
  XNOR2_X1   g18218(.A1(new_n18470_), .A2(new_n18475_), .ZN(new_n18476_));
  NOR2_X1    g18219(.A1(new_n18476_), .A2(new_n18469_), .ZN(new_n18477_));
  INV_X1     g18220(.I(new_n18469_), .ZN(new_n18478_));
  NOR2_X1    g18221(.A1(new_n18470_), .A2(new_n18475_), .ZN(new_n18479_));
  INV_X1     g18222(.I(new_n18479_), .ZN(new_n18480_));
  NAND2_X1   g18223(.A1(new_n18470_), .A2(new_n18475_), .ZN(new_n18481_));
  AOI21_X1   g18224(.A1(new_n18480_), .A2(new_n18481_), .B(new_n18478_), .ZN(new_n18482_));
  NOR2_X1    g18225(.A1(new_n18477_), .A2(new_n18482_), .ZN(new_n18483_));
  NOR3_X1    g18226(.A1(new_n18483_), .A2(new_n18315_), .A3(new_n18343_), .ZN(new_n18484_));
  NOR2_X1    g18227(.A1(new_n18343_), .A2(new_n18315_), .ZN(new_n18485_));
  INV_X1     g18228(.I(new_n18483_), .ZN(new_n18486_));
  NOR2_X1    g18229(.A1(new_n18486_), .A2(new_n18485_), .ZN(new_n18487_));
  NOR2_X1    g18230(.A1(new_n18487_), .A2(new_n18484_), .ZN(new_n18488_));
  NOR2_X1    g18231(.A1(new_n18488_), .A2(new_n18342_), .ZN(new_n18489_));
  INV_X1     g18232(.I(new_n18342_), .ZN(new_n18490_));
  XOR2_X1    g18233(.A1(new_n18485_), .A2(new_n18483_), .Z(new_n18491_));
  NOR2_X1    g18234(.A1(new_n18491_), .A2(new_n18490_), .ZN(new_n18492_));
  NOR2_X1    g18235(.A1(new_n18489_), .A2(new_n18492_), .ZN(new_n18493_));
  NOR2_X1    g18236(.A1(new_n18325_), .A2(new_n18175_), .ZN(new_n18494_));
  NOR2_X1    g18237(.A1(new_n18494_), .A2(new_n18326_), .ZN(new_n18495_));
  NOR3_X1    g18238(.A1(new_n18336_), .A2(new_n18166_), .A3(new_n18333_), .ZN(new_n18496_));
  NOR2_X1    g18239(.A1(new_n18329_), .A2(new_n18173_), .ZN(new_n18497_));
  NOR2_X1    g18240(.A1(new_n18496_), .A2(new_n18497_), .ZN(new_n18498_));
  XNOR2_X1   g18241(.A1(new_n18498_), .A2(new_n18495_), .ZN(new_n18499_));
  XOR2_X1    g18242(.A1(new_n18499_), .A2(new_n18493_), .Z(\f[97] ));
  XNOR2_X1   g18243(.A1(new_n18493_), .A2(new_n18495_), .ZN(new_n18501_));
  INV_X1     g18244(.I(new_n18501_), .ZN(new_n18502_));
  NAND2_X1   g18245(.A1(new_n18502_), .A2(new_n18495_), .ZN(new_n18503_));
  INV_X1     g18246(.I(new_n18503_), .ZN(new_n18504_));
  NOR2_X1    g18247(.A1(new_n18501_), .A2(new_n18497_), .ZN(new_n18505_));
  AOI21_X1   g18248(.A1(new_n18332_), .A2(new_n18505_), .B(new_n18504_), .ZN(new_n18506_));
  INV_X1     g18249(.I(new_n18484_), .ZN(new_n18507_));
  AOI21_X1   g18250(.A1(new_n18507_), .A2(new_n18490_), .B(new_n18487_), .ZN(new_n18508_));
  INV_X1     g18251(.I(new_n18508_), .ZN(new_n18509_));
  AOI21_X1   g18252(.A1(new_n18478_), .A2(new_n18481_), .B(new_n18479_), .ZN(new_n18510_));
  OAI22_X1   g18253(.A1(new_n9595_), .A2(new_n2849_), .B1(new_n8956_), .B2(new_n3015_), .ZN(new_n18511_));
  OAI22_X1   g18254(.A1(new_n3298_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n3293_), .ZN(new_n18512_));
  NAND2_X1   g18255(.A1(new_n4227_), .A2(\b[60] ), .ZN(new_n18513_));
  AOI21_X1   g18256(.A1(new_n18512_), .A2(new_n18513_), .B(new_n3301_), .ZN(new_n18514_));
  NAND2_X1   g18257(.A1(new_n8935_), .A2(new_n18514_), .ZN(new_n18515_));
  XOR2_X1    g18258(.A1(new_n18515_), .A2(\a[38] ), .Z(new_n18516_));
  OAI22_X1   g18259(.A1(new_n4208_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n4203_), .ZN(new_n18517_));
  NAND2_X1   g18260(.A1(new_n5244_), .A2(\b[54] ), .ZN(new_n18518_));
  AOI21_X1   g18261(.A1(new_n18517_), .A2(new_n18518_), .B(new_n4211_), .ZN(new_n18519_));
  NAND2_X1   g18262(.A1(new_n6994_), .A2(new_n18519_), .ZN(new_n18520_));
  XOR2_X1    g18263(.A1(new_n18520_), .A2(\a[44] ), .Z(new_n18521_));
  INV_X1     g18264(.I(new_n18441_), .ZN(new_n18522_));
  OAI21_X1   g18265(.A1(new_n18357_), .A2(new_n18444_), .B(new_n18522_), .ZN(new_n18523_));
  OAI22_X1   g18266(.A1(new_n4711_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n4706_), .ZN(new_n18524_));
  NAND2_X1   g18267(.A1(new_n5814_), .A2(\b[51] ), .ZN(new_n18525_));
  AOI21_X1   g18268(.A1(new_n18524_), .A2(new_n18525_), .B(new_n4714_), .ZN(new_n18526_));
  NAND2_X1   g18269(.A1(new_n6219_), .A2(new_n18526_), .ZN(new_n18527_));
  XOR2_X1    g18270(.A1(new_n18527_), .A2(\a[47] ), .Z(new_n18528_));
  OAI22_X1   g18271(.A1(new_n5228_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n5225_), .ZN(new_n18529_));
  NAND2_X1   g18272(.A1(new_n5387_), .A2(\b[48] ), .ZN(new_n18530_));
  AOI21_X1   g18273(.A1(new_n18529_), .A2(new_n18530_), .B(new_n5231_), .ZN(new_n18531_));
  NAND2_X1   g18274(.A1(new_n5537_), .A2(new_n18531_), .ZN(new_n18532_));
  XOR2_X1    g18275(.A1(new_n18532_), .A2(\a[50] ), .Z(new_n18533_));
  OAI22_X1   g18276(.A1(new_n6721_), .A2(new_n4316_), .B1(new_n6723_), .B2(new_n4501_), .ZN(new_n18534_));
  NAND2_X1   g18277(.A1(new_n7617_), .A2(\b[42] ), .ZN(new_n18535_));
  AOI21_X1   g18278(.A1(new_n18535_), .A2(new_n18534_), .B(new_n6731_), .ZN(new_n18536_));
  NAND2_X1   g18279(.A1(new_n4500_), .A2(new_n18536_), .ZN(new_n18537_));
  XOR2_X1    g18280(.A1(new_n18537_), .A2(\a[56] ), .Z(new_n18538_));
  OAI21_X1   g18281(.A1(new_n18368_), .A2(new_n18394_), .B(new_n18396_), .ZN(new_n18539_));
  OAI21_X1   g18282(.A1(new_n18375_), .A2(new_n18385_), .B(new_n18387_), .ZN(new_n18540_));
  NOR3_X1    g18283(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n2964_), .ZN(new_n18541_));
  NOR2_X1    g18284(.A1(new_n9364_), .A2(new_n2964_), .ZN(new_n18542_));
  NOR3_X1    g18285(.A1(new_n18542_), .A2(new_n3097_), .A3(new_n8985_), .ZN(new_n18543_));
  NOR2_X1    g18286(.A1(new_n18543_), .A2(new_n18541_), .ZN(new_n18544_));
  NOR2_X1    g18287(.A1(new_n18382_), .A2(new_n18544_), .ZN(new_n18545_));
  INV_X1     g18288(.I(new_n18544_), .ZN(new_n18546_));
  NOR2_X1    g18289(.A1(new_n18546_), .A2(new_n18381_), .ZN(new_n18547_));
  OAI21_X1   g18290(.A1(new_n18545_), .A2(new_n18547_), .B(new_n18540_), .ZN(new_n18548_));
  XOR2_X1    g18291(.A1(new_n18381_), .A2(new_n18544_), .Z(new_n18549_));
  OR2_X2     g18292(.A1(new_n18540_), .A2(new_n18549_), .Z(new_n18550_));
  NAND2_X1   g18293(.A1(new_n18550_), .A2(new_n18548_), .ZN(new_n18551_));
  OAI22_X1   g18294(.A1(new_n3997_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n3845_), .ZN(new_n18552_));
  NAND2_X1   g18295(.A1(new_n8628_), .A2(\b[39] ), .ZN(new_n18553_));
  AOI21_X1   g18296(.A1(new_n18553_), .A2(new_n18552_), .B(new_n7354_), .ZN(new_n18554_));
  NAND2_X1   g18297(.A1(new_n3996_), .A2(new_n18554_), .ZN(new_n18555_));
  XOR2_X1    g18298(.A1(new_n18555_), .A2(\a[59] ), .Z(new_n18556_));
  OAI22_X1   g18299(.A1(new_n3566_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n3408_), .ZN(new_n18557_));
  NAND2_X1   g18300(.A1(new_n9644_), .A2(\b[36] ), .ZN(new_n18558_));
  AOI21_X1   g18301(.A1(new_n18558_), .A2(new_n18557_), .B(new_n8321_), .ZN(new_n18559_));
  NAND2_X1   g18302(.A1(new_n3565_), .A2(new_n18559_), .ZN(new_n18560_));
  XOR2_X1    g18303(.A1(new_n18560_), .A2(\a[62] ), .Z(new_n18561_));
  NOR2_X1    g18304(.A1(new_n18556_), .A2(new_n18561_), .ZN(new_n18562_));
  INV_X1     g18305(.I(new_n18562_), .ZN(new_n18563_));
  NAND2_X1   g18306(.A1(new_n18556_), .A2(new_n18561_), .ZN(new_n18564_));
  NAND2_X1   g18307(.A1(new_n18563_), .A2(new_n18564_), .ZN(new_n18565_));
  XNOR2_X1   g18308(.A1(new_n18556_), .A2(new_n18561_), .ZN(new_n18566_));
  NOR2_X1    g18309(.A1(new_n18566_), .A2(new_n18551_), .ZN(new_n18567_));
  AOI21_X1   g18310(.A1(new_n18551_), .A2(new_n18565_), .B(new_n18567_), .ZN(new_n18568_));
  XOR2_X1    g18311(.A1(new_n18568_), .A2(new_n18539_), .Z(new_n18569_));
  INV_X1     g18312(.I(new_n18539_), .ZN(new_n18570_));
  NOR2_X1    g18313(.A1(new_n18568_), .A2(new_n18570_), .ZN(new_n18571_));
  NAND2_X1   g18314(.A1(new_n18568_), .A2(new_n18570_), .ZN(new_n18572_));
  INV_X1     g18315(.I(new_n18572_), .ZN(new_n18573_));
  OAI21_X1   g18316(.A1(new_n18573_), .A2(new_n18571_), .B(new_n18538_), .ZN(new_n18574_));
  OAI21_X1   g18317(.A1(new_n18538_), .A2(new_n18569_), .B(new_n18574_), .ZN(new_n18575_));
  OAI22_X1   g18318(.A1(new_n5786_), .A2(new_n4997_), .B1(new_n4834_), .B2(new_n5792_), .ZN(new_n18576_));
  NAND2_X1   g18319(.A1(new_n6745_), .A2(\b[45] ), .ZN(new_n18577_));
  AOI21_X1   g18320(.A1(new_n18577_), .A2(new_n18576_), .B(new_n5796_), .ZN(new_n18578_));
  NAND2_X1   g18321(.A1(new_n5004_), .A2(new_n18578_), .ZN(new_n18579_));
  XOR2_X1    g18322(.A1(new_n18579_), .A2(\a[53] ), .Z(new_n18580_));
  NOR2_X1    g18323(.A1(new_n18407_), .A2(new_n18363_), .ZN(new_n18581_));
  NOR2_X1    g18324(.A1(new_n18581_), .A2(new_n18405_), .ZN(new_n18582_));
  XOR2_X1    g18325(.A1(new_n18580_), .A2(new_n18582_), .Z(new_n18583_));
  NOR2_X1    g18326(.A1(new_n18580_), .A2(new_n18582_), .ZN(new_n18584_));
  INV_X1     g18327(.I(new_n18584_), .ZN(new_n18585_));
  NAND2_X1   g18328(.A1(new_n18580_), .A2(new_n18582_), .ZN(new_n18586_));
  AOI21_X1   g18329(.A1(new_n18585_), .A2(new_n18586_), .B(new_n18575_), .ZN(new_n18587_));
  AOI21_X1   g18330(.A1(new_n18575_), .A2(new_n18583_), .B(new_n18587_), .ZN(new_n18588_));
  NAND2_X1   g18331(.A1(new_n18418_), .A2(new_n18420_), .ZN(new_n18589_));
  NAND2_X1   g18332(.A1(new_n18589_), .A2(new_n18417_), .ZN(new_n18590_));
  XOR2_X1    g18333(.A1(new_n18588_), .A2(new_n18590_), .Z(new_n18591_));
  NOR2_X1    g18334(.A1(new_n18591_), .A2(new_n18533_), .ZN(new_n18592_));
  INV_X1     g18335(.I(new_n18533_), .ZN(new_n18593_));
  INV_X1     g18336(.I(new_n18590_), .ZN(new_n18594_));
  NOR2_X1    g18337(.A1(new_n18588_), .A2(new_n18594_), .ZN(new_n18595_));
  INV_X1     g18338(.I(new_n18595_), .ZN(new_n18596_));
  NAND2_X1   g18339(.A1(new_n18588_), .A2(new_n18594_), .ZN(new_n18597_));
  AOI21_X1   g18340(.A1(new_n18596_), .A2(new_n18597_), .B(new_n18593_), .ZN(new_n18598_));
  NOR2_X1    g18341(.A1(new_n18592_), .A2(new_n18598_), .ZN(new_n18599_));
  OAI21_X1   g18342(.A1(new_n18423_), .A2(new_n18433_), .B(new_n18432_), .ZN(new_n18600_));
  INV_X1     g18343(.I(new_n18600_), .ZN(new_n18601_));
  XOR2_X1    g18344(.A1(new_n18599_), .A2(new_n18601_), .Z(new_n18602_));
  NOR2_X1    g18345(.A1(new_n18602_), .A2(new_n18528_), .ZN(new_n18603_));
  INV_X1     g18346(.I(new_n18528_), .ZN(new_n18604_));
  INV_X1     g18347(.I(new_n18599_), .ZN(new_n18605_));
  NOR2_X1    g18348(.A1(new_n18605_), .A2(new_n18601_), .ZN(new_n18606_));
  NOR2_X1    g18349(.A1(new_n18599_), .A2(new_n18600_), .ZN(new_n18607_));
  NOR2_X1    g18350(.A1(new_n18606_), .A2(new_n18607_), .ZN(new_n18608_));
  NOR2_X1    g18351(.A1(new_n18608_), .A2(new_n18604_), .ZN(new_n18609_));
  NOR2_X1    g18352(.A1(new_n18609_), .A2(new_n18603_), .ZN(new_n18610_));
  XNOR2_X1   g18353(.A1(new_n18610_), .A2(new_n18523_), .ZN(new_n18611_));
  NOR2_X1    g18354(.A1(new_n18610_), .A2(new_n18523_), .ZN(new_n18612_));
  NAND2_X1   g18355(.A1(new_n18610_), .A2(new_n18523_), .ZN(new_n18613_));
  INV_X1     g18356(.I(new_n18613_), .ZN(new_n18614_));
  OAI21_X1   g18357(.A1(new_n18614_), .A2(new_n18612_), .B(new_n18521_), .ZN(new_n18615_));
  OAI21_X1   g18358(.A1(new_n18521_), .A2(new_n18611_), .B(new_n18615_), .ZN(new_n18616_));
  OAI22_X1   g18359(.A1(new_n3736_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n3731_), .ZN(new_n18617_));
  NAND2_X1   g18360(.A1(new_n4730_), .A2(\b[57] ), .ZN(new_n18618_));
  AOI21_X1   g18361(.A1(new_n18617_), .A2(new_n18618_), .B(new_n3739_), .ZN(new_n18619_));
  NAND2_X1   g18362(.A1(new_n7895_), .A2(new_n18619_), .ZN(new_n18620_));
  XOR2_X1    g18363(.A1(new_n18620_), .A2(\a[41] ), .Z(new_n18621_));
  INV_X1     g18364(.I(new_n18621_), .ZN(new_n18622_));
  NAND2_X1   g18365(.A1(new_n18459_), .A2(new_n18456_), .ZN(new_n18623_));
  NAND2_X1   g18366(.A1(new_n18623_), .A2(new_n18458_), .ZN(new_n18624_));
  XOR2_X1    g18367(.A1(new_n18624_), .A2(new_n18622_), .Z(new_n18625_));
  NAND2_X1   g18368(.A1(new_n18616_), .A2(new_n18625_), .ZN(new_n18626_));
  AOI21_X1   g18369(.A1(new_n18623_), .A2(new_n18458_), .B(new_n18621_), .ZN(new_n18627_));
  NOR2_X1    g18370(.A1(new_n18624_), .A2(new_n18622_), .ZN(new_n18628_));
  NOR2_X1    g18371(.A1(new_n18628_), .A2(new_n18627_), .ZN(new_n18629_));
  OAI21_X1   g18372(.A1(new_n18616_), .A2(new_n18629_), .B(new_n18626_), .ZN(new_n18630_));
  OAI21_X1   g18373(.A1(new_n18348_), .A2(new_n18462_), .B(new_n18464_), .ZN(new_n18631_));
  AND2_X2    g18374(.A1(new_n18630_), .A2(new_n18631_), .Z(new_n18632_));
  NOR2_X1    g18375(.A1(new_n18630_), .A2(new_n18631_), .ZN(new_n18633_));
  NOR2_X1    g18376(.A1(new_n18632_), .A2(new_n18633_), .ZN(new_n18634_));
  NOR2_X1    g18377(.A1(new_n18634_), .A2(new_n18516_), .ZN(new_n18635_));
  XOR2_X1    g18378(.A1(new_n18630_), .A2(new_n18631_), .Z(new_n18636_));
  AOI21_X1   g18379(.A1(new_n18516_), .A2(new_n18636_), .B(new_n18635_), .ZN(new_n18637_));
  XOR2_X1    g18380(.A1(new_n18637_), .A2(new_n18511_), .Z(new_n18638_));
  XOR2_X1    g18381(.A1(new_n18638_), .A2(\a[35] ), .Z(new_n18639_));
  XNOR2_X1   g18382(.A1(new_n18639_), .A2(new_n18510_), .ZN(new_n18640_));
  XOR2_X1    g18383(.A1(new_n18640_), .A2(new_n18509_), .Z(new_n18641_));
  XOR2_X1    g18384(.A1(new_n18640_), .A2(new_n18509_), .Z(new_n18642_));
  NAND2_X1   g18385(.A1(new_n18506_), .A2(new_n18642_), .ZN(new_n18643_));
  OAI21_X1   g18386(.A1(new_n18506_), .A2(new_n18641_), .B(new_n18643_), .ZN(\f[98] ));
  OAI22_X1   g18387(.A1(new_n3298_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n3293_), .ZN(new_n18645_));
  NAND2_X1   g18388(.A1(new_n4227_), .A2(\b[61] ), .ZN(new_n18646_));
  AOI21_X1   g18389(.A1(new_n18645_), .A2(new_n18646_), .B(new_n3301_), .ZN(new_n18647_));
  NAND2_X1   g18390(.A1(new_n8963_), .A2(new_n18647_), .ZN(new_n18648_));
  XOR2_X1    g18391(.A1(new_n18648_), .A2(\a[38] ), .Z(new_n18649_));
  INV_X1     g18392(.I(new_n18649_), .ZN(new_n18650_));
  INV_X1     g18393(.I(new_n18632_), .ZN(new_n18651_));
  OAI21_X1   g18394(.A1(new_n18516_), .A2(new_n18633_), .B(new_n18651_), .ZN(new_n18652_));
  OAI21_X1   g18395(.A1(new_n18521_), .A2(new_n18612_), .B(new_n18613_), .ZN(new_n18653_));
  INV_X1     g18396(.I(new_n18653_), .ZN(new_n18654_));
  INV_X1     g18397(.I(new_n18607_), .ZN(new_n18655_));
  AOI21_X1   g18398(.A1(new_n18604_), .A2(new_n18655_), .B(new_n18606_), .ZN(new_n18656_));
  OAI22_X1   g18399(.A1(new_n4711_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n4706_), .ZN(new_n18657_));
  NAND2_X1   g18400(.A1(new_n5814_), .A2(\b[52] ), .ZN(new_n18658_));
  AOI21_X1   g18401(.A1(new_n18657_), .A2(new_n18658_), .B(new_n4714_), .ZN(new_n18659_));
  NAND2_X1   g18402(.A1(new_n6237_), .A2(new_n18659_), .ZN(new_n18660_));
  XOR2_X1    g18403(.A1(new_n18660_), .A2(\a[47] ), .Z(new_n18661_));
  AOI21_X1   g18404(.A1(new_n18593_), .A2(new_n18597_), .B(new_n18595_), .ZN(new_n18662_));
  INV_X1     g18405(.I(new_n18538_), .ZN(new_n18663_));
  AOI21_X1   g18406(.A1(new_n18663_), .A2(new_n18572_), .B(new_n18571_), .ZN(new_n18664_));
  INV_X1     g18407(.I(new_n18545_), .ZN(new_n18665_));
  AOI21_X1   g18408(.A1(new_n18540_), .A2(new_n18665_), .B(new_n18547_), .ZN(new_n18666_));
  OAI22_X1   g18409(.A1(new_n3696_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n3566_), .ZN(new_n18667_));
  NAND2_X1   g18410(.A1(new_n9644_), .A2(\b[37] ), .ZN(new_n18668_));
  AOI21_X1   g18411(.A1(new_n18668_), .A2(new_n18667_), .B(new_n8321_), .ZN(new_n18669_));
  NAND2_X1   g18412(.A1(new_n3700_), .A2(new_n18669_), .ZN(new_n18670_));
  XOR2_X1    g18413(.A1(new_n18670_), .A2(\a[62] ), .Z(new_n18671_));
  NOR2_X1    g18414(.A1(new_n8985_), .A2(new_n3247_), .ZN(new_n18672_));
  NOR2_X1    g18415(.A1(new_n9364_), .A2(new_n3097_), .ZN(new_n18673_));
  XNOR2_X1   g18416(.A1(new_n18672_), .A2(new_n18673_), .ZN(new_n18674_));
  XOR2_X1    g18417(.A1(new_n18674_), .A2(\a[35] ), .Z(new_n18675_));
  NOR2_X1    g18418(.A1(new_n18675_), .A2(new_n18544_), .ZN(new_n18676_));
  NOR2_X1    g18419(.A1(new_n18674_), .A2(new_n2836_), .ZN(new_n18677_));
  INV_X1     g18420(.I(new_n18677_), .ZN(new_n18678_));
  NAND2_X1   g18421(.A1(new_n18674_), .A2(new_n2836_), .ZN(new_n18679_));
  AOI21_X1   g18422(.A1(new_n18678_), .A2(new_n18679_), .B(new_n18546_), .ZN(new_n18680_));
  NOR2_X1    g18423(.A1(new_n18676_), .A2(new_n18680_), .ZN(new_n18681_));
  XOR2_X1    g18424(.A1(new_n18671_), .A2(new_n18681_), .Z(new_n18682_));
  NOR2_X1    g18425(.A1(new_n18682_), .A2(new_n18666_), .ZN(new_n18683_));
  OAI21_X1   g18426(.A1(new_n18676_), .A2(new_n18680_), .B(new_n18671_), .ZN(new_n18684_));
  INV_X1     g18427(.I(new_n18671_), .ZN(new_n18685_));
  NAND2_X1   g18428(.A1(new_n18685_), .A2(new_n18681_), .ZN(new_n18686_));
  NAND2_X1   g18429(.A1(new_n18686_), .A2(new_n18684_), .ZN(new_n18687_));
  AOI21_X1   g18430(.A1(new_n18666_), .A2(new_n18687_), .B(new_n18683_), .ZN(new_n18688_));
  OAI22_X1   g18431(.A1(new_n4018_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n3997_), .ZN(new_n18689_));
  NAND2_X1   g18432(.A1(new_n8628_), .A2(\b[40] ), .ZN(new_n18690_));
  AOI21_X1   g18433(.A1(new_n18690_), .A2(new_n18689_), .B(new_n7354_), .ZN(new_n18691_));
  NAND2_X1   g18434(.A1(new_n4017_), .A2(new_n18691_), .ZN(new_n18692_));
  XOR2_X1    g18435(.A1(new_n18692_), .A2(\a[59] ), .Z(new_n18693_));
  NAND2_X1   g18436(.A1(new_n18564_), .A2(new_n18551_), .ZN(new_n18694_));
  NAND2_X1   g18437(.A1(new_n18694_), .A2(new_n18563_), .ZN(new_n18695_));
  XOR2_X1    g18438(.A1(new_n18695_), .A2(new_n18693_), .Z(new_n18696_));
  NOR2_X1    g18439(.A1(new_n18696_), .A2(new_n18688_), .ZN(new_n18697_));
  INV_X1     g18440(.I(new_n18695_), .ZN(new_n18698_));
  NOR2_X1    g18441(.A1(new_n18698_), .A2(new_n18693_), .ZN(new_n18699_));
  INV_X1     g18442(.I(new_n18699_), .ZN(new_n18700_));
  NAND2_X1   g18443(.A1(new_n18698_), .A2(new_n18693_), .ZN(new_n18701_));
  NAND2_X1   g18444(.A1(new_n18700_), .A2(new_n18701_), .ZN(new_n18702_));
  AOI21_X1   g18445(.A1(new_n18688_), .A2(new_n18702_), .B(new_n18697_), .ZN(new_n18703_));
  OAI22_X1   g18446(.A1(new_n6721_), .A2(new_n4501_), .B1(new_n6723_), .B2(new_n4509_), .ZN(new_n18704_));
  NAND2_X1   g18447(.A1(new_n7617_), .A2(\b[43] ), .ZN(new_n18705_));
  AOI21_X1   g18448(.A1(new_n18705_), .A2(new_n18704_), .B(new_n6731_), .ZN(new_n18706_));
  NAND2_X1   g18449(.A1(new_n4513_), .A2(new_n18706_), .ZN(new_n18707_));
  XOR2_X1    g18450(.A1(new_n18707_), .A2(\a[56] ), .Z(new_n18708_));
  XNOR2_X1   g18451(.A1(new_n18703_), .A2(new_n18708_), .ZN(new_n18709_));
  NOR2_X1    g18452(.A1(new_n18709_), .A2(new_n18664_), .ZN(new_n18710_));
  INV_X1     g18453(.I(new_n18664_), .ZN(new_n18711_));
  NOR2_X1    g18454(.A1(new_n18703_), .A2(new_n18708_), .ZN(new_n18712_));
  INV_X1     g18455(.I(new_n18712_), .ZN(new_n18713_));
  NAND2_X1   g18456(.A1(new_n18703_), .A2(new_n18708_), .ZN(new_n18714_));
  AOI21_X1   g18457(.A1(new_n18713_), .A2(new_n18714_), .B(new_n18711_), .ZN(new_n18715_));
  NOR2_X1    g18458(.A1(new_n18710_), .A2(new_n18715_), .ZN(new_n18716_));
  OAI22_X1   g18459(.A1(new_n5786_), .A2(new_n5178_), .B1(new_n4997_), .B2(new_n5792_), .ZN(new_n18717_));
  NAND2_X1   g18460(.A1(new_n6745_), .A2(\b[46] ), .ZN(new_n18718_));
  AOI21_X1   g18461(.A1(new_n18718_), .A2(new_n18717_), .B(new_n5796_), .ZN(new_n18719_));
  NAND2_X1   g18462(.A1(new_n5177_), .A2(new_n18719_), .ZN(new_n18720_));
  XOR2_X1    g18463(.A1(new_n18720_), .A2(\a[53] ), .Z(new_n18721_));
  INV_X1     g18464(.I(new_n18575_), .ZN(new_n18722_));
  AOI21_X1   g18465(.A1(new_n18722_), .A2(new_n18586_), .B(new_n18584_), .ZN(new_n18723_));
  NOR2_X1    g18466(.A1(new_n18723_), .A2(new_n18721_), .ZN(new_n18724_));
  INV_X1     g18467(.I(new_n18724_), .ZN(new_n18725_));
  NAND2_X1   g18468(.A1(new_n18723_), .A2(new_n18721_), .ZN(new_n18726_));
  AOI21_X1   g18469(.A1(new_n18725_), .A2(new_n18726_), .B(new_n18716_), .ZN(new_n18727_));
  XNOR2_X1   g18470(.A1(new_n18723_), .A2(new_n18721_), .ZN(new_n18728_));
  NOR3_X1    g18471(.A1(new_n18728_), .A2(new_n18710_), .A3(new_n18715_), .ZN(new_n18729_));
  NOR2_X1    g18472(.A1(new_n18729_), .A2(new_n18727_), .ZN(new_n18730_));
  OAI22_X1   g18473(.A1(new_n5228_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n5225_), .ZN(new_n18731_));
  NAND2_X1   g18474(.A1(new_n5387_), .A2(\b[49] ), .ZN(new_n18732_));
  AOI21_X1   g18475(.A1(new_n18731_), .A2(new_n18732_), .B(new_n5231_), .ZN(new_n18733_));
  NAND2_X1   g18476(.A1(new_n5741_), .A2(new_n18733_), .ZN(new_n18734_));
  XOR2_X1    g18477(.A1(new_n18734_), .A2(\a[50] ), .Z(new_n18735_));
  XOR2_X1    g18478(.A1(new_n18730_), .A2(new_n18735_), .Z(new_n18736_));
  NOR2_X1    g18479(.A1(new_n18736_), .A2(new_n18662_), .ZN(new_n18737_));
  INV_X1     g18480(.I(new_n18662_), .ZN(new_n18738_));
  INV_X1     g18481(.I(new_n18730_), .ZN(new_n18739_));
  NOR2_X1    g18482(.A1(new_n18739_), .A2(new_n18735_), .ZN(new_n18740_));
  INV_X1     g18483(.I(new_n18740_), .ZN(new_n18741_));
  NAND2_X1   g18484(.A1(new_n18739_), .A2(new_n18735_), .ZN(new_n18742_));
  AOI21_X1   g18485(.A1(new_n18741_), .A2(new_n18742_), .B(new_n18738_), .ZN(new_n18743_));
  NOR2_X1    g18486(.A1(new_n18743_), .A2(new_n18737_), .ZN(new_n18744_));
  XOR2_X1    g18487(.A1(new_n18744_), .A2(new_n18661_), .Z(new_n18745_));
  INV_X1     g18488(.I(new_n18661_), .ZN(new_n18746_));
  NOR2_X1    g18489(.A1(new_n18744_), .A2(new_n18746_), .ZN(new_n18747_));
  NAND2_X1   g18490(.A1(new_n18744_), .A2(new_n18746_), .ZN(new_n18748_));
  INV_X1     g18491(.I(new_n18748_), .ZN(new_n18749_));
  OAI21_X1   g18492(.A1(new_n18749_), .A2(new_n18747_), .B(new_n18656_), .ZN(new_n18750_));
  OAI21_X1   g18493(.A1(new_n18656_), .A2(new_n18745_), .B(new_n18750_), .ZN(new_n18751_));
  OAI22_X1   g18494(.A1(new_n4208_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n4203_), .ZN(new_n18752_));
  NAND2_X1   g18495(.A1(new_n5244_), .A2(\b[55] ), .ZN(new_n18753_));
  AOI21_X1   g18496(.A1(new_n18752_), .A2(new_n18753_), .B(new_n4211_), .ZN(new_n18754_));
  NAND2_X1   g18497(.A1(new_n7308_), .A2(new_n18754_), .ZN(new_n18755_));
  XOR2_X1    g18498(.A1(new_n18755_), .A2(\a[44] ), .Z(new_n18756_));
  XNOR2_X1   g18499(.A1(new_n18751_), .A2(new_n18756_), .ZN(new_n18757_));
  NOR2_X1    g18500(.A1(new_n18757_), .A2(new_n18654_), .ZN(new_n18758_));
  NOR2_X1    g18501(.A1(new_n18751_), .A2(new_n18756_), .ZN(new_n18759_));
  INV_X1     g18502(.I(new_n18759_), .ZN(new_n18760_));
  NAND2_X1   g18503(.A1(new_n18751_), .A2(new_n18756_), .ZN(new_n18761_));
  AOI21_X1   g18504(.A1(new_n18760_), .A2(new_n18761_), .B(new_n18653_), .ZN(new_n18762_));
  NOR2_X1    g18505(.A1(new_n18758_), .A2(new_n18762_), .ZN(new_n18763_));
  OAI22_X1   g18506(.A1(new_n3736_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n3731_), .ZN(new_n18764_));
  NAND2_X1   g18507(.A1(new_n4730_), .A2(\b[58] ), .ZN(new_n18765_));
  AOI21_X1   g18508(.A1(new_n18764_), .A2(new_n18765_), .B(new_n3739_), .ZN(new_n18766_));
  NAND2_X1   g18509(.A1(new_n7929_), .A2(new_n18766_), .ZN(new_n18767_));
  XOR2_X1    g18510(.A1(new_n18767_), .A2(\a[41] ), .Z(new_n18768_));
  NOR2_X1    g18511(.A1(new_n18616_), .A2(new_n18628_), .ZN(new_n18769_));
  NOR2_X1    g18512(.A1(new_n18769_), .A2(new_n18627_), .ZN(new_n18770_));
  NOR2_X1    g18513(.A1(new_n18770_), .A2(new_n18768_), .ZN(new_n18771_));
  NAND2_X1   g18514(.A1(new_n18770_), .A2(new_n18768_), .ZN(new_n18772_));
  INV_X1     g18515(.I(new_n18772_), .ZN(new_n18773_));
  NOR2_X1    g18516(.A1(new_n18773_), .A2(new_n18771_), .ZN(new_n18774_));
  XOR2_X1    g18517(.A1(new_n18770_), .A2(new_n18768_), .Z(new_n18775_));
  NAND2_X1   g18518(.A1(new_n18775_), .A2(new_n18763_), .ZN(new_n18776_));
  OAI21_X1   g18519(.A1(new_n18763_), .A2(new_n18774_), .B(new_n18776_), .ZN(new_n18777_));
  XNOR2_X1   g18520(.A1(new_n18777_), .A2(new_n18652_), .ZN(new_n18778_));
  NAND2_X1   g18521(.A1(new_n18778_), .A2(new_n18650_), .ZN(new_n18779_));
  INV_X1     g18522(.I(new_n18652_), .ZN(new_n18780_));
  NAND2_X1   g18523(.A1(new_n18780_), .A2(new_n18777_), .ZN(new_n18781_));
  NOR2_X1    g18524(.A1(new_n18780_), .A2(new_n18777_), .ZN(new_n18782_));
  INV_X1     g18525(.I(new_n18782_), .ZN(new_n18783_));
  NAND2_X1   g18526(.A1(new_n18783_), .A2(new_n18781_), .ZN(new_n18784_));
  NAND2_X1   g18527(.A1(new_n18784_), .A2(new_n18649_), .ZN(new_n18785_));
  NAND2_X1   g18528(.A1(new_n18785_), .A2(new_n18779_), .ZN(new_n18786_));
  NAND2_X1   g18529(.A1(new_n18637_), .A2(new_n18510_), .ZN(new_n18787_));
  XOR2_X1    g18530(.A1(new_n18511_), .A2(\a[35] ), .Z(new_n18788_));
  NAND2_X1   g18531(.A1(new_n18787_), .A2(new_n18788_), .ZN(new_n18789_));
  OAI21_X1   g18532(.A1(new_n18510_), .A2(new_n18637_), .B(new_n18789_), .ZN(new_n18790_));
  XOR2_X1    g18533(.A1(new_n18786_), .A2(new_n18790_), .Z(new_n18791_));
  NOR2_X1    g18534(.A1(new_n18506_), .A2(new_n18508_), .ZN(new_n18792_));
  XOR2_X1    g18535(.A1(new_n18792_), .A2(new_n18791_), .Z(new_n18793_));
  INV_X1     g18536(.I(new_n18640_), .ZN(new_n18794_));
  XOR2_X1    g18537(.A1(new_n18506_), .A2(new_n18508_), .Z(new_n18795_));
  NAND2_X1   g18538(.A1(new_n18795_), .A2(new_n18794_), .ZN(new_n18796_));
  XOR2_X1    g18539(.A1(new_n18793_), .A2(new_n18796_), .Z(\f[99] ));
  NOR2_X1    g18540(.A1(new_n3447_), .A2(new_n8932_), .ZN(new_n18798_));
  NOR2_X1    g18541(.A1(new_n3293_), .A2(new_n8956_), .ZN(new_n18799_));
  NOR4_X1    g18542(.A1(new_n9323_), .A2(new_n3301_), .A3(new_n18798_), .A4(new_n18799_), .ZN(new_n18800_));
  XOR2_X1    g18543(.A1(new_n18800_), .A2(new_n3288_), .Z(new_n18801_));
  AOI21_X1   g18544(.A1(new_n18763_), .A2(new_n18772_), .B(new_n18771_), .ZN(new_n18802_));
  INV_X1     g18545(.I(new_n18802_), .ZN(new_n18803_));
  OAI22_X1   g18546(.A1(new_n4208_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n4203_), .ZN(new_n18804_));
  NAND2_X1   g18547(.A1(new_n5244_), .A2(\b[56] ), .ZN(new_n18805_));
  AOI21_X1   g18548(.A1(new_n18804_), .A2(new_n18805_), .B(new_n4211_), .ZN(new_n18806_));
  NAND2_X1   g18549(.A1(new_n7559_), .A2(new_n18806_), .ZN(new_n18807_));
  XOR2_X1    g18550(.A1(new_n18807_), .A2(\a[44] ), .Z(new_n18808_));
  OAI22_X1   g18551(.A1(new_n5228_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n5225_), .ZN(new_n18809_));
  NAND2_X1   g18552(.A1(new_n5387_), .A2(\b[50] ), .ZN(new_n18810_));
  AOI21_X1   g18553(.A1(new_n18809_), .A2(new_n18810_), .B(new_n5231_), .ZN(new_n18811_));
  NAND2_X1   g18554(.A1(new_n5954_), .A2(new_n18811_), .ZN(new_n18812_));
  XOR2_X1    g18555(.A1(new_n18812_), .A2(\a[50] ), .Z(new_n18813_));
  OAI22_X1   g18556(.A1(new_n6721_), .A2(new_n4509_), .B1(new_n6723_), .B2(new_n4834_), .ZN(new_n18814_));
  NAND2_X1   g18557(.A1(new_n7617_), .A2(\b[44] ), .ZN(new_n18815_));
  AOI21_X1   g18558(.A1(new_n18815_), .A2(new_n18814_), .B(new_n6731_), .ZN(new_n18816_));
  NAND2_X1   g18559(.A1(new_n4833_), .A2(new_n18816_), .ZN(new_n18817_));
  XOR2_X1    g18560(.A1(new_n18817_), .A2(\a[56] ), .Z(new_n18818_));
  OAI22_X1   g18561(.A1(new_n3845_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n3696_), .ZN(new_n18819_));
  NAND2_X1   g18562(.A1(new_n9644_), .A2(\b[38] ), .ZN(new_n18820_));
  AOI21_X1   g18563(.A1(new_n18820_), .A2(new_n18819_), .B(new_n8321_), .ZN(new_n18821_));
  NAND2_X1   g18564(.A1(new_n3844_), .A2(new_n18821_), .ZN(new_n18822_));
  XOR2_X1    g18565(.A1(new_n18822_), .A2(\a[62] ), .Z(new_n18823_));
  NAND2_X1   g18566(.A1(new_n18679_), .A2(new_n18546_), .ZN(new_n18824_));
  NAND2_X1   g18567(.A1(new_n18824_), .A2(new_n18678_), .ZN(new_n18825_));
  NOR3_X1    g18568(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n3247_), .ZN(new_n18826_));
  NOR2_X1    g18569(.A1(new_n9364_), .A2(new_n3247_), .ZN(new_n18827_));
  NOR3_X1    g18570(.A1(new_n18827_), .A2(new_n3408_), .A3(new_n8985_), .ZN(new_n18828_));
  NOR2_X1    g18571(.A1(new_n18828_), .A2(new_n18826_), .ZN(new_n18829_));
  NOR2_X1    g18572(.A1(new_n18825_), .A2(new_n18829_), .ZN(new_n18830_));
  INV_X1     g18573(.I(new_n18830_), .ZN(new_n18831_));
  NAND2_X1   g18574(.A1(new_n18825_), .A2(new_n18829_), .ZN(new_n18832_));
  AOI21_X1   g18575(.A1(new_n18831_), .A2(new_n18832_), .B(new_n18823_), .ZN(new_n18833_));
  INV_X1     g18576(.I(new_n18829_), .ZN(new_n18834_));
  XOR2_X1    g18577(.A1(new_n18825_), .A2(new_n18834_), .Z(new_n18835_));
  INV_X1     g18578(.I(new_n18835_), .ZN(new_n18836_));
  AOI21_X1   g18579(.A1(new_n18823_), .A2(new_n18836_), .B(new_n18833_), .ZN(new_n18837_));
  INV_X1     g18580(.I(new_n18837_), .ZN(new_n18838_));
  INV_X1     g18581(.I(new_n18666_), .ZN(new_n18839_));
  NAND2_X1   g18582(.A1(new_n18839_), .A2(new_n18684_), .ZN(new_n18840_));
  NAND2_X1   g18583(.A1(new_n18840_), .A2(new_n18686_), .ZN(new_n18841_));
  INV_X1     g18584(.I(new_n18841_), .ZN(new_n18842_));
  OAI22_X1   g18585(.A1(new_n4316_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n4018_), .ZN(new_n18843_));
  NAND2_X1   g18586(.A1(new_n8628_), .A2(\b[41] ), .ZN(new_n18844_));
  AOI21_X1   g18587(.A1(new_n18844_), .A2(new_n18843_), .B(new_n7354_), .ZN(new_n18845_));
  NAND2_X1   g18588(.A1(new_n4320_), .A2(new_n18845_), .ZN(new_n18846_));
  XOR2_X1    g18589(.A1(new_n18846_), .A2(\a[59] ), .Z(new_n18847_));
  NOR2_X1    g18590(.A1(new_n18842_), .A2(new_n18847_), .ZN(new_n18848_));
  INV_X1     g18591(.I(new_n18847_), .ZN(new_n18849_));
  NOR2_X1    g18592(.A1(new_n18849_), .A2(new_n18841_), .ZN(new_n18850_));
  OAI21_X1   g18593(.A1(new_n18850_), .A2(new_n18848_), .B(new_n18838_), .ZN(new_n18851_));
  XNOR2_X1   g18594(.A1(new_n18847_), .A2(new_n18841_), .ZN(new_n18852_));
  NAND2_X1   g18595(.A1(new_n18852_), .A2(new_n18837_), .ZN(new_n18853_));
  NAND2_X1   g18596(.A1(new_n18853_), .A2(new_n18851_), .ZN(new_n18854_));
  INV_X1     g18597(.I(new_n18854_), .ZN(new_n18855_));
  NAND2_X1   g18598(.A1(new_n18701_), .A2(new_n18688_), .ZN(new_n18856_));
  NAND2_X1   g18599(.A1(new_n18856_), .A2(new_n18700_), .ZN(new_n18857_));
  INV_X1     g18600(.I(new_n18857_), .ZN(new_n18858_));
  NOR2_X1    g18601(.A1(new_n18858_), .A2(new_n18855_), .ZN(new_n18859_));
  NOR2_X1    g18602(.A1(new_n18857_), .A2(new_n18854_), .ZN(new_n18860_));
  NOR2_X1    g18603(.A1(new_n18859_), .A2(new_n18860_), .ZN(new_n18861_));
  NOR2_X1    g18604(.A1(new_n18861_), .A2(new_n18818_), .ZN(new_n18862_));
  INV_X1     g18605(.I(new_n18818_), .ZN(new_n18863_));
  XOR2_X1    g18606(.A1(new_n18857_), .A2(new_n18855_), .Z(new_n18864_));
  NOR2_X1    g18607(.A1(new_n18864_), .A2(new_n18863_), .ZN(new_n18865_));
  NOR2_X1    g18608(.A1(new_n18862_), .A2(new_n18865_), .ZN(new_n18866_));
  NAND2_X1   g18609(.A1(new_n18714_), .A2(new_n18711_), .ZN(new_n18867_));
  NAND2_X1   g18610(.A1(new_n18867_), .A2(new_n18713_), .ZN(new_n18868_));
  INV_X1     g18611(.I(new_n18868_), .ZN(new_n18869_));
  OAI22_X1   g18612(.A1(new_n5786_), .A2(new_n5197_), .B1(new_n5178_), .B2(new_n5792_), .ZN(new_n18870_));
  NAND2_X1   g18613(.A1(new_n6745_), .A2(\b[47] ), .ZN(new_n18871_));
  AOI21_X1   g18614(.A1(new_n18871_), .A2(new_n18870_), .B(new_n5796_), .ZN(new_n18872_));
  NAND2_X1   g18615(.A1(new_n5196_), .A2(new_n18872_), .ZN(new_n18873_));
  XOR2_X1    g18616(.A1(new_n18873_), .A2(\a[53] ), .Z(new_n18874_));
  NOR2_X1    g18617(.A1(new_n18869_), .A2(new_n18874_), .ZN(new_n18875_));
  INV_X1     g18618(.I(new_n18874_), .ZN(new_n18876_));
  NOR2_X1    g18619(.A1(new_n18868_), .A2(new_n18876_), .ZN(new_n18877_));
  NOR2_X1    g18620(.A1(new_n18875_), .A2(new_n18877_), .ZN(new_n18878_));
  NOR2_X1    g18621(.A1(new_n18878_), .A2(new_n18866_), .ZN(new_n18879_));
  INV_X1     g18622(.I(new_n18866_), .ZN(new_n18880_));
  XOR2_X1    g18623(.A1(new_n18868_), .A2(new_n18874_), .Z(new_n18881_));
  NOR2_X1    g18624(.A1(new_n18881_), .A2(new_n18880_), .ZN(new_n18882_));
  NOR2_X1    g18625(.A1(new_n18879_), .A2(new_n18882_), .ZN(new_n18883_));
  AOI21_X1   g18626(.A1(new_n18716_), .A2(new_n18726_), .B(new_n18724_), .ZN(new_n18884_));
  NOR2_X1    g18627(.A1(new_n18883_), .A2(new_n18884_), .ZN(new_n18885_));
  INV_X1     g18628(.I(new_n18885_), .ZN(new_n18886_));
  NAND2_X1   g18629(.A1(new_n18883_), .A2(new_n18884_), .ZN(new_n18887_));
  AOI21_X1   g18630(.A1(new_n18886_), .A2(new_n18887_), .B(new_n18813_), .ZN(new_n18888_));
  INV_X1     g18631(.I(new_n18813_), .ZN(new_n18889_));
  XNOR2_X1   g18632(.A1(new_n18883_), .A2(new_n18884_), .ZN(new_n18890_));
  NOR2_X1    g18633(.A1(new_n18890_), .A2(new_n18889_), .ZN(new_n18891_));
  NAND2_X1   g18634(.A1(new_n18742_), .A2(new_n18738_), .ZN(new_n18892_));
  OAI22_X1   g18635(.A1(new_n4711_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n4706_), .ZN(new_n18893_));
  NAND2_X1   g18636(.A1(new_n5814_), .A2(\b[53] ), .ZN(new_n18894_));
  AOI21_X1   g18637(.A1(new_n18893_), .A2(new_n18894_), .B(new_n4714_), .ZN(new_n18895_));
  NAND2_X1   g18638(.A1(new_n6471_), .A2(new_n18895_), .ZN(new_n18896_));
  XOR2_X1    g18639(.A1(new_n18896_), .A2(\a[47] ), .Z(new_n18897_));
  AOI21_X1   g18640(.A1(new_n18892_), .A2(new_n18741_), .B(new_n18897_), .ZN(new_n18898_));
  NAND2_X1   g18641(.A1(new_n18892_), .A2(new_n18741_), .ZN(new_n18899_));
  INV_X1     g18642(.I(new_n18897_), .ZN(new_n18900_));
  NOR2_X1    g18643(.A1(new_n18899_), .A2(new_n18900_), .ZN(new_n18901_));
  OAI22_X1   g18644(.A1(new_n18901_), .A2(new_n18898_), .B1(new_n18888_), .B2(new_n18891_), .ZN(new_n18902_));
  NOR2_X1    g18645(.A1(new_n18891_), .A2(new_n18888_), .ZN(new_n18903_));
  XOR2_X1    g18646(.A1(new_n18899_), .A2(new_n18900_), .Z(new_n18904_));
  NAND2_X1   g18647(.A1(new_n18904_), .A2(new_n18903_), .ZN(new_n18905_));
  NAND2_X1   g18648(.A1(new_n18905_), .A2(new_n18902_), .ZN(new_n18906_));
  INV_X1     g18649(.I(new_n18906_), .ZN(new_n18907_));
  OAI21_X1   g18650(.A1(new_n18656_), .A2(new_n18747_), .B(new_n18748_), .ZN(new_n18908_));
  INV_X1     g18651(.I(new_n18908_), .ZN(new_n18909_));
  NOR2_X1    g18652(.A1(new_n18907_), .A2(new_n18909_), .ZN(new_n18910_));
  NOR2_X1    g18653(.A1(new_n18906_), .A2(new_n18908_), .ZN(new_n18911_));
  NOR2_X1    g18654(.A1(new_n18910_), .A2(new_n18911_), .ZN(new_n18912_));
  NOR2_X1    g18655(.A1(new_n18912_), .A2(new_n18808_), .ZN(new_n18913_));
  INV_X1     g18656(.I(new_n18808_), .ZN(new_n18914_));
  XOR2_X1    g18657(.A1(new_n18906_), .A2(new_n18909_), .Z(new_n18915_));
  NOR2_X1    g18658(.A1(new_n18915_), .A2(new_n18914_), .ZN(new_n18916_));
  NOR2_X1    g18659(.A1(new_n18913_), .A2(new_n18916_), .ZN(new_n18917_));
  NAND2_X1   g18660(.A1(new_n18761_), .A2(new_n18653_), .ZN(new_n18918_));
  NAND2_X1   g18661(.A1(new_n18918_), .A2(new_n18760_), .ZN(new_n18919_));
  OAI22_X1   g18662(.A1(new_n3736_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n3731_), .ZN(new_n18920_));
  NAND2_X1   g18663(.A1(new_n4730_), .A2(\b[59] ), .ZN(new_n18921_));
  AOI21_X1   g18664(.A1(new_n18920_), .A2(new_n18921_), .B(new_n3739_), .ZN(new_n18922_));
  NAND2_X1   g18665(.A1(new_n8550_), .A2(new_n18922_), .ZN(new_n18923_));
  XOR2_X1    g18666(.A1(new_n18923_), .A2(\a[41] ), .Z(new_n18924_));
  XOR2_X1    g18667(.A1(new_n18919_), .A2(new_n18924_), .Z(new_n18925_));
  NOR2_X1    g18668(.A1(new_n18925_), .A2(new_n18917_), .ZN(new_n18926_));
  INV_X1     g18669(.I(new_n18917_), .ZN(new_n18927_));
  INV_X1     g18670(.I(new_n18919_), .ZN(new_n18928_));
  NOR2_X1    g18671(.A1(new_n18928_), .A2(new_n18924_), .ZN(new_n18929_));
  INV_X1     g18672(.I(new_n18929_), .ZN(new_n18930_));
  NAND2_X1   g18673(.A1(new_n18928_), .A2(new_n18924_), .ZN(new_n18931_));
  AOI21_X1   g18674(.A1(new_n18930_), .A2(new_n18931_), .B(new_n18927_), .ZN(new_n18932_));
  NOR2_X1    g18675(.A1(new_n18932_), .A2(new_n18926_), .ZN(new_n18933_));
  NOR2_X1    g18676(.A1(new_n18933_), .A2(new_n18803_), .ZN(new_n18934_));
  INV_X1     g18677(.I(new_n18933_), .ZN(new_n18935_));
  NOR2_X1    g18678(.A1(new_n18935_), .A2(new_n18802_), .ZN(new_n18936_));
  NOR2_X1    g18679(.A1(new_n18936_), .A2(new_n18934_), .ZN(new_n18937_));
  NOR2_X1    g18680(.A1(new_n18937_), .A2(new_n18801_), .ZN(new_n18938_));
  INV_X1     g18681(.I(new_n18801_), .ZN(new_n18939_));
  XOR2_X1    g18682(.A1(new_n18933_), .A2(new_n18802_), .Z(new_n18940_));
  NOR2_X1    g18683(.A1(new_n18940_), .A2(new_n18939_), .ZN(new_n18941_));
  NOR2_X1    g18684(.A1(new_n18938_), .A2(new_n18941_), .ZN(new_n18942_));
  AOI21_X1   g18685(.A1(new_n18650_), .A2(new_n18781_), .B(new_n18782_), .ZN(new_n18943_));
  INV_X1     g18686(.I(new_n18943_), .ZN(new_n18944_));
  NAND2_X1   g18687(.A1(new_n18794_), .A2(new_n18791_), .ZN(new_n18945_));
  INV_X1     g18688(.I(new_n18945_), .ZN(new_n18946_));
  NOR3_X1    g18689(.A1(new_n18506_), .A2(new_n18508_), .A3(new_n18946_), .ZN(new_n18947_));
  AOI21_X1   g18690(.A1(new_n18785_), .A2(new_n18779_), .B(new_n18790_), .ZN(new_n18948_));
  NOR2_X1    g18691(.A1(new_n18947_), .A2(new_n18948_), .ZN(new_n18949_));
  XOR2_X1    g18692(.A1(new_n18949_), .A2(new_n18944_), .Z(new_n18950_));
  XOR2_X1    g18693(.A1(new_n18950_), .A2(new_n18942_), .Z(\f[100] ));
  NOR2_X1    g18694(.A1(new_n18942_), .A2(new_n18944_), .ZN(new_n18952_));
  INV_X1     g18695(.I(new_n18952_), .ZN(new_n18953_));
  XOR2_X1    g18696(.A1(new_n18942_), .A2(new_n18944_), .Z(new_n18954_));
  NOR2_X1    g18697(.A1(new_n18954_), .A2(new_n18948_), .ZN(new_n18955_));
  INV_X1     g18698(.I(new_n18955_), .ZN(new_n18956_));
  OAI21_X1   g18699(.A1(new_n18947_), .A2(new_n18956_), .B(new_n18953_), .ZN(new_n18957_));
  INV_X1     g18700(.I(new_n18934_), .ZN(new_n18958_));
  AOI21_X1   g18701(.A1(new_n18939_), .A2(new_n18958_), .B(new_n18936_), .ZN(new_n18959_));
  AOI21_X1   g18702(.A1(new_n18927_), .A2(new_n18931_), .B(new_n18929_), .ZN(new_n18960_));
  OAI22_X1   g18703(.A1(new_n9595_), .A2(new_n3301_), .B1(new_n8956_), .B2(new_n3447_), .ZN(new_n18961_));
  OAI22_X1   g18704(.A1(new_n3736_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n3731_), .ZN(new_n18962_));
  NAND2_X1   g18705(.A1(new_n4730_), .A2(\b[60] ), .ZN(new_n18963_));
  AOI21_X1   g18706(.A1(new_n18962_), .A2(new_n18963_), .B(new_n3739_), .ZN(new_n18964_));
  NAND2_X1   g18707(.A1(new_n8935_), .A2(new_n18964_), .ZN(new_n18965_));
  XOR2_X1    g18708(.A1(new_n18965_), .A2(\a[41] ), .Z(new_n18966_));
  OAI22_X1   g18709(.A1(new_n4711_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n4706_), .ZN(new_n18967_));
  NAND2_X1   g18710(.A1(new_n5814_), .A2(\b[54] ), .ZN(new_n18968_));
  AOI21_X1   g18711(.A1(new_n18967_), .A2(new_n18968_), .B(new_n4714_), .ZN(new_n18969_));
  NAND2_X1   g18712(.A1(new_n6994_), .A2(new_n18969_), .ZN(new_n18970_));
  XOR2_X1    g18713(.A1(new_n18970_), .A2(\a[47] ), .Z(new_n18971_));
  INV_X1     g18714(.I(new_n18971_), .ZN(new_n18972_));
  NAND2_X1   g18715(.A1(new_n18887_), .A2(new_n18889_), .ZN(new_n18973_));
  NAND2_X1   g18716(.A1(new_n18973_), .A2(new_n18886_), .ZN(new_n18974_));
  OAI22_X1   g18717(.A1(new_n5228_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n5225_), .ZN(new_n18975_));
  NAND2_X1   g18718(.A1(new_n5387_), .A2(\b[51] ), .ZN(new_n18976_));
  AOI21_X1   g18719(.A1(new_n18975_), .A2(new_n18976_), .B(new_n5231_), .ZN(new_n18977_));
  NAND2_X1   g18720(.A1(new_n6219_), .A2(new_n18977_), .ZN(new_n18978_));
  XOR2_X1    g18721(.A1(new_n18978_), .A2(\a[50] ), .Z(new_n18979_));
  INV_X1     g18722(.I(new_n18979_), .ZN(new_n18980_));
  OAI22_X1   g18723(.A1(new_n5786_), .A2(new_n5538_), .B1(new_n5197_), .B2(new_n5792_), .ZN(new_n18981_));
  NAND2_X1   g18724(.A1(new_n6745_), .A2(\b[48] ), .ZN(new_n18982_));
  AOI21_X1   g18725(.A1(new_n18982_), .A2(new_n18981_), .B(new_n5796_), .ZN(new_n18983_));
  NAND2_X1   g18726(.A1(new_n5537_), .A2(new_n18983_), .ZN(new_n18984_));
  XOR2_X1    g18727(.A1(new_n18984_), .A2(\a[53] ), .Z(new_n18985_));
  OAI21_X1   g18728(.A1(new_n18823_), .A2(new_n18830_), .B(new_n18832_), .ZN(new_n18986_));
  NOR3_X1    g18729(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n3408_), .ZN(new_n18987_));
  NOR2_X1    g18730(.A1(new_n9364_), .A2(new_n3408_), .ZN(new_n18988_));
  NOR3_X1    g18731(.A1(new_n18988_), .A2(new_n3566_), .A3(new_n8985_), .ZN(new_n18989_));
  NOR2_X1    g18732(.A1(new_n18989_), .A2(new_n18987_), .ZN(new_n18990_));
  NOR2_X1    g18733(.A1(new_n18834_), .A2(new_n18990_), .ZN(new_n18991_));
  INV_X1     g18734(.I(new_n18990_), .ZN(new_n18992_));
  NOR2_X1    g18735(.A1(new_n18992_), .A2(new_n18829_), .ZN(new_n18993_));
  OAI21_X1   g18736(.A1(new_n18991_), .A2(new_n18993_), .B(new_n18986_), .ZN(new_n18994_));
  XOR2_X1    g18737(.A1(new_n18829_), .A2(new_n18990_), .Z(new_n18995_));
  OR2_X2     g18738(.A1(new_n18986_), .A2(new_n18995_), .Z(new_n18996_));
  NAND2_X1   g18739(.A1(new_n18996_), .A2(new_n18994_), .ZN(new_n18997_));
  INV_X1     g18740(.I(new_n18997_), .ZN(new_n18998_));
  OAI22_X1   g18741(.A1(new_n4501_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n4316_), .ZN(new_n18999_));
  NAND2_X1   g18742(.A1(new_n8628_), .A2(\b[42] ), .ZN(new_n19000_));
  AOI21_X1   g18743(.A1(new_n19000_), .A2(new_n18999_), .B(new_n7354_), .ZN(new_n19001_));
  NAND2_X1   g18744(.A1(new_n4500_), .A2(new_n19001_), .ZN(new_n19002_));
  XOR2_X1    g18745(.A1(new_n19002_), .A2(\a[59] ), .Z(new_n19003_));
  OAI22_X1   g18746(.A1(new_n3997_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n3845_), .ZN(new_n19004_));
  NAND2_X1   g18747(.A1(new_n9644_), .A2(\b[39] ), .ZN(new_n19005_));
  AOI21_X1   g18748(.A1(new_n19005_), .A2(new_n19004_), .B(new_n8321_), .ZN(new_n19006_));
  NAND2_X1   g18749(.A1(new_n3996_), .A2(new_n19006_), .ZN(new_n19007_));
  XOR2_X1    g18750(.A1(new_n19007_), .A2(\a[62] ), .Z(new_n19008_));
  NOR2_X1    g18751(.A1(new_n19003_), .A2(new_n19008_), .ZN(new_n19009_));
  INV_X1     g18752(.I(new_n19009_), .ZN(new_n19010_));
  NAND2_X1   g18753(.A1(new_n19003_), .A2(new_n19008_), .ZN(new_n19011_));
  AOI21_X1   g18754(.A1(new_n19010_), .A2(new_n19011_), .B(new_n18998_), .ZN(new_n19012_));
  XNOR2_X1   g18755(.A1(new_n19003_), .A2(new_n19008_), .ZN(new_n19013_));
  NOR2_X1    g18756(.A1(new_n19013_), .A2(new_n18997_), .ZN(new_n19014_));
  NOR2_X1    g18757(.A1(new_n19014_), .A2(new_n19012_), .ZN(new_n19015_));
  INV_X1     g18758(.I(new_n19015_), .ZN(new_n19016_));
  OAI22_X1   g18759(.A1(new_n6721_), .A2(new_n4834_), .B1(new_n6723_), .B2(new_n4997_), .ZN(new_n19017_));
  NAND2_X1   g18760(.A1(new_n7617_), .A2(\b[45] ), .ZN(new_n19018_));
  AOI21_X1   g18761(.A1(new_n19018_), .A2(new_n19017_), .B(new_n6731_), .ZN(new_n19019_));
  NAND2_X1   g18762(.A1(new_n5004_), .A2(new_n19019_), .ZN(new_n19020_));
  XOR2_X1    g18763(.A1(new_n19020_), .A2(\a[56] ), .Z(new_n19021_));
  NOR2_X1    g18764(.A1(new_n18850_), .A2(new_n18837_), .ZN(new_n19022_));
  NOR2_X1    g18765(.A1(new_n19022_), .A2(new_n18848_), .ZN(new_n19023_));
  NOR2_X1    g18766(.A1(new_n19021_), .A2(new_n19023_), .ZN(new_n19024_));
  INV_X1     g18767(.I(new_n19024_), .ZN(new_n19025_));
  NAND2_X1   g18768(.A1(new_n19021_), .A2(new_n19023_), .ZN(new_n19026_));
  NAND2_X1   g18769(.A1(new_n19025_), .A2(new_n19026_), .ZN(new_n19027_));
  NAND2_X1   g18770(.A1(new_n19027_), .A2(new_n19016_), .ZN(new_n19028_));
  XOR2_X1    g18771(.A1(new_n19021_), .A2(new_n19023_), .Z(new_n19029_));
  NAND2_X1   g18772(.A1(new_n19029_), .A2(new_n19015_), .ZN(new_n19030_));
  NAND2_X1   g18773(.A1(new_n19028_), .A2(new_n19030_), .ZN(new_n19031_));
  NOR2_X1    g18774(.A1(new_n18860_), .A2(new_n18818_), .ZN(new_n19032_));
  NOR2_X1    g18775(.A1(new_n19032_), .A2(new_n18859_), .ZN(new_n19033_));
  XOR2_X1    g18776(.A1(new_n19031_), .A2(new_n19033_), .Z(new_n19034_));
  NOR2_X1    g18777(.A1(new_n19034_), .A2(new_n18985_), .ZN(new_n19035_));
  INV_X1     g18778(.I(new_n18985_), .ZN(new_n19036_));
  INV_X1     g18779(.I(new_n19031_), .ZN(new_n19037_));
  NOR2_X1    g18780(.A1(new_n19037_), .A2(new_n19033_), .ZN(new_n19038_));
  INV_X1     g18781(.I(new_n19038_), .ZN(new_n19039_));
  NAND2_X1   g18782(.A1(new_n19037_), .A2(new_n19033_), .ZN(new_n19040_));
  AOI21_X1   g18783(.A1(new_n19039_), .A2(new_n19040_), .B(new_n19036_), .ZN(new_n19041_));
  NOR2_X1    g18784(.A1(new_n19041_), .A2(new_n19035_), .ZN(new_n19042_));
  NOR2_X1    g18785(.A1(new_n18877_), .A2(new_n18866_), .ZN(new_n19043_));
  NOR2_X1    g18786(.A1(new_n19043_), .A2(new_n18875_), .ZN(new_n19044_));
  XNOR2_X1   g18787(.A1(new_n19042_), .A2(new_n19044_), .ZN(new_n19045_));
  INV_X1     g18788(.I(new_n19042_), .ZN(new_n19046_));
  NOR2_X1    g18789(.A1(new_n19046_), .A2(new_n19044_), .ZN(new_n19047_));
  INV_X1     g18790(.I(new_n19047_), .ZN(new_n19048_));
  NAND2_X1   g18791(.A1(new_n19046_), .A2(new_n19044_), .ZN(new_n19049_));
  AOI21_X1   g18792(.A1(new_n19048_), .A2(new_n19049_), .B(new_n18980_), .ZN(new_n19050_));
  AOI21_X1   g18793(.A1(new_n18980_), .A2(new_n19045_), .B(new_n19050_), .ZN(new_n19051_));
  XOR2_X1    g18794(.A1(new_n19051_), .A2(new_n18974_), .Z(new_n19052_));
  NAND2_X1   g18795(.A1(new_n19052_), .A2(new_n18972_), .ZN(new_n19053_));
  NOR2_X1    g18796(.A1(new_n19051_), .A2(new_n18974_), .ZN(new_n19054_));
  NAND2_X1   g18797(.A1(new_n19051_), .A2(new_n18974_), .ZN(new_n19055_));
  INV_X1     g18798(.I(new_n19055_), .ZN(new_n19056_));
  OAI21_X1   g18799(.A1(new_n19056_), .A2(new_n19054_), .B(new_n18971_), .ZN(new_n19057_));
  NAND2_X1   g18800(.A1(new_n19053_), .A2(new_n19057_), .ZN(new_n19058_));
  OAI22_X1   g18801(.A1(new_n4208_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n4203_), .ZN(new_n19059_));
  NAND2_X1   g18802(.A1(new_n5244_), .A2(\b[57] ), .ZN(new_n19060_));
  AOI21_X1   g18803(.A1(new_n19059_), .A2(new_n19060_), .B(new_n4211_), .ZN(new_n19061_));
  NAND2_X1   g18804(.A1(new_n7895_), .A2(new_n19061_), .ZN(new_n19062_));
  XOR2_X1    g18805(.A1(new_n19062_), .A2(\a[44] ), .Z(new_n19063_));
  NOR2_X1    g18806(.A1(new_n18901_), .A2(new_n18903_), .ZN(new_n19064_));
  NOR2_X1    g18807(.A1(new_n19064_), .A2(new_n18898_), .ZN(new_n19065_));
  XOR2_X1    g18808(.A1(new_n19065_), .A2(new_n19063_), .Z(new_n19066_));
  NAND2_X1   g18809(.A1(new_n19066_), .A2(new_n19058_), .ZN(new_n19067_));
  INV_X1     g18810(.I(new_n19058_), .ZN(new_n19068_));
  NOR2_X1    g18811(.A1(new_n19065_), .A2(new_n19063_), .ZN(new_n19069_));
  NAND2_X1   g18812(.A1(new_n19065_), .A2(new_n19063_), .ZN(new_n19070_));
  INV_X1     g18813(.I(new_n19070_), .ZN(new_n19071_));
  OAI21_X1   g18814(.A1(new_n19069_), .A2(new_n19071_), .B(new_n19068_), .ZN(new_n19072_));
  NAND2_X1   g18815(.A1(new_n19072_), .A2(new_n19067_), .ZN(new_n19073_));
  INV_X1     g18816(.I(new_n19073_), .ZN(new_n19074_));
  NOR2_X1    g18817(.A1(new_n18911_), .A2(new_n18808_), .ZN(new_n19075_));
  NOR2_X1    g18818(.A1(new_n19075_), .A2(new_n18910_), .ZN(new_n19076_));
  NOR2_X1    g18819(.A1(new_n19074_), .A2(new_n19076_), .ZN(new_n19077_));
  INV_X1     g18820(.I(new_n19077_), .ZN(new_n19078_));
  NAND2_X1   g18821(.A1(new_n19074_), .A2(new_n19076_), .ZN(new_n19079_));
  AOI21_X1   g18822(.A1(new_n19078_), .A2(new_n19079_), .B(new_n18966_), .ZN(new_n19080_));
  XNOR2_X1   g18823(.A1(new_n19073_), .A2(new_n19076_), .ZN(new_n19081_));
  AOI21_X1   g18824(.A1(new_n18966_), .A2(new_n19081_), .B(new_n19080_), .ZN(new_n19082_));
  XOR2_X1    g18825(.A1(new_n19082_), .A2(new_n18961_), .Z(new_n19083_));
  XOR2_X1    g18826(.A1(new_n19083_), .A2(\a[38] ), .Z(new_n19084_));
  XNOR2_X1   g18827(.A1(new_n19084_), .A2(new_n18960_), .ZN(new_n19085_));
  XOR2_X1    g18828(.A1(new_n19085_), .A2(new_n18959_), .Z(new_n19086_));
  NAND2_X1   g18829(.A1(new_n18957_), .A2(new_n19086_), .ZN(new_n19087_));
  XOR2_X1    g18830(.A1(new_n19085_), .A2(new_n18959_), .Z(new_n19088_));
  OAI21_X1   g18831(.A1(new_n18957_), .A2(new_n19088_), .B(new_n19087_), .ZN(\f[101] ));
  OAI22_X1   g18832(.A1(new_n3736_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n3731_), .ZN(new_n19090_));
  NAND2_X1   g18833(.A1(new_n4730_), .A2(\b[61] ), .ZN(new_n19091_));
  AOI21_X1   g18834(.A1(new_n19090_), .A2(new_n19091_), .B(new_n3739_), .ZN(new_n19092_));
  NAND2_X1   g18835(.A1(new_n8963_), .A2(new_n19092_), .ZN(new_n19093_));
  XOR2_X1    g18836(.A1(new_n19093_), .A2(\a[41] ), .Z(new_n19094_));
  INV_X1     g18837(.I(new_n19094_), .ZN(new_n19095_));
  INV_X1     g18838(.I(new_n18966_), .ZN(new_n19096_));
  AOI21_X1   g18839(.A1(new_n19096_), .A2(new_n19079_), .B(new_n19077_), .ZN(new_n19097_));
  OAI21_X1   g18840(.A1(new_n18971_), .A2(new_n19054_), .B(new_n19055_), .ZN(new_n19098_));
  AOI21_X1   g18841(.A1(new_n18980_), .A2(new_n19049_), .B(new_n19047_), .ZN(new_n19099_));
  OAI22_X1   g18842(.A1(new_n5228_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n5225_), .ZN(new_n19100_));
  NAND2_X1   g18843(.A1(new_n5387_), .A2(\b[52] ), .ZN(new_n19101_));
  AOI21_X1   g18844(.A1(new_n19100_), .A2(new_n19101_), .B(new_n5231_), .ZN(new_n19102_));
  NAND2_X1   g18845(.A1(new_n6237_), .A2(new_n19102_), .ZN(new_n19103_));
  XOR2_X1    g18846(.A1(new_n19103_), .A2(\a[50] ), .Z(new_n19104_));
  NAND2_X1   g18847(.A1(new_n19040_), .A2(new_n19036_), .ZN(new_n19105_));
  NAND2_X1   g18848(.A1(new_n19105_), .A2(new_n19039_), .ZN(new_n19106_));
  INV_X1     g18849(.I(new_n18993_), .ZN(new_n19107_));
  AOI21_X1   g18850(.A1(new_n18986_), .A2(new_n19107_), .B(new_n18991_), .ZN(new_n19108_));
  OAI22_X1   g18851(.A1(new_n4018_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n3997_), .ZN(new_n19109_));
  NAND2_X1   g18852(.A1(new_n9644_), .A2(\b[40] ), .ZN(new_n19110_));
  AOI21_X1   g18853(.A1(new_n19110_), .A2(new_n19109_), .B(new_n8321_), .ZN(new_n19111_));
  NAND2_X1   g18854(.A1(new_n4017_), .A2(new_n19111_), .ZN(new_n19112_));
  XOR2_X1    g18855(.A1(new_n19112_), .A2(\a[62] ), .Z(new_n19113_));
  INV_X1     g18856(.I(new_n19113_), .ZN(new_n19114_));
  NOR2_X1    g18857(.A1(new_n8985_), .A2(new_n3696_), .ZN(new_n19115_));
  NOR2_X1    g18858(.A1(new_n9364_), .A2(new_n3566_), .ZN(new_n19116_));
  XNOR2_X1   g18859(.A1(new_n19115_), .A2(new_n19116_), .ZN(new_n19117_));
  XOR2_X1    g18860(.A1(new_n19117_), .A2(\a[38] ), .Z(new_n19118_));
  NOR2_X1    g18861(.A1(new_n19118_), .A2(new_n18829_), .ZN(new_n19119_));
  NOR2_X1    g18862(.A1(new_n19117_), .A2(new_n3288_), .ZN(new_n19120_));
  INV_X1     g18863(.I(new_n19120_), .ZN(new_n19121_));
  NAND2_X1   g18864(.A1(new_n19117_), .A2(new_n3288_), .ZN(new_n19122_));
  AOI21_X1   g18865(.A1(new_n19121_), .A2(new_n19122_), .B(new_n18834_), .ZN(new_n19123_));
  NOR2_X1    g18866(.A1(new_n19119_), .A2(new_n19123_), .ZN(new_n19124_));
  NOR2_X1    g18867(.A1(new_n19114_), .A2(new_n19124_), .ZN(new_n19125_));
  INV_X1     g18868(.I(new_n19125_), .ZN(new_n19126_));
  NAND2_X1   g18869(.A1(new_n19114_), .A2(new_n19124_), .ZN(new_n19127_));
  AOI21_X1   g18870(.A1(new_n19126_), .A2(new_n19127_), .B(new_n19108_), .ZN(new_n19128_));
  XNOR2_X1   g18871(.A1(new_n19113_), .A2(new_n19124_), .ZN(new_n19129_));
  AOI21_X1   g18872(.A1(new_n19129_), .A2(new_n19108_), .B(new_n19128_), .ZN(new_n19130_));
  INV_X1     g18873(.I(new_n19130_), .ZN(new_n19131_));
  NAND2_X1   g18874(.A1(new_n19011_), .A2(new_n18997_), .ZN(new_n19132_));
  OAI22_X1   g18875(.A1(new_n4509_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n4501_), .ZN(new_n19133_));
  NAND2_X1   g18876(.A1(new_n8628_), .A2(\b[43] ), .ZN(new_n19134_));
  AOI21_X1   g18877(.A1(new_n19134_), .A2(new_n19133_), .B(new_n7354_), .ZN(new_n19135_));
  NAND2_X1   g18878(.A1(new_n4513_), .A2(new_n19135_), .ZN(new_n19136_));
  XOR2_X1    g18879(.A1(new_n19136_), .A2(\a[59] ), .Z(new_n19137_));
  AOI21_X1   g18880(.A1(new_n19132_), .A2(new_n19010_), .B(new_n19137_), .ZN(new_n19138_));
  NAND2_X1   g18881(.A1(new_n19132_), .A2(new_n19010_), .ZN(new_n19139_));
  INV_X1     g18882(.I(new_n19137_), .ZN(new_n19140_));
  NOR2_X1    g18883(.A1(new_n19139_), .A2(new_n19140_), .ZN(new_n19141_));
  OAI21_X1   g18884(.A1(new_n19141_), .A2(new_n19138_), .B(new_n19131_), .ZN(new_n19142_));
  XOR2_X1    g18885(.A1(new_n19139_), .A2(new_n19140_), .Z(new_n19143_));
  NAND2_X1   g18886(.A1(new_n19143_), .A2(new_n19130_), .ZN(new_n19144_));
  NAND2_X1   g18887(.A1(new_n19144_), .A2(new_n19142_), .ZN(new_n19145_));
  INV_X1     g18888(.I(new_n19145_), .ZN(new_n19146_));
  OAI22_X1   g18889(.A1(new_n6721_), .A2(new_n4997_), .B1(new_n6723_), .B2(new_n5178_), .ZN(new_n19147_));
  NAND2_X1   g18890(.A1(new_n7617_), .A2(\b[46] ), .ZN(new_n19148_));
  AOI21_X1   g18891(.A1(new_n19148_), .A2(new_n19147_), .B(new_n6731_), .ZN(new_n19149_));
  NAND2_X1   g18892(.A1(new_n5177_), .A2(new_n19149_), .ZN(new_n19150_));
  XOR2_X1    g18893(.A1(new_n19150_), .A2(\a[56] ), .Z(new_n19151_));
  NAND2_X1   g18894(.A1(new_n19026_), .A2(new_n19016_), .ZN(new_n19152_));
  NAND2_X1   g18895(.A1(new_n19152_), .A2(new_n19025_), .ZN(new_n19153_));
  XOR2_X1    g18896(.A1(new_n19153_), .A2(new_n19151_), .Z(new_n19154_));
  AOI21_X1   g18897(.A1(new_n19152_), .A2(new_n19025_), .B(new_n19151_), .ZN(new_n19155_));
  INV_X1     g18898(.I(new_n19151_), .ZN(new_n19156_));
  NOR2_X1    g18899(.A1(new_n19153_), .A2(new_n19156_), .ZN(new_n19157_));
  OAI21_X1   g18900(.A1(new_n19157_), .A2(new_n19155_), .B(new_n19146_), .ZN(new_n19158_));
  OAI21_X1   g18901(.A1(new_n19146_), .A2(new_n19154_), .B(new_n19158_), .ZN(new_n19159_));
  OAI22_X1   g18902(.A1(new_n5786_), .A2(new_n5738_), .B1(new_n5538_), .B2(new_n5792_), .ZN(new_n19160_));
  NAND2_X1   g18903(.A1(new_n6745_), .A2(\b[49] ), .ZN(new_n19161_));
  AOI21_X1   g18904(.A1(new_n19161_), .A2(new_n19160_), .B(new_n5796_), .ZN(new_n19162_));
  NAND2_X1   g18905(.A1(new_n5741_), .A2(new_n19162_), .ZN(new_n19163_));
  XOR2_X1    g18906(.A1(new_n19163_), .A2(\a[53] ), .Z(new_n19164_));
  XNOR2_X1   g18907(.A1(new_n19159_), .A2(new_n19164_), .ZN(new_n19165_));
  INV_X1     g18908(.I(new_n19165_), .ZN(new_n19166_));
  NOR2_X1    g18909(.A1(new_n19159_), .A2(new_n19164_), .ZN(new_n19167_));
  INV_X1     g18910(.I(new_n19167_), .ZN(new_n19168_));
  NAND2_X1   g18911(.A1(new_n19159_), .A2(new_n19164_), .ZN(new_n19169_));
  AOI21_X1   g18912(.A1(new_n19168_), .A2(new_n19169_), .B(new_n19106_), .ZN(new_n19170_));
  AOI21_X1   g18913(.A1(new_n19166_), .A2(new_n19106_), .B(new_n19170_), .ZN(new_n19171_));
  XOR2_X1    g18914(.A1(new_n19171_), .A2(new_n19104_), .Z(new_n19172_));
  NOR2_X1    g18915(.A1(new_n19172_), .A2(new_n19099_), .ZN(new_n19173_));
  INV_X1     g18916(.I(new_n19099_), .ZN(new_n19174_));
  INV_X1     g18917(.I(new_n19104_), .ZN(new_n19175_));
  NOR2_X1    g18918(.A1(new_n19171_), .A2(new_n19175_), .ZN(new_n19176_));
  INV_X1     g18919(.I(new_n19176_), .ZN(new_n19177_));
  NAND2_X1   g18920(.A1(new_n19171_), .A2(new_n19175_), .ZN(new_n19178_));
  AOI21_X1   g18921(.A1(new_n19177_), .A2(new_n19178_), .B(new_n19174_), .ZN(new_n19179_));
  NOR2_X1    g18922(.A1(new_n19179_), .A2(new_n19173_), .ZN(new_n19180_));
  OAI22_X1   g18923(.A1(new_n4711_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n4706_), .ZN(new_n19181_));
  NAND2_X1   g18924(.A1(new_n5814_), .A2(\b[55] ), .ZN(new_n19182_));
  AOI21_X1   g18925(.A1(new_n19181_), .A2(new_n19182_), .B(new_n4714_), .ZN(new_n19183_));
  NAND2_X1   g18926(.A1(new_n7308_), .A2(new_n19183_), .ZN(new_n19184_));
  XOR2_X1    g18927(.A1(new_n19184_), .A2(\a[47] ), .Z(new_n19185_));
  INV_X1     g18928(.I(new_n19185_), .ZN(new_n19186_));
  XOR2_X1    g18929(.A1(new_n19180_), .A2(new_n19186_), .Z(new_n19187_));
  NAND2_X1   g18930(.A1(new_n19187_), .A2(new_n19098_), .ZN(new_n19188_));
  INV_X1     g18931(.I(new_n19180_), .ZN(new_n19189_));
  NOR2_X1    g18932(.A1(new_n19189_), .A2(new_n19185_), .ZN(new_n19190_));
  NOR2_X1    g18933(.A1(new_n19180_), .A2(new_n19186_), .ZN(new_n19191_));
  NOR2_X1    g18934(.A1(new_n19190_), .A2(new_n19191_), .ZN(new_n19192_));
  OAI21_X1   g18935(.A1(new_n19098_), .A2(new_n19192_), .B(new_n19188_), .ZN(new_n19193_));
  OAI22_X1   g18936(.A1(new_n4208_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n4203_), .ZN(new_n19194_));
  NAND2_X1   g18937(.A1(new_n5244_), .A2(\b[58] ), .ZN(new_n19195_));
  AOI21_X1   g18938(.A1(new_n19194_), .A2(new_n19195_), .B(new_n4211_), .ZN(new_n19196_));
  NAND2_X1   g18939(.A1(new_n7929_), .A2(new_n19196_), .ZN(new_n19197_));
  XOR2_X1    g18940(.A1(new_n19197_), .A2(\a[44] ), .Z(new_n19198_));
  NOR2_X1    g18941(.A1(new_n19058_), .A2(new_n19071_), .ZN(new_n19199_));
  NOR2_X1    g18942(.A1(new_n19199_), .A2(new_n19069_), .ZN(new_n19200_));
  NOR2_X1    g18943(.A1(new_n19200_), .A2(new_n19198_), .ZN(new_n19201_));
  INV_X1     g18944(.I(new_n19198_), .ZN(new_n19202_));
  NOR3_X1    g18945(.A1(new_n19199_), .A2(new_n19069_), .A3(new_n19202_), .ZN(new_n19203_));
  OAI21_X1   g18946(.A1(new_n19201_), .A2(new_n19203_), .B(new_n19193_), .ZN(new_n19204_));
  XOR2_X1    g18947(.A1(new_n19200_), .A2(new_n19202_), .Z(new_n19205_));
  OAI21_X1   g18948(.A1(new_n19205_), .A2(new_n19193_), .B(new_n19204_), .ZN(new_n19206_));
  XOR2_X1    g18949(.A1(new_n19097_), .A2(new_n19206_), .Z(new_n19207_));
  NAND2_X1   g18950(.A1(new_n19207_), .A2(new_n19095_), .ZN(new_n19208_));
  NAND2_X1   g18951(.A1(new_n19097_), .A2(new_n19206_), .ZN(new_n19209_));
  NOR2_X1    g18952(.A1(new_n19097_), .A2(new_n19206_), .ZN(new_n19210_));
  INV_X1     g18953(.I(new_n19210_), .ZN(new_n19211_));
  NAND2_X1   g18954(.A1(new_n19211_), .A2(new_n19209_), .ZN(new_n19212_));
  NAND2_X1   g18955(.A1(new_n19212_), .A2(new_n19094_), .ZN(new_n19213_));
  NAND2_X1   g18956(.A1(new_n19213_), .A2(new_n19208_), .ZN(new_n19214_));
  NAND2_X1   g18957(.A1(new_n19082_), .A2(new_n18960_), .ZN(new_n19215_));
  XOR2_X1    g18958(.A1(new_n18961_), .A2(\a[38] ), .Z(new_n19216_));
  NAND2_X1   g18959(.A1(new_n19215_), .A2(new_n19216_), .ZN(new_n19217_));
  OAI21_X1   g18960(.A1(new_n18960_), .A2(new_n19082_), .B(new_n19217_), .ZN(new_n19218_));
  XOR2_X1    g18961(.A1(new_n19218_), .A2(new_n19214_), .Z(new_n19219_));
  INV_X1     g18962(.I(new_n19219_), .ZN(new_n19220_));
  INV_X1     g18963(.I(new_n18959_), .ZN(new_n19221_));
  NAND2_X1   g18964(.A1(new_n18957_), .A2(new_n19221_), .ZN(new_n19222_));
  XOR2_X1    g18965(.A1(new_n19222_), .A2(new_n19220_), .Z(new_n19223_));
  INV_X1     g18966(.I(new_n19085_), .ZN(new_n19224_));
  XOR2_X1    g18967(.A1(new_n18957_), .A2(new_n19221_), .Z(new_n19225_));
  NAND2_X1   g18968(.A1(new_n19225_), .A2(new_n19224_), .ZN(new_n19226_));
  XOR2_X1    g18969(.A1(new_n19223_), .A2(new_n19226_), .Z(\f[102] ));
  NOR2_X1    g18970(.A1(new_n3889_), .A2(new_n8932_), .ZN(new_n19228_));
  NOR2_X1    g18971(.A1(new_n3731_), .A2(new_n8956_), .ZN(new_n19229_));
  NOR4_X1    g18972(.A1(new_n9323_), .A2(new_n3739_), .A3(new_n19228_), .A4(new_n19229_), .ZN(new_n19230_));
  XOR2_X1    g18973(.A1(new_n19230_), .A2(new_n3726_), .Z(new_n19231_));
  NOR2_X1    g18974(.A1(new_n19203_), .A2(new_n19193_), .ZN(new_n19232_));
  OAI22_X1   g18975(.A1(new_n4711_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n4706_), .ZN(new_n19233_));
  NAND2_X1   g18976(.A1(new_n5814_), .A2(\b[56] ), .ZN(new_n19234_));
  AOI21_X1   g18977(.A1(new_n19233_), .A2(new_n19234_), .B(new_n4714_), .ZN(new_n19235_));
  NAND2_X1   g18978(.A1(new_n7559_), .A2(new_n19235_), .ZN(new_n19236_));
  XOR2_X1    g18979(.A1(new_n19236_), .A2(\a[47] ), .Z(new_n19237_));
  INV_X1     g18980(.I(new_n19237_), .ZN(new_n19238_));
  OAI22_X1   g18981(.A1(new_n5786_), .A2(new_n5955_), .B1(new_n5738_), .B2(new_n5792_), .ZN(new_n19239_));
  NAND2_X1   g18982(.A1(new_n6745_), .A2(\b[50] ), .ZN(new_n19240_));
  AOI21_X1   g18983(.A1(new_n19240_), .A2(new_n19239_), .B(new_n5796_), .ZN(new_n19241_));
  NAND2_X1   g18984(.A1(new_n5954_), .A2(new_n19241_), .ZN(new_n19242_));
  XOR2_X1    g18985(.A1(new_n19242_), .A2(\a[53] ), .Z(new_n19243_));
  OAI21_X1   g18986(.A1(new_n19108_), .A2(new_n19125_), .B(new_n19127_), .ZN(new_n19244_));
  INV_X1     g18987(.I(new_n19244_), .ZN(new_n19245_));
  OAI22_X1   g18988(.A1(new_n4834_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n4509_), .ZN(new_n19246_));
  NAND2_X1   g18989(.A1(new_n8628_), .A2(\b[44] ), .ZN(new_n19247_));
  AOI21_X1   g18990(.A1(new_n19247_), .A2(new_n19246_), .B(new_n7354_), .ZN(new_n19248_));
  NAND2_X1   g18991(.A1(new_n4833_), .A2(new_n19248_), .ZN(new_n19249_));
  XOR2_X1    g18992(.A1(new_n19249_), .A2(\a[59] ), .Z(new_n19250_));
  INV_X1     g18993(.I(new_n19250_), .ZN(new_n19251_));
  OAI22_X1   g18994(.A1(new_n4316_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n4018_), .ZN(new_n19252_));
  NAND2_X1   g18995(.A1(new_n9644_), .A2(\b[41] ), .ZN(new_n19253_));
  AOI21_X1   g18996(.A1(new_n19253_), .A2(new_n19252_), .B(new_n8321_), .ZN(new_n19254_));
  NAND2_X1   g18997(.A1(new_n4320_), .A2(new_n19254_), .ZN(new_n19255_));
  XOR2_X1    g18998(.A1(new_n19255_), .A2(\a[62] ), .Z(new_n19256_));
  NAND2_X1   g18999(.A1(new_n19122_), .A2(new_n18834_), .ZN(new_n19257_));
  NAND2_X1   g19000(.A1(new_n19257_), .A2(new_n19121_), .ZN(new_n19258_));
  NOR3_X1    g19001(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n3696_), .ZN(new_n19259_));
  NOR2_X1    g19002(.A1(new_n9364_), .A2(new_n3696_), .ZN(new_n19260_));
  NOR3_X1    g19003(.A1(new_n19260_), .A2(new_n3845_), .A3(new_n8985_), .ZN(new_n19261_));
  NOR2_X1    g19004(.A1(new_n19261_), .A2(new_n19259_), .ZN(new_n19262_));
  INV_X1     g19005(.I(new_n19262_), .ZN(new_n19263_));
  XOR2_X1    g19006(.A1(new_n19258_), .A2(new_n19263_), .Z(new_n19264_));
  NOR2_X1    g19007(.A1(new_n19256_), .A2(new_n19264_), .ZN(new_n19265_));
  NOR2_X1    g19008(.A1(new_n19258_), .A2(new_n19262_), .ZN(new_n19266_));
  INV_X1     g19009(.I(new_n19266_), .ZN(new_n19267_));
  NAND2_X1   g19010(.A1(new_n19258_), .A2(new_n19262_), .ZN(new_n19268_));
  NAND2_X1   g19011(.A1(new_n19267_), .A2(new_n19268_), .ZN(new_n19269_));
  AOI21_X1   g19012(.A1(new_n19256_), .A2(new_n19269_), .B(new_n19265_), .ZN(new_n19270_));
  NOR2_X1    g19013(.A1(new_n19270_), .A2(new_n19251_), .ZN(new_n19271_));
  INV_X1     g19014(.I(new_n19271_), .ZN(new_n19272_));
  NAND2_X1   g19015(.A1(new_n19270_), .A2(new_n19251_), .ZN(new_n19273_));
  AOI21_X1   g19016(.A1(new_n19272_), .A2(new_n19273_), .B(new_n19245_), .ZN(new_n19274_));
  XOR2_X1    g19017(.A1(new_n19270_), .A2(new_n19250_), .Z(new_n19275_));
  NOR2_X1    g19018(.A1(new_n19275_), .A2(new_n19244_), .ZN(new_n19276_));
  NOR2_X1    g19019(.A1(new_n19276_), .A2(new_n19274_), .ZN(new_n19277_));
  NOR2_X1    g19020(.A1(new_n19141_), .A2(new_n19130_), .ZN(new_n19278_));
  NOR2_X1    g19021(.A1(new_n19278_), .A2(new_n19138_), .ZN(new_n19279_));
  OAI22_X1   g19022(.A1(new_n6721_), .A2(new_n5178_), .B1(new_n6723_), .B2(new_n5197_), .ZN(new_n19280_));
  NAND2_X1   g19023(.A1(new_n7617_), .A2(\b[47] ), .ZN(new_n19281_));
  AOI21_X1   g19024(.A1(new_n19281_), .A2(new_n19280_), .B(new_n6731_), .ZN(new_n19282_));
  NAND2_X1   g19025(.A1(new_n5196_), .A2(new_n19282_), .ZN(new_n19283_));
  XOR2_X1    g19026(.A1(new_n19283_), .A2(\a[56] ), .Z(new_n19284_));
  NOR2_X1    g19027(.A1(new_n19284_), .A2(new_n19279_), .ZN(new_n19285_));
  INV_X1     g19028(.I(new_n19285_), .ZN(new_n19286_));
  NAND2_X1   g19029(.A1(new_n19284_), .A2(new_n19279_), .ZN(new_n19287_));
  AOI21_X1   g19030(.A1(new_n19286_), .A2(new_n19287_), .B(new_n19277_), .ZN(new_n19288_));
  INV_X1     g19031(.I(new_n19277_), .ZN(new_n19289_));
  XNOR2_X1   g19032(.A1(new_n19284_), .A2(new_n19279_), .ZN(new_n19290_));
  NOR2_X1    g19033(.A1(new_n19290_), .A2(new_n19289_), .ZN(new_n19291_));
  NOR2_X1    g19034(.A1(new_n19291_), .A2(new_n19288_), .ZN(new_n19292_));
  NOR2_X1    g19035(.A1(new_n19157_), .A2(new_n19146_), .ZN(new_n19293_));
  NOR2_X1    g19036(.A1(new_n19293_), .A2(new_n19155_), .ZN(new_n19294_));
  NOR2_X1    g19037(.A1(new_n19294_), .A2(new_n19292_), .ZN(new_n19295_));
  INV_X1     g19038(.I(new_n19294_), .ZN(new_n19296_));
  NOR3_X1    g19039(.A1(new_n19296_), .A2(new_n19288_), .A3(new_n19291_), .ZN(new_n19297_));
  NOR2_X1    g19040(.A1(new_n19297_), .A2(new_n19295_), .ZN(new_n19298_));
  NOR2_X1    g19041(.A1(new_n19298_), .A2(new_n19243_), .ZN(new_n19299_));
  INV_X1     g19042(.I(new_n19243_), .ZN(new_n19300_));
  XNOR2_X1   g19043(.A1(new_n19294_), .A2(new_n19292_), .ZN(new_n19301_));
  NOR2_X1    g19044(.A1(new_n19301_), .A2(new_n19300_), .ZN(new_n19302_));
  NOR2_X1    g19045(.A1(new_n19299_), .A2(new_n19302_), .ZN(new_n19303_));
  NAND2_X1   g19046(.A1(new_n19106_), .A2(new_n19169_), .ZN(new_n19304_));
  NAND2_X1   g19047(.A1(new_n19304_), .A2(new_n19168_), .ZN(new_n19305_));
  INV_X1     g19048(.I(new_n19305_), .ZN(new_n19306_));
  OAI22_X1   g19049(.A1(new_n5228_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n5225_), .ZN(new_n19307_));
  NAND2_X1   g19050(.A1(new_n5387_), .A2(\b[53] ), .ZN(new_n19308_));
  AOI21_X1   g19051(.A1(new_n19307_), .A2(new_n19308_), .B(new_n5231_), .ZN(new_n19309_));
  NAND2_X1   g19052(.A1(new_n6471_), .A2(new_n19309_), .ZN(new_n19310_));
  XOR2_X1    g19053(.A1(new_n19310_), .A2(\a[50] ), .Z(new_n19311_));
  NOR2_X1    g19054(.A1(new_n19306_), .A2(new_n19311_), .ZN(new_n19312_));
  INV_X1     g19055(.I(new_n19311_), .ZN(new_n19313_));
  NOR2_X1    g19056(.A1(new_n19305_), .A2(new_n19313_), .ZN(new_n19314_));
  NOR2_X1    g19057(.A1(new_n19312_), .A2(new_n19314_), .ZN(new_n19315_));
  NOR2_X1    g19058(.A1(new_n19315_), .A2(new_n19303_), .ZN(new_n19316_));
  INV_X1     g19059(.I(new_n19303_), .ZN(new_n19317_));
  XOR2_X1    g19060(.A1(new_n19305_), .A2(new_n19311_), .Z(new_n19318_));
  NOR2_X1    g19061(.A1(new_n19318_), .A2(new_n19317_), .ZN(new_n19319_));
  NOR2_X1    g19062(.A1(new_n19316_), .A2(new_n19319_), .ZN(new_n19320_));
  NAND2_X1   g19063(.A1(new_n19174_), .A2(new_n19177_), .ZN(new_n19321_));
  AOI21_X1   g19064(.A1(new_n19178_), .A2(new_n19321_), .B(new_n19320_), .ZN(new_n19322_));
  NAND2_X1   g19065(.A1(new_n19321_), .A2(new_n19178_), .ZN(new_n19323_));
  NOR3_X1    g19066(.A1(new_n19323_), .A2(new_n19316_), .A3(new_n19319_), .ZN(new_n19324_));
  OAI21_X1   g19067(.A1(new_n19324_), .A2(new_n19322_), .B(new_n19238_), .ZN(new_n19325_));
  XNOR2_X1   g19068(.A1(new_n19323_), .A2(new_n19320_), .ZN(new_n19326_));
  NAND2_X1   g19069(.A1(new_n19326_), .A2(new_n19237_), .ZN(new_n19327_));
  INV_X1     g19070(.I(new_n19190_), .ZN(new_n19328_));
  OAI21_X1   g19071(.A1(new_n19180_), .A2(new_n19186_), .B(new_n19098_), .ZN(new_n19329_));
  NAND2_X1   g19072(.A1(new_n19328_), .A2(new_n19329_), .ZN(new_n19330_));
  OAI22_X1   g19073(.A1(new_n4208_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n4203_), .ZN(new_n19331_));
  NAND2_X1   g19074(.A1(new_n5244_), .A2(\b[59] ), .ZN(new_n19332_));
  AOI21_X1   g19075(.A1(new_n19331_), .A2(new_n19332_), .B(new_n4211_), .ZN(new_n19333_));
  NAND2_X1   g19076(.A1(new_n8550_), .A2(new_n19333_), .ZN(new_n19334_));
  XOR2_X1    g19077(.A1(new_n19334_), .A2(\a[44] ), .Z(new_n19335_));
  XOR2_X1    g19078(.A1(new_n19330_), .A2(new_n19335_), .Z(new_n19336_));
  AOI21_X1   g19079(.A1(new_n19325_), .A2(new_n19327_), .B(new_n19336_), .ZN(new_n19337_));
  NAND2_X1   g19080(.A1(new_n19327_), .A2(new_n19325_), .ZN(new_n19338_));
  INV_X1     g19081(.I(new_n19330_), .ZN(new_n19339_));
  NOR2_X1    g19082(.A1(new_n19339_), .A2(new_n19335_), .ZN(new_n19340_));
  INV_X1     g19083(.I(new_n19340_), .ZN(new_n19341_));
  NAND2_X1   g19084(.A1(new_n19339_), .A2(new_n19335_), .ZN(new_n19342_));
  AOI21_X1   g19085(.A1(new_n19341_), .A2(new_n19342_), .B(new_n19338_), .ZN(new_n19343_));
  NOR2_X1    g19086(.A1(new_n19337_), .A2(new_n19343_), .ZN(new_n19344_));
  NOR3_X1    g19087(.A1(new_n19344_), .A2(new_n19201_), .A3(new_n19232_), .ZN(new_n19345_));
  NOR2_X1    g19088(.A1(new_n19232_), .A2(new_n19201_), .ZN(new_n19346_));
  INV_X1     g19089(.I(new_n19344_), .ZN(new_n19347_));
  NOR2_X1    g19090(.A1(new_n19347_), .A2(new_n19346_), .ZN(new_n19348_));
  NOR2_X1    g19091(.A1(new_n19348_), .A2(new_n19345_), .ZN(new_n19349_));
  NOR2_X1    g19092(.A1(new_n19349_), .A2(new_n19231_), .ZN(new_n19350_));
  INV_X1     g19093(.I(new_n19231_), .ZN(new_n19351_));
  XOR2_X1    g19094(.A1(new_n19344_), .A2(new_n19346_), .Z(new_n19352_));
  NOR2_X1    g19095(.A1(new_n19352_), .A2(new_n19351_), .ZN(new_n19353_));
  NOR2_X1    g19096(.A1(new_n19350_), .A2(new_n19353_), .ZN(new_n19354_));
  AOI21_X1   g19097(.A1(new_n19095_), .A2(new_n19209_), .B(new_n19210_), .ZN(new_n19355_));
  INV_X1     g19098(.I(new_n19355_), .ZN(new_n19356_));
  INV_X1     g19099(.I(new_n18505_), .ZN(new_n19357_));
  OAI21_X1   g19100(.A1(new_n18496_), .A2(new_n19357_), .B(new_n18503_), .ZN(new_n19358_));
  NAND3_X1   g19101(.A1(new_n19358_), .A2(new_n18509_), .A3(new_n18945_), .ZN(new_n19359_));
  AOI21_X1   g19102(.A1(new_n19359_), .A2(new_n18955_), .B(new_n18952_), .ZN(new_n19360_));
  NOR2_X1    g19103(.A1(new_n19085_), .A2(new_n19220_), .ZN(new_n19361_));
  NOR3_X1    g19104(.A1(new_n19360_), .A2(new_n18959_), .A3(new_n19361_), .ZN(new_n19362_));
  AOI21_X1   g19105(.A1(new_n19208_), .A2(new_n19213_), .B(new_n19218_), .ZN(new_n19363_));
  NOR2_X1    g19106(.A1(new_n19362_), .A2(new_n19363_), .ZN(new_n19364_));
  XOR2_X1    g19107(.A1(new_n19364_), .A2(new_n19356_), .Z(new_n19365_));
  XOR2_X1    g19108(.A1(new_n19365_), .A2(new_n19354_), .Z(\f[103] ));
  INV_X1     g19109(.I(new_n19361_), .ZN(new_n19367_));
  NAND3_X1   g19110(.A1(new_n18957_), .A2(new_n19221_), .A3(new_n19367_), .ZN(new_n19368_));
  NOR2_X1    g19111(.A1(new_n19354_), .A2(new_n19356_), .ZN(new_n19369_));
  XOR2_X1    g19112(.A1(new_n19354_), .A2(new_n19356_), .Z(new_n19370_));
  NOR2_X1    g19113(.A1(new_n19363_), .A2(new_n19370_), .ZN(new_n19371_));
  AOI21_X1   g19114(.A1(new_n19368_), .A2(new_n19371_), .B(new_n19369_), .ZN(new_n19372_));
  INV_X1     g19115(.I(new_n19345_), .ZN(new_n19373_));
  AOI21_X1   g19116(.A1(new_n19373_), .A2(new_n19351_), .B(new_n19348_), .ZN(new_n19374_));
  INV_X1     g19117(.I(new_n19374_), .ZN(new_n19375_));
  AOI21_X1   g19118(.A1(new_n19338_), .A2(new_n19342_), .B(new_n19340_), .ZN(new_n19376_));
  INV_X1     g19119(.I(new_n19376_), .ZN(new_n19377_));
  OAI22_X1   g19120(.A1(new_n9595_), .A2(new_n3739_), .B1(new_n8956_), .B2(new_n3889_), .ZN(new_n19378_));
  OAI22_X1   g19121(.A1(new_n4208_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n4203_), .ZN(new_n19379_));
  NAND2_X1   g19122(.A1(new_n5244_), .A2(\b[60] ), .ZN(new_n19380_));
  AOI21_X1   g19123(.A1(new_n19379_), .A2(new_n19380_), .B(new_n4211_), .ZN(new_n19381_));
  NAND2_X1   g19124(.A1(new_n8935_), .A2(new_n19381_), .ZN(new_n19382_));
  XOR2_X1    g19125(.A1(new_n19382_), .A2(\a[44] ), .Z(new_n19383_));
  OAI22_X1   g19126(.A1(new_n5228_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n5225_), .ZN(new_n19384_));
  NAND2_X1   g19127(.A1(new_n5387_), .A2(\b[54] ), .ZN(new_n19385_));
  AOI21_X1   g19128(.A1(new_n19384_), .A2(new_n19385_), .B(new_n5231_), .ZN(new_n19386_));
  NAND2_X1   g19129(.A1(new_n6994_), .A2(new_n19386_), .ZN(new_n19387_));
  XOR2_X1    g19130(.A1(new_n19387_), .A2(\a[50] ), .Z(new_n19388_));
  INV_X1     g19131(.I(new_n19388_), .ZN(new_n19389_));
  NOR2_X1    g19132(.A1(new_n19297_), .A2(new_n19243_), .ZN(new_n19390_));
  NOR2_X1    g19133(.A1(new_n19390_), .A2(new_n19295_), .ZN(new_n19391_));
  INV_X1     g19134(.I(new_n19391_), .ZN(new_n19392_));
  OAI22_X1   g19135(.A1(new_n5786_), .A2(new_n6215_), .B1(new_n5955_), .B2(new_n5792_), .ZN(new_n19393_));
  NAND2_X1   g19136(.A1(new_n6745_), .A2(\b[51] ), .ZN(new_n19394_));
  AOI21_X1   g19137(.A1(new_n19394_), .A2(new_n19393_), .B(new_n5796_), .ZN(new_n19395_));
  NAND2_X1   g19138(.A1(new_n6219_), .A2(new_n19395_), .ZN(new_n19396_));
  XOR2_X1    g19139(.A1(new_n19396_), .A2(\a[53] ), .Z(new_n19397_));
  OAI22_X1   g19140(.A1(new_n6721_), .A2(new_n5197_), .B1(new_n6723_), .B2(new_n5538_), .ZN(new_n19398_));
  NAND2_X1   g19141(.A1(new_n7617_), .A2(\b[48] ), .ZN(new_n19399_));
  AOI21_X1   g19142(.A1(new_n19399_), .A2(new_n19398_), .B(new_n6731_), .ZN(new_n19400_));
  NAND2_X1   g19143(.A1(new_n5537_), .A2(new_n19400_), .ZN(new_n19401_));
  XOR2_X1    g19144(.A1(new_n19401_), .A2(\a[56] ), .Z(new_n19402_));
  OAI21_X1   g19145(.A1(new_n19245_), .A2(new_n19271_), .B(new_n19273_), .ZN(new_n19403_));
  OAI21_X1   g19146(.A1(new_n19256_), .A2(new_n19266_), .B(new_n19268_), .ZN(new_n19404_));
  NOR3_X1    g19147(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n3845_), .ZN(new_n19405_));
  NOR2_X1    g19148(.A1(new_n9364_), .A2(new_n3845_), .ZN(new_n19406_));
  NOR3_X1    g19149(.A1(new_n19406_), .A2(new_n3997_), .A3(new_n8985_), .ZN(new_n19407_));
  NOR2_X1    g19150(.A1(new_n19407_), .A2(new_n19405_), .ZN(new_n19408_));
  NOR2_X1    g19151(.A1(new_n19263_), .A2(new_n19408_), .ZN(new_n19409_));
  INV_X1     g19152(.I(new_n19408_), .ZN(new_n19410_));
  NOR2_X1    g19153(.A1(new_n19410_), .A2(new_n19262_), .ZN(new_n19411_));
  OAI21_X1   g19154(.A1(new_n19409_), .A2(new_n19411_), .B(new_n19404_), .ZN(new_n19412_));
  XOR2_X1    g19155(.A1(new_n19262_), .A2(new_n19408_), .Z(new_n19413_));
  OR2_X2     g19156(.A1(new_n19404_), .A2(new_n19413_), .Z(new_n19414_));
  NAND2_X1   g19157(.A1(new_n19414_), .A2(new_n19412_), .ZN(new_n19415_));
  OAI22_X1   g19158(.A1(new_n4997_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n4834_), .ZN(new_n19416_));
  NAND2_X1   g19159(.A1(new_n8628_), .A2(\b[45] ), .ZN(new_n19417_));
  AOI21_X1   g19160(.A1(new_n19417_), .A2(new_n19416_), .B(new_n7354_), .ZN(new_n19418_));
  NAND2_X1   g19161(.A1(new_n5004_), .A2(new_n19418_), .ZN(new_n19419_));
  XOR2_X1    g19162(.A1(new_n19419_), .A2(\a[59] ), .Z(new_n19420_));
  OAI22_X1   g19163(.A1(new_n4501_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n4316_), .ZN(new_n19421_));
  NAND2_X1   g19164(.A1(new_n9644_), .A2(\b[42] ), .ZN(new_n19422_));
  AOI21_X1   g19165(.A1(new_n19422_), .A2(new_n19421_), .B(new_n8321_), .ZN(new_n19423_));
  NAND2_X1   g19166(.A1(new_n4500_), .A2(new_n19423_), .ZN(new_n19424_));
  XOR2_X1    g19167(.A1(new_n19424_), .A2(\a[62] ), .Z(new_n19425_));
  XNOR2_X1   g19168(.A1(new_n19420_), .A2(new_n19425_), .ZN(new_n19426_));
  INV_X1     g19169(.I(new_n19426_), .ZN(new_n19427_));
  NOR2_X1    g19170(.A1(new_n19420_), .A2(new_n19425_), .ZN(new_n19428_));
  INV_X1     g19171(.I(new_n19428_), .ZN(new_n19429_));
  NAND2_X1   g19172(.A1(new_n19420_), .A2(new_n19425_), .ZN(new_n19430_));
  AOI21_X1   g19173(.A1(new_n19429_), .A2(new_n19430_), .B(new_n19415_), .ZN(new_n19431_));
  AOI21_X1   g19174(.A1(new_n19427_), .A2(new_n19415_), .B(new_n19431_), .ZN(new_n19432_));
  XNOR2_X1   g19175(.A1(new_n19432_), .A2(new_n19403_), .ZN(new_n19433_));
  NOR2_X1    g19176(.A1(new_n19433_), .A2(new_n19402_), .ZN(new_n19434_));
  INV_X1     g19177(.I(new_n19402_), .ZN(new_n19435_));
  NOR2_X1    g19178(.A1(new_n19432_), .A2(new_n19403_), .ZN(new_n19436_));
  INV_X1     g19179(.I(new_n19436_), .ZN(new_n19437_));
  NAND2_X1   g19180(.A1(new_n19432_), .A2(new_n19403_), .ZN(new_n19438_));
  AOI21_X1   g19181(.A1(new_n19437_), .A2(new_n19438_), .B(new_n19435_), .ZN(new_n19439_));
  NOR2_X1    g19182(.A1(new_n19434_), .A2(new_n19439_), .ZN(new_n19440_));
  AOI21_X1   g19183(.A1(new_n19289_), .A2(new_n19287_), .B(new_n19285_), .ZN(new_n19441_));
  XOR2_X1    g19184(.A1(new_n19440_), .A2(new_n19441_), .Z(new_n19442_));
  NOR2_X1    g19185(.A1(new_n19442_), .A2(new_n19397_), .ZN(new_n19443_));
  INV_X1     g19186(.I(new_n19397_), .ZN(new_n19444_));
  INV_X1     g19187(.I(new_n19440_), .ZN(new_n19445_));
  NOR2_X1    g19188(.A1(new_n19445_), .A2(new_n19441_), .ZN(new_n19446_));
  INV_X1     g19189(.I(new_n19446_), .ZN(new_n19447_));
  NAND2_X1   g19190(.A1(new_n19445_), .A2(new_n19441_), .ZN(new_n19448_));
  AOI21_X1   g19191(.A1(new_n19447_), .A2(new_n19448_), .B(new_n19444_), .ZN(new_n19449_));
  NOR2_X1    g19192(.A1(new_n19449_), .A2(new_n19443_), .ZN(new_n19450_));
  XOR2_X1    g19193(.A1(new_n19450_), .A2(new_n19392_), .Z(new_n19451_));
  NOR2_X1    g19194(.A1(new_n19450_), .A2(new_n19392_), .ZN(new_n19452_));
  INV_X1     g19195(.I(new_n19452_), .ZN(new_n19453_));
  NAND2_X1   g19196(.A1(new_n19450_), .A2(new_n19392_), .ZN(new_n19454_));
  AOI21_X1   g19197(.A1(new_n19453_), .A2(new_n19454_), .B(new_n19389_), .ZN(new_n19455_));
  AOI21_X1   g19198(.A1(new_n19389_), .A2(new_n19451_), .B(new_n19455_), .ZN(new_n19456_));
  OAI22_X1   g19199(.A1(new_n4711_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n4706_), .ZN(new_n19457_));
  NAND2_X1   g19200(.A1(new_n5814_), .A2(\b[57] ), .ZN(new_n19458_));
  AOI21_X1   g19201(.A1(new_n19457_), .A2(new_n19458_), .B(new_n4714_), .ZN(new_n19459_));
  NAND2_X1   g19202(.A1(new_n7895_), .A2(new_n19459_), .ZN(new_n19460_));
  XOR2_X1    g19203(.A1(new_n19460_), .A2(\a[47] ), .Z(new_n19461_));
  NOR2_X1    g19204(.A1(new_n19314_), .A2(new_n19303_), .ZN(new_n19462_));
  NOR2_X1    g19205(.A1(new_n19462_), .A2(new_n19312_), .ZN(new_n19463_));
  XNOR2_X1   g19206(.A1(new_n19463_), .A2(new_n19461_), .ZN(new_n19464_));
  OR2_X2     g19207(.A1(new_n19456_), .A2(new_n19464_), .Z(new_n19465_));
  NOR2_X1    g19208(.A1(new_n19463_), .A2(new_n19461_), .ZN(new_n19466_));
  INV_X1     g19209(.I(new_n19466_), .ZN(new_n19467_));
  NAND2_X1   g19210(.A1(new_n19463_), .A2(new_n19461_), .ZN(new_n19468_));
  NAND2_X1   g19211(.A1(new_n19467_), .A2(new_n19468_), .ZN(new_n19469_));
  NAND2_X1   g19212(.A1(new_n19456_), .A2(new_n19469_), .ZN(new_n19470_));
  NAND2_X1   g19213(.A1(new_n19465_), .A2(new_n19470_), .ZN(new_n19471_));
  INV_X1     g19214(.I(new_n19471_), .ZN(new_n19472_));
  NOR2_X1    g19215(.A1(new_n19324_), .A2(new_n19237_), .ZN(new_n19473_));
  NOR2_X1    g19216(.A1(new_n19473_), .A2(new_n19322_), .ZN(new_n19474_));
  NOR2_X1    g19217(.A1(new_n19472_), .A2(new_n19474_), .ZN(new_n19475_));
  NOR3_X1    g19218(.A1(new_n19471_), .A2(new_n19322_), .A3(new_n19473_), .ZN(new_n19476_));
  NOR2_X1    g19219(.A1(new_n19475_), .A2(new_n19476_), .ZN(new_n19477_));
  NOR2_X1    g19220(.A1(new_n19477_), .A2(new_n19383_), .ZN(new_n19478_));
  INV_X1     g19221(.I(new_n19383_), .ZN(new_n19479_));
  XOR2_X1    g19222(.A1(new_n19471_), .A2(new_n19474_), .Z(new_n19480_));
  NOR2_X1    g19223(.A1(new_n19480_), .A2(new_n19479_), .ZN(new_n19481_));
  NOR2_X1    g19224(.A1(new_n19478_), .A2(new_n19481_), .ZN(new_n19482_));
  XOR2_X1    g19225(.A1(new_n19482_), .A2(new_n19378_), .Z(new_n19483_));
  XOR2_X1    g19226(.A1(new_n19483_), .A2(\a[41] ), .Z(new_n19484_));
  XOR2_X1    g19227(.A1(new_n19484_), .A2(new_n19377_), .Z(new_n19485_));
  XOR2_X1    g19228(.A1(new_n19485_), .A2(new_n19375_), .Z(new_n19486_));
  XOR2_X1    g19229(.A1(new_n19485_), .A2(new_n19375_), .Z(new_n19487_));
  NAND2_X1   g19230(.A1(new_n19372_), .A2(new_n19487_), .ZN(new_n19488_));
  OAI21_X1   g19231(.A1(new_n19372_), .A2(new_n19486_), .B(new_n19488_), .ZN(\f[104] ));
  OAI22_X1   g19232(.A1(new_n4208_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n4203_), .ZN(new_n19490_));
  NAND2_X1   g19233(.A1(new_n5244_), .A2(\b[61] ), .ZN(new_n19491_));
  AOI21_X1   g19234(.A1(new_n19490_), .A2(new_n19491_), .B(new_n4211_), .ZN(new_n19492_));
  NAND2_X1   g19235(.A1(new_n8963_), .A2(new_n19492_), .ZN(new_n19493_));
  XOR2_X1    g19236(.A1(new_n19493_), .A2(\a[44] ), .Z(new_n19494_));
  INV_X1     g19237(.I(new_n19476_), .ZN(new_n19495_));
  AOI21_X1   g19238(.A1(new_n19495_), .A2(new_n19479_), .B(new_n19475_), .ZN(new_n19496_));
  OAI21_X1   g19239(.A1(new_n19388_), .A2(new_n19452_), .B(new_n19454_), .ZN(new_n19497_));
  INV_X1     g19240(.I(new_n19497_), .ZN(new_n19498_));
  OAI22_X1   g19241(.A1(new_n5228_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n5225_), .ZN(new_n19499_));
  NAND2_X1   g19242(.A1(new_n5387_), .A2(\b[55] ), .ZN(new_n19500_));
  AOI21_X1   g19243(.A1(new_n19499_), .A2(new_n19500_), .B(new_n5231_), .ZN(new_n19501_));
  NAND2_X1   g19244(.A1(new_n7308_), .A2(new_n19501_), .ZN(new_n19502_));
  XOR2_X1    g19245(.A1(new_n19502_), .A2(\a[50] ), .Z(new_n19503_));
  AOI21_X1   g19246(.A1(new_n19444_), .A2(new_n19448_), .B(new_n19446_), .ZN(new_n19504_));
  OAI21_X1   g19247(.A1(new_n19402_), .A2(new_n19436_), .B(new_n19438_), .ZN(new_n19505_));
  OAI22_X1   g19248(.A1(new_n6721_), .A2(new_n5538_), .B1(new_n6723_), .B2(new_n5738_), .ZN(new_n19506_));
  NAND2_X1   g19249(.A1(new_n7617_), .A2(\b[49] ), .ZN(new_n19507_));
  AOI21_X1   g19250(.A1(new_n19507_), .A2(new_n19506_), .B(new_n6731_), .ZN(new_n19508_));
  NAND2_X1   g19251(.A1(new_n5741_), .A2(new_n19508_), .ZN(new_n19509_));
  XOR2_X1    g19252(.A1(new_n19509_), .A2(\a[56] ), .Z(new_n19510_));
  INV_X1     g19253(.I(new_n19510_), .ZN(new_n19511_));
  INV_X1     g19254(.I(new_n19411_), .ZN(new_n19512_));
  AOI21_X1   g19255(.A1(new_n19404_), .A2(new_n19512_), .B(new_n19409_), .ZN(new_n19513_));
  OAI22_X1   g19256(.A1(new_n4509_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n4501_), .ZN(new_n19514_));
  NAND2_X1   g19257(.A1(new_n9644_), .A2(\b[43] ), .ZN(new_n19515_));
  AOI21_X1   g19258(.A1(new_n19515_), .A2(new_n19514_), .B(new_n8321_), .ZN(new_n19516_));
  NAND2_X1   g19259(.A1(new_n4513_), .A2(new_n19516_), .ZN(new_n19517_));
  XOR2_X1    g19260(.A1(new_n19517_), .A2(\a[62] ), .Z(new_n19518_));
  NOR2_X1    g19261(.A1(new_n8985_), .A2(new_n4018_), .ZN(new_n19519_));
  NOR2_X1    g19262(.A1(new_n9364_), .A2(new_n3997_), .ZN(new_n19520_));
  XNOR2_X1   g19263(.A1(new_n19519_), .A2(new_n19520_), .ZN(new_n19521_));
  XOR2_X1    g19264(.A1(new_n19521_), .A2(\a[41] ), .Z(new_n19522_));
  NOR2_X1    g19265(.A1(new_n19522_), .A2(new_n19262_), .ZN(new_n19523_));
  NOR2_X1    g19266(.A1(new_n19521_), .A2(new_n3726_), .ZN(new_n19524_));
  INV_X1     g19267(.I(new_n19524_), .ZN(new_n19525_));
  NAND2_X1   g19268(.A1(new_n19521_), .A2(new_n3726_), .ZN(new_n19526_));
  AOI21_X1   g19269(.A1(new_n19525_), .A2(new_n19526_), .B(new_n19263_), .ZN(new_n19527_));
  NOR2_X1    g19270(.A1(new_n19523_), .A2(new_n19527_), .ZN(new_n19528_));
  XOR2_X1    g19271(.A1(new_n19518_), .A2(new_n19528_), .Z(new_n19529_));
  NOR2_X1    g19272(.A1(new_n19529_), .A2(new_n19513_), .ZN(new_n19530_));
  INV_X1     g19273(.I(new_n19518_), .ZN(new_n19531_));
  NOR2_X1    g19274(.A1(new_n19531_), .A2(new_n19528_), .ZN(new_n19532_));
  INV_X1     g19275(.I(new_n19532_), .ZN(new_n19533_));
  NAND2_X1   g19276(.A1(new_n19531_), .A2(new_n19528_), .ZN(new_n19534_));
  NAND2_X1   g19277(.A1(new_n19533_), .A2(new_n19534_), .ZN(new_n19535_));
  AOI21_X1   g19278(.A1(new_n19513_), .A2(new_n19535_), .B(new_n19530_), .ZN(new_n19536_));
  INV_X1     g19279(.I(new_n19536_), .ZN(new_n19537_));
  OAI22_X1   g19280(.A1(new_n5178_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n4997_), .ZN(new_n19538_));
  NAND2_X1   g19281(.A1(new_n8628_), .A2(\b[46] ), .ZN(new_n19539_));
  AOI21_X1   g19282(.A1(new_n19539_), .A2(new_n19538_), .B(new_n7354_), .ZN(new_n19540_));
  NAND2_X1   g19283(.A1(new_n5177_), .A2(new_n19540_), .ZN(new_n19541_));
  XOR2_X1    g19284(.A1(new_n19541_), .A2(\a[59] ), .Z(new_n19542_));
  NAND2_X1   g19285(.A1(new_n19430_), .A2(new_n19415_), .ZN(new_n19543_));
  NAND2_X1   g19286(.A1(new_n19543_), .A2(new_n19429_), .ZN(new_n19544_));
  INV_X1     g19287(.I(new_n19544_), .ZN(new_n19545_));
  NOR2_X1    g19288(.A1(new_n19545_), .A2(new_n19542_), .ZN(new_n19546_));
  INV_X1     g19289(.I(new_n19542_), .ZN(new_n19547_));
  NOR2_X1    g19290(.A1(new_n19544_), .A2(new_n19547_), .ZN(new_n19548_));
  OAI21_X1   g19291(.A1(new_n19546_), .A2(new_n19548_), .B(new_n19537_), .ZN(new_n19549_));
  XOR2_X1    g19292(.A1(new_n19544_), .A2(new_n19547_), .Z(new_n19550_));
  NAND2_X1   g19293(.A1(new_n19550_), .A2(new_n19536_), .ZN(new_n19551_));
  AOI21_X1   g19294(.A1(new_n19551_), .A2(new_n19549_), .B(new_n19511_), .ZN(new_n19552_));
  NAND2_X1   g19295(.A1(new_n19551_), .A2(new_n19549_), .ZN(new_n19553_));
  NOR2_X1    g19296(.A1(new_n19553_), .A2(new_n19510_), .ZN(new_n19554_));
  NOR2_X1    g19297(.A1(new_n19554_), .A2(new_n19552_), .ZN(new_n19555_));
  XOR2_X1    g19298(.A1(new_n19553_), .A2(new_n19511_), .Z(new_n19556_));
  MUX2_X1    g19299(.I0(new_n19556_), .I1(new_n19555_), .S(new_n19505_), .Z(new_n19557_));
  OAI22_X1   g19300(.A1(new_n5786_), .A2(new_n6238_), .B1(new_n6215_), .B2(new_n5792_), .ZN(new_n19558_));
  NAND2_X1   g19301(.A1(new_n6745_), .A2(\b[52] ), .ZN(new_n19559_));
  AOI21_X1   g19302(.A1(new_n19559_), .A2(new_n19558_), .B(new_n5796_), .ZN(new_n19560_));
  NAND2_X1   g19303(.A1(new_n6237_), .A2(new_n19560_), .ZN(new_n19561_));
  XOR2_X1    g19304(.A1(new_n19561_), .A2(\a[53] ), .Z(new_n19562_));
  XNOR2_X1   g19305(.A1(new_n19557_), .A2(new_n19562_), .ZN(new_n19563_));
  NOR2_X1    g19306(.A1(new_n19563_), .A2(new_n19504_), .ZN(new_n19564_));
  INV_X1     g19307(.I(new_n19504_), .ZN(new_n19565_));
  NOR2_X1    g19308(.A1(new_n19557_), .A2(new_n19562_), .ZN(new_n19566_));
  INV_X1     g19309(.I(new_n19566_), .ZN(new_n19567_));
  NAND2_X1   g19310(.A1(new_n19557_), .A2(new_n19562_), .ZN(new_n19568_));
  AOI21_X1   g19311(.A1(new_n19567_), .A2(new_n19568_), .B(new_n19565_), .ZN(new_n19569_));
  NOR2_X1    g19312(.A1(new_n19564_), .A2(new_n19569_), .ZN(new_n19570_));
  XOR2_X1    g19313(.A1(new_n19570_), .A2(new_n19503_), .Z(new_n19571_));
  NOR2_X1    g19314(.A1(new_n19571_), .A2(new_n19498_), .ZN(new_n19572_));
  INV_X1     g19315(.I(new_n19503_), .ZN(new_n19573_));
  NOR2_X1    g19316(.A1(new_n19570_), .A2(new_n19573_), .ZN(new_n19574_));
  INV_X1     g19317(.I(new_n19574_), .ZN(new_n19575_));
  NAND2_X1   g19318(.A1(new_n19570_), .A2(new_n19573_), .ZN(new_n19576_));
  AOI21_X1   g19319(.A1(new_n19575_), .A2(new_n19576_), .B(new_n19497_), .ZN(new_n19577_));
  NOR2_X1    g19320(.A1(new_n19572_), .A2(new_n19577_), .ZN(new_n19578_));
  OAI22_X1   g19321(.A1(new_n4711_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n4706_), .ZN(new_n19579_));
  NAND2_X1   g19322(.A1(new_n5814_), .A2(\b[58] ), .ZN(new_n19580_));
  AOI21_X1   g19323(.A1(new_n19579_), .A2(new_n19580_), .B(new_n4714_), .ZN(new_n19581_));
  NAND2_X1   g19324(.A1(new_n7929_), .A2(new_n19581_), .ZN(new_n19582_));
  XOR2_X1    g19325(.A1(new_n19582_), .A2(\a[47] ), .Z(new_n19583_));
  NAND2_X1   g19326(.A1(new_n19456_), .A2(new_n19468_), .ZN(new_n19584_));
  NAND2_X1   g19327(.A1(new_n19584_), .A2(new_n19467_), .ZN(new_n19585_));
  INV_X1     g19328(.I(new_n19585_), .ZN(new_n19586_));
  NOR2_X1    g19329(.A1(new_n19586_), .A2(new_n19583_), .ZN(new_n19587_));
  INV_X1     g19330(.I(new_n19583_), .ZN(new_n19588_));
  NOR2_X1    g19331(.A1(new_n19585_), .A2(new_n19588_), .ZN(new_n19589_));
  NOR2_X1    g19332(.A1(new_n19587_), .A2(new_n19589_), .ZN(new_n19590_));
  NOR2_X1    g19333(.A1(new_n19590_), .A2(new_n19578_), .ZN(new_n19591_));
  XOR2_X1    g19334(.A1(new_n19585_), .A2(new_n19583_), .Z(new_n19592_));
  INV_X1     g19335(.I(new_n19592_), .ZN(new_n19593_));
  AOI21_X1   g19336(.A1(new_n19578_), .A2(new_n19593_), .B(new_n19591_), .ZN(new_n19594_));
  XOR2_X1    g19337(.A1(new_n19594_), .A2(new_n19496_), .Z(new_n19595_));
  NOR2_X1    g19338(.A1(new_n19595_), .A2(new_n19494_), .ZN(new_n19596_));
  INV_X1     g19339(.I(new_n19496_), .ZN(new_n19597_));
  NOR2_X1    g19340(.A1(new_n19594_), .A2(new_n19597_), .ZN(new_n19598_));
  INV_X1     g19341(.I(new_n19598_), .ZN(new_n19599_));
  NAND2_X1   g19342(.A1(new_n19594_), .A2(new_n19597_), .ZN(new_n19600_));
  NAND2_X1   g19343(.A1(new_n19599_), .A2(new_n19600_), .ZN(new_n19601_));
  AOI21_X1   g19344(.A1(new_n19494_), .A2(new_n19601_), .B(new_n19596_), .ZN(new_n19602_));
  NOR2_X1    g19345(.A1(new_n19482_), .A2(new_n19376_), .ZN(new_n19603_));
  XOR2_X1    g19346(.A1(new_n19378_), .A2(new_n3726_), .Z(new_n19604_));
  AOI21_X1   g19347(.A1(new_n19482_), .A2(new_n19376_), .B(new_n19604_), .ZN(new_n19605_));
  NOR2_X1    g19348(.A1(new_n19605_), .A2(new_n19603_), .ZN(new_n19606_));
  XOR2_X1    g19349(.A1(new_n19602_), .A2(new_n19606_), .Z(new_n19607_));
  NOR2_X1    g19350(.A1(new_n19372_), .A2(new_n19374_), .ZN(new_n19608_));
  XOR2_X1    g19351(.A1(new_n19608_), .A2(new_n19607_), .Z(new_n19609_));
  INV_X1     g19352(.I(new_n19485_), .ZN(new_n19610_));
  XOR2_X1    g19353(.A1(new_n19372_), .A2(new_n19374_), .Z(new_n19611_));
  NAND2_X1   g19354(.A1(new_n19611_), .A2(new_n19610_), .ZN(new_n19612_));
  XOR2_X1    g19355(.A1(new_n19609_), .A2(new_n19612_), .Z(\f[105] ));
  NOR2_X1    g19356(.A1(new_n4362_), .A2(new_n8932_), .ZN(new_n19614_));
  NOR2_X1    g19357(.A1(new_n4203_), .A2(new_n8956_), .ZN(new_n19615_));
  NOR4_X1    g19358(.A1(new_n9323_), .A2(new_n4211_), .A3(new_n19614_), .A4(new_n19615_), .ZN(new_n19616_));
  XOR2_X1    g19359(.A1(new_n19616_), .A2(new_n4198_), .Z(new_n19617_));
  INV_X1     g19360(.I(new_n19589_), .ZN(new_n19618_));
  AOI21_X1   g19361(.A1(new_n19578_), .A2(new_n19618_), .B(new_n19587_), .ZN(new_n19619_));
  OAI22_X1   g19362(.A1(new_n4711_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n4706_), .ZN(new_n19620_));
  NAND2_X1   g19363(.A1(new_n5814_), .A2(\b[59] ), .ZN(new_n19621_));
  AOI21_X1   g19364(.A1(new_n19620_), .A2(new_n19621_), .B(new_n4714_), .ZN(new_n19622_));
  NAND2_X1   g19365(.A1(new_n8550_), .A2(new_n19622_), .ZN(new_n19623_));
  XOR2_X1    g19366(.A1(new_n19623_), .A2(\a[47] ), .Z(new_n19624_));
  OAI21_X1   g19367(.A1(new_n19498_), .A2(new_n19574_), .B(new_n19576_), .ZN(new_n19625_));
  OAI22_X1   g19368(.A1(new_n5228_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n5225_), .ZN(new_n19626_));
  NAND2_X1   g19369(.A1(new_n5387_), .A2(\b[56] ), .ZN(new_n19627_));
  AOI21_X1   g19370(.A1(new_n19626_), .A2(new_n19627_), .B(new_n5231_), .ZN(new_n19628_));
  NAND2_X1   g19371(.A1(new_n7559_), .A2(new_n19628_), .ZN(new_n19629_));
  XOR2_X1    g19372(.A1(new_n19629_), .A2(\a[50] ), .Z(new_n19630_));
  NAND2_X1   g19373(.A1(new_n19565_), .A2(new_n19568_), .ZN(new_n19631_));
  NAND2_X1   g19374(.A1(new_n19631_), .A2(new_n19567_), .ZN(new_n19632_));
  OAI22_X1   g19375(.A1(new_n6721_), .A2(new_n5738_), .B1(new_n6723_), .B2(new_n5955_), .ZN(new_n19633_));
  NAND2_X1   g19376(.A1(new_n7617_), .A2(\b[50] ), .ZN(new_n19634_));
  AOI21_X1   g19377(.A1(new_n19634_), .A2(new_n19633_), .B(new_n6731_), .ZN(new_n19635_));
  NAND2_X1   g19378(.A1(new_n5954_), .A2(new_n19635_), .ZN(new_n19636_));
  XOR2_X1    g19379(.A1(new_n19636_), .A2(\a[56] ), .Z(new_n19637_));
  OAI21_X1   g19380(.A1(new_n19513_), .A2(new_n19532_), .B(new_n19534_), .ZN(new_n19638_));
  INV_X1     g19381(.I(new_n19638_), .ZN(new_n19639_));
  OAI22_X1   g19382(.A1(new_n4834_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n4509_), .ZN(new_n19640_));
  NAND2_X1   g19383(.A1(new_n9644_), .A2(\b[44] ), .ZN(new_n19641_));
  AOI21_X1   g19384(.A1(new_n19641_), .A2(new_n19640_), .B(new_n8321_), .ZN(new_n19642_));
  NAND2_X1   g19385(.A1(new_n4833_), .A2(new_n19642_), .ZN(new_n19643_));
  XOR2_X1    g19386(.A1(new_n19643_), .A2(new_n8309_), .Z(new_n19644_));
  NAND2_X1   g19387(.A1(new_n19526_), .A2(new_n19263_), .ZN(new_n19645_));
  NAND2_X1   g19388(.A1(new_n19645_), .A2(new_n19525_), .ZN(new_n19646_));
  NOR3_X1    g19389(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n4018_), .ZN(new_n19647_));
  NOR2_X1    g19390(.A1(new_n9364_), .A2(new_n4018_), .ZN(new_n19648_));
  NOR3_X1    g19391(.A1(new_n19648_), .A2(new_n4316_), .A3(new_n8985_), .ZN(new_n19649_));
  NOR2_X1    g19392(.A1(new_n19649_), .A2(new_n19647_), .ZN(new_n19650_));
  INV_X1     g19393(.I(new_n19650_), .ZN(new_n19651_));
  XOR2_X1    g19394(.A1(new_n19646_), .A2(new_n19651_), .Z(new_n19652_));
  INV_X1     g19395(.I(new_n19652_), .ZN(new_n19653_));
  NOR2_X1    g19396(.A1(new_n19646_), .A2(new_n19650_), .ZN(new_n19654_));
  INV_X1     g19397(.I(new_n19654_), .ZN(new_n19655_));
  NAND2_X1   g19398(.A1(new_n19646_), .A2(new_n19650_), .ZN(new_n19656_));
  AOI21_X1   g19399(.A1(new_n19655_), .A2(new_n19656_), .B(new_n19644_), .ZN(new_n19657_));
  AOI21_X1   g19400(.A1(new_n19644_), .A2(new_n19653_), .B(new_n19657_), .ZN(new_n19658_));
  INV_X1     g19401(.I(new_n19658_), .ZN(new_n19659_));
  OAI22_X1   g19402(.A1(new_n5197_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n5178_), .ZN(new_n19660_));
  NAND2_X1   g19403(.A1(new_n8628_), .A2(\b[47] ), .ZN(new_n19661_));
  AOI21_X1   g19404(.A1(new_n19661_), .A2(new_n19660_), .B(new_n7354_), .ZN(new_n19662_));
  NAND2_X1   g19405(.A1(new_n5196_), .A2(new_n19662_), .ZN(new_n19663_));
  XOR2_X1    g19406(.A1(new_n19663_), .A2(\a[59] ), .Z(new_n19664_));
  NOR2_X1    g19407(.A1(new_n19664_), .A2(new_n19659_), .ZN(new_n19665_));
  AND2_X2    g19408(.A1(new_n19664_), .A2(new_n19659_), .Z(new_n19666_));
  NOR2_X1    g19409(.A1(new_n19666_), .A2(new_n19665_), .ZN(new_n19667_));
  NOR2_X1    g19410(.A1(new_n19667_), .A2(new_n19639_), .ZN(new_n19668_));
  XOR2_X1    g19411(.A1(new_n19664_), .A2(new_n19658_), .Z(new_n19669_));
  NOR2_X1    g19412(.A1(new_n19669_), .A2(new_n19638_), .ZN(new_n19670_));
  NOR2_X1    g19413(.A1(new_n19668_), .A2(new_n19670_), .ZN(new_n19671_));
  INV_X1     g19414(.I(new_n19546_), .ZN(new_n19672_));
  OAI21_X1   g19415(.A1(new_n19544_), .A2(new_n19547_), .B(new_n19536_), .ZN(new_n19673_));
  NAND2_X1   g19416(.A1(new_n19672_), .A2(new_n19673_), .ZN(new_n19674_));
  INV_X1     g19417(.I(new_n19674_), .ZN(new_n19675_));
  NOR2_X1    g19418(.A1(new_n19675_), .A2(new_n19671_), .ZN(new_n19676_));
  NOR3_X1    g19419(.A1(new_n19674_), .A2(new_n19668_), .A3(new_n19670_), .ZN(new_n19677_));
  NOR2_X1    g19420(.A1(new_n19676_), .A2(new_n19677_), .ZN(new_n19678_));
  NOR2_X1    g19421(.A1(new_n19678_), .A2(new_n19637_), .ZN(new_n19679_));
  INV_X1     g19422(.I(new_n19637_), .ZN(new_n19680_));
  XOR2_X1    g19423(.A1(new_n19674_), .A2(new_n19671_), .Z(new_n19681_));
  NOR2_X1    g19424(.A1(new_n19681_), .A2(new_n19680_), .ZN(new_n19682_));
  NOR2_X1    g19425(.A1(new_n19679_), .A2(new_n19682_), .ZN(new_n19683_));
  INV_X1     g19426(.I(new_n19552_), .ZN(new_n19684_));
  AOI21_X1   g19427(.A1(new_n19684_), .A2(new_n19505_), .B(new_n19554_), .ZN(new_n19685_));
  OAI22_X1   g19428(.A1(new_n5786_), .A2(new_n6467_), .B1(new_n6238_), .B2(new_n5792_), .ZN(new_n19686_));
  NAND2_X1   g19429(.A1(new_n6745_), .A2(\b[53] ), .ZN(new_n19687_));
  AOI21_X1   g19430(.A1(new_n19687_), .A2(new_n19686_), .B(new_n5796_), .ZN(new_n19688_));
  NAND2_X1   g19431(.A1(new_n6471_), .A2(new_n19688_), .ZN(new_n19689_));
  XOR2_X1    g19432(.A1(new_n19689_), .A2(\a[53] ), .Z(new_n19690_));
  NOR2_X1    g19433(.A1(new_n19685_), .A2(new_n19690_), .ZN(new_n19691_));
  AND2_X2    g19434(.A1(new_n19685_), .A2(new_n19690_), .Z(new_n19692_));
  NOR2_X1    g19435(.A1(new_n19692_), .A2(new_n19691_), .ZN(new_n19693_));
  NOR2_X1    g19436(.A1(new_n19693_), .A2(new_n19683_), .ZN(new_n19694_));
  INV_X1     g19437(.I(new_n19683_), .ZN(new_n19695_));
  XNOR2_X1   g19438(.A1(new_n19685_), .A2(new_n19690_), .ZN(new_n19696_));
  NOR2_X1    g19439(.A1(new_n19696_), .A2(new_n19695_), .ZN(new_n19697_));
  NOR2_X1    g19440(.A1(new_n19694_), .A2(new_n19697_), .ZN(new_n19698_));
  XOR2_X1    g19441(.A1(new_n19632_), .A2(new_n19698_), .Z(new_n19699_));
  NOR2_X1    g19442(.A1(new_n19699_), .A2(new_n19630_), .ZN(new_n19700_));
  INV_X1     g19443(.I(new_n19630_), .ZN(new_n19701_));
  INV_X1     g19444(.I(new_n19632_), .ZN(new_n19702_));
  NOR2_X1    g19445(.A1(new_n19702_), .A2(new_n19698_), .ZN(new_n19703_));
  INV_X1     g19446(.I(new_n19703_), .ZN(new_n19704_));
  NAND2_X1   g19447(.A1(new_n19702_), .A2(new_n19698_), .ZN(new_n19705_));
  AOI21_X1   g19448(.A1(new_n19704_), .A2(new_n19705_), .B(new_n19701_), .ZN(new_n19706_));
  NOR2_X1    g19449(.A1(new_n19706_), .A2(new_n19700_), .ZN(new_n19707_));
  NOR2_X1    g19450(.A1(new_n19707_), .A2(new_n19625_), .ZN(new_n19708_));
  INV_X1     g19451(.I(new_n19708_), .ZN(new_n19709_));
  NAND2_X1   g19452(.A1(new_n19707_), .A2(new_n19625_), .ZN(new_n19710_));
  AOI21_X1   g19453(.A1(new_n19709_), .A2(new_n19710_), .B(new_n19624_), .ZN(new_n19711_));
  XNOR2_X1   g19454(.A1(new_n19707_), .A2(new_n19625_), .ZN(new_n19712_));
  INV_X1     g19455(.I(new_n19712_), .ZN(new_n19713_));
  AOI21_X1   g19456(.A1(new_n19713_), .A2(new_n19624_), .B(new_n19711_), .ZN(new_n19714_));
  NOR2_X1    g19457(.A1(new_n19714_), .A2(new_n19619_), .ZN(new_n19715_));
  INV_X1     g19458(.I(new_n19715_), .ZN(new_n19716_));
  NAND2_X1   g19459(.A1(new_n19714_), .A2(new_n19619_), .ZN(new_n19717_));
  AOI21_X1   g19460(.A1(new_n19716_), .A2(new_n19717_), .B(new_n19617_), .ZN(new_n19718_));
  INV_X1     g19461(.I(new_n19617_), .ZN(new_n19719_));
  XNOR2_X1   g19462(.A1(new_n19714_), .A2(new_n19619_), .ZN(new_n19720_));
  NOR2_X1    g19463(.A1(new_n19720_), .A2(new_n19719_), .ZN(new_n19721_));
  NOR2_X1    g19464(.A1(new_n19721_), .A2(new_n19718_), .ZN(new_n19722_));
  OAI21_X1   g19465(.A1(new_n19494_), .A2(new_n19598_), .B(new_n19600_), .ZN(new_n19723_));
  NAND2_X1   g19466(.A1(new_n19610_), .A2(new_n19607_), .ZN(new_n19724_));
  INV_X1     g19467(.I(new_n19724_), .ZN(new_n19725_));
  NOR3_X1    g19468(.A1(new_n19372_), .A2(new_n19374_), .A3(new_n19725_), .ZN(new_n19726_));
  NOR3_X1    g19469(.A1(new_n19602_), .A2(new_n19603_), .A3(new_n19605_), .ZN(new_n19727_));
  NOR2_X1    g19470(.A1(new_n19726_), .A2(new_n19727_), .ZN(new_n19728_));
  XOR2_X1    g19471(.A1(new_n19728_), .A2(new_n19723_), .Z(new_n19729_));
  XOR2_X1    g19472(.A1(new_n19729_), .A2(new_n19722_), .Z(\f[106] ));
  NOR2_X1    g19473(.A1(new_n19722_), .A2(new_n19723_), .ZN(new_n19731_));
  INV_X1     g19474(.I(new_n19731_), .ZN(new_n19732_));
  XOR2_X1    g19475(.A1(new_n19722_), .A2(new_n19723_), .Z(new_n19733_));
  NOR2_X1    g19476(.A1(new_n19727_), .A2(new_n19733_), .ZN(new_n19734_));
  INV_X1     g19477(.I(new_n19734_), .ZN(new_n19735_));
  OAI21_X1   g19478(.A1(new_n19726_), .A2(new_n19735_), .B(new_n19732_), .ZN(new_n19736_));
  AOI21_X1   g19479(.A1(new_n19719_), .A2(new_n19717_), .B(new_n19715_), .ZN(new_n19737_));
  OAI21_X1   g19480(.A1(new_n19624_), .A2(new_n19708_), .B(new_n19710_), .ZN(new_n19738_));
  OAI22_X1   g19481(.A1(new_n9595_), .A2(new_n4211_), .B1(new_n8956_), .B2(new_n4362_), .ZN(new_n19739_));
  OAI22_X1   g19482(.A1(new_n4711_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n4706_), .ZN(new_n19740_));
  NAND2_X1   g19483(.A1(new_n5814_), .A2(\b[60] ), .ZN(new_n19741_));
  AOI21_X1   g19484(.A1(new_n19740_), .A2(new_n19741_), .B(new_n4714_), .ZN(new_n19742_));
  NAND2_X1   g19485(.A1(new_n8935_), .A2(new_n19742_), .ZN(new_n19743_));
  XOR2_X1    g19486(.A1(new_n19743_), .A2(\a[47] ), .Z(new_n19744_));
  OAI22_X1   g19487(.A1(new_n5786_), .A2(new_n6995_), .B1(new_n6467_), .B2(new_n5792_), .ZN(new_n19745_));
  NAND2_X1   g19488(.A1(new_n6745_), .A2(\b[54] ), .ZN(new_n19746_));
  AOI21_X1   g19489(.A1(new_n19746_), .A2(new_n19745_), .B(new_n5796_), .ZN(new_n19747_));
  NAND2_X1   g19490(.A1(new_n6994_), .A2(new_n19747_), .ZN(new_n19748_));
  XOR2_X1    g19491(.A1(new_n19748_), .A2(\a[53] ), .Z(new_n19749_));
  INV_X1     g19492(.I(new_n19677_), .ZN(new_n19750_));
  AOI21_X1   g19493(.A1(new_n19750_), .A2(new_n19680_), .B(new_n19676_), .ZN(new_n19751_));
  OAI22_X1   g19494(.A1(new_n6721_), .A2(new_n5955_), .B1(new_n6723_), .B2(new_n6215_), .ZN(new_n19752_));
  NAND2_X1   g19495(.A1(new_n7617_), .A2(\b[51] ), .ZN(new_n19753_));
  AOI21_X1   g19496(.A1(new_n19753_), .A2(new_n19752_), .B(new_n6731_), .ZN(new_n19754_));
  NAND2_X1   g19497(.A1(new_n6219_), .A2(new_n19754_), .ZN(new_n19755_));
  XOR2_X1    g19498(.A1(new_n19755_), .A2(\a[56] ), .Z(new_n19756_));
  OAI22_X1   g19499(.A1(new_n5538_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n5197_), .ZN(new_n19757_));
  NAND2_X1   g19500(.A1(new_n8628_), .A2(\b[48] ), .ZN(new_n19758_));
  AOI21_X1   g19501(.A1(new_n19758_), .A2(new_n19757_), .B(new_n7354_), .ZN(new_n19759_));
  NAND2_X1   g19502(.A1(new_n5537_), .A2(new_n19759_), .ZN(new_n19760_));
  XOR2_X1    g19503(.A1(new_n19760_), .A2(\a[59] ), .Z(new_n19761_));
  INV_X1     g19504(.I(new_n19656_), .ZN(new_n19762_));
  AOI21_X1   g19505(.A1(new_n19644_), .A2(new_n19655_), .B(new_n19762_), .ZN(new_n19763_));
  OAI22_X1   g19506(.A1(new_n4997_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n4834_), .ZN(new_n19764_));
  NAND2_X1   g19507(.A1(new_n9644_), .A2(\b[45] ), .ZN(new_n19765_));
  AOI21_X1   g19508(.A1(new_n19765_), .A2(new_n19764_), .B(new_n8321_), .ZN(new_n19766_));
  NAND2_X1   g19509(.A1(new_n5004_), .A2(new_n19766_), .ZN(new_n19767_));
  XOR2_X1    g19510(.A1(new_n19767_), .A2(\a[62] ), .Z(new_n19768_));
  NOR2_X1    g19511(.A1(new_n8985_), .A2(new_n4501_), .ZN(new_n19769_));
  NOR2_X1    g19512(.A1(new_n9364_), .A2(new_n4316_), .ZN(new_n19770_));
  XNOR2_X1   g19513(.A1(new_n19769_), .A2(new_n19770_), .ZN(new_n19771_));
  XOR2_X1    g19514(.A1(new_n19771_), .A2(new_n19650_), .Z(new_n19772_));
  NOR2_X1    g19515(.A1(new_n19768_), .A2(new_n19772_), .ZN(new_n19773_));
  NOR2_X1    g19516(.A1(new_n19651_), .A2(new_n19771_), .ZN(new_n19774_));
  INV_X1     g19517(.I(new_n19774_), .ZN(new_n19775_));
  NAND2_X1   g19518(.A1(new_n19651_), .A2(new_n19771_), .ZN(new_n19776_));
  NAND2_X1   g19519(.A1(new_n19775_), .A2(new_n19776_), .ZN(new_n19777_));
  AOI21_X1   g19520(.A1(new_n19768_), .A2(new_n19777_), .B(new_n19773_), .ZN(new_n19778_));
  XOR2_X1    g19521(.A1(new_n19778_), .A2(new_n19763_), .Z(new_n19779_));
  NOR2_X1    g19522(.A1(new_n19779_), .A2(new_n19761_), .ZN(new_n19780_));
  INV_X1     g19523(.I(new_n19761_), .ZN(new_n19781_));
  INV_X1     g19524(.I(new_n19763_), .ZN(new_n19782_));
  NOR2_X1    g19525(.A1(new_n19778_), .A2(new_n19782_), .ZN(new_n19783_));
  INV_X1     g19526(.I(new_n19783_), .ZN(new_n19784_));
  NAND2_X1   g19527(.A1(new_n19778_), .A2(new_n19782_), .ZN(new_n19785_));
  AOI21_X1   g19528(.A1(new_n19784_), .A2(new_n19785_), .B(new_n19781_), .ZN(new_n19786_));
  NOR2_X1    g19529(.A1(new_n19780_), .A2(new_n19786_), .ZN(new_n19787_));
  NOR2_X1    g19530(.A1(new_n19666_), .A2(new_n19639_), .ZN(new_n19788_));
  NOR2_X1    g19531(.A1(new_n19788_), .A2(new_n19665_), .ZN(new_n19789_));
  XOR2_X1    g19532(.A1(new_n19787_), .A2(new_n19789_), .Z(new_n19790_));
  NOR2_X1    g19533(.A1(new_n19790_), .A2(new_n19756_), .ZN(new_n19791_));
  INV_X1     g19534(.I(new_n19756_), .ZN(new_n19792_));
  INV_X1     g19535(.I(new_n19787_), .ZN(new_n19793_));
  NOR2_X1    g19536(.A1(new_n19793_), .A2(new_n19789_), .ZN(new_n19794_));
  INV_X1     g19537(.I(new_n19794_), .ZN(new_n19795_));
  NAND2_X1   g19538(.A1(new_n19793_), .A2(new_n19789_), .ZN(new_n19796_));
  AOI21_X1   g19539(.A1(new_n19795_), .A2(new_n19796_), .B(new_n19792_), .ZN(new_n19797_));
  NOR2_X1    g19540(.A1(new_n19797_), .A2(new_n19791_), .ZN(new_n19798_));
  XOR2_X1    g19541(.A1(new_n19798_), .A2(new_n19751_), .Z(new_n19799_));
  NOR2_X1    g19542(.A1(new_n19799_), .A2(new_n19749_), .ZN(new_n19800_));
  INV_X1     g19543(.I(new_n19749_), .ZN(new_n19801_));
  INV_X1     g19544(.I(new_n19751_), .ZN(new_n19802_));
  NOR2_X1    g19545(.A1(new_n19798_), .A2(new_n19802_), .ZN(new_n19803_));
  INV_X1     g19546(.I(new_n19803_), .ZN(new_n19804_));
  NAND2_X1   g19547(.A1(new_n19798_), .A2(new_n19802_), .ZN(new_n19805_));
  AOI21_X1   g19548(.A1(new_n19804_), .A2(new_n19805_), .B(new_n19801_), .ZN(new_n19806_));
  NOR2_X1    g19549(.A1(new_n19800_), .A2(new_n19806_), .ZN(new_n19807_));
  OAI22_X1   g19550(.A1(new_n5228_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n5225_), .ZN(new_n19808_));
  NAND2_X1   g19551(.A1(new_n5387_), .A2(\b[57] ), .ZN(new_n19809_));
  AOI21_X1   g19552(.A1(new_n19808_), .A2(new_n19809_), .B(new_n5231_), .ZN(new_n19810_));
  NAND2_X1   g19553(.A1(new_n7895_), .A2(new_n19810_), .ZN(new_n19811_));
  XOR2_X1    g19554(.A1(new_n19811_), .A2(\a[50] ), .Z(new_n19812_));
  NOR2_X1    g19555(.A1(new_n19692_), .A2(new_n19683_), .ZN(new_n19813_));
  NOR2_X1    g19556(.A1(new_n19813_), .A2(new_n19691_), .ZN(new_n19814_));
  XNOR2_X1   g19557(.A1(new_n19814_), .A2(new_n19812_), .ZN(new_n19815_));
  NOR2_X1    g19558(.A1(new_n19815_), .A2(new_n19807_), .ZN(new_n19816_));
  INV_X1     g19559(.I(new_n19807_), .ZN(new_n19817_));
  NOR2_X1    g19560(.A1(new_n19814_), .A2(new_n19812_), .ZN(new_n19818_));
  INV_X1     g19561(.I(new_n19818_), .ZN(new_n19819_));
  NAND2_X1   g19562(.A1(new_n19814_), .A2(new_n19812_), .ZN(new_n19820_));
  AOI21_X1   g19563(.A1(new_n19819_), .A2(new_n19820_), .B(new_n19817_), .ZN(new_n19821_));
  NOR2_X1    g19564(.A1(new_n19821_), .A2(new_n19816_), .ZN(new_n19822_));
  NAND2_X1   g19565(.A1(new_n19705_), .A2(new_n19701_), .ZN(new_n19823_));
  NAND2_X1   g19566(.A1(new_n19823_), .A2(new_n19704_), .ZN(new_n19824_));
  INV_X1     g19567(.I(new_n19824_), .ZN(new_n19825_));
  NOR2_X1    g19568(.A1(new_n19825_), .A2(new_n19822_), .ZN(new_n19826_));
  NOR3_X1    g19569(.A1(new_n19824_), .A2(new_n19816_), .A3(new_n19821_), .ZN(new_n19827_));
  NOR2_X1    g19570(.A1(new_n19826_), .A2(new_n19827_), .ZN(new_n19828_));
  NOR2_X1    g19571(.A1(new_n19828_), .A2(new_n19744_), .ZN(new_n19829_));
  INV_X1     g19572(.I(new_n19744_), .ZN(new_n19830_));
  XOR2_X1    g19573(.A1(new_n19822_), .A2(new_n19824_), .Z(new_n19831_));
  NOR2_X1    g19574(.A1(new_n19831_), .A2(new_n19830_), .ZN(new_n19832_));
  NOR2_X1    g19575(.A1(new_n19832_), .A2(new_n19829_), .ZN(new_n19833_));
  XOR2_X1    g19576(.A1(new_n19833_), .A2(new_n19739_), .Z(new_n19834_));
  XOR2_X1    g19577(.A1(new_n19834_), .A2(\a[44] ), .Z(new_n19835_));
  XOR2_X1    g19578(.A1(new_n19835_), .A2(new_n19738_), .Z(new_n19836_));
  XOR2_X1    g19579(.A1(new_n19836_), .A2(new_n19737_), .Z(new_n19837_));
  NAND2_X1   g19580(.A1(new_n19736_), .A2(new_n19837_), .ZN(new_n19838_));
  XOR2_X1    g19581(.A1(new_n19836_), .A2(new_n19737_), .Z(new_n19839_));
  OAI21_X1   g19582(.A1(new_n19736_), .A2(new_n19839_), .B(new_n19838_), .ZN(\f[107] ));
  OAI22_X1   g19583(.A1(new_n4711_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n4706_), .ZN(new_n19841_));
  NAND2_X1   g19584(.A1(new_n5814_), .A2(\b[61] ), .ZN(new_n19842_));
  AOI21_X1   g19585(.A1(new_n19841_), .A2(new_n19842_), .B(new_n4714_), .ZN(new_n19843_));
  NAND2_X1   g19586(.A1(new_n8963_), .A2(new_n19843_), .ZN(new_n19844_));
  XOR2_X1    g19587(.A1(new_n19844_), .A2(\a[47] ), .Z(new_n19845_));
  INV_X1     g19588(.I(new_n19827_), .ZN(new_n19846_));
  AOI21_X1   g19589(.A1(new_n19846_), .A2(new_n19830_), .B(new_n19826_), .ZN(new_n19847_));
  AOI21_X1   g19590(.A1(new_n19807_), .A2(new_n19820_), .B(new_n19818_), .ZN(new_n19848_));
  OAI22_X1   g19591(.A1(new_n5228_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n5225_), .ZN(new_n19849_));
  NAND2_X1   g19592(.A1(new_n5387_), .A2(\b[58] ), .ZN(new_n19850_));
  AOI21_X1   g19593(.A1(new_n19849_), .A2(new_n19850_), .B(new_n5231_), .ZN(new_n19851_));
  NAND2_X1   g19594(.A1(new_n7929_), .A2(new_n19851_), .ZN(new_n19852_));
  XOR2_X1    g19595(.A1(new_n19852_), .A2(\a[50] ), .Z(new_n19853_));
  OAI21_X1   g19596(.A1(new_n19749_), .A2(new_n19803_), .B(new_n19805_), .ZN(new_n19854_));
  INV_X1     g19597(.I(new_n19854_), .ZN(new_n19855_));
  OAI22_X1   g19598(.A1(new_n5786_), .A2(new_n7305_), .B1(new_n6995_), .B2(new_n5792_), .ZN(new_n19856_));
  NAND2_X1   g19599(.A1(new_n6745_), .A2(\b[55] ), .ZN(new_n19857_));
  AOI21_X1   g19600(.A1(new_n19857_), .A2(new_n19856_), .B(new_n5796_), .ZN(new_n19858_));
  NAND2_X1   g19601(.A1(new_n7308_), .A2(new_n19858_), .ZN(new_n19859_));
  XOR2_X1    g19602(.A1(new_n19859_), .A2(\a[53] ), .Z(new_n19860_));
  AOI21_X1   g19603(.A1(new_n19792_), .A2(new_n19796_), .B(new_n19794_), .ZN(new_n19861_));
  OAI22_X1   g19604(.A1(new_n6721_), .A2(new_n6215_), .B1(new_n6723_), .B2(new_n6238_), .ZN(new_n19862_));
  NAND2_X1   g19605(.A1(new_n7617_), .A2(\b[52] ), .ZN(new_n19863_));
  AOI21_X1   g19606(.A1(new_n19863_), .A2(new_n19862_), .B(new_n6731_), .ZN(new_n19864_));
  NAND2_X1   g19607(.A1(new_n6237_), .A2(new_n19864_), .ZN(new_n19865_));
  XOR2_X1    g19608(.A1(new_n19865_), .A2(\a[56] ), .Z(new_n19866_));
  OAI21_X1   g19609(.A1(new_n19761_), .A2(new_n19783_), .B(new_n19785_), .ZN(new_n19867_));
  INV_X1     g19610(.I(new_n19768_), .ZN(new_n19868_));
  NAND2_X1   g19611(.A1(new_n19868_), .A2(new_n19776_), .ZN(new_n19869_));
  NAND2_X1   g19612(.A1(new_n19869_), .A2(new_n19775_), .ZN(new_n19870_));
  OAI22_X1   g19613(.A1(new_n5178_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n4997_), .ZN(new_n19871_));
  NAND2_X1   g19614(.A1(new_n9644_), .A2(\b[46] ), .ZN(new_n19872_));
  AOI21_X1   g19615(.A1(new_n19872_), .A2(new_n19871_), .B(new_n8321_), .ZN(new_n19873_));
  NAND2_X1   g19616(.A1(new_n5177_), .A2(new_n19873_), .ZN(new_n19874_));
  XOR2_X1    g19617(.A1(new_n19874_), .A2(\a[62] ), .Z(new_n19875_));
  NOR2_X1    g19618(.A1(new_n8985_), .A2(new_n4509_), .ZN(new_n19876_));
  NOR2_X1    g19619(.A1(new_n9364_), .A2(new_n4501_), .ZN(new_n19877_));
  XNOR2_X1   g19620(.A1(new_n19876_), .A2(new_n19877_), .ZN(new_n19878_));
  NOR2_X1    g19621(.A1(new_n19878_), .A2(new_n4198_), .ZN(new_n19879_));
  INV_X1     g19622(.I(new_n19879_), .ZN(new_n19880_));
  NAND2_X1   g19623(.A1(new_n19878_), .A2(new_n4198_), .ZN(new_n19881_));
  AOI21_X1   g19624(.A1(new_n19880_), .A2(new_n19881_), .B(new_n19650_), .ZN(new_n19882_));
  XOR2_X1    g19625(.A1(new_n19878_), .A2(\a[44] ), .Z(new_n19883_));
  NOR2_X1    g19626(.A1(new_n19883_), .A2(new_n19651_), .ZN(new_n19884_));
  NOR2_X1    g19627(.A1(new_n19884_), .A2(new_n19882_), .ZN(new_n19885_));
  OR2_X2     g19628(.A1(new_n19875_), .A2(new_n19885_), .Z(new_n19886_));
  NAND2_X1   g19629(.A1(new_n19875_), .A2(new_n19885_), .ZN(new_n19887_));
  NAND2_X1   g19630(.A1(new_n19886_), .A2(new_n19887_), .ZN(new_n19888_));
  XNOR2_X1   g19631(.A1(new_n19875_), .A2(new_n19885_), .ZN(new_n19889_));
  NOR2_X1    g19632(.A1(new_n19870_), .A2(new_n19889_), .ZN(new_n19890_));
  AOI21_X1   g19633(.A1(new_n19870_), .A2(new_n19888_), .B(new_n19890_), .ZN(new_n19891_));
  OAI22_X1   g19634(.A1(new_n5738_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n5538_), .ZN(new_n19892_));
  NAND2_X1   g19635(.A1(new_n8628_), .A2(\b[49] ), .ZN(new_n19893_));
  AOI21_X1   g19636(.A1(new_n19893_), .A2(new_n19892_), .B(new_n7354_), .ZN(new_n19894_));
  NAND2_X1   g19637(.A1(new_n5741_), .A2(new_n19894_), .ZN(new_n19895_));
  XOR2_X1    g19638(.A1(new_n19895_), .A2(\a[59] ), .Z(new_n19896_));
  XNOR2_X1   g19639(.A1(new_n19891_), .A2(new_n19896_), .ZN(new_n19897_));
  INV_X1     g19640(.I(new_n19897_), .ZN(new_n19898_));
  NOR2_X1    g19641(.A1(new_n19891_), .A2(new_n19896_), .ZN(new_n19899_));
  INV_X1     g19642(.I(new_n19899_), .ZN(new_n19900_));
  NAND2_X1   g19643(.A1(new_n19891_), .A2(new_n19896_), .ZN(new_n19901_));
  AOI21_X1   g19644(.A1(new_n19900_), .A2(new_n19901_), .B(new_n19867_), .ZN(new_n19902_));
  AOI21_X1   g19645(.A1(new_n19898_), .A2(new_n19867_), .B(new_n19902_), .ZN(new_n19903_));
  XOR2_X1    g19646(.A1(new_n19903_), .A2(new_n19866_), .Z(new_n19904_));
  NOR2_X1    g19647(.A1(new_n19904_), .A2(new_n19861_), .ZN(new_n19905_));
  INV_X1     g19648(.I(new_n19866_), .ZN(new_n19906_));
  NOR2_X1    g19649(.A1(new_n19903_), .A2(new_n19906_), .ZN(new_n19907_));
  INV_X1     g19650(.I(new_n19907_), .ZN(new_n19908_));
  NAND2_X1   g19651(.A1(new_n19903_), .A2(new_n19906_), .ZN(new_n19909_));
  NAND2_X1   g19652(.A1(new_n19908_), .A2(new_n19909_), .ZN(new_n19910_));
  AOI21_X1   g19653(.A1(new_n19861_), .A2(new_n19910_), .B(new_n19905_), .ZN(new_n19911_));
  XOR2_X1    g19654(.A1(new_n19911_), .A2(new_n19860_), .Z(new_n19912_));
  NOR2_X1    g19655(.A1(new_n19912_), .A2(new_n19855_), .ZN(new_n19913_));
  INV_X1     g19656(.I(new_n19860_), .ZN(new_n19914_));
  NOR2_X1    g19657(.A1(new_n19911_), .A2(new_n19914_), .ZN(new_n19915_));
  INV_X1     g19658(.I(new_n19915_), .ZN(new_n19916_));
  NAND2_X1   g19659(.A1(new_n19911_), .A2(new_n19914_), .ZN(new_n19917_));
  AOI21_X1   g19660(.A1(new_n19916_), .A2(new_n19917_), .B(new_n19854_), .ZN(new_n19918_));
  NOR2_X1    g19661(.A1(new_n19913_), .A2(new_n19918_), .ZN(new_n19919_));
  XOR2_X1    g19662(.A1(new_n19919_), .A2(new_n19853_), .Z(new_n19920_));
  NOR2_X1    g19663(.A1(new_n19920_), .A2(new_n19848_), .ZN(new_n19921_));
  INV_X1     g19664(.I(new_n19853_), .ZN(new_n19922_));
  NOR2_X1    g19665(.A1(new_n19919_), .A2(new_n19922_), .ZN(new_n19923_));
  INV_X1     g19666(.I(new_n19923_), .ZN(new_n19924_));
  NAND2_X1   g19667(.A1(new_n19919_), .A2(new_n19922_), .ZN(new_n19925_));
  NAND2_X1   g19668(.A1(new_n19924_), .A2(new_n19925_), .ZN(new_n19926_));
  AOI21_X1   g19669(.A1(new_n19848_), .A2(new_n19926_), .B(new_n19921_), .ZN(new_n19927_));
  XOR2_X1    g19670(.A1(new_n19927_), .A2(new_n19847_), .Z(new_n19928_));
  NOR2_X1    g19671(.A1(new_n19928_), .A2(new_n19845_), .ZN(new_n19929_));
  INV_X1     g19672(.I(new_n19847_), .ZN(new_n19930_));
  NOR2_X1    g19673(.A1(new_n19927_), .A2(new_n19930_), .ZN(new_n19931_));
  INV_X1     g19674(.I(new_n19931_), .ZN(new_n19932_));
  NAND2_X1   g19675(.A1(new_n19927_), .A2(new_n19930_), .ZN(new_n19933_));
  NAND2_X1   g19676(.A1(new_n19932_), .A2(new_n19933_), .ZN(new_n19934_));
  AOI21_X1   g19677(.A1(new_n19845_), .A2(new_n19934_), .B(new_n19929_), .ZN(new_n19935_));
  INV_X1     g19678(.I(new_n19738_), .ZN(new_n19936_));
  NOR2_X1    g19679(.A1(new_n19833_), .A2(new_n19936_), .ZN(new_n19937_));
  XOR2_X1    g19680(.A1(new_n19739_), .A2(new_n4198_), .Z(new_n19938_));
  AOI21_X1   g19681(.A1(new_n19833_), .A2(new_n19936_), .B(new_n19938_), .ZN(new_n19939_));
  NOR2_X1    g19682(.A1(new_n19939_), .A2(new_n19937_), .ZN(new_n19940_));
  XOR2_X1    g19683(.A1(new_n19935_), .A2(new_n19940_), .Z(new_n19941_));
  INV_X1     g19684(.I(new_n19941_), .ZN(new_n19942_));
  INV_X1     g19685(.I(new_n19737_), .ZN(new_n19943_));
  NAND2_X1   g19686(.A1(new_n19736_), .A2(new_n19943_), .ZN(new_n19944_));
  XOR2_X1    g19687(.A1(new_n19944_), .A2(new_n19942_), .Z(new_n19945_));
  INV_X1     g19688(.I(new_n19836_), .ZN(new_n19946_));
  XOR2_X1    g19689(.A1(new_n19736_), .A2(new_n19943_), .Z(new_n19947_));
  NAND2_X1   g19690(.A1(new_n19947_), .A2(new_n19946_), .ZN(new_n19948_));
  XOR2_X1    g19691(.A1(new_n19945_), .A2(new_n19948_), .Z(\f[108] ));
  NOR2_X1    g19692(.A1(new_n4873_), .A2(new_n8932_), .ZN(new_n19950_));
  NOR2_X1    g19693(.A1(new_n4706_), .A2(new_n8956_), .ZN(new_n19951_));
  NOR4_X1    g19694(.A1(new_n9323_), .A2(new_n4714_), .A3(new_n19950_), .A4(new_n19951_), .ZN(new_n19952_));
  XOR2_X1    g19695(.A1(new_n19952_), .A2(new_n4701_), .Z(new_n19953_));
  OAI21_X1   g19696(.A1(new_n19848_), .A2(new_n19923_), .B(new_n19925_), .ZN(new_n19954_));
  INV_X1     g19697(.I(new_n19954_), .ZN(new_n19955_));
  OAI22_X1   g19698(.A1(new_n5228_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n5225_), .ZN(new_n19956_));
  NAND2_X1   g19699(.A1(new_n5387_), .A2(\b[59] ), .ZN(new_n19957_));
  AOI21_X1   g19700(.A1(new_n19956_), .A2(new_n19957_), .B(new_n5231_), .ZN(new_n19958_));
  NAND2_X1   g19701(.A1(new_n8550_), .A2(new_n19958_), .ZN(new_n19959_));
  XOR2_X1    g19702(.A1(new_n19959_), .A2(\a[50] ), .Z(new_n19960_));
  OAI21_X1   g19703(.A1(new_n19855_), .A2(new_n19915_), .B(new_n19917_), .ZN(new_n19961_));
  OAI22_X1   g19704(.A1(new_n5786_), .A2(new_n7560_), .B1(new_n7305_), .B2(new_n5792_), .ZN(new_n19962_));
  NAND2_X1   g19705(.A1(new_n6745_), .A2(\b[56] ), .ZN(new_n19963_));
  AOI21_X1   g19706(.A1(new_n19963_), .A2(new_n19962_), .B(new_n5796_), .ZN(new_n19964_));
  NAND2_X1   g19707(.A1(new_n7559_), .A2(new_n19964_), .ZN(new_n19965_));
  XOR2_X1    g19708(.A1(new_n19965_), .A2(\a[53] ), .Z(new_n19966_));
  OAI21_X1   g19709(.A1(new_n19861_), .A2(new_n19907_), .B(new_n19909_), .ZN(new_n19967_));
  AOI21_X1   g19710(.A1(new_n19867_), .A2(new_n19901_), .B(new_n19899_), .ZN(new_n19968_));
  OAI22_X1   g19711(.A1(new_n5955_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n5738_), .ZN(new_n19969_));
  NAND2_X1   g19712(.A1(new_n8628_), .A2(\b[50] ), .ZN(new_n19970_));
  AOI21_X1   g19713(.A1(new_n19970_), .A2(new_n19969_), .B(new_n7354_), .ZN(new_n19971_));
  NAND2_X1   g19714(.A1(new_n5954_), .A2(new_n19971_), .ZN(new_n19972_));
  XOR2_X1    g19715(.A1(new_n19972_), .A2(\a[59] ), .Z(new_n19973_));
  NAND2_X1   g19716(.A1(new_n19870_), .A2(new_n19887_), .ZN(new_n19974_));
  NAND2_X1   g19717(.A1(new_n19974_), .A2(new_n19886_), .ZN(new_n19975_));
  OAI22_X1   g19718(.A1(new_n5197_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n5178_), .ZN(new_n19976_));
  NAND2_X1   g19719(.A1(new_n9644_), .A2(\b[47] ), .ZN(new_n19977_));
  AOI21_X1   g19720(.A1(new_n19977_), .A2(new_n19976_), .B(new_n8321_), .ZN(new_n19978_));
  NAND2_X1   g19721(.A1(new_n5196_), .A2(new_n19978_), .ZN(new_n19979_));
  XOR2_X1    g19722(.A1(new_n19979_), .A2(\a[62] ), .Z(new_n19980_));
  NAND2_X1   g19723(.A1(new_n19881_), .A2(new_n19651_), .ZN(new_n19981_));
  NAND2_X1   g19724(.A1(new_n19981_), .A2(new_n19880_), .ZN(new_n19982_));
  NOR3_X1    g19725(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n4509_), .ZN(new_n19983_));
  NOR2_X1    g19726(.A1(new_n9364_), .A2(new_n4509_), .ZN(new_n19984_));
  NOR3_X1    g19727(.A1(new_n19984_), .A2(new_n4834_), .A3(new_n8985_), .ZN(new_n19985_));
  NOR2_X1    g19728(.A1(new_n19985_), .A2(new_n19983_), .ZN(new_n19986_));
  INV_X1     g19729(.I(new_n19986_), .ZN(new_n19987_));
  XOR2_X1    g19730(.A1(new_n19982_), .A2(new_n19987_), .Z(new_n19988_));
  OR2_X2     g19731(.A1(new_n19980_), .A2(new_n19988_), .Z(new_n19989_));
  NOR2_X1    g19732(.A1(new_n19982_), .A2(new_n19986_), .ZN(new_n19990_));
  NAND2_X1   g19733(.A1(new_n19982_), .A2(new_n19986_), .ZN(new_n19991_));
  INV_X1     g19734(.I(new_n19991_), .ZN(new_n19992_));
  OAI21_X1   g19735(.A1(new_n19990_), .A2(new_n19992_), .B(new_n19980_), .ZN(new_n19993_));
  NAND2_X1   g19736(.A1(new_n19989_), .A2(new_n19993_), .ZN(new_n19994_));
  XOR2_X1    g19737(.A1(new_n19975_), .A2(new_n19994_), .Z(new_n19995_));
  NOR2_X1    g19738(.A1(new_n19995_), .A2(new_n19973_), .ZN(new_n19996_));
  INV_X1     g19739(.I(new_n19973_), .ZN(new_n19997_));
  INV_X1     g19740(.I(new_n19994_), .ZN(new_n19998_));
  NOR2_X1    g19741(.A1(new_n19998_), .A2(new_n19975_), .ZN(new_n19999_));
  INV_X1     g19742(.I(new_n19999_), .ZN(new_n20000_));
  NAND2_X1   g19743(.A1(new_n19998_), .A2(new_n19975_), .ZN(new_n20001_));
  AOI21_X1   g19744(.A1(new_n20000_), .A2(new_n20001_), .B(new_n19997_), .ZN(new_n20002_));
  NOR2_X1    g19745(.A1(new_n19996_), .A2(new_n20002_), .ZN(new_n20003_));
  INV_X1     g19746(.I(new_n20003_), .ZN(new_n20004_));
  OAI22_X1   g19747(.A1(new_n6721_), .A2(new_n6238_), .B1(new_n6723_), .B2(new_n6467_), .ZN(new_n20005_));
  NAND2_X1   g19748(.A1(new_n7617_), .A2(\b[53] ), .ZN(new_n20006_));
  AOI21_X1   g19749(.A1(new_n20006_), .A2(new_n20005_), .B(new_n6731_), .ZN(new_n20007_));
  NAND2_X1   g19750(.A1(new_n6471_), .A2(new_n20007_), .ZN(new_n20008_));
  XOR2_X1    g19751(.A1(new_n20008_), .A2(\a[56] ), .Z(new_n20009_));
  NOR2_X1    g19752(.A1(new_n20004_), .A2(new_n20009_), .ZN(new_n20010_));
  INV_X1     g19753(.I(new_n20009_), .ZN(new_n20011_));
  NOR2_X1    g19754(.A1(new_n20003_), .A2(new_n20011_), .ZN(new_n20012_));
  NOR2_X1    g19755(.A1(new_n20010_), .A2(new_n20012_), .ZN(new_n20013_));
  NOR2_X1    g19756(.A1(new_n20013_), .A2(new_n19968_), .ZN(new_n20014_));
  INV_X1     g19757(.I(new_n19968_), .ZN(new_n20015_));
  XOR2_X1    g19758(.A1(new_n20003_), .A2(new_n20009_), .Z(new_n20016_));
  NOR2_X1    g19759(.A1(new_n20016_), .A2(new_n20015_), .ZN(new_n20017_));
  NOR2_X1    g19760(.A1(new_n20014_), .A2(new_n20017_), .ZN(new_n20018_));
  XOR2_X1    g19761(.A1(new_n20018_), .A2(new_n19967_), .Z(new_n20019_));
  NOR2_X1    g19762(.A1(new_n20019_), .A2(new_n19966_), .ZN(new_n20020_));
  INV_X1     g19763(.I(new_n19966_), .ZN(new_n20021_));
  INV_X1     g19764(.I(new_n19967_), .ZN(new_n20022_));
  NOR2_X1    g19765(.A1(new_n20018_), .A2(new_n20022_), .ZN(new_n20023_));
  INV_X1     g19766(.I(new_n20023_), .ZN(new_n20024_));
  NAND2_X1   g19767(.A1(new_n20018_), .A2(new_n20022_), .ZN(new_n20025_));
  AOI21_X1   g19768(.A1(new_n20024_), .A2(new_n20025_), .B(new_n20021_), .ZN(new_n20026_));
  NOR2_X1    g19769(.A1(new_n20020_), .A2(new_n20026_), .ZN(new_n20027_));
  NOR2_X1    g19770(.A1(new_n20027_), .A2(new_n19961_), .ZN(new_n20028_));
  INV_X1     g19771(.I(new_n20028_), .ZN(new_n20029_));
  NAND2_X1   g19772(.A1(new_n20027_), .A2(new_n19961_), .ZN(new_n20030_));
  AOI21_X1   g19773(.A1(new_n20029_), .A2(new_n20030_), .B(new_n19960_), .ZN(new_n20031_));
  INV_X1     g19774(.I(new_n19960_), .ZN(new_n20032_));
  XNOR2_X1   g19775(.A1(new_n20027_), .A2(new_n19961_), .ZN(new_n20033_));
  NOR2_X1    g19776(.A1(new_n20033_), .A2(new_n20032_), .ZN(new_n20034_));
  NOR2_X1    g19777(.A1(new_n20034_), .A2(new_n20031_), .ZN(new_n20035_));
  NOR2_X1    g19778(.A1(new_n20035_), .A2(new_n19955_), .ZN(new_n20036_));
  NOR3_X1    g19779(.A1(new_n20034_), .A2(new_n19954_), .A3(new_n20031_), .ZN(new_n20037_));
  NOR2_X1    g19780(.A1(new_n20036_), .A2(new_n20037_), .ZN(new_n20038_));
  NOR2_X1    g19781(.A1(new_n20038_), .A2(new_n19953_), .ZN(new_n20039_));
  INV_X1     g19782(.I(new_n19953_), .ZN(new_n20040_));
  XOR2_X1    g19783(.A1(new_n20035_), .A2(new_n19954_), .Z(new_n20041_));
  NOR2_X1    g19784(.A1(new_n20041_), .A2(new_n20040_), .ZN(new_n20042_));
  NOR2_X1    g19785(.A1(new_n20042_), .A2(new_n20039_), .ZN(new_n20043_));
  OAI21_X1   g19786(.A1(new_n19845_), .A2(new_n19931_), .B(new_n19933_), .ZN(new_n20044_));
  INV_X1     g19787(.I(new_n19369_), .ZN(new_n20045_));
  INV_X1     g19788(.I(new_n19371_), .ZN(new_n20046_));
  OAI21_X1   g19789(.A1(new_n19362_), .A2(new_n20046_), .B(new_n20045_), .ZN(new_n20047_));
  NAND3_X1   g19790(.A1(new_n20047_), .A2(new_n19375_), .A3(new_n19724_), .ZN(new_n20048_));
  AOI21_X1   g19791(.A1(new_n20048_), .A2(new_n19734_), .B(new_n19731_), .ZN(new_n20049_));
  NOR2_X1    g19792(.A1(new_n19942_), .A2(new_n19836_), .ZN(new_n20050_));
  NOR3_X1    g19793(.A1(new_n20049_), .A2(new_n19737_), .A3(new_n20050_), .ZN(new_n20051_));
  NOR3_X1    g19794(.A1(new_n19935_), .A2(new_n19937_), .A3(new_n19939_), .ZN(new_n20052_));
  NOR2_X1    g19795(.A1(new_n20051_), .A2(new_n20052_), .ZN(new_n20053_));
  XOR2_X1    g19796(.A1(new_n20053_), .A2(new_n20044_), .Z(new_n20054_));
  XOR2_X1    g19797(.A1(new_n20054_), .A2(new_n20043_), .Z(\f[109] ));
  INV_X1     g19798(.I(new_n20050_), .ZN(new_n20056_));
  NAND3_X1   g19799(.A1(new_n19736_), .A2(new_n19943_), .A3(new_n20056_), .ZN(new_n20057_));
  NOR2_X1    g19800(.A1(new_n20043_), .A2(new_n20044_), .ZN(new_n20058_));
  XOR2_X1    g19801(.A1(new_n20043_), .A2(new_n20044_), .Z(new_n20059_));
  NOR2_X1    g19802(.A1(new_n20052_), .A2(new_n20059_), .ZN(new_n20060_));
  AOI21_X1   g19803(.A1(new_n20057_), .A2(new_n20060_), .B(new_n20058_), .ZN(new_n20061_));
  OAI21_X1   g19804(.A1(new_n19960_), .A2(new_n20028_), .B(new_n20030_), .ZN(new_n20062_));
  OAI22_X1   g19805(.A1(new_n5228_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n5225_), .ZN(new_n20063_));
  NAND2_X1   g19806(.A1(new_n5387_), .A2(\b[60] ), .ZN(new_n20064_));
  AOI21_X1   g19807(.A1(new_n20063_), .A2(new_n20064_), .B(new_n5231_), .ZN(new_n20065_));
  NAND2_X1   g19808(.A1(new_n8935_), .A2(new_n20065_), .ZN(new_n20066_));
  XOR2_X1    g19809(.A1(new_n20066_), .A2(\a[50] ), .Z(new_n20067_));
  INV_X1     g19810(.I(new_n20067_), .ZN(new_n20068_));
  OAI22_X1   g19811(.A1(new_n6721_), .A2(new_n6467_), .B1(new_n6723_), .B2(new_n6995_), .ZN(new_n20069_));
  NAND2_X1   g19812(.A1(new_n7617_), .A2(\b[54] ), .ZN(new_n20070_));
  AOI21_X1   g19813(.A1(new_n20070_), .A2(new_n20069_), .B(new_n6731_), .ZN(new_n20071_));
  NAND2_X1   g19814(.A1(new_n6994_), .A2(new_n20071_), .ZN(new_n20072_));
  XOR2_X1    g19815(.A1(new_n20072_), .A2(\a[56] ), .Z(new_n20073_));
  OAI21_X1   g19816(.A1(new_n19973_), .A2(new_n19999_), .B(new_n20001_), .ZN(new_n20074_));
  OAI22_X1   g19817(.A1(new_n6215_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n5955_), .ZN(new_n20075_));
  NAND2_X1   g19818(.A1(new_n8628_), .A2(\b[51] ), .ZN(new_n20076_));
  AOI21_X1   g19819(.A1(new_n20076_), .A2(new_n20075_), .B(new_n7354_), .ZN(new_n20077_));
  NAND2_X1   g19820(.A1(new_n6219_), .A2(new_n20077_), .ZN(new_n20078_));
  XOR2_X1    g19821(.A1(new_n20078_), .A2(\a[59] ), .Z(new_n20079_));
  OAI21_X1   g19822(.A1(new_n19980_), .A2(new_n19990_), .B(new_n19991_), .ZN(new_n20080_));
  NOR3_X1    g19823(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n4834_), .ZN(new_n20081_));
  NOR2_X1    g19824(.A1(new_n9364_), .A2(new_n4834_), .ZN(new_n20082_));
  NOR3_X1    g19825(.A1(new_n20082_), .A2(new_n4997_), .A3(new_n8985_), .ZN(new_n20083_));
  NOR2_X1    g19826(.A1(new_n20083_), .A2(new_n20081_), .ZN(new_n20084_));
  NOR2_X1    g19827(.A1(new_n19987_), .A2(new_n20084_), .ZN(new_n20085_));
  INV_X1     g19828(.I(new_n20085_), .ZN(new_n20086_));
  INV_X1     g19829(.I(new_n20084_), .ZN(new_n20087_));
  NOR2_X1    g19830(.A1(new_n20087_), .A2(new_n19986_), .ZN(new_n20088_));
  INV_X1     g19831(.I(new_n20088_), .ZN(new_n20089_));
  NAND2_X1   g19832(.A1(new_n20086_), .A2(new_n20089_), .ZN(new_n20090_));
  XOR2_X1    g19833(.A1(new_n19986_), .A2(new_n20084_), .Z(new_n20091_));
  NOR2_X1    g19834(.A1(new_n20080_), .A2(new_n20091_), .ZN(new_n20092_));
  AOI21_X1   g19835(.A1(new_n20080_), .A2(new_n20090_), .B(new_n20092_), .ZN(new_n20093_));
  OAI22_X1   g19836(.A1(new_n5538_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n5197_), .ZN(new_n20094_));
  NAND2_X1   g19837(.A1(new_n9644_), .A2(\b[48] ), .ZN(new_n20095_));
  AOI21_X1   g19838(.A1(new_n20095_), .A2(new_n20094_), .B(new_n8321_), .ZN(new_n20096_));
  NAND2_X1   g19839(.A1(new_n5537_), .A2(new_n20096_), .ZN(new_n20097_));
  XOR2_X1    g19840(.A1(new_n20097_), .A2(\a[62] ), .Z(new_n20098_));
  XNOR2_X1   g19841(.A1(new_n20093_), .A2(new_n20098_), .ZN(new_n20099_));
  NOR2_X1    g19842(.A1(new_n20099_), .A2(new_n20079_), .ZN(new_n20100_));
  INV_X1     g19843(.I(new_n20079_), .ZN(new_n20101_));
  NOR2_X1    g19844(.A1(new_n20093_), .A2(new_n20098_), .ZN(new_n20102_));
  INV_X1     g19845(.I(new_n20102_), .ZN(new_n20103_));
  NAND2_X1   g19846(.A1(new_n20093_), .A2(new_n20098_), .ZN(new_n20104_));
  AOI21_X1   g19847(.A1(new_n20103_), .A2(new_n20104_), .B(new_n20101_), .ZN(new_n20105_));
  NOR2_X1    g19848(.A1(new_n20100_), .A2(new_n20105_), .ZN(new_n20106_));
  XNOR2_X1   g19849(.A1(new_n20106_), .A2(new_n20074_), .ZN(new_n20107_));
  NOR2_X1    g19850(.A1(new_n20107_), .A2(new_n20073_), .ZN(new_n20108_));
  INV_X1     g19851(.I(new_n20073_), .ZN(new_n20109_));
  NOR2_X1    g19852(.A1(new_n20106_), .A2(new_n20074_), .ZN(new_n20110_));
  INV_X1     g19853(.I(new_n20110_), .ZN(new_n20111_));
  NAND2_X1   g19854(.A1(new_n20106_), .A2(new_n20074_), .ZN(new_n20112_));
  AOI21_X1   g19855(.A1(new_n20111_), .A2(new_n20112_), .B(new_n20109_), .ZN(new_n20113_));
  NOR2_X1    g19856(.A1(new_n20108_), .A2(new_n20113_), .ZN(new_n20114_));
  OAI22_X1   g19857(.A1(new_n5786_), .A2(new_n7890_), .B1(new_n7560_), .B2(new_n5792_), .ZN(new_n20115_));
  NAND2_X1   g19858(.A1(new_n6745_), .A2(\b[57] ), .ZN(new_n20116_));
  AOI21_X1   g19859(.A1(new_n20116_), .A2(new_n20115_), .B(new_n5796_), .ZN(new_n20117_));
  NAND2_X1   g19860(.A1(new_n7895_), .A2(new_n20117_), .ZN(new_n20118_));
  XOR2_X1    g19861(.A1(new_n20118_), .A2(\a[53] ), .Z(new_n20119_));
  NOR2_X1    g19862(.A1(new_n20012_), .A2(new_n19968_), .ZN(new_n20120_));
  NOR2_X1    g19863(.A1(new_n20120_), .A2(new_n20010_), .ZN(new_n20121_));
  XNOR2_X1   g19864(.A1(new_n20121_), .A2(new_n20119_), .ZN(new_n20122_));
  NOR2_X1    g19865(.A1(new_n20122_), .A2(new_n20114_), .ZN(new_n20123_));
  INV_X1     g19866(.I(new_n20114_), .ZN(new_n20124_));
  NOR2_X1    g19867(.A1(new_n20121_), .A2(new_n20119_), .ZN(new_n20125_));
  INV_X1     g19868(.I(new_n20125_), .ZN(new_n20126_));
  NAND2_X1   g19869(.A1(new_n20121_), .A2(new_n20119_), .ZN(new_n20127_));
  AOI21_X1   g19870(.A1(new_n20126_), .A2(new_n20127_), .B(new_n20124_), .ZN(new_n20128_));
  NOR2_X1    g19871(.A1(new_n20128_), .A2(new_n20123_), .ZN(new_n20129_));
  AOI21_X1   g19872(.A1(new_n20021_), .A2(new_n20025_), .B(new_n20023_), .ZN(new_n20130_));
  NOR2_X1    g19873(.A1(new_n20129_), .A2(new_n20130_), .ZN(new_n20131_));
  INV_X1     g19874(.I(new_n20130_), .ZN(new_n20132_));
  NOR3_X1    g19875(.A1(new_n20132_), .A2(new_n20123_), .A3(new_n20128_), .ZN(new_n20133_));
  OAI21_X1   g19876(.A1(new_n20131_), .A2(new_n20133_), .B(new_n20068_), .ZN(new_n20134_));
  XOR2_X1    g19877(.A1(new_n20129_), .A2(new_n20132_), .Z(new_n20135_));
  OAI21_X1   g19878(.A1(new_n20135_), .A2(new_n20068_), .B(new_n20134_), .ZN(new_n20136_));
  OAI22_X1   g19879(.A1(new_n9595_), .A2(new_n4714_), .B1(new_n8956_), .B2(new_n4873_), .ZN(new_n20137_));
  XOR2_X1    g19880(.A1(new_n20136_), .A2(new_n20137_), .Z(new_n20138_));
  XOR2_X1    g19881(.A1(new_n20138_), .A2(new_n4701_), .Z(new_n20139_));
  XOR2_X1    g19882(.A1(new_n20139_), .A2(new_n20062_), .Z(new_n20140_));
  NOR2_X1    g19883(.A1(new_n20037_), .A2(new_n19953_), .ZN(new_n20141_));
  NOR2_X1    g19884(.A1(new_n20141_), .A2(new_n20036_), .ZN(new_n20142_));
  INV_X1     g19885(.I(new_n20142_), .ZN(new_n20143_));
  XOR2_X1    g19886(.A1(new_n20140_), .A2(new_n20143_), .Z(new_n20144_));
  XOR2_X1    g19887(.A1(new_n20140_), .A2(new_n20143_), .Z(new_n20145_));
  NAND2_X1   g19888(.A1(new_n20061_), .A2(new_n20145_), .ZN(new_n20146_));
  OAI21_X1   g19889(.A1(new_n20061_), .A2(new_n20144_), .B(new_n20146_), .ZN(\f[110] ));
  OAI22_X1   g19890(.A1(new_n5228_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n5225_), .ZN(new_n20148_));
  NAND2_X1   g19891(.A1(new_n5387_), .A2(\b[61] ), .ZN(new_n20149_));
  AOI21_X1   g19892(.A1(new_n20148_), .A2(new_n20149_), .B(new_n5231_), .ZN(new_n20150_));
  NAND2_X1   g19893(.A1(new_n8963_), .A2(new_n20150_), .ZN(new_n20151_));
  XOR2_X1    g19894(.A1(new_n20151_), .A2(\a[50] ), .Z(new_n20152_));
  INV_X1     g19895(.I(new_n20131_), .ZN(new_n20153_));
  OAI21_X1   g19896(.A1(new_n20067_), .A2(new_n20133_), .B(new_n20153_), .ZN(new_n20154_));
  AOI21_X1   g19897(.A1(new_n20114_), .A2(new_n20127_), .B(new_n20125_), .ZN(new_n20155_));
  INV_X1     g19898(.I(new_n20155_), .ZN(new_n20156_));
  OAI22_X1   g19899(.A1(new_n5786_), .A2(new_n7930_), .B1(new_n7890_), .B2(new_n5792_), .ZN(new_n20157_));
  NAND2_X1   g19900(.A1(new_n6745_), .A2(\b[58] ), .ZN(new_n20158_));
  AOI21_X1   g19901(.A1(new_n20158_), .A2(new_n20157_), .B(new_n5796_), .ZN(new_n20159_));
  NAND2_X1   g19902(.A1(new_n7929_), .A2(new_n20159_), .ZN(new_n20160_));
  XOR2_X1    g19903(.A1(new_n20160_), .A2(\a[53] ), .Z(new_n20161_));
  OAI21_X1   g19904(.A1(new_n20073_), .A2(new_n20110_), .B(new_n20112_), .ZN(new_n20162_));
  INV_X1     g19905(.I(new_n20162_), .ZN(new_n20163_));
  OAI22_X1   g19906(.A1(new_n6721_), .A2(new_n6995_), .B1(new_n6723_), .B2(new_n7305_), .ZN(new_n20164_));
  NAND2_X1   g19907(.A1(new_n7617_), .A2(\b[55] ), .ZN(new_n20165_));
  AOI21_X1   g19908(.A1(new_n20165_), .A2(new_n20164_), .B(new_n6731_), .ZN(new_n20166_));
  NAND2_X1   g19909(.A1(new_n7308_), .A2(new_n20166_), .ZN(new_n20167_));
  XOR2_X1    g19910(.A1(new_n20167_), .A2(\a[56] ), .Z(new_n20168_));
  INV_X1     g19911(.I(new_n20168_), .ZN(new_n20169_));
  AOI21_X1   g19912(.A1(new_n20101_), .A2(new_n20104_), .B(new_n20102_), .ZN(new_n20170_));
  INV_X1     g19913(.I(new_n20170_), .ZN(new_n20171_));
  AOI21_X1   g19914(.A1(new_n20080_), .A2(new_n20086_), .B(new_n20088_), .ZN(new_n20172_));
  OAI22_X1   g19915(.A1(new_n5738_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n5538_), .ZN(new_n20173_));
  NAND2_X1   g19916(.A1(new_n9644_), .A2(\b[49] ), .ZN(new_n20174_));
  AOI21_X1   g19917(.A1(new_n20174_), .A2(new_n20173_), .B(new_n8321_), .ZN(new_n20175_));
  NAND2_X1   g19918(.A1(new_n5741_), .A2(new_n20175_), .ZN(new_n20176_));
  XOR2_X1    g19919(.A1(new_n20176_), .A2(\a[62] ), .Z(new_n20177_));
  INV_X1     g19920(.I(new_n20177_), .ZN(new_n20178_));
  NOR2_X1    g19921(.A1(new_n8985_), .A2(new_n5178_), .ZN(new_n20179_));
  NOR2_X1    g19922(.A1(new_n9364_), .A2(new_n4997_), .ZN(new_n20180_));
  XNOR2_X1   g19923(.A1(new_n20179_), .A2(new_n20180_), .ZN(new_n20181_));
  XOR2_X1    g19924(.A1(new_n20181_), .A2(\a[47] ), .Z(new_n20182_));
  NOR2_X1    g19925(.A1(new_n20182_), .A2(new_n20084_), .ZN(new_n20183_));
  NOR2_X1    g19926(.A1(new_n20181_), .A2(new_n4701_), .ZN(new_n20184_));
  INV_X1     g19927(.I(new_n20184_), .ZN(new_n20185_));
  NAND2_X1   g19928(.A1(new_n20181_), .A2(new_n4701_), .ZN(new_n20186_));
  AOI21_X1   g19929(.A1(new_n20185_), .A2(new_n20186_), .B(new_n20087_), .ZN(new_n20187_));
  NOR2_X1    g19930(.A1(new_n20183_), .A2(new_n20187_), .ZN(new_n20188_));
  NOR2_X1    g19931(.A1(new_n20178_), .A2(new_n20188_), .ZN(new_n20189_));
  INV_X1     g19932(.I(new_n20189_), .ZN(new_n20190_));
  NAND2_X1   g19933(.A1(new_n20178_), .A2(new_n20188_), .ZN(new_n20191_));
  AOI21_X1   g19934(.A1(new_n20190_), .A2(new_n20191_), .B(new_n20172_), .ZN(new_n20192_));
  XNOR2_X1   g19935(.A1(new_n20177_), .A2(new_n20188_), .ZN(new_n20193_));
  AOI21_X1   g19936(.A1(new_n20172_), .A2(new_n20193_), .B(new_n20192_), .ZN(new_n20194_));
  OAI22_X1   g19937(.A1(new_n6238_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n6215_), .ZN(new_n20195_));
  NAND2_X1   g19938(.A1(new_n8628_), .A2(\b[52] ), .ZN(new_n20196_));
  AOI21_X1   g19939(.A1(new_n20196_), .A2(new_n20195_), .B(new_n7354_), .ZN(new_n20197_));
  NAND2_X1   g19940(.A1(new_n6237_), .A2(new_n20197_), .ZN(new_n20198_));
  XOR2_X1    g19941(.A1(new_n20198_), .A2(\a[59] ), .Z(new_n20199_));
  XOR2_X1    g19942(.A1(new_n20194_), .A2(new_n20199_), .Z(new_n20200_));
  NAND2_X1   g19943(.A1(new_n20200_), .A2(new_n20171_), .ZN(new_n20201_));
  NOR2_X1    g19944(.A1(new_n20194_), .A2(new_n20199_), .ZN(new_n20202_));
  NAND2_X1   g19945(.A1(new_n20194_), .A2(new_n20199_), .ZN(new_n20203_));
  INV_X1     g19946(.I(new_n20203_), .ZN(new_n20204_));
  OAI21_X1   g19947(.A1(new_n20204_), .A2(new_n20202_), .B(new_n20170_), .ZN(new_n20205_));
  NAND2_X1   g19948(.A1(new_n20201_), .A2(new_n20205_), .ZN(new_n20206_));
  XOR2_X1    g19949(.A1(new_n20206_), .A2(new_n20169_), .Z(new_n20207_));
  NOR2_X1    g19950(.A1(new_n20207_), .A2(new_n20163_), .ZN(new_n20208_));
  AOI21_X1   g19951(.A1(new_n20201_), .A2(new_n20205_), .B(new_n20169_), .ZN(new_n20209_));
  NOR2_X1    g19952(.A1(new_n20206_), .A2(new_n20168_), .ZN(new_n20210_));
  NOR2_X1    g19953(.A1(new_n20210_), .A2(new_n20209_), .ZN(new_n20211_));
  NOR2_X1    g19954(.A1(new_n20211_), .A2(new_n20162_), .ZN(new_n20212_));
  NOR2_X1    g19955(.A1(new_n20208_), .A2(new_n20212_), .ZN(new_n20213_));
  XNOR2_X1   g19956(.A1(new_n20213_), .A2(new_n20161_), .ZN(new_n20214_));
  INV_X1     g19957(.I(new_n20213_), .ZN(new_n20215_));
  NAND2_X1   g19958(.A1(new_n20215_), .A2(new_n20161_), .ZN(new_n20216_));
  NOR2_X1    g19959(.A1(new_n20215_), .A2(new_n20161_), .ZN(new_n20217_));
  INV_X1     g19960(.I(new_n20217_), .ZN(new_n20218_));
  AOI21_X1   g19961(.A1(new_n20218_), .A2(new_n20216_), .B(new_n20156_), .ZN(new_n20219_));
  AOI21_X1   g19962(.A1(new_n20156_), .A2(new_n20214_), .B(new_n20219_), .ZN(new_n20220_));
  XNOR2_X1   g19963(.A1(new_n20220_), .A2(new_n20154_), .ZN(new_n20221_));
  NOR2_X1    g19964(.A1(new_n20221_), .A2(new_n20152_), .ZN(new_n20222_));
  INV_X1     g19965(.I(new_n20152_), .ZN(new_n20223_));
  NOR2_X1    g19966(.A1(new_n20220_), .A2(new_n20154_), .ZN(new_n20224_));
  INV_X1     g19967(.I(new_n20224_), .ZN(new_n20225_));
  NAND2_X1   g19968(.A1(new_n20220_), .A2(new_n20154_), .ZN(new_n20226_));
  AOI21_X1   g19969(.A1(new_n20225_), .A2(new_n20226_), .B(new_n20223_), .ZN(new_n20227_));
  NOR2_X1    g19970(.A1(new_n20222_), .A2(new_n20227_), .ZN(new_n20228_));
  XOR2_X1    g19971(.A1(new_n20137_), .A2(new_n4701_), .Z(new_n20229_));
  NOR3_X1    g19972(.A1(new_n20136_), .A2(new_n20062_), .A3(new_n20229_), .ZN(new_n20230_));
  AOI21_X1   g19973(.A1(new_n20062_), .A2(new_n20136_), .B(new_n20230_), .ZN(new_n20231_));
  XOR2_X1    g19974(.A1(new_n20228_), .A2(new_n20231_), .Z(new_n20232_));
  NOR2_X1    g19975(.A1(new_n20061_), .A2(new_n20140_), .ZN(new_n20233_));
  XOR2_X1    g19976(.A1(new_n20233_), .A2(new_n20232_), .Z(new_n20234_));
  XOR2_X1    g19977(.A1(new_n20061_), .A2(new_n20140_), .Z(new_n20235_));
  NAND2_X1   g19978(.A1(new_n20235_), .A2(new_n20143_), .ZN(new_n20236_));
  XOR2_X1    g19979(.A1(new_n20234_), .A2(new_n20236_), .Z(\f[111] ));
  NOR2_X1    g19980(.A1(new_n5378_), .A2(new_n8932_), .ZN(new_n20238_));
  NOR2_X1    g19981(.A1(new_n5225_), .A2(new_n8956_), .ZN(new_n20239_));
  NOR4_X1    g19982(.A1(new_n9323_), .A2(new_n5231_), .A3(new_n20238_), .A4(new_n20239_), .ZN(new_n20240_));
  XOR2_X1    g19983(.A1(new_n20240_), .A2(new_n5220_), .Z(new_n20241_));
  AOI21_X1   g19984(.A1(new_n20156_), .A2(new_n20216_), .B(new_n20217_), .ZN(new_n20242_));
  INV_X1     g19985(.I(new_n20242_), .ZN(new_n20243_));
  OAI22_X1   g19986(.A1(new_n5786_), .A2(new_n8548_), .B1(new_n7930_), .B2(new_n5792_), .ZN(new_n20244_));
  NAND2_X1   g19987(.A1(new_n6745_), .A2(\b[59] ), .ZN(new_n20245_));
  AOI21_X1   g19988(.A1(new_n20245_), .A2(new_n20244_), .B(new_n5796_), .ZN(new_n20246_));
  NAND2_X1   g19989(.A1(new_n8550_), .A2(new_n20246_), .ZN(new_n20247_));
  XOR2_X1    g19990(.A1(new_n20247_), .A2(\a[53] ), .Z(new_n20248_));
  INV_X1     g19991(.I(new_n20209_), .ZN(new_n20249_));
  AOI21_X1   g19992(.A1(new_n20249_), .A2(new_n20162_), .B(new_n20210_), .ZN(new_n20250_));
  OAI22_X1   g19993(.A1(new_n6721_), .A2(new_n7305_), .B1(new_n6723_), .B2(new_n7560_), .ZN(new_n20251_));
  NAND2_X1   g19994(.A1(new_n7617_), .A2(\b[56] ), .ZN(new_n20252_));
  AOI21_X1   g19995(.A1(new_n20252_), .A2(new_n20251_), .B(new_n6731_), .ZN(new_n20253_));
  NAND2_X1   g19996(.A1(new_n7559_), .A2(new_n20253_), .ZN(new_n20254_));
  XOR2_X1    g19997(.A1(new_n20254_), .A2(\a[56] ), .Z(new_n20255_));
  NOR2_X1    g19998(.A1(new_n20204_), .A2(new_n20170_), .ZN(new_n20256_));
  NOR2_X1    g19999(.A1(new_n20256_), .A2(new_n20202_), .ZN(new_n20257_));
  OAI22_X1   g20000(.A1(new_n6467_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n6238_), .ZN(new_n20258_));
  NAND2_X1   g20001(.A1(new_n8628_), .A2(\b[53] ), .ZN(new_n20259_));
  AOI21_X1   g20002(.A1(new_n20259_), .A2(new_n20258_), .B(new_n7354_), .ZN(new_n20260_));
  NAND2_X1   g20003(.A1(new_n6471_), .A2(new_n20260_), .ZN(new_n20261_));
  XOR2_X1    g20004(.A1(new_n20261_), .A2(\a[59] ), .Z(new_n20262_));
  OAI21_X1   g20005(.A1(new_n20172_), .A2(new_n20189_), .B(new_n20191_), .ZN(new_n20263_));
  OAI22_X1   g20006(.A1(new_n5955_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n5738_), .ZN(new_n20264_));
  NAND2_X1   g20007(.A1(new_n9644_), .A2(\b[50] ), .ZN(new_n20265_));
  AOI21_X1   g20008(.A1(new_n20265_), .A2(new_n20264_), .B(new_n8321_), .ZN(new_n20266_));
  NAND2_X1   g20009(.A1(new_n5954_), .A2(new_n20266_), .ZN(new_n20267_));
  XOR2_X1    g20010(.A1(new_n20267_), .A2(new_n8309_), .Z(new_n20268_));
  NAND2_X1   g20011(.A1(new_n20186_), .A2(new_n20087_), .ZN(new_n20269_));
  NAND2_X1   g20012(.A1(new_n20269_), .A2(new_n20185_), .ZN(new_n20270_));
  NOR3_X1    g20013(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n5178_), .ZN(new_n20271_));
  NOR2_X1    g20014(.A1(new_n9364_), .A2(new_n5178_), .ZN(new_n20272_));
  NOR3_X1    g20015(.A1(new_n20272_), .A2(new_n5197_), .A3(new_n8985_), .ZN(new_n20273_));
  NOR2_X1    g20016(.A1(new_n20273_), .A2(new_n20271_), .ZN(new_n20274_));
  INV_X1     g20017(.I(new_n20274_), .ZN(new_n20275_));
  XOR2_X1    g20018(.A1(new_n20270_), .A2(new_n20275_), .Z(new_n20276_));
  INV_X1     g20019(.I(new_n20276_), .ZN(new_n20277_));
  NOR2_X1    g20020(.A1(new_n20270_), .A2(new_n20274_), .ZN(new_n20278_));
  INV_X1     g20021(.I(new_n20278_), .ZN(new_n20279_));
  NAND2_X1   g20022(.A1(new_n20270_), .A2(new_n20274_), .ZN(new_n20280_));
  AOI21_X1   g20023(.A1(new_n20279_), .A2(new_n20280_), .B(new_n20268_), .ZN(new_n20281_));
  AOI21_X1   g20024(.A1(new_n20268_), .A2(new_n20277_), .B(new_n20281_), .ZN(new_n20282_));
  XNOR2_X1   g20025(.A1(new_n20263_), .A2(new_n20282_), .ZN(new_n20283_));
  NOR2_X1    g20026(.A1(new_n20283_), .A2(new_n20262_), .ZN(new_n20284_));
  NOR2_X1    g20027(.A1(new_n20263_), .A2(new_n20282_), .ZN(new_n20285_));
  INV_X1     g20028(.I(new_n20285_), .ZN(new_n20286_));
  NAND2_X1   g20029(.A1(new_n20263_), .A2(new_n20282_), .ZN(new_n20287_));
  NAND2_X1   g20030(.A1(new_n20286_), .A2(new_n20287_), .ZN(new_n20288_));
  AOI21_X1   g20031(.A1(new_n20262_), .A2(new_n20288_), .B(new_n20284_), .ZN(new_n20289_));
  XOR2_X1    g20032(.A1(new_n20257_), .A2(new_n20289_), .Z(new_n20290_));
  NOR2_X1    g20033(.A1(new_n20290_), .A2(new_n20255_), .ZN(new_n20291_));
  INV_X1     g20034(.I(new_n20257_), .ZN(new_n20292_));
  NOR2_X1    g20035(.A1(new_n20292_), .A2(new_n20289_), .ZN(new_n20293_));
  INV_X1     g20036(.I(new_n20293_), .ZN(new_n20294_));
  NAND2_X1   g20037(.A1(new_n20292_), .A2(new_n20289_), .ZN(new_n20295_));
  NAND2_X1   g20038(.A1(new_n20294_), .A2(new_n20295_), .ZN(new_n20296_));
  AOI21_X1   g20039(.A1(new_n20255_), .A2(new_n20296_), .B(new_n20291_), .ZN(new_n20297_));
  XOR2_X1    g20040(.A1(new_n20297_), .A2(new_n20250_), .Z(new_n20298_));
  NOR2_X1    g20041(.A1(new_n20298_), .A2(new_n20248_), .ZN(new_n20299_));
  INV_X1     g20042(.I(new_n20250_), .ZN(new_n20300_));
  NOR2_X1    g20043(.A1(new_n20297_), .A2(new_n20300_), .ZN(new_n20301_));
  INV_X1     g20044(.I(new_n20301_), .ZN(new_n20302_));
  NAND2_X1   g20045(.A1(new_n20297_), .A2(new_n20300_), .ZN(new_n20303_));
  NAND2_X1   g20046(.A1(new_n20302_), .A2(new_n20303_), .ZN(new_n20304_));
  AOI21_X1   g20047(.A1(new_n20248_), .A2(new_n20304_), .B(new_n20299_), .ZN(new_n20305_));
  NOR2_X1    g20048(.A1(new_n20305_), .A2(new_n20243_), .ZN(new_n20306_));
  INV_X1     g20049(.I(new_n20306_), .ZN(new_n20307_));
  NAND2_X1   g20050(.A1(new_n20305_), .A2(new_n20243_), .ZN(new_n20308_));
  AOI21_X1   g20051(.A1(new_n20307_), .A2(new_n20308_), .B(new_n20241_), .ZN(new_n20309_));
  XOR2_X1    g20052(.A1(new_n20305_), .A2(new_n20242_), .Z(new_n20310_));
  INV_X1     g20053(.I(new_n20310_), .ZN(new_n20311_));
  AOI21_X1   g20054(.A1(new_n20311_), .A2(new_n20241_), .B(new_n20309_), .ZN(new_n20312_));
  OAI21_X1   g20055(.A1(new_n20152_), .A2(new_n20224_), .B(new_n20226_), .ZN(new_n20313_));
  NAND2_X1   g20056(.A1(new_n20232_), .A2(new_n20143_), .ZN(new_n20314_));
  INV_X1     g20057(.I(new_n20314_), .ZN(new_n20315_));
  NOR3_X1    g20058(.A1(new_n20061_), .A2(new_n20140_), .A3(new_n20315_), .ZN(new_n20316_));
  OAI21_X1   g20059(.A1(new_n20222_), .A2(new_n20227_), .B(new_n20231_), .ZN(new_n20317_));
  INV_X1     g20060(.I(new_n20317_), .ZN(new_n20318_));
  NOR2_X1    g20061(.A1(new_n20316_), .A2(new_n20318_), .ZN(new_n20319_));
  XOR2_X1    g20062(.A1(new_n20319_), .A2(new_n20313_), .Z(new_n20320_));
  XOR2_X1    g20063(.A1(new_n20320_), .A2(new_n20312_), .Z(\f[112] ));
  NOR2_X1    g20064(.A1(new_n20312_), .A2(new_n20313_), .ZN(new_n20322_));
  INV_X1     g20065(.I(new_n20322_), .ZN(new_n20323_));
  XOR2_X1    g20066(.A1(new_n20312_), .A2(new_n20313_), .Z(new_n20324_));
  NOR2_X1    g20067(.A1(new_n20324_), .A2(new_n20318_), .ZN(new_n20325_));
  INV_X1     g20068(.I(new_n20325_), .ZN(new_n20326_));
  OAI21_X1   g20069(.A1(new_n20316_), .A2(new_n20326_), .B(new_n20323_), .ZN(new_n20327_));
  OAI21_X1   g20070(.A1(new_n20248_), .A2(new_n20301_), .B(new_n20303_), .ZN(new_n20328_));
  OAI22_X1   g20071(.A1(new_n5786_), .A2(new_n8932_), .B1(new_n8548_), .B2(new_n5792_), .ZN(new_n20329_));
  NAND2_X1   g20072(.A1(new_n6745_), .A2(\b[60] ), .ZN(new_n20330_));
  AOI21_X1   g20073(.A1(new_n20330_), .A2(new_n20329_), .B(new_n5796_), .ZN(new_n20331_));
  NAND2_X1   g20074(.A1(new_n8935_), .A2(new_n20331_), .ZN(new_n20332_));
  XOR2_X1    g20075(.A1(new_n20332_), .A2(\a[53] ), .Z(new_n20333_));
  OAI22_X1   g20076(.A1(new_n6995_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n6467_), .ZN(new_n20334_));
  NAND2_X1   g20077(.A1(new_n8628_), .A2(\b[54] ), .ZN(new_n20335_));
  AOI21_X1   g20078(.A1(new_n20335_), .A2(new_n20334_), .B(new_n7354_), .ZN(new_n20336_));
  NAND2_X1   g20079(.A1(new_n6994_), .A2(new_n20336_), .ZN(new_n20337_));
  XOR2_X1    g20080(.A1(new_n20337_), .A2(\a[59] ), .Z(new_n20338_));
  OAI22_X1   g20081(.A1(new_n6215_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n5955_), .ZN(new_n20339_));
  NAND2_X1   g20082(.A1(new_n9644_), .A2(\b[51] ), .ZN(new_n20340_));
  AOI21_X1   g20083(.A1(new_n20340_), .A2(new_n20339_), .B(new_n8321_), .ZN(new_n20341_));
  NAND2_X1   g20084(.A1(new_n6219_), .A2(new_n20341_), .ZN(new_n20342_));
  XOR2_X1    g20085(.A1(new_n20342_), .A2(\a[62] ), .Z(new_n20343_));
  NOR3_X1    g20086(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n5197_), .ZN(new_n20344_));
  NOR2_X1    g20087(.A1(new_n9364_), .A2(new_n5197_), .ZN(new_n20345_));
  NOR3_X1    g20088(.A1(new_n20345_), .A2(new_n5538_), .A3(new_n8985_), .ZN(new_n20346_));
  NOR2_X1    g20089(.A1(new_n20346_), .A2(new_n20344_), .ZN(new_n20347_));
  NOR2_X1    g20090(.A1(new_n20275_), .A2(new_n20347_), .ZN(new_n20348_));
  NOR3_X1    g20091(.A1(new_n20274_), .A2(new_n20344_), .A3(new_n20346_), .ZN(new_n20349_));
  NOR2_X1    g20092(.A1(new_n20348_), .A2(new_n20349_), .ZN(new_n20350_));
  NOR2_X1    g20093(.A1(new_n20343_), .A2(new_n20350_), .ZN(new_n20351_));
  INV_X1     g20094(.I(new_n20343_), .ZN(new_n20352_));
  XOR2_X1    g20095(.A1(new_n20274_), .A2(new_n20347_), .Z(new_n20353_));
  NOR2_X1    g20096(.A1(new_n20352_), .A2(new_n20353_), .ZN(new_n20354_));
  NOR2_X1    g20097(.A1(new_n20354_), .A2(new_n20351_), .ZN(new_n20355_));
  INV_X1     g20098(.I(new_n20280_), .ZN(new_n20356_));
  AOI21_X1   g20099(.A1(new_n20268_), .A2(new_n20279_), .B(new_n20356_), .ZN(new_n20357_));
  XNOR2_X1   g20100(.A1(new_n20355_), .A2(new_n20357_), .ZN(new_n20358_));
  NOR2_X1    g20101(.A1(new_n20358_), .A2(new_n20338_), .ZN(new_n20359_));
  INV_X1     g20102(.I(new_n20338_), .ZN(new_n20360_));
  NOR2_X1    g20103(.A1(new_n20355_), .A2(new_n20357_), .ZN(new_n20361_));
  INV_X1     g20104(.I(new_n20361_), .ZN(new_n20362_));
  NAND2_X1   g20105(.A1(new_n20355_), .A2(new_n20357_), .ZN(new_n20363_));
  AOI21_X1   g20106(.A1(new_n20362_), .A2(new_n20363_), .B(new_n20360_), .ZN(new_n20364_));
  NOR2_X1    g20107(.A1(new_n20359_), .A2(new_n20364_), .ZN(new_n20365_));
  OAI22_X1   g20108(.A1(new_n6721_), .A2(new_n7560_), .B1(new_n6723_), .B2(new_n7890_), .ZN(new_n20366_));
  NAND2_X1   g20109(.A1(new_n7617_), .A2(\b[57] ), .ZN(new_n20367_));
  AOI21_X1   g20110(.A1(new_n20367_), .A2(new_n20366_), .B(new_n6731_), .ZN(new_n20368_));
  NAND2_X1   g20111(.A1(new_n7895_), .A2(new_n20368_), .ZN(new_n20369_));
  XOR2_X1    g20112(.A1(new_n20369_), .A2(\a[56] ), .Z(new_n20370_));
  OAI21_X1   g20113(.A1(new_n20262_), .A2(new_n20285_), .B(new_n20287_), .ZN(new_n20371_));
  XOR2_X1    g20114(.A1(new_n20371_), .A2(new_n20370_), .Z(new_n20372_));
  NOR2_X1    g20115(.A1(new_n20365_), .A2(new_n20372_), .ZN(new_n20373_));
  INV_X1     g20116(.I(new_n20365_), .ZN(new_n20374_));
  INV_X1     g20117(.I(new_n20371_), .ZN(new_n20375_));
  NOR2_X1    g20118(.A1(new_n20375_), .A2(new_n20370_), .ZN(new_n20376_));
  INV_X1     g20119(.I(new_n20376_), .ZN(new_n20377_));
  NAND2_X1   g20120(.A1(new_n20375_), .A2(new_n20370_), .ZN(new_n20378_));
  AOI21_X1   g20121(.A1(new_n20377_), .A2(new_n20378_), .B(new_n20374_), .ZN(new_n20379_));
  NOR2_X1    g20122(.A1(new_n20379_), .A2(new_n20373_), .ZN(new_n20380_));
  OAI21_X1   g20123(.A1(new_n20255_), .A2(new_n20293_), .B(new_n20295_), .ZN(new_n20381_));
  INV_X1     g20124(.I(new_n20381_), .ZN(new_n20382_));
  NOR2_X1    g20125(.A1(new_n20382_), .A2(new_n20380_), .ZN(new_n20383_));
  NOR3_X1    g20126(.A1(new_n20381_), .A2(new_n20373_), .A3(new_n20379_), .ZN(new_n20384_));
  NOR2_X1    g20127(.A1(new_n20383_), .A2(new_n20384_), .ZN(new_n20385_));
  NOR2_X1    g20128(.A1(new_n20385_), .A2(new_n20333_), .ZN(new_n20386_));
  INV_X1     g20129(.I(new_n20333_), .ZN(new_n20387_));
  XOR2_X1    g20130(.A1(new_n20381_), .A2(new_n20380_), .Z(new_n20388_));
  NOR2_X1    g20131(.A1(new_n20388_), .A2(new_n20387_), .ZN(new_n20389_));
  NOR2_X1    g20132(.A1(new_n20386_), .A2(new_n20389_), .ZN(new_n20390_));
  OAI22_X1   g20133(.A1(new_n9595_), .A2(new_n5231_), .B1(new_n8956_), .B2(new_n5378_), .ZN(new_n20391_));
  XOR2_X1    g20134(.A1(new_n20390_), .A2(new_n20391_), .Z(new_n20392_));
  XOR2_X1    g20135(.A1(new_n20392_), .A2(\a[50] ), .Z(new_n20393_));
  XOR2_X1    g20136(.A1(new_n20393_), .A2(new_n20328_), .Z(new_n20394_));
  OAI21_X1   g20137(.A1(new_n20241_), .A2(new_n20306_), .B(new_n20308_), .ZN(new_n20395_));
  INV_X1     g20138(.I(new_n20395_), .ZN(new_n20396_));
  XOR2_X1    g20139(.A1(new_n20394_), .A2(new_n20396_), .Z(new_n20397_));
  NAND2_X1   g20140(.A1(new_n20327_), .A2(new_n20397_), .ZN(new_n20398_));
  XOR2_X1    g20141(.A1(new_n20394_), .A2(new_n20396_), .Z(new_n20399_));
  OAI21_X1   g20142(.A1(new_n20327_), .A2(new_n20399_), .B(new_n20398_), .ZN(\f[113] ));
  OAI22_X1   g20143(.A1(new_n5786_), .A2(new_n8956_), .B1(new_n8932_), .B2(new_n5792_), .ZN(new_n20401_));
  NAND2_X1   g20144(.A1(new_n6745_), .A2(\b[61] ), .ZN(new_n20402_));
  AOI21_X1   g20145(.A1(new_n20402_), .A2(new_n20401_), .B(new_n5796_), .ZN(new_n20403_));
  NAND2_X1   g20146(.A1(new_n8963_), .A2(new_n20403_), .ZN(new_n20404_));
  XOR2_X1    g20147(.A1(new_n20404_), .A2(\a[53] ), .Z(new_n20405_));
  INV_X1     g20148(.I(new_n20384_), .ZN(new_n20406_));
  AOI21_X1   g20149(.A1(new_n20406_), .A2(new_n20387_), .B(new_n20383_), .ZN(new_n20407_));
  AOI21_X1   g20150(.A1(new_n20365_), .A2(new_n20378_), .B(new_n20376_), .ZN(new_n20408_));
  OAI22_X1   g20151(.A1(new_n6721_), .A2(new_n7890_), .B1(new_n6723_), .B2(new_n7930_), .ZN(new_n20409_));
  NAND2_X1   g20152(.A1(new_n7617_), .A2(\b[58] ), .ZN(new_n20410_));
  AOI21_X1   g20153(.A1(new_n20410_), .A2(new_n20409_), .B(new_n6731_), .ZN(new_n20411_));
  NAND2_X1   g20154(.A1(new_n7929_), .A2(new_n20411_), .ZN(new_n20412_));
  XOR2_X1    g20155(.A1(new_n20412_), .A2(\a[56] ), .Z(new_n20413_));
  INV_X1     g20156(.I(new_n20413_), .ZN(new_n20414_));
  AOI21_X1   g20157(.A1(new_n20360_), .A2(new_n20363_), .B(new_n20361_), .ZN(new_n20415_));
  INV_X1     g20158(.I(new_n20415_), .ZN(new_n20416_));
  OAI22_X1   g20159(.A1(new_n7305_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n6995_), .ZN(new_n20417_));
  NAND2_X1   g20160(.A1(new_n8628_), .A2(\b[55] ), .ZN(new_n20418_));
  AOI21_X1   g20161(.A1(new_n20418_), .A2(new_n20417_), .B(new_n7354_), .ZN(new_n20419_));
  NAND2_X1   g20162(.A1(new_n7308_), .A2(new_n20419_), .ZN(new_n20420_));
  XOR2_X1    g20163(.A1(new_n20420_), .A2(\a[59] ), .Z(new_n20421_));
  OAI22_X1   g20164(.A1(new_n6238_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n6215_), .ZN(new_n20422_));
  NAND2_X1   g20165(.A1(new_n9644_), .A2(\b[52] ), .ZN(new_n20423_));
  AOI21_X1   g20166(.A1(new_n20423_), .A2(new_n20422_), .B(new_n8321_), .ZN(new_n20424_));
  NAND2_X1   g20167(.A1(new_n6237_), .A2(new_n20424_), .ZN(new_n20425_));
  XOR2_X1    g20168(.A1(new_n20425_), .A2(\a[62] ), .Z(new_n20426_));
  INV_X1     g20169(.I(new_n20426_), .ZN(new_n20427_));
  INV_X1     g20170(.I(new_n20349_), .ZN(new_n20428_));
  AOI21_X1   g20171(.A1(new_n20352_), .A2(new_n20428_), .B(new_n20348_), .ZN(new_n20429_));
  NOR2_X1    g20172(.A1(new_n8985_), .A2(new_n5738_), .ZN(new_n20430_));
  NOR2_X1    g20173(.A1(new_n9364_), .A2(new_n5538_), .ZN(new_n20431_));
  XNOR2_X1   g20174(.A1(new_n20430_), .A2(new_n20431_), .ZN(new_n20432_));
  XOR2_X1    g20175(.A1(new_n20432_), .A2(\a[50] ), .Z(new_n20433_));
  NOR2_X1    g20176(.A1(new_n20433_), .A2(new_n20274_), .ZN(new_n20434_));
  NOR2_X1    g20177(.A1(new_n20432_), .A2(new_n5220_), .ZN(new_n20435_));
  INV_X1     g20178(.I(new_n20435_), .ZN(new_n20436_));
  NAND2_X1   g20179(.A1(new_n20432_), .A2(new_n5220_), .ZN(new_n20437_));
  AOI21_X1   g20180(.A1(new_n20436_), .A2(new_n20437_), .B(new_n20275_), .ZN(new_n20438_));
  NOR2_X1    g20181(.A1(new_n20434_), .A2(new_n20438_), .ZN(new_n20439_));
  INV_X1     g20182(.I(new_n20439_), .ZN(new_n20440_));
  XOR2_X1    g20183(.A1(new_n20429_), .A2(new_n20440_), .Z(new_n20441_));
  NAND2_X1   g20184(.A1(new_n20441_), .A2(new_n20427_), .ZN(new_n20442_));
  AND2_X2    g20185(.A1(new_n20429_), .A2(new_n20440_), .Z(new_n20443_));
  NOR2_X1    g20186(.A1(new_n20429_), .A2(new_n20440_), .ZN(new_n20444_));
  OAI21_X1   g20187(.A1(new_n20443_), .A2(new_n20444_), .B(new_n20426_), .ZN(new_n20445_));
  NAND2_X1   g20188(.A1(new_n20442_), .A2(new_n20445_), .ZN(new_n20446_));
  XOR2_X1    g20189(.A1(new_n20446_), .A2(new_n20421_), .Z(new_n20447_));
  NAND2_X1   g20190(.A1(new_n20447_), .A2(new_n20416_), .ZN(new_n20448_));
  AND2_X2    g20191(.A1(new_n20446_), .A2(new_n20421_), .Z(new_n20449_));
  NOR2_X1    g20192(.A1(new_n20446_), .A2(new_n20421_), .ZN(new_n20450_));
  OAI21_X1   g20193(.A1(new_n20449_), .A2(new_n20450_), .B(new_n20415_), .ZN(new_n20451_));
  NAND2_X1   g20194(.A1(new_n20448_), .A2(new_n20451_), .ZN(new_n20452_));
  XOR2_X1    g20195(.A1(new_n20452_), .A2(new_n20414_), .Z(new_n20453_));
  NOR2_X1    g20196(.A1(new_n20453_), .A2(new_n20408_), .ZN(new_n20454_));
  INV_X1     g20197(.I(new_n20408_), .ZN(new_n20455_));
  AOI21_X1   g20198(.A1(new_n20448_), .A2(new_n20451_), .B(new_n20414_), .ZN(new_n20456_));
  NOR2_X1    g20199(.A1(new_n20452_), .A2(new_n20413_), .ZN(new_n20457_));
  NOR2_X1    g20200(.A1(new_n20457_), .A2(new_n20456_), .ZN(new_n20458_));
  NOR2_X1    g20201(.A1(new_n20458_), .A2(new_n20455_), .ZN(new_n20459_));
  NOR2_X1    g20202(.A1(new_n20454_), .A2(new_n20459_), .ZN(new_n20460_));
  XOR2_X1    g20203(.A1(new_n20460_), .A2(new_n20407_), .Z(new_n20461_));
  NOR2_X1    g20204(.A1(new_n20461_), .A2(new_n20405_), .ZN(new_n20462_));
  INV_X1     g20205(.I(new_n20407_), .ZN(new_n20463_));
  NOR2_X1    g20206(.A1(new_n20460_), .A2(new_n20463_), .ZN(new_n20464_));
  INV_X1     g20207(.I(new_n20464_), .ZN(new_n20465_));
  NAND2_X1   g20208(.A1(new_n20460_), .A2(new_n20463_), .ZN(new_n20466_));
  NAND2_X1   g20209(.A1(new_n20465_), .A2(new_n20466_), .ZN(new_n20467_));
  AOI21_X1   g20210(.A1(new_n20405_), .A2(new_n20467_), .B(new_n20462_), .ZN(new_n20468_));
  INV_X1     g20211(.I(new_n20328_), .ZN(new_n20469_));
  NOR2_X1    g20212(.A1(new_n20469_), .A2(new_n20390_), .ZN(new_n20470_));
  XOR2_X1    g20213(.A1(new_n20391_), .A2(new_n5220_), .Z(new_n20471_));
  NOR4_X1    g20214(.A1(new_n20386_), .A2(new_n20328_), .A3(new_n20389_), .A4(new_n20471_), .ZN(new_n20472_));
  NOR2_X1    g20215(.A1(new_n20470_), .A2(new_n20472_), .ZN(new_n20473_));
  XOR2_X1    g20216(.A1(new_n20468_), .A2(new_n20473_), .Z(new_n20474_));
  INV_X1     g20217(.I(new_n20474_), .ZN(new_n20475_));
  INV_X1     g20218(.I(new_n20394_), .ZN(new_n20476_));
  NAND2_X1   g20219(.A1(new_n20327_), .A2(new_n20476_), .ZN(new_n20477_));
  XOR2_X1    g20220(.A1(new_n20477_), .A2(new_n20475_), .Z(new_n20478_));
  XOR2_X1    g20221(.A1(new_n20327_), .A2(new_n20476_), .Z(new_n20479_));
  NAND2_X1   g20222(.A1(new_n20479_), .A2(new_n20395_), .ZN(new_n20480_));
  XOR2_X1    g20223(.A1(new_n20478_), .A2(new_n20480_), .Z(\f[114] ));
  NOR2_X1    g20224(.A1(new_n6012_), .A2(new_n8932_), .ZN(new_n20482_));
  NOR2_X1    g20225(.A1(new_n5792_), .A2(new_n8956_), .ZN(new_n20483_));
  NOR4_X1    g20226(.A1(new_n9323_), .A2(new_n5796_), .A3(new_n20482_), .A4(new_n20483_), .ZN(new_n20484_));
  XOR2_X1    g20227(.A1(new_n20484_), .A2(new_n5783_), .Z(new_n20485_));
  INV_X1     g20228(.I(new_n20456_), .ZN(new_n20486_));
  AOI21_X1   g20229(.A1(new_n20486_), .A2(new_n20455_), .B(new_n20457_), .ZN(new_n20487_));
  INV_X1     g20230(.I(new_n20487_), .ZN(new_n20488_));
  OAI22_X1   g20231(.A1(new_n6721_), .A2(new_n7930_), .B1(new_n6723_), .B2(new_n8548_), .ZN(new_n20489_));
  NAND2_X1   g20232(.A1(new_n7617_), .A2(\b[59] ), .ZN(new_n20490_));
  AOI21_X1   g20233(.A1(new_n20490_), .A2(new_n20489_), .B(new_n6731_), .ZN(new_n20491_));
  NAND2_X1   g20234(.A1(new_n8550_), .A2(new_n20491_), .ZN(new_n20492_));
  XOR2_X1    g20235(.A1(new_n20492_), .A2(\a[56] ), .Z(new_n20493_));
  NOR2_X1    g20236(.A1(new_n20449_), .A2(new_n20415_), .ZN(new_n20494_));
  NOR2_X1    g20237(.A1(new_n20494_), .A2(new_n20450_), .ZN(new_n20495_));
  OAI22_X1   g20238(.A1(new_n7560_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n7305_), .ZN(new_n20496_));
  NAND2_X1   g20239(.A1(new_n8628_), .A2(\b[56] ), .ZN(new_n20497_));
  AOI21_X1   g20240(.A1(new_n20497_), .A2(new_n20496_), .B(new_n7354_), .ZN(new_n20498_));
  NAND2_X1   g20241(.A1(new_n7559_), .A2(new_n20498_), .ZN(new_n20499_));
  XOR2_X1    g20242(.A1(new_n20499_), .A2(\a[59] ), .Z(new_n20500_));
  NOR2_X1    g20243(.A1(new_n20443_), .A2(new_n20426_), .ZN(new_n20501_));
  NOR2_X1    g20244(.A1(new_n20501_), .A2(new_n20444_), .ZN(new_n20502_));
  OAI22_X1   g20245(.A1(new_n6467_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n6238_), .ZN(new_n20503_));
  NAND2_X1   g20246(.A1(new_n9644_), .A2(\b[53] ), .ZN(new_n20504_));
  AOI21_X1   g20247(.A1(new_n20504_), .A2(new_n20503_), .B(new_n8321_), .ZN(new_n20505_));
  NAND2_X1   g20248(.A1(new_n6471_), .A2(new_n20505_), .ZN(new_n20506_));
  XOR2_X1    g20249(.A1(new_n20506_), .A2(\a[62] ), .Z(new_n20507_));
  NAND2_X1   g20250(.A1(new_n20437_), .A2(new_n20275_), .ZN(new_n20508_));
  NAND2_X1   g20251(.A1(new_n20508_), .A2(new_n20436_), .ZN(new_n20509_));
  NOR3_X1    g20252(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n5738_), .ZN(new_n20510_));
  NOR2_X1    g20253(.A1(new_n9364_), .A2(new_n5738_), .ZN(new_n20511_));
  NOR3_X1    g20254(.A1(new_n20511_), .A2(new_n5955_), .A3(new_n8985_), .ZN(new_n20512_));
  NOR2_X1    g20255(.A1(new_n20512_), .A2(new_n20510_), .ZN(new_n20513_));
  INV_X1     g20256(.I(new_n20513_), .ZN(new_n20514_));
  XOR2_X1    g20257(.A1(new_n20509_), .A2(new_n20514_), .Z(new_n20515_));
  NOR2_X1    g20258(.A1(new_n20507_), .A2(new_n20515_), .ZN(new_n20516_));
  NOR2_X1    g20259(.A1(new_n20509_), .A2(new_n20513_), .ZN(new_n20517_));
  INV_X1     g20260(.I(new_n20517_), .ZN(new_n20518_));
  NAND2_X1   g20261(.A1(new_n20509_), .A2(new_n20513_), .ZN(new_n20519_));
  NAND2_X1   g20262(.A1(new_n20518_), .A2(new_n20519_), .ZN(new_n20520_));
  AOI21_X1   g20263(.A1(new_n20507_), .A2(new_n20520_), .B(new_n20516_), .ZN(new_n20521_));
  XOR2_X1    g20264(.A1(new_n20502_), .A2(new_n20521_), .Z(new_n20522_));
  NOR2_X1    g20265(.A1(new_n20522_), .A2(new_n20500_), .ZN(new_n20523_));
  INV_X1     g20266(.I(new_n20502_), .ZN(new_n20524_));
  NOR2_X1    g20267(.A1(new_n20524_), .A2(new_n20521_), .ZN(new_n20525_));
  INV_X1     g20268(.I(new_n20525_), .ZN(new_n20526_));
  NAND2_X1   g20269(.A1(new_n20524_), .A2(new_n20521_), .ZN(new_n20527_));
  NAND2_X1   g20270(.A1(new_n20526_), .A2(new_n20527_), .ZN(new_n20528_));
  AOI21_X1   g20271(.A1(new_n20500_), .A2(new_n20528_), .B(new_n20523_), .ZN(new_n20529_));
  XOR2_X1    g20272(.A1(new_n20529_), .A2(new_n20495_), .Z(new_n20530_));
  NOR2_X1    g20273(.A1(new_n20530_), .A2(new_n20493_), .ZN(new_n20531_));
  INV_X1     g20274(.I(new_n20493_), .ZN(new_n20532_));
  INV_X1     g20275(.I(new_n20495_), .ZN(new_n20533_));
  NOR2_X1    g20276(.A1(new_n20533_), .A2(new_n20529_), .ZN(new_n20534_));
  INV_X1     g20277(.I(new_n20534_), .ZN(new_n20535_));
  NAND2_X1   g20278(.A1(new_n20533_), .A2(new_n20529_), .ZN(new_n20536_));
  AOI21_X1   g20279(.A1(new_n20535_), .A2(new_n20536_), .B(new_n20532_), .ZN(new_n20537_));
  NOR2_X1    g20280(.A1(new_n20531_), .A2(new_n20537_), .ZN(new_n20538_));
  NOR2_X1    g20281(.A1(new_n20538_), .A2(new_n20488_), .ZN(new_n20539_));
  INV_X1     g20282(.I(new_n20538_), .ZN(new_n20540_));
  NOR2_X1    g20283(.A1(new_n20540_), .A2(new_n20487_), .ZN(new_n20541_));
  NOR2_X1    g20284(.A1(new_n20541_), .A2(new_n20539_), .ZN(new_n20542_));
  NOR2_X1    g20285(.A1(new_n20542_), .A2(new_n20485_), .ZN(new_n20543_));
  INV_X1     g20286(.I(new_n20485_), .ZN(new_n20544_));
  XOR2_X1    g20287(.A1(new_n20538_), .A2(new_n20487_), .Z(new_n20545_));
  NOR2_X1    g20288(.A1(new_n20545_), .A2(new_n20544_), .ZN(new_n20546_));
  NOR2_X1    g20289(.A1(new_n20543_), .A2(new_n20546_), .ZN(new_n20547_));
  OAI21_X1   g20290(.A1(new_n20405_), .A2(new_n20464_), .B(new_n20466_), .ZN(new_n20548_));
  INV_X1     g20291(.I(new_n20058_), .ZN(new_n20549_));
  INV_X1     g20292(.I(new_n20060_), .ZN(new_n20550_));
  OAI21_X1   g20293(.A1(new_n20051_), .A2(new_n20550_), .B(new_n20549_), .ZN(new_n20551_));
  INV_X1     g20294(.I(new_n20140_), .ZN(new_n20552_));
  NAND3_X1   g20295(.A1(new_n20551_), .A2(new_n20552_), .A3(new_n20314_), .ZN(new_n20553_));
  AOI21_X1   g20296(.A1(new_n20553_), .A2(new_n20325_), .B(new_n20322_), .ZN(new_n20554_));
  NOR2_X1    g20297(.A1(new_n20475_), .A2(new_n20396_), .ZN(new_n20555_));
  NOR3_X1    g20298(.A1(new_n20554_), .A2(new_n20394_), .A3(new_n20555_), .ZN(new_n20556_));
  NOR3_X1    g20299(.A1(new_n20468_), .A2(new_n20470_), .A3(new_n20472_), .ZN(new_n20557_));
  NOR2_X1    g20300(.A1(new_n20556_), .A2(new_n20557_), .ZN(new_n20558_));
  XOR2_X1    g20301(.A1(new_n20558_), .A2(new_n20548_), .Z(new_n20559_));
  XOR2_X1    g20302(.A1(new_n20559_), .A2(new_n20547_), .Z(\f[115] ));
  INV_X1     g20303(.I(new_n20555_), .ZN(new_n20561_));
  NAND3_X1   g20304(.A1(new_n20327_), .A2(new_n20476_), .A3(new_n20561_), .ZN(new_n20562_));
  NOR2_X1    g20305(.A1(new_n20547_), .A2(new_n20548_), .ZN(new_n20563_));
  XOR2_X1    g20306(.A1(new_n20547_), .A2(new_n20548_), .Z(new_n20564_));
  NOR2_X1    g20307(.A1(new_n20564_), .A2(new_n20557_), .ZN(new_n20565_));
  AOI21_X1   g20308(.A1(new_n20562_), .A2(new_n20565_), .B(new_n20563_), .ZN(new_n20566_));
  OAI21_X1   g20309(.A1(new_n20493_), .A2(new_n20534_), .B(new_n20536_), .ZN(new_n20567_));
  OAI22_X1   g20310(.A1(new_n6721_), .A2(new_n8548_), .B1(new_n6723_), .B2(new_n8932_), .ZN(new_n20568_));
  NAND2_X1   g20311(.A1(new_n7617_), .A2(\b[60] ), .ZN(new_n20569_));
  AOI21_X1   g20312(.A1(new_n20569_), .A2(new_n20568_), .B(new_n6731_), .ZN(new_n20570_));
  NAND2_X1   g20313(.A1(new_n8935_), .A2(new_n20570_), .ZN(new_n20571_));
  XOR2_X1    g20314(.A1(new_n20571_), .A2(\a[56] ), .Z(new_n20572_));
  OAI21_X1   g20315(.A1(new_n20500_), .A2(new_n20525_), .B(new_n20527_), .ZN(new_n20573_));
  OAI21_X1   g20316(.A1(new_n20507_), .A2(new_n20517_), .B(new_n20519_), .ZN(new_n20574_));
  NOR3_X1    g20317(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n5955_), .ZN(new_n20575_));
  NOR2_X1    g20318(.A1(new_n9364_), .A2(new_n5955_), .ZN(new_n20576_));
  NOR3_X1    g20319(.A1(new_n20576_), .A2(new_n6215_), .A3(new_n8985_), .ZN(new_n20577_));
  NOR2_X1    g20320(.A1(new_n20577_), .A2(new_n20575_), .ZN(new_n20578_));
  NOR2_X1    g20321(.A1(new_n20514_), .A2(new_n20578_), .ZN(new_n20579_));
  INV_X1     g20322(.I(new_n20578_), .ZN(new_n20580_));
  NOR2_X1    g20323(.A1(new_n20580_), .A2(new_n20513_), .ZN(new_n20581_));
  OAI21_X1   g20324(.A1(new_n20579_), .A2(new_n20581_), .B(new_n20574_), .ZN(new_n20582_));
  XOR2_X1    g20325(.A1(new_n20513_), .A2(new_n20578_), .Z(new_n20583_));
  OR2_X2     g20326(.A1(new_n20574_), .A2(new_n20583_), .Z(new_n20584_));
  NAND2_X1   g20327(.A1(new_n20584_), .A2(new_n20582_), .ZN(new_n20585_));
  OAI22_X1   g20328(.A1(new_n7890_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n7560_), .ZN(new_n20586_));
  NAND2_X1   g20329(.A1(new_n8628_), .A2(\b[57] ), .ZN(new_n20587_));
  AOI21_X1   g20330(.A1(new_n20587_), .A2(new_n20586_), .B(new_n7354_), .ZN(new_n20588_));
  NAND2_X1   g20331(.A1(new_n7895_), .A2(new_n20588_), .ZN(new_n20589_));
  XOR2_X1    g20332(.A1(new_n20589_), .A2(\a[59] ), .Z(new_n20590_));
  OAI22_X1   g20333(.A1(new_n6995_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n6467_), .ZN(new_n20591_));
  NAND2_X1   g20334(.A1(new_n9644_), .A2(\b[54] ), .ZN(new_n20592_));
  AOI21_X1   g20335(.A1(new_n20592_), .A2(new_n20591_), .B(new_n8321_), .ZN(new_n20593_));
  NAND2_X1   g20336(.A1(new_n6994_), .A2(new_n20593_), .ZN(new_n20594_));
  XOR2_X1    g20337(.A1(new_n20594_), .A2(\a[62] ), .Z(new_n20595_));
  XNOR2_X1   g20338(.A1(new_n20590_), .A2(new_n20595_), .ZN(new_n20596_));
  INV_X1     g20339(.I(new_n20596_), .ZN(new_n20597_));
  NOR2_X1    g20340(.A1(new_n20590_), .A2(new_n20595_), .ZN(new_n20598_));
  INV_X1     g20341(.I(new_n20598_), .ZN(new_n20599_));
  NAND2_X1   g20342(.A1(new_n20590_), .A2(new_n20595_), .ZN(new_n20600_));
  AOI21_X1   g20343(.A1(new_n20599_), .A2(new_n20600_), .B(new_n20585_), .ZN(new_n20601_));
  AOI21_X1   g20344(.A1(new_n20597_), .A2(new_n20585_), .B(new_n20601_), .ZN(new_n20602_));
  NOR2_X1    g20345(.A1(new_n20573_), .A2(new_n20602_), .ZN(new_n20603_));
  INV_X1     g20346(.I(new_n20603_), .ZN(new_n20604_));
  NAND2_X1   g20347(.A1(new_n20573_), .A2(new_n20602_), .ZN(new_n20605_));
  AOI21_X1   g20348(.A1(new_n20604_), .A2(new_n20605_), .B(new_n20572_), .ZN(new_n20606_));
  INV_X1     g20349(.I(new_n20572_), .ZN(new_n20607_));
  XNOR2_X1   g20350(.A1(new_n20573_), .A2(new_n20602_), .ZN(new_n20608_));
  NOR2_X1    g20351(.A1(new_n20608_), .A2(new_n20607_), .ZN(new_n20609_));
  NOR2_X1    g20352(.A1(new_n20609_), .A2(new_n20606_), .ZN(new_n20610_));
  OAI22_X1   g20353(.A1(new_n9595_), .A2(new_n5796_), .B1(new_n8956_), .B2(new_n6012_), .ZN(new_n20611_));
  XOR2_X1    g20354(.A1(new_n20610_), .A2(new_n20611_), .Z(new_n20612_));
  XOR2_X1    g20355(.A1(new_n20612_), .A2(\a[53] ), .Z(new_n20613_));
  XOR2_X1    g20356(.A1(new_n20613_), .A2(new_n20567_), .Z(new_n20614_));
  NOR2_X1    g20357(.A1(new_n20539_), .A2(new_n20485_), .ZN(new_n20615_));
  NOR2_X1    g20358(.A1(new_n20615_), .A2(new_n20541_), .ZN(new_n20616_));
  INV_X1     g20359(.I(new_n20616_), .ZN(new_n20617_));
  XOR2_X1    g20360(.A1(new_n20614_), .A2(new_n20617_), .Z(new_n20618_));
  XOR2_X1    g20361(.A1(new_n20614_), .A2(new_n20617_), .Z(new_n20619_));
  NAND2_X1   g20362(.A1(new_n20566_), .A2(new_n20619_), .ZN(new_n20620_));
  OAI21_X1   g20363(.A1(new_n20566_), .A2(new_n20618_), .B(new_n20620_), .ZN(\f[116] ));
  INV_X1     g20364(.I(new_n20567_), .ZN(new_n20622_));
  NOR2_X1    g20365(.A1(new_n20622_), .A2(new_n20610_), .ZN(new_n20623_));
  XOR2_X1    g20366(.A1(new_n20611_), .A2(new_n5783_), .Z(new_n20624_));
  NOR4_X1    g20367(.A1(new_n20567_), .A2(new_n20606_), .A3(new_n20609_), .A4(new_n20624_), .ZN(new_n20625_));
  NOR2_X1    g20368(.A1(new_n20623_), .A2(new_n20625_), .ZN(new_n20626_));
  OAI21_X1   g20369(.A1(new_n20572_), .A2(new_n20603_), .B(new_n20605_), .ZN(new_n20627_));
  OAI22_X1   g20370(.A1(new_n6721_), .A2(new_n8932_), .B1(new_n6723_), .B2(new_n8956_), .ZN(new_n20628_));
  NAND2_X1   g20371(.A1(new_n7617_), .A2(\b[61] ), .ZN(new_n20629_));
  AOI21_X1   g20372(.A1(new_n20629_), .A2(new_n20628_), .B(new_n6731_), .ZN(new_n20630_));
  NAND2_X1   g20373(.A1(new_n8963_), .A2(new_n20630_), .ZN(new_n20631_));
  XOR2_X1    g20374(.A1(new_n20631_), .A2(\a[56] ), .Z(new_n20632_));
  AOI21_X1   g20375(.A1(new_n20585_), .A2(new_n20600_), .B(new_n20598_), .ZN(new_n20633_));
  OAI22_X1   g20376(.A1(new_n7930_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n7890_), .ZN(new_n20634_));
  NAND2_X1   g20377(.A1(new_n8628_), .A2(\b[58] ), .ZN(new_n20635_));
  AOI21_X1   g20378(.A1(new_n20635_), .A2(new_n20634_), .B(new_n7354_), .ZN(new_n20636_));
  NAND2_X1   g20379(.A1(new_n7929_), .A2(new_n20636_), .ZN(new_n20637_));
  XOR2_X1    g20380(.A1(new_n20637_), .A2(\a[59] ), .Z(new_n20638_));
  INV_X1     g20381(.I(new_n20638_), .ZN(new_n20639_));
  INV_X1     g20382(.I(new_n20579_), .ZN(new_n20640_));
  AOI21_X1   g20383(.A1(new_n20574_), .A2(new_n20640_), .B(new_n20581_), .ZN(new_n20641_));
  INV_X1     g20384(.I(new_n20641_), .ZN(new_n20642_));
  OAI22_X1   g20385(.A1(new_n7305_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n6995_), .ZN(new_n20643_));
  NAND2_X1   g20386(.A1(new_n9644_), .A2(\b[55] ), .ZN(new_n20644_));
  AOI21_X1   g20387(.A1(new_n20644_), .A2(new_n20643_), .B(new_n8321_), .ZN(new_n20645_));
  NAND2_X1   g20388(.A1(new_n7308_), .A2(new_n20645_), .ZN(new_n20646_));
  XOR2_X1    g20389(.A1(new_n20646_), .A2(\a[62] ), .Z(new_n20647_));
  NOR2_X1    g20390(.A1(new_n8985_), .A2(new_n6238_), .ZN(new_n20648_));
  NOR2_X1    g20391(.A1(new_n9364_), .A2(new_n6215_), .ZN(new_n20649_));
  XNOR2_X1   g20392(.A1(new_n20648_), .A2(new_n20649_), .ZN(new_n20650_));
  XOR2_X1    g20393(.A1(new_n20650_), .A2(\a[53] ), .Z(new_n20651_));
  NOR2_X1    g20394(.A1(new_n20651_), .A2(new_n20578_), .ZN(new_n20652_));
  NOR2_X1    g20395(.A1(new_n20650_), .A2(new_n5783_), .ZN(new_n20653_));
  INV_X1     g20396(.I(new_n20653_), .ZN(new_n20654_));
  NAND2_X1   g20397(.A1(new_n20650_), .A2(new_n5783_), .ZN(new_n20655_));
  AOI21_X1   g20398(.A1(new_n20654_), .A2(new_n20655_), .B(new_n20580_), .ZN(new_n20656_));
  NOR2_X1    g20399(.A1(new_n20652_), .A2(new_n20656_), .ZN(new_n20657_));
  INV_X1     g20400(.I(new_n20657_), .ZN(new_n20658_));
  XOR2_X1    g20401(.A1(new_n20647_), .A2(new_n20658_), .Z(new_n20659_));
  NAND2_X1   g20402(.A1(new_n20659_), .A2(new_n20642_), .ZN(new_n20660_));
  AND2_X2    g20403(.A1(new_n20647_), .A2(new_n20658_), .Z(new_n20661_));
  NOR2_X1    g20404(.A1(new_n20647_), .A2(new_n20658_), .ZN(new_n20662_));
  OAI21_X1   g20405(.A1(new_n20661_), .A2(new_n20662_), .B(new_n20641_), .ZN(new_n20663_));
  AOI21_X1   g20406(.A1(new_n20660_), .A2(new_n20663_), .B(new_n20639_), .ZN(new_n20664_));
  NAND2_X1   g20407(.A1(new_n20660_), .A2(new_n20663_), .ZN(new_n20665_));
  NOR2_X1    g20408(.A1(new_n20665_), .A2(new_n20638_), .ZN(new_n20666_));
  NOR2_X1    g20409(.A1(new_n20666_), .A2(new_n20664_), .ZN(new_n20667_));
  NOR2_X1    g20410(.A1(new_n20667_), .A2(new_n20633_), .ZN(new_n20668_));
  INV_X1     g20411(.I(new_n20633_), .ZN(new_n20669_));
  XOR2_X1    g20412(.A1(new_n20665_), .A2(new_n20639_), .Z(new_n20670_));
  NOR2_X1    g20413(.A1(new_n20670_), .A2(new_n20669_), .ZN(new_n20671_));
  NOR2_X1    g20414(.A1(new_n20671_), .A2(new_n20668_), .ZN(new_n20672_));
  NOR2_X1    g20415(.A1(new_n20672_), .A2(new_n20632_), .ZN(new_n20673_));
  NAND2_X1   g20416(.A1(new_n20672_), .A2(new_n20632_), .ZN(new_n20674_));
  INV_X1     g20417(.I(new_n20674_), .ZN(new_n20675_));
  OAI21_X1   g20418(.A1(new_n20675_), .A2(new_n20673_), .B(new_n20627_), .ZN(new_n20676_));
  XNOR2_X1   g20419(.A1(new_n20672_), .A2(new_n20632_), .ZN(new_n20677_));
  OAI21_X1   g20420(.A1(new_n20627_), .A2(new_n20677_), .B(new_n20676_), .ZN(new_n20678_));
  XOR2_X1    g20421(.A1(new_n20626_), .A2(new_n20678_), .Z(new_n20679_));
  NOR2_X1    g20422(.A1(new_n20566_), .A2(new_n20614_), .ZN(new_n20680_));
  XOR2_X1    g20423(.A1(new_n20680_), .A2(new_n20679_), .Z(new_n20681_));
  XOR2_X1    g20424(.A1(new_n20566_), .A2(new_n20614_), .Z(new_n20682_));
  NAND2_X1   g20425(.A1(new_n20682_), .A2(new_n20617_), .ZN(new_n20683_));
  XOR2_X1    g20426(.A1(new_n20681_), .A2(new_n20683_), .Z(\f[117] ));
  NOR2_X1    g20427(.A1(new_n6729_), .A2(new_n8932_), .ZN(new_n20685_));
  NOR2_X1    g20428(.A1(new_n6721_), .A2(new_n8956_), .ZN(new_n20686_));
  NOR4_X1    g20429(.A1(new_n9323_), .A2(new_n6731_), .A3(new_n20685_), .A4(new_n20686_), .ZN(new_n20687_));
  XOR2_X1    g20430(.A1(new_n20687_), .A2(new_n6516_), .Z(new_n20688_));
  INV_X1     g20431(.I(new_n20664_), .ZN(new_n20689_));
  AOI21_X1   g20432(.A1(new_n20689_), .A2(new_n20669_), .B(new_n20666_), .ZN(new_n20690_));
  INV_X1     g20433(.I(new_n20690_), .ZN(new_n20691_));
  OAI22_X1   g20434(.A1(new_n8548_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n7930_), .ZN(new_n20692_));
  NAND2_X1   g20435(.A1(new_n8628_), .A2(\b[59] ), .ZN(new_n20693_));
  AOI21_X1   g20436(.A1(new_n20693_), .A2(new_n20692_), .B(new_n7354_), .ZN(new_n20694_));
  NAND2_X1   g20437(.A1(new_n8550_), .A2(new_n20694_), .ZN(new_n20695_));
  XOR2_X1    g20438(.A1(new_n20695_), .A2(\a[59] ), .Z(new_n20696_));
  NOR2_X1    g20439(.A1(new_n20661_), .A2(new_n20641_), .ZN(new_n20697_));
  NOR2_X1    g20440(.A1(new_n20697_), .A2(new_n20662_), .ZN(new_n20698_));
  OAI22_X1   g20441(.A1(new_n7560_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n7305_), .ZN(new_n20699_));
  NAND2_X1   g20442(.A1(new_n9644_), .A2(\b[56] ), .ZN(new_n20700_));
  AOI21_X1   g20443(.A1(new_n20700_), .A2(new_n20699_), .B(new_n8321_), .ZN(new_n20701_));
  NAND2_X1   g20444(.A1(new_n7559_), .A2(new_n20701_), .ZN(new_n20702_));
  XOR2_X1    g20445(.A1(new_n20702_), .A2(new_n8309_), .Z(new_n20703_));
  NAND2_X1   g20446(.A1(new_n20655_), .A2(new_n20580_), .ZN(new_n20704_));
  NAND2_X1   g20447(.A1(new_n20704_), .A2(new_n20654_), .ZN(new_n20705_));
  NOR3_X1    g20448(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n6238_), .ZN(new_n20706_));
  NOR2_X1    g20449(.A1(new_n9364_), .A2(new_n6238_), .ZN(new_n20707_));
  NOR3_X1    g20450(.A1(new_n20707_), .A2(new_n6467_), .A3(new_n8985_), .ZN(new_n20708_));
  NOR2_X1    g20451(.A1(new_n20708_), .A2(new_n20706_), .ZN(new_n20709_));
  INV_X1     g20452(.I(new_n20709_), .ZN(new_n20710_));
  XOR2_X1    g20453(.A1(new_n20705_), .A2(new_n20710_), .Z(new_n20711_));
  INV_X1     g20454(.I(new_n20711_), .ZN(new_n20712_));
  NOR2_X1    g20455(.A1(new_n20705_), .A2(new_n20709_), .ZN(new_n20713_));
  INV_X1     g20456(.I(new_n20713_), .ZN(new_n20714_));
  NAND2_X1   g20457(.A1(new_n20705_), .A2(new_n20709_), .ZN(new_n20715_));
  AOI21_X1   g20458(.A1(new_n20714_), .A2(new_n20715_), .B(new_n20703_), .ZN(new_n20716_));
  AOI21_X1   g20459(.A1(new_n20703_), .A2(new_n20712_), .B(new_n20716_), .ZN(new_n20717_));
  XOR2_X1    g20460(.A1(new_n20698_), .A2(new_n20717_), .Z(new_n20718_));
  NOR2_X1    g20461(.A1(new_n20718_), .A2(new_n20696_), .ZN(new_n20719_));
  INV_X1     g20462(.I(new_n20698_), .ZN(new_n20720_));
  NOR2_X1    g20463(.A1(new_n20720_), .A2(new_n20717_), .ZN(new_n20721_));
  INV_X1     g20464(.I(new_n20721_), .ZN(new_n20722_));
  NAND2_X1   g20465(.A1(new_n20720_), .A2(new_n20717_), .ZN(new_n20723_));
  NAND2_X1   g20466(.A1(new_n20722_), .A2(new_n20723_), .ZN(new_n20724_));
  AOI21_X1   g20467(.A1(new_n20696_), .A2(new_n20724_), .B(new_n20719_), .ZN(new_n20725_));
  NOR2_X1    g20468(.A1(new_n20725_), .A2(new_n20691_), .ZN(new_n20726_));
  INV_X1     g20469(.I(new_n20726_), .ZN(new_n20727_));
  NAND2_X1   g20470(.A1(new_n20725_), .A2(new_n20691_), .ZN(new_n20728_));
  AOI21_X1   g20471(.A1(new_n20727_), .A2(new_n20728_), .B(new_n20688_), .ZN(new_n20729_));
  INV_X1     g20472(.I(new_n20688_), .ZN(new_n20730_));
  XOR2_X1    g20473(.A1(new_n20725_), .A2(new_n20690_), .Z(new_n20731_));
  NOR2_X1    g20474(.A1(new_n20731_), .A2(new_n20730_), .ZN(new_n20732_));
  NOR2_X1    g20475(.A1(new_n20732_), .A2(new_n20729_), .ZN(new_n20733_));
  AOI21_X1   g20476(.A1(new_n20627_), .A2(new_n20674_), .B(new_n20673_), .ZN(new_n20734_));
  INV_X1     g20477(.I(new_n20734_), .ZN(new_n20735_));
  NAND2_X1   g20478(.A1(new_n20617_), .A2(new_n20679_), .ZN(new_n20736_));
  INV_X1     g20479(.I(new_n20736_), .ZN(new_n20737_));
  NOR3_X1    g20480(.A1(new_n20566_), .A2(new_n20614_), .A3(new_n20737_), .ZN(new_n20738_));
  NOR3_X1    g20481(.A1(new_n20678_), .A2(new_n20623_), .A3(new_n20625_), .ZN(new_n20739_));
  NOR2_X1    g20482(.A1(new_n20738_), .A2(new_n20739_), .ZN(new_n20740_));
  XOR2_X1    g20483(.A1(new_n20740_), .A2(new_n20735_), .Z(new_n20741_));
  XOR2_X1    g20484(.A1(new_n20741_), .A2(new_n20733_), .Z(\f[118] ));
  NOR2_X1    g20485(.A1(new_n20733_), .A2(new_n20735_), .ZN(new_n20743_));
  INV_X1     g20486(.I(new_n20743_), .ZN(new_n20744_));
  XOR2_X1    g20487(.A1(new_n20733_), .A2(new_n20735_), .Z(new_n20745_));
  NOR2_X1    g20488(.A1(new_n20745_), .A2(new_n20739_), .ZN(new_n20746_));
  INV_X1     g20489(.I(new_n20746_), .ZN(new_n20747_));
  OAI21_X1   g20490(.A1(new_n20738_), .A2(new_n20747_), .B(new_n20744_), .ZN(new_n20748_));
  OAI21_X1   g20491(.A1(new_n20696_), .A2(new_n20721_), .B(new_n20723_), .ZN(new_n20749_));
  OAI22_X1   g20492(.A1(new_n8932_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n8548_), .ZN(new_n20750_));
  NAND2_X1   g20493(.A1(new_n8628_), .A2(\b[60] ), .ZN(new_n20751_));
  AOI21_X1   g20494(.A1(new_n20751_), .A2(new_n20750_), .B(new_n7354_), .ZN(new_n20752_));
  NAND2_X1   g20495(.A1(new_n8935_), .A2(new_n20752_), .ZN(new_n20753_));
  XOR2_X1    g20496(.A1(new_n20753_), .A2(\a[59] ), .Z(new_n20754_));
  OAI22_X1   g20497(.A1(new_n7890_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n7560_), .ZN(new_n20755_));
  NAND2_X1   g20498(.A1(new_n9644_), .A2(\b[57] ), .ZN(new_n20756_));
  AOI21_X1   g20499(.A1(new_n20756_), .A2(new_n20755_), .B(new_n8321_), .ZN(new_n20757_));
  NAND2_X1   g20500(.A1(new_n7895_), .A2(new_n20757_), .ZN(new_n20758_));
  XOR2_X1    g20501(.A1(new_n20758_), .A2(\a[62] ), .Z(new_n20759_));
  NOR3_X1    g20502(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n6467_), .ZN(new_n20760_));
  NOR2_X1    g20503(.A1(new_n9364_), .A2(new_n6467_), .ZN(new_n20761_));
  NOR3_X1    g20504(.A1(new_n20761_), .A2(new_n6995_), .A3(new_n8985_), .ZN(new_n20762_));
  NOR2_X1    g20505(.A1(new_n20762_), .A2(new_n20760_), .ZN(new_n20763_));
  NOR2_X1    g20506(.A1(new_n20710_), .A2(new_n20763_), .ZN(new_n20764_));
  NOR3_X1    g20507(.A1(new_n20709_), .A2(new_n20760_), .A3(new_n20762_), .ZN(new_n20765_));
  NOR2_X1    g20508(.A1(new_n20764_), .A2(new_n20765_), .ZN(new_n20766_));
  NOR2_X1    g20509(.A1(new_n20759_), .A2(new_n20766_), .ZN(new_n20767_));
  INV_X1     g20510(.I(new_n20759_), .ZN(new_n20768_));
  XOR2_X1    g20511(.A1(new_n20709_), .A2(new_n20763_), .Z(new_n20769_));
  NOR2_X1    g20512(.A1(new_n20768_), .A2(new_n20769_), .ZN(new_n20770_));
  NOR2_X1    g20513(.A1(new_n20770_), .A2(new_n20767_), .ZN(new_n20771_));
  INV_X1     g20514(.I(new_n20715_), .ZN(new_n20772_));
  AOI21_X1   g20515(.A1(new_n20703_), .A2(new_n20714_), .B(new_n20772_), .ZN(new_n20773_));
  NOR2_X1    g20516(.A1(new_n20771_), .A2(new_n20773_), .ZN(new_n20774_));
  INV_X1     g20517(.I(new_n20774_), .ZN(new_n20775_));
  NAND2_X1   g20518(.A1(new_n20771_), .A2(new_n20773_), .ZN(new_n20776_));
  AOI21_X1   g20519(.A1(new_n20775_), .A2(new_n20776_), .B(new_n20754_), .ZN(new_n20777_));
  INV_X1     g20520(.I(new_n20754_), .ZN(new_n20778_));
  XNOR2_X1   g20521(.A1(new_n20771_), .A2(new_n20773_), .ZN(new_n20779_));
  NOR2_X1    g20522(.A1(new_n20779_), .A2(new_n20778_), .ZN(new_n20780_));
  NOR2_X1    g20523(.A1(new_n20780_), .A2(new_n20777_), .ZN(new_n20781_));
  OAI22_X1   g20524(.A1(new_n9595_), .A2(new_n6731_), .B1(new_n8956_), .B2(new_n6729_), .ZN(new_n20782_));
  XOR2_X1    g20525(.A1(new_n20781_), .A2(new_n20782_), .Z(new_n20783_));
  XOR2_X1    g20526(.A1(new_n20783_), .A2(\a[56] ), .Z(new_n20784_));
  XOR2_X1    g20527(.A1(new_n20784_), .A2(new_n20749_), .Z(new_n20785_));
  OAI21_X1   g20528(.A1(new_n20688_), .A2(new_n20726_), .B(new_n20728_), .ZN(new_n20786_));
  INV_X1     g20529(.I(new_n20786_), .ZN(new_n20787_));
  XOR2_X1    g20530(.A1(new_n20785_), .A2(new_n20787_), .Z(new_n20788_));
  NAND2_X1   g20531(.A1(new_n20748_), .A2(new_n20788_), .ZN(new_n20789_));
  XOR2_X1    g20532(.A1(new_n20785_), .A2(new_n20787_), .Z(new_n20790_));
  OAI21_X1   g20533(.A1(new_n20748_), .A2(new_n20790_), .B(new_n20789_), .ZN(\f[119] ));
  AOI21_X1   g20534(.A1(new_n20778_), .A2(new_n20776_), .B(new_n20774_), .ZN(new_n20792_));
  INV_X1     g20535(.I(new_n20792_), .ZN(new_n20793_));
  OAI22_X1   g20536(.A1(new_n8956_), .A2(new_n7346_), .B1(new_n7351_), .B2(new_n8932_), .ZN(new_n20794_));
  NAND2_X1   g20537(.A1(new_n8628_), .A2(\b[61] ), .ZN(new_n20795_));
  AOI21_X1   g20538(.A1(new_n20795_), .A2(new_n20794_), .B(new_n7354_), .ZN(new_n20796_));
  NAND2_X1   g20539(.A1(new_n8963_), .A2(new_n20796_), .ZN(new_n20797_));
  XOR2_X1    g20540(.A1(new_n20797_), .A2(\a[59] ), .Z(new_n20798_));
  INV_X1     g20541(.I(new_n20798_), .ZN(new_n20799_));
  NOR2_X1    g20542(.A1(new_n20759_), .A2(new_n20765_), .ZN(new_n20800_));
  NOR2_X1    g20543(.A1(new_n20800_), .A2(new_n20764_), .ZN(new_n20801_));
  INV_X1     g20544(.I(new_n20801_), .ZN(new_n20802_));
  OAI22_X1   g20545(.A1(new_n7930_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n7890_), .ZN(new_n20803_));
  NAND2_X1   g20546(.A1(new_n9644_), .A2(\b[58] ), .ZN(new_n20804_));
  AOI21_X1   g20547(.A1(new_n20804_), .A2(new_n20803_), .B(new_n8321_), .ZN(new_n20805_));
  NAND2_X1   g20548(.A1(new_n7929_), .A2(new_n20805_), .ZN(new_n20806_));
  XOR2_X1    g20549(.A1(new_n20806_), .A2(\a[62] ), .Z(new_n20807_));
  NOR2_X1    g20550(.A1(new_n8985_), .A2(new_n7305_), .ZN(new_n20808_));
  NOR2_X1    g20551(.A1(new_n9364_), .A2(new_n6995_), .ZN(new_n20809_));
  XNOR2_X1   g20552(.A1(new_n20808_), .A2(new_n20809_), .ZN(new_n20810_));
  NOR2_X1    g20553(.A1(new_n20810_), .A2(new_n6516_), .ZN(new_n20811_));
  INV_X1     g20554(.I(new_n20811_), .ZN(new_n20812_));
  NAND2_X1   g20555(.A1(new_n20810_), .A2(new_n6516_), .ZN(new_n20813_));
  AOI21_X1   g20556(.A1(new_n20812_), .A2(new_n20813_), .B(new_n20709_), .ZN(new_n20814_));
  XOR2_X1    g20557(.A1(new_n20810_), .A2(\a[56] ), .Z(new_n20815_));
  NOR2_X1    g20558(.A1(new_n20815_), .A2(new_n20710_), .ZN(new_n20816_));
  NOR2_X1    g20559(.A1(new_n20816_), .A2(new_n20814_), .ZN(new_n20817_));
  XOR2_X1    g20560(.A1(new_n20807_), .A2(new_n20817_), .Z(new_n20818_));
  NOR2_X1    g20561(.A1(new_n20807_), .A2(new_n20817_), .ZN(new_n20819_));
  INV_X1     g20562(.I(new_n20819_), .ZN(new_n20820_));
  NAND2_X1   g20563(.A1(new_n20807_), .A2(new_n20817_), .ZN(new_n20821_));
  AOI21_X1   g20564(.A1(new_n20820_), .A2(new_n20821_), .B(new_n20802_), .ZN(new_n20822_));
  AOI21_X1   g20565(.A1(new_n20802_), .A2(new_n20818_), .B(new_n20822_), .ZN(new_n20823_));
  NOR2_X1    g20566(.A1(new_n20823_), .A2(new_n20799_), .ZN(new_n20824_));
  AND2_X2    g20567(.A1(new_n20823_), .A2(new_n20799_), .Z(new_n20825_));
  OAI21_X1   g20568(.A1(new_n20825_), .A2(new_n20824_), .B(new_n20793_), .ZN(new_n20826_));
  XOR2_X1    g20569(.A1(new_n20823_), .A2(new_n20798_), .Z(new_n20827_));
  OAI21_X1   g20570(.A1(new_n20793_), .A2(new_n20827_), .B(new_n20826_), .ZN(new_n20828_));
  INV_X1     g20571(.I(new_n20749_), .ZN(new_n20829_));
  XOR2_X1    g20572(.A1(new_n20782_), .A2(\a[56] ), .Z(new_n20830_));
  NAND3_X1   g20573(.A1(new_n20781_), .A2(new_n20829_), .A3(new_n20830_), .ZN(new_n20831_));
  OAI21_X1   g20574(.A1(new_n20829_), .A2(new_n20781_), .B(new_n20831_), .ZN(new_n20832_));
  XNOR2_X1   g20575(.A1(new_n20828_), .A2(new_n20832_), .ZN(new_n20833_));
  INV_X1     g20576(.I(new_n20833_), .ZN(new_n20834_));
  INV_X1     g20577(.I(new_n20785_), .ZN(new_n20835_));
  NAND2_X1   g20578(.A1(new_n20748_), .A2(new_n20835_), .ZN(new_n20836_));
  XOR2_X1    g20579(.A1(new_n20836_), .A2(new_n20834_), .Z(new_n20837_));
  XOR2_X1    g20580(.A1(new_n20748_), .A2(new_n20835_), .Z(new_n20838_));
  NAND2_X1   g20581(.A1(new_n20838_), .A2(new_n20786_), .ZN(new_n20839_));
  XOR2_X1    g20582(.A1(new_n20837_), .A2(new_n20839_), .Z(\f[120] ));
  NOR2_X1    g20583(.A1(new_n7611_), .A2(new_n8932_), .ZN(new_n20841_));
  NOR2_X1    g20584(.A1(new_n7351_), .A2(new_n8956_), .ZN(new_n20842_));
  NOR4_X1    g20585(.A1(new_n9323_), .A2(new_n7354_), .A3(new_n20841_), .A4(new_n20842_), .ZN(new_n20843_));
  XOR2_X1    g20586(.A1(new_n20843_), .A2(new_n7343_), .Z(new_n20844_));
  NAND2_X1   g20587(.A1(new_n20802_), .A2(new_n20821_), .ZN(new_n20845_));
  NAND2_X1   g20588(.A1(new_n20845_), .A2(new_n20820_), .ZN(new_n20846_));
  INV_X1     g20589(.I(new_n20846_), .ZN(new_n20847_));
  OAI22_X1   g20590(.A1(new_n8548_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n7930_), .ZN(new_n20848_));
  NAND2_X1   g20591(.A1(new_n9644_), .A2(\b[59] ), .ZN(new_n20849_));
  AOI21_X1   g20592(.A1(new_n20849_), .A2(new_n20848_), .B(new_n8321_), .ZN(new_n20850_));
  NAND2_X1   g20593(.A1(new_n8550_), .A2(new_n20850_), .ZN(new_n20851_));
  XOR2_X1    g20594(.A1(new_n20851_), .A2(\a[62] ), .Z(new_n20852_));
  NAND2_X1   g20595(.A1(new_n20813_), .A2(new_n20710_), .ZN(new_n20853_));
  NAND2_X1   g20596(.A1(new_n20853_), .A2(new_n20812_), .ZN(new_n20854_));
  NOR3_X1    g20597(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n7305_), .ZN(new_n20855_));
  NOR2_X1    g20598(.A1(new_n9364_), .A2(new_n7305_), .ZN(new_n20856_));
  NOR3_X1    g20599(.A1(new_n20856_), .A2(new_n7560_), .A3(new_n8985_), .ZN(new_n20857_));
  NOR2_X1    g20600(.A1(new_n20857_), .A2(new_n20855_), .ZN(new_n20858_));
  INV_X1     g20601(.I(new_n20858_), .ZN(new_n20859_));
  XOR2_X1    g20602(.A1(new_n20854_), .A2(new_n20859_), .Z(new_n20860_));
  NOR2_X1    g20603(.A1(new_n20854_), .A2(new_n20858_), .ZN(new_n20861_));
  NAND2_X1   g20604(.A1(new_n20854_), .A2(new_n20858_), .ZN(new_n20862_));
  INV_X1     g20605(.I(new_n20862_), .ZN(new_n20863_));
  OAI21_X1   g20606(.A1(new_n20861_), .A2(new_n20863_), .B(new_n20852_), .ZN(new_n20864_));
  OAI21_X1   g20607(.A1(new_n20852_), .A2(new_n20860_), .B(new_n20864_), .ZN(new_n20865_));
  NAND2_X1   g20608(.A1(new_n20865_), .A2(new_n20847_), .ZN(new_n20866_));
  NOR2_X1    g20609(.A1(new_n20865_), .A2(new_n20847_), .ZN(new_n20867_));
  INV_X1     g20610(.I(new_n20867_), .ZN(new_n20868_));
  AOI21_X1   g20611(.A1(new_n20868_), .A2(new_n20866_), .B(new_n20844_), .ZN(new_n20869_));
  INV_X1     g20612(.I(new_n20844_), .ZN(new_n20870_));
  XOR2_X1    g20613(.A1(new_n20865_), .A2(new_n20846_), .Z(new_n20871_));
  NOR2_X1    g20614(.A1(new_n20871_), .A2(new_n20870_), .ZN(new_n20872_));
  NOR2_X1    g20615(.A1(new_n20872_), .A2(new_n20869_), .ZN(new_n20873_));
  NOR2_X1    g20616(.A1(new_n20824_), .A2(new_n20792_), .ZN(new_n20874_));
  NOR2_X1    g20617(.A1(new_n20874_), .A2(new_n20825_), .ZN(new_n20875_));
  INV_X1     g20618(.I(new_n20875_), .ZN(new_n20876_));
  INV_X1     g20619(.I(new_n20563_), .ZN(new_n20877_));
  INV_X1     g20620(.I(new_n20565_), .ZN(new_n20878_));
  OAI21_X1   g20621(.A1(new_n20556_), .A2(new_n20878_), .B(new_n20877_), .ZN(new_n20879_));
  INV_X1     g20622(.I(new_n20614_), .ZN(new_n20880_));
  NAND3_X1   g20623(.A1(new_n20879_), .A2(new_n20880_), .A3(new_n20736_), .ZN(new_n20881_));
  AOI21_X1   g20624(.A1(new_n20881_), .A2(new_n20746_), .B(new_n20743_), .ZN(new_n20882_));
  NOR2_X1    g20625(.A1(new_n20834_), .A2(new_n20787_), .ZN(new_n20883_));
  NOR3_X1    g20626(.A1(new_n20882_), .A2(new_n20785_), .A3(new_n20883_), .ZN(new_n20884_));
  NOR2_X1    g20627(.A1(new_n20828_), .A2(new_n20832_), .ZN(new_n20885_));
  NOR2_X1    g20628(.A1(new_n20884_), .A2(new_n20885_), .ZN(new_n20886_));
  XOR2_X1    g20629(.A1(new_n20886_), .A2(new_n20876_), .Z(new_n20887_));
  XOR2_X1    g20630(.A1(new_n20887_), .A2(new_n20873_), .Z(\f[121] ));
  INV_X1     g20631(.I(new_n20883_), .ZN(new_n20889_));
  NAND3_X1   g20632(.A1(new_n20748_), .A2(new_n20835_), .A3(new_n20889_), .ZN(new_n20890_));
  NOR2_X1    g20633(.A1(new_n20873_), .A2(new_n20876_), .ZN(new_n20891_));
  XOR2_X1    g20634(.A1(new_n20873_), .A2(new_n20876_), .Z(new_n20892_));
  NOR2_X1    g20635(.A1(new_n20892_), .A2(new_n20885_), .ZN(new_n20893_));
  AOI21_X1   g20636(.A1(new_n20890_), .A2(new_n20893_), .B(new_n20891_), .ZN(new_n20894_));
  AOI21_X1   g20637(.A1(new_n20870_), .A2(new_n20866_), .B(new_n20867_), .ZN(new_n20895_));
  OAI22_X1   g20638(.A1(new_n8932_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n8548_), .ZN(new_n20896_));
  NAND2_X1   g20639(.A1(new_n9644_), .A2(\b[60] ), .ZN(new_n20897_));
  AOI21_X1   g20640(.A1(new_n20897_), .A2(new_n20896_), .B(new_n8321_), .ZN(new_n20898_));
  NAND2_X1   g20641(.A1(new_n8935_), .A2(new_n20898_), .ZN(new_n20899_));
  XOR2_X1    g20642(.A1(new_n20899_), .A2(\a[62] ), .Z(new_n20900_));
  INV_X1     g20643(.I(new_n20900_), .ZN(new_n20901_));
  OAI21_X1   g20644(.A1(new_n20852_), .A2(new_n20861_), .B(new_n20862_), .ZN(new_n20902_));
  INV_X1     g20645(.I(new_n20902_), .ZN(new_n20903_));
  NOR3_X1    g20646(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n7560_), .ZN(new_n20904_));
  NOR2_X1    g20647(.A1(new_n9364_), .A2(new_n7560_), .ZN(new_n20905_));
  NOR3_X1    g20648(.A1(new_n20905_), .A2(new_n7890_), .A3(new_n8985_), .ZN(new_n20906_));
  NOR2_X1    g20649(.A1(new_n20906_), .A2(new_n20904_), .ZN(new_n20907_));
  NOR2_X1    g20650(.A1(new_n20859_), .A2(new_n20907_), .ZN(new_n20908_));
  INV_X1     g20651(.I(new_n20907_), .ZN(new_n20909_));
  NOR2_X1    g20652(.A1(new_n20909_), .A2(new_n20858_), .ZN(new_n20910_));
  NOR2_X1    g20653(.A1(new_n20908_), .A2(new_n20910_), .ZN(new_n20911_));
  NOR2_X1    g20654(.A1(new_n20903_), .A2(new_n20911_), .ZN(new_n20912_));
  XOR2_X1    g20655(.A1(new_n20858_), .A2(new_n20907_), .Z(new_n20913_));
  NOR2_X1    g20656(.A1(new_n20902_), .A2(new_n20913_), .ZN(new_n20914_));
  NOR2_X1    g20657(.A1(new_n20912_), .A2(new_n20914_), .ZN(new_n20915_));
  OAI22_X1   g20658(.A1(new_n9595_), .A2(new_n7354_), .B1(new_n8956_), .B2(new_n7611_), .ZN(new_n20916_));
  XOR2_X1    g20659(.A1(new_n20915_), .A2(new_n20916_), .Z(new_n20917_));
  XOR2_X1    g20660(.A1(new_n20917_), .A2(\a[59] ), .Z(new_n20918_));
  XOR2_X1    g20661(.A1(new_n20918_), .A2(new_n20901_), .Z(new_n20919_));
  NOR2_X1    g20662(.A1(new_n20919_), .A2(new_n20895_), .ZN(new_n20920_));
  NAND2_X1   g20663(.A1(new_n20919_), .A2(new_n20895_), .ZN(new_n20921_));
  INV_X1     g20664(.I(new_n20921_), .ZN(new_n20922_));
  NOR2_X1    g20665(.A1(new_n20922_), .A2(new_n20920_), .ZN(new_n20923_));
  XOR2_X1    g20666(.A1(new_n20894_), .A2(new_n20923_), .Z(\f[122] ));
  NAND2_X1   g20667(.A1(new_n20915_), .A2(new_n20900_), .ZN(new_n20925_));
  XOR2_X1    g20668(.A1(new_n20916_), .A2(\a[59] ), .Z(new_n20926_));
  NAND2_X1   g20669(.A1(new_n20925_), .A2(new_n20926_), .ZN(new_n20927_));
  OAI21_X1   g20670(.A1(new_n20900_), .A2(new_n20915_), .B(new_n20927_), .ZN(new_n20928_));
  NOR2_X1    g20671(.A1(new_n20903_), .A2(new_n20908_), .ZN(new_n20929_));
  NOR2_X1    g20672(.A1(new_n20929_), .A2(new_n20910_), .ZN(new_n20930_));
  INV_X1     g20673(.I(new_n20930_), .ZN(new_n20931_));
  OAI22_X1   g20674(.A1(new_n8956_), .A2(new_n8312_), .B1(new_n8317_), .B2(new_n8932_), .ZN(new_n20932_));
  NAND2_X1   g20675(.A1(new_n9644_), .A2(\b[61] ), .ZN(new_n20933_));
  AOI21_X1   g20676(.A1(new_n20933_), .A2(new_n20932_), .B(new_n8321_), .ZN(new_n20934_));
  NAND2_X1   g20677(.A1(new_n8963_), .A2(new_n20934_), .ZN(new_n20935_));
  XOR2_X1    g20678(.A1(new_n20935_), .A2(\a[62] ), .Z(new_n20936_));
  NOR2_X1    g20679(.A1(new_n8985_), .A2(new_n7930_), .ZN(new_n20937_));
  NOR2_X1    g20680(.A1(new_n9364_), .A2(new_n7890_), .ZN(new_n20938_));
  XNOR2_X1   g20681(.A1(new_n20937_), .A2(new_n20938_), .ZN(new_n20939_));
  XOR2_X1    g20682(.A1(new_n20939_), .A2(\a[59] ), .Z(new_n20940_));
  NOR2_X1    g20683(.A1(new_n20940_), .A2(new_n20907_), .ZN(new_n20941_));
  NOR2_X1    g20684(.A1(new_n20939_), .A2(new_n7343_), .ZN(new_n20942_));
  INV_X1     g20685(.I(new_n20942_), .ZN(new_n20943_));
  NAND2_X1   g20686(.A1(new_n20939_), .A2(new_n7343_), .ZN(new_n20944_));
  AOI21_X1   g20687(.A1(new_n20943_), .A2(new_n20944_), .B(new_n20909_), .ZN(new_n20945_));
  NOR2_X1    g20688(.A1(new_n20941_), .A2(new_n20945_), .ZN(new_n20946_));
  INV_X1     g20689(.I(new_n20946_), .ZN(new_n20947_));
  XOR2_X1    g20690(.A1(new_n20936_), .A2(new_n20947_), .Z(new_n20948_));
  AND2_X2    g20691(.A1(new_n20936_), .A2(new_n20947_), .Z(new_n20949_));
  INV_X1     g20692(.I(new_n20949_), .ZN(new_n20950_));
  NOR2_X1    g20693(.A1(new_n20936_), .A2(new_n20947_), .ZN(new_n20951_));
  INV_X1     g20694(.I(new_n20951_), .ZN(new_n20952_));
  AOI21_X1   g20695(.A1(new_n20950_), .A2(new_n20952_), .B(new_n20931_), .ZN(new_n20953_));
  AOI21_X1   g20696(.A1(new_n20931_), .A2(new_n20948_), .B(new_n20953_), .ZN(new_n20954_));
  XOR2_X1    g20697(.A1(new_n20954_), .A2(new_n20928_), .Z(new_n20955_));
  INV_X1     g20698(.I(new_n20955_), .ZN(new_n20956_));
  AOI21_X1   g20699(.A1(new_n20894_), .A2(new_n20923_), .B(new_n20922_), .ZN(new_n20957_));
  XOR2_X1    g20700(.A1(new_n20957_), .A2(new_n20956_), .Z(\f[123] ));
  AOI21_X1   g20701(.A1(new_n20931_), .A2(new_n20950_), .B(new_n20951_), .ZN(new_n20959_));
  INV_X1     g20702(.I(new_n20959_), .ZN(new_n20960_));
  NOR2_X1    g20703(.A1(new_n8622_), .A2(new_n8932_), .ZN(new_n20961_));
  NOR2_X1    g20704(.A1(new_n8317_), .A2(new_n8956_), .ZN(new_n20962_));
  NOR4_X1    g20705(.A1(new_n9323_), .A2(new_n8321_), .A3(new_n20961_), .A4(new_n20962_), .ZN(new_n20963_));
  XOR2_X1    g20706(.A1(new_n20963_), .A2(\a[62] ), .Z(new_n20964_));
  NAND2_X1   g20707(.A1(new_n20944_), .A2(new_n20909_), .ZN(new_n20965_));
  NAND2_X1   g20708(.A1(new_n20965_), .A2(new_n20943_), .ZN(new_n20966_));
  NAND2_X1   g20709(.A1(new_n9649_), .A2(\b[61] ), .ZN(new_n20967_));
  NOR2_X1    g20710(.A1(new_n9364_), .A2(new_n7930_), .ZN(new_n20968_));
  XOR2_X1    g20711(.A1(new_n20967_), .A2(new_n20968_), .Z(new_n20969_));
  INV_X1     g20712(.I(new_n20969_), .ZN(new_n20970_));
  XOR2_X1    g20713(.A1(new_n20966_), .A2(new_n20970_), .Z(new_n20971_));
  INV_X1     g20714(.I(new_n20971_), .ZN(new_n20972_));
  NOR2_X1    g20715(.A1(new_n20966_), .A2(new_n20969_), .ZN(new_n20973_));
  INV_X1     g20716(.I(new_n20973_), .ZN(new_n20974_));
  NAND2_X1   g20717(.A1(new_n20966_), .A2(new_n20969_), .ZN(new_n20975_));
  AOI21_X1   g20718(.A1(new_n20974_), .A2(new_n20975_), .B(new_n20964_), .ZN(new_n20976_));
  AOI21_X1   g20719(.A1(new_n20964_), .A2(new_n20972_), .B(new_n20976_), .ZN(new_n20977_));
  NOR2_X1    g20720(.A1(new_n20954_), .A2(new_n20928_), .ZN(new_n20978_));
  NOR2_X1    g20721(.A1(new_n20956_), .A2(new_n20978_), .ZN(new_n20979_));
  INV_X1     g20722(.I(new_n20979_), .ZN(new_n20980_));
  OAI21_X1   g20723(.A1(new_n20957_), .A2(new_n20980_), .B(new_n20977_), .ZN(new_n20981_));
  INV_X1     g20724(.I(new_n20891_), .ZN(new_n20982_));
  INV_X1     g20725(.I(new_n20893_), .ZN(new_n20983_));
  OAI21_X1   g20726(.A1(new_n20884_), .A2(new_n20983_), .B(new_n20982_), .ZN(new_n20984_));
  OAI21_X1   g20727(.A1(new_n20984_), .A2(new_n20920_), .B(new_n20921_), .ZN(new_n20985_));
  INV_X1     g20728(.I(new_n20977_), .ZN(new_n20986_));
  NAND3_X1   g20729(.A1(new_n20985_), .A2(new_n20986_), .A3(new_n20979_), .ZN(new_n20987_));
  NAND2_X1   g20730(.A1(new_n20987_), .A2(new_n20981_), .ZN(new_n20988_));
  XOR2_X1    g20731(.A1(new_n20988_), .A2(new_n20960_), .Z(\f[124] ));
  NOR2_X1    g20732(.A1(new_n20957_), .A2(new_n20980_), .ZN(new_n20990_));
  AOI21_X1   g20733(.A1(new_n20985_), .A2(new_n20979_), .B(new_n20986_), .ZN(new_n20991_));
  NOR3_X1    g20734(.A1(new_n20957_), .A2(new_n20977_), .A3(new_n20980_), .ZN(new_n20992_));
  OAI22_X1   g20735(.A1(new_n20991_), .A2(new_n20992_), .B1(new_n20990_), .B2(new_n20959_), .ZN(new_n20993_));
  INV_X1     g20736(.I(new_n20975_), .ZN(new_n20994_));
  AOI21_X1   g20737(.A1(new_n20964_), .A2(new_n20974_), .B(new_n20994_), .ZN(new_n20995_));
  NAND2_X1   g20738(.A1(new_n9649_), .A2(\b[62] ), .ZN(new_n20996_));
  NOR2_X1    g20739(.A1(new_n9364_), .A2(new_n8548_), .ZN(new_n20997_));
  XOR2_X1    g20740(.A1(new_n20996_), .A2(new_n20997_), .Z(new_n20998_));
  OAI22_X1   g20741(.A1(new_n9595_), .A2(new_n8321_), .B1(new_n8956_), .B2(new_n8622_), .ZN(new_n20999_));
  XOR2_X1    g20742(.A1(new_n20999_), .A2(new_n20970_), .Z(new_n21000_));
  XOR2_X1    g20743(.A1(new_n21000_), .A2(new_n8309_), .Z(new_n21001_));
  XNOR2_X1   g20744(.A1(new_n21001_), .A2(new_n20998_), .ZN(new_n21002_));
  XOR2_X1    g20745(.A1(new_n21002_), .A2(new_n20995_), .Z(new_n21003_));
  INV_X1     g20746(.I(new_n20995_), .ZN(new_n21004_));
  NOR2_X1    g20747(.A1(new_n21002_), .A2(new_n21004_), .ZN(new_n21005_));
  INV_X1     g20748(.I(new_n21005_), .ZN(new_n21006_));
  NAND2_X1   g20749(.A1(new_n21002_), .A2(new_n21004_), .ZN(new_n21007_));
  NAND2_X1   g20750(.A1(new_n21006_), .A2(new_n21007_), .ZN(new_n21008_));
  NAND2_X1   g20751(.A1(new_n20993_), .A2(new_n21008_), .ZN(new_n21009_));
  OAI21_X1   g20752(.A1(new_n20993_), .A2(new_n21003_), .B(new_n21009_), .ZN(\f[125] ));
  OAI21_X1   g20753(.A1(new_n20993_), .A2(new_n21005_), .B(new_n21007_), .ZN(new_n21011_));
  XOR2_X1    g20754(.A1(new_n20999_), .A2(new_n8309_), .Z(new_n21012_));
  XOR2_X1    g20755(.A1(new_n21012_), .A2(new_n20970_), .Z(new_n21013_));
  INV_X1     g20756(.I(new_n21013_), .ZN(new_n21014_));
  OAI21_X1   g20757(.A1(new_n20998_), .A2(new_n21012_), .B(new_n21014_), .ZN(new_n21015_));
  NOR3_X1    g20758(.A1(new_n8309_), .A2(new_n9362_), .A3(new_n8932_), .ZN(new_n21016_));
  NOR2_X1    g20759(.A1(new_n9364_), .A2(new_n8932_), .ZN(new_n21017_));
  NOR3_X1    g20760(.A1(new_n21017_), .A2(new_n8956_), .A3(new_n8985_), .ZN(new_n21018_));
  NOR2_X1    g20761(.A1(new_n21018_), .A2(new_n21016_), .ZN(new_n21019_));
  XOR2_X1    g20762(.A1(new_n21019_), .A2(new_n8309_), .Z(new_n21020_));
  OAI21_X1   g20763(.A1(new_n21018_), .A2(new_n21016_), .B(\a[62] ), .ZN(new_n21021_));
  NAND2_X1   g20764(.A1(new_n21019_), .A2(new_n8309_), .ZN(new_n21022_));
  AOI21_X1   g20765(.A1(new_n21021_), .A2(new_n21022_), .B(new_n20970_), .ZN(new_n21023_));
  AOI21_X1   g20766(.A1(new_n20970_), .A2(new_n21020_), .B(new_n21023_), .ZN(new_n21024_));
  XNOR2_X1   g20767(.A1(new_n21015_), .A2(new_n21024_), .ZN(new_n21025_));
  NAND2_X1   g20768(.A1(new_n21011_), .A2(new_n21025_), .ZN(new_n21026_));
  XNOR2_X1   g20769(.A1(new_n21015_), .A2(new_n21024_), .ZN(new_n21027_));
  OAI21_X1   g20770(.A1(new_n21011_), .A2(new_n21027_), .B(new_n21026_), .ZN(\f[126] ));
  NOR2_X1    g20771(.A1(new_n9364_), .A2(new_n8956_), .ZN(new_n21029_));
  NOR2_X1    g20772(.A1(new_n20969_), .A2(new_n21019_), .ZN(new_n21030_));
  XOR2_X1    g20773(.A1(new_n21030_), .A2(new_n21029_), .Z(new_n21031_));
  XOR2_X1    g20774(.A1(new_n20969_), .A2(new_n21019_), .Z(new_n21032_));
  NAND2_X1   g20775(.A1(new_n21032_), .A2(\a[62] ), .ZN(new_n21033_));
  XOR2_X1    g20776(.A1(new_n21031_), .A2(new_n21033_), .Z(new_n21034_));
  AOI21_X1   g20777(.A1(new_n20987_), .A2(new_n20981_), .B(new_n20960_), .ZN(new_n21035_));
  NOR3_X1    g20778(.A1(new_n20957_), .A2(new_n20977_), .A3(new_n20980_), .ZN(new_n21036_));
  OAI21_X1   g20779(.A1(new_n21035_), .A2(new_n21036_), .B(new_n21006_), .ZN(new_n21037_));
  INV_X1     g20780(.I(new_n21015_), .ZN(new_n21038_));
  NAND3_X1   g20781(.A1(new_n21037_), .A2(new_n21007_), .A3(new_n21038_), .ZN(new_n21039_));
  NAND2_X1   g20782(.A1(new_n21011_), .A2(new_n21015_), .ZN(new_n21040_));
  NAND2_X1   g20783(.A1(new_n21040_), .A2(new_n21039_), .ZN(new_n21041_));
  NAND3_X1   g20784(.A1(new_n21041_), .A2(new_n21024_), .A3(new_n21034_), .ZN(new_n21042_));
  INV_X1     g20785(.I(new_n21034_), .ZN(new_n21043_));
  NOR2_X1    g20786(.A1(new_n21011_), .A2(new_n21015_), .ZN(new_n21044_));
  AOI21_X1   g20787(.A1(new_n21037_), .A2(new_n21007_), .B(new_n21038_), .ZN(new_n21045_));
  OAI21_X1   g20788(.A1(new_n21044_), .A2(new_n21045_), .B(new_n21024_), .ZN(new_n21046_));
  NAND2_X1   g20789(.A1(new_n21046_), .A2(new_n21043_), .ZN(new_n21047_));
  NAND2_X1   g20790(.A1(new_n21011_), .A2(new_n21038_), .ZN(new_n21048_));
  INV_X1     g20791(.I(new_n21048_), .ZN(new_n21049_));
  NAND3_X1   g20792(.A1(new_n21047_), .A2(new_n21042_), .A3(new_n21049_), .ZN(new_n21050_));
  NOR2_X1    g20793(.A1(new_n21046_), .A2(new_n21043_), .ZN(new_n21051_));
  AOI21_X1   g20794(.A1(new_n21041_), .A2(new_n21024_), .B(new_n21034_), .ZN(new_n21052_));
  OAI21_X1   g20795(.A1(new_n21051_), .A2(new_n21052_), .B(new_n21048_), .ZN(new_n21053_));
  NAND2_X1   g20796(.A1(new_n21053_), .A2(new_n21050_), .ZN(\f[127] ));
endmodule


