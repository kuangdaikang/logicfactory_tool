// Benchmark "max" written by ABC on Fri Sep 15 11:23:28 2023

module max ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_,
    new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_,
    new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_,
    new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_,
    new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_,
    new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_,
    new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3413_, new_n3415_, new_n3417_, new_n3419_,
    new_n3421_, new_n3423_, new_n3425_, new_n3427_, new_n3429_, new_n3431_,
    new_n3433_, new_n3435_, new_n3437_, new_n3439_, new_n3441_, new_n3443_,
    new_n3445_, new_n3447_, new_n3449_, new_n3451_, new_n3453_, new_n3455_,
    new_n3457_, new_n3459_, new_n3461_, new_n3463_, new_n3465_, new_n3467_,
    new_n3469_, new_n3471_, new_n3473_, new_n3475_, new_n3476_, new_n3478_,
    new_n3479_, new_n3481_, new_n3483_, new_n3484_, new_n3486_, new_n3487_,
    new_n3489_, new_n3490_, new_n3492_, new_n3494_, new_n3496_, new_n3498_,
    new_n3499_, new_n3501_, new_n3503_, new_n3505_, new_n3507_, new_n3508_,
    new_n3510_, new_n3512_, new_n3513_, new_n3515_, new_n3516_, new_n3518_,
    new_n3519_, new_n3521_, new_n3523_, new_n3525_, new_n3526_, new_n3528_,
    new_n3529_, new_n3531_, new_n3533_, new_n3535_, new_n3537_, new_n3538_,
    new_n3540_, new_n3542_, new_n3544_, new_n3546_, new_n3547_, new_n3549_,
    new_n3551_, new_n3552_, new_n3554_, new_n3555_, new_n3557_, new_n3558_,
    new_n3560_, new_n3562_, new_n3564_, new_n3566_, new_n3568_, new_n3570_,
    new_n3572_, new_n3573_, new_n3575_, new_n3576_, new_n3578_, new_n3580_,
    new_n3582_, new_n3584_, new_n3586_, new_n3588_, new_n3590_, new_n3591_,
    new_n3593_, new_n3594_, new_n3596_, new_n3598_, new_n3600_, new_n3601_,
    new_n3603_, new_n3604_, new_n3606_, new_n3608_, new_n3610_, new_n3611_,
    new_n3613_, new_n3614_, new_n3616_, new_n3618_, new_n3620_, new_n3622_,
    new_n3624_, new_n3626_, new_n3628_, new_n3629_, new_n3631_, new_n3632_,
    new_n3634_, new_n3636_, new_n3638_, new_n3640_, new_n3642_, new_n3644_,
    new_n3646_, new_n3647_, new_n3649_, new_n3650_, new_n3652_, new_n3654_,
    new_n3656_, new_n3657_, new_n3659_, new_n3660_, new_n3662_, new_n3664_,
    new_n3666_, new_n3667_, new_n3669_, new_n3670_, new_n3672_, new_n3674_,
    new_n3676_, new_n3678_, new_n3680_, new_n3682_, new_n3684_, new_n3685_,
    new_n3687_, new_n3688_, new_n3690_, new_n3692_, new_n3694_, new_n3696_,
    new_n3698_, new_n3702_;
  INV_X1     g0000(.I(\in1[0] ), .ZN(new_n643_));
  INV_X1     g0001(.I(\in0[127] ), .ZN(new_n644_));
  NOR2_X1    g0002(.A1(new_n644_), .A2(\in1[127] ), .ZN(new_n645_));
  INV_X1     g0003(.I(\in0[125] ), .ZN(new_n646_));
  INV_X1     g0004(.I(\in0[126] ), .ZN(new_n647_));
  AOI22_X1   g0005(.A1(new_n646_), .A2(\in1[125] ), .B1(new_n647_), .B2(\in1[126] ), .ZN(new_n648_));
  INV_X1     g0006(.I(\in1[124] ), .ZN(new_n649_));
  INV_X1     g0007(.I(\in1[125] ), .ZN(new_n650_));
  AOI22_X1   g0008(.A1(\in0[124] ), .A2(new_n649_), .B1(new_n650_), .B2(\in0[125] ), .ZN(new_n651_));
  INV_X1     g0009(.I(new_n651_), .ZN(new_n652_));
  NAND2_X1   g0010(.A1(new_n652_), .A2(new_n648_), .ZN(new_n653_));
  INV_X1     g0011(.I(\in1[126] ), .ZN(new_n654_));
  NAND2_X1   g0012(.A1(new_n654_), .A2(\in0[126] ), .ZN(new_n655_));
  AOI21_X1   g0013(.A1(new_n653_), .A2(new_n655_), .B(new_n645_), .ZN(new_n656_));
  INV_X1     g0014(.I(new_n656_), .ZN(new_n657_));
  INV_X1     g0015(.I(new_n648_), .ZN(new_n658_));
  NOR2_X1    g0016(.A1(new_n649_), .A2(\in0[124] ), .ZN(new_n659_));
  NOR3_X1    g0017(.A1(new_n658_), .A2(new_n645_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1     g0018(.I(new_n660_), .ZN(new_n661_));
  INV_X1     g0019(.I(\in1[121] ), .ZN(new_n662_));
  NOR2_X1    g0020(.A1(new_n662_), .A2(\in0[121] ), .ZN(new_n663_));
  INV_X1     g0021(.I(\in0[122] ), .ZN(new_n664_));
  INV_X1     g0022(.I(\in0[123] ), .ZN(new_n665_));
  AOI22_X1   g0023(.A1(new_n664_), .A2(\in1[122] ), .B1(new_n665_), .B2(\in1[123] ), .ZN(new_n666_));
  INV_X1     g0024(.I(new_n666_), .ZN(new_n667_));
  INV_X1     g0025(.I(\in1[120] ), .ZN(new_n668_));
  NOR2_X1    g0026(.A1(new_n668_), .A2(\in0[120] ), .ZN(new_n669_));
  NOR3_X1    g0027(.A1(new_n667_), .A2(new_n663_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1     g0028(.I(\in1[119] ), .ZN(new_n671_));
  NOR2_X1    g0029(.A1(new_n671_), .A2(\in0[119] ), .ZN(new_n672_));
  INV_X1     g0030(.I(\in0[118] ), .ZN(new_n673_));
  AOI21_X1   g0031(.A1(new_n673_), .A2(\in1[118] ), .B(new_n672_), .ZN(new_n674_));
  INV_X1     g0032(.I(new_n674_), .ZN(new_n675_));
  INV_X1     g0033(.I(\in1[117] ), .ZN(new_n676_));
  NOR2_X1    g0034(.A1(new_n676_), .A2(\in0[117] ), .ZN(new_n677_));
  INV_X1     g0035(.I(\in1[116] ), .ZN(new_n678_));
  AOI22_X1   g0036(.A1(\in0[116] ), .A2(new_n678_), .B1(new_n676_), .B2(\in0[117] ), .ZN(new_n679_));
  NOR2_X1    g0037(.A1(new_n679_), .A2(new_n677_), .ZN(new_n680_));
  INV_X1     g0038(.I(new_n680_), .ZN(new_n681_));
  INV_X1     g0039(.I(\in1[118] ), .ZN(new_n682_));
  AOI22_X1   g0040(.A1(\in0[118] ), .A2(new_n682_), .B1(new_n671_), .B2(\in0[119] ), .ZN(new_n683_));
  OAI22_X1   g0041(.A1(new_n681_), .A2(new_n675_), .B1(new_n672_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1     g0042(.I(new_n684_), .ZN(new_n685_));
  INV_X1     g0043(.I(\in1[115] ), .ZN(new_n686_));
  INV_X1     g0044(.I(\in0[114] ), .ZN(new_n687_));
  INV_X1     g0045(.I(\in0[115] ), .ZN(new_n688_));
  AOI22_X1   g0046(.A1(new_n687_), .A2(\in1[114] ), .B1(new_n688_), .B2(\in1[115] ), .ZN(new_n689_));
  INV_X1     g0047(.I(\in1[113] ), .ZN(new_n690_));
  INV_X1     g0048(.I(\in1[114] ), .ZN(new_n691_));
  AOI22_X1   g0049(.A1(\in0[113] ), .A2(new_n690_), .B1(new_n691_), .B2(\in0[114] ), .ZN(new_n692_));
  NOR2_X1    g0050(.A1(new_n690_), .A2(\in0[113] ), .ZN(new_n693_));
  INV_X1     g0051(.I(\in1[112] ), .ZN(new_n694_));
  NAND2_X1   g0052(.A1(new_n694_), .A2(\in0[112] ), .ZN(new_n695_));
  OAI21_X1   g0053(.A1(new_n693_), .A2(new_n695_), .B(new_n692_), .ZN(new_n696_));
  AOI22_X1   g0054(.A1(new_n696_), .A2(new_n689_), .B1(\in0[115] ), .B2(new_n686_), .ZN(new_n697_));
  INV_X1     g0055(.I(new_n697_), .ZN(new_n698_));
  INV_X1     g0056(.I(new_n689_), .ZN(new_n699_));
  NOR2_X1    g0057(.A1(new_n694_), .A2(\in0[112] ), .ZN(new_n700_));
  NOR3_X1    g0058(.A1(new_n699_), .A2(new_n693_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1     g0059(.I(\in0[110] ), .ZN(new_n702_));
  INV_X1     g0060(.I(\in1[111] ), .ZN(new_n703_));
  NOR2_X1    g0061(.A1(new_n703_), .A2(\in0[111] ), .ZN(new_n704_));
  AOI21_X1   g0062(.A1(new_n702_), .A2(\in1[110] ), .B(new_n704_), .ZN(new_n705_));
  INV_X1     g0063(.I(new_n705_), .ZN(new_n706_));
  INV_X1     g0064(.I(\in1[108] ), .ZN(new_n707_));
  NOR2_X1    g0065(.A1(new_n707_), .A2(\in0[108] ), .ZN(new_n708_));
  INV_X1     g0066(.I(\in1[109] ), .ZN(new_n709_));
  NOR2_X1    g0067(.A1(new_n709_), .A2(\in0[109] ), .ZN(new_n710_));
  NOR3_X1    g0068(.A1(new_n706_), .A2(new_n708_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1     g0069(.I(new_n711_), .ZN(new_n712_));
  INV_X1     g0070(.I(\in1[107] ), .ZN(new_n713_));
  INV_X1     g0071(.I(\in0[106] ), .ZN(new_n714_));
  INV_X1     g0072(.I(\in0[107] ), .ZN(new_n715_));
  AOI22_X1   g0073(.A1(new_n714_), .A2(\in1[106] ), .B1(new_n715_), .B2(\in1[107] ), .ZN(new_n716_));
  INV_X1     g0074(.I(\in1[105] ), .ZN(new_n717_));
  INV_X1     g0075(.I(\in1[106] ), .ZN(new_n718_));
  AOI22_X1   g0076(.A1(\in0[105] ), .A2(new_n717_), .B1(new_n718_), .B2(\in0[106] ), .ZN(new_n719_));
  NOR2_X1    g0077(.A1(new_n717_), .A2(\in0[105] ), .ZN(new_n720_));
  INV_X1     g0078(.I(\in1[104] ), .ZN(new_n721_));
  NAND2_X1   g0079(.A1(new_n721_), .A2(\in0[104] ), .ZN(new_n722_));
  OAI21_X1   g0080(.A1(new_n720_), .A2(new_n722_), .B(new_n719_), .ZN(new_n723_));
  AOI22_X1   g0081(.A1(new_n723_), .A2(new_n716_), .B1(\in0[107] ), .B2(new_n713_), .ZN(new_n724_));
  INV_X1     g0082(.I(new_n724_), .ZN(new_n725_));
  INV_X1     g0083(.I(\in1[103] ), .ZN(new_n726_));
  NOR2_X1    g0084(.A1(new_n726_), .A2(\in0[103] ), .ZN(new_n727_));
  INV_X1     g0085(.I(\in0[102] ), .ZN(new_n728_));
  AOI21_X1   g0086(.A1(new_n728_), .A2(\in1[102] ), .B(new_n727_), .ZN(new_n729_));
  INV_X1     g0087(.I(new_n729_), .ZN(new_n730_));
  INV_X1     g0088(.I(\in1[101] ), .ZN(new_n731_));
  NOR2_X1    g0089(.A1(new_n731_), .A2(\in0[101] ), .ZN(new_n732_));
  INV_X1     g0090(.I(\in1[100] ), .ZN(new_n733_));
  AOI22_X1   g0091(.A1(\in0[100] ), .A2(new_n733_), .B1(new_n731_), .B2(\in0[101] ), .ZN(new_n734_));
  NOR2_X1    g0092(.A1(new_n734_), .A2(new_n732_), .ZN(new_n735_));
  INV_X1     g0093(.I(new_n735_), .ZN(new_n736_));
  INV_X1     g0094(.I(\in1[102] ), .ZN(new_n737_));
  AOI22_X1   g0095(.A1(\in0[102] ), .A2(new_n737_), .B1(new_n726_), .B2(\in0[103] ), .ZN(new_n738_));
  OAI22_X1   g0096(.A1(new_n736_), .A2(new_n730_), .B1(new_n727_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1     g0097(.I(new_n739_), .ZN(new_n740_));
  NOR2_X1    g0098(.A1(new_n733_), .A2(\in0[100] ), .ZN(new_n741_));
  NOR3_X1    g0099(.A1(new_n730_), .A2(new_n732_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1     g0100(.I(new_n742_), .ZN(new_n743_));
  INV_X1     g0101(.I(\in1[97] ), .ZN(new_n744_));
  NOR2_X1    g0102(.A1(new_n744_), .A2(\in0[97] ), .ZN(new_n745_));
  INV_X1     g0103(.I(\in0[98] ), .ZN(new_n746_));
  INV_X1     g0104(.I(\in0[99] ), .ZN(new_n747_));
  AOI22_X1   g0105(.A1(new_n746_), .A2(\in1[98] ), .B1(new_n747_), .B2(\in1[99] ), .ZN(new_n748_));
  INV_X1     g0106(.I(new_n748_), .ZN(new_n749_));
  INV_X1     g0107(.I(\in1[96] ), .ZN(new_n750_));
  NOR2_X1    g0108(.A1(new_n750_), .A2(\in0[96] ), .ZN(new_n751_));
  NOR3_X1    g0109(.A1(new_n749_), .A2(new_n745_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1     g0110(.I(\in1[95] ), .ZN(new_n753_));
  NOR2_X1    g0111(.A1(new_n753_), .A2(\in0[95] ), .ZN(new_n754_));
  INV_X1     g0112(.I(\in0[94] ), .ZN(new_n755_));
  AOI21_X1   g0113(.A1(new_n755_), .A2(\in1[94] ), .B(new_n754_), .ZN(new_n756_));
  INV_X1     g0114(.I(new_n756_), .ZN(new_n757_));
  INV_X1     g0115(.I(\in1[93] ), .ZN(new_n758_));
  NOR2_X1    g0116(.A1(new_n758_), .A2(\in0[93] ), .ZN(new_n759_));
  INV_X1     g0117(.I(\in1[92] ), .ZN(new_n760_));
  AOI22_X1   g0118(.A1(\in0[92] ), .A2(new_n760_), .B1(new_n758_), .B2(\in0[93] ), .ZN(new_n761_));
  NOR2_X1    g0119(.A1(new_n761_), .A2(new_n759_), .ZN(new_n762_));
  INV_X1     g0120(.I(new_n762_), .ZN(new_n763_));
  INV_X1     g0121(.I(\in1[94] ), .ZN(new_n764_));
  AOI22_X1   g0122(.A1(\in0[94] ), .A2(new_n764_), .B1(new_n753_), .B2(\in0[95] ), .ZN(new_n765_));
  OAI22_X1   g0123(.A1(new_n763_), .A2(new_n757_), .B1(new_n754_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1     g0124(.I(new_n766_), .ZN(new_n767_));
  INV_X1     g0125(.I(\in1[91] ), .ZN(new_n768_));
  INV_X1     g0126(.I(\in0[90] ), .ZN(new_n769_));
  INV_X1     g0127(.I(\in0[91] ), .ZN(new_n770_));
  AOI22_X1   g0128(.A1(new_n769_), .A2(\in1[90] ), .B1(new_n770_), .B2(\in1[91] ), .ZN(new_n771_));
  INV_X1     g0129(.I(\in1[89] ), .ZN(new_n772_));
  INV_X1     g0130(.I(\in1[90] ), .ZN(new_n773_));
  AOI22_X1   g0131(.A1(\in0[89] ), .A2(new_n772_), .B1(new_n773_), .B2(\in0[90] ), .ZN(new_n774_));
  NOR2_X1    g0132(.A1(new_n772_), .A2(\in0[89] ), .ZN(new_n775_));
  INV_X1     g0133(.I(\in1[88] ), .ZN(new_n776_));
  NAND2_X1   g0134(.A1(new_n776_), .A2(\in0[88] ), .ZN(new_n777_));
  OAI21_X1   g0135(.A1(new_n775_), .A2(new_n777_), .B(new_n774_), .ZN(new_n778_));
  AOI22_X1   g0136(.A1(new_n778_), .A2(new_n771_), .B1(\in0[91] ), .B2(new_n768_), .ZN(new_n779_));
  INV_X1     g0137(.I(new_n779_), .ZN(new_n780_));
  INV_X1     g0138(.I(new_n771_), .ZN(new_n781_));
  NOR2_X1    g0139(.A1(new_n776_), .A2(\in0[88] ), .ZN(new_n782_));
  NOR3_X1    g0140(.A1(new_n781_), .A2(new_n775_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1     g0141(.I(\in0[86] ), .ZN(new_n784_));
  INV_X1     g0142(.I(\in1[87] ), .ZN(new_n785_));
  NOR2_X1    g0143(.A1(new_n785_), .A2(\in0[87] ), .ZN(new_n786_));
  AOI21_X1   g0144(.A1(new_n784_), .A2(\in1[86] ), .B(new_n786_), .ZN(new_n787_));
  INV_X1     g0145(.I(new_n787_), .ZN(new_n788_));
  INV_X1     g0146(.I(\in1[84] ), .ZN(new_n789_));
  NOR2_X1    g0147(.A1(new_n789_), .A2(\in0[84] ), .ZN(new_n790_));
  INV_X1     g0148(.I(\in1[85] ), .ZN(new_n791_));
  NOR2_X1    g0149(.A1(new_n791_), .A2(\in0[85] ), .ZN(new_n792_));
  NOR3_X1    g0150(.A1(new_n788_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1     g0151(.I(new_n793_), .ZN(new_n794_));
  INV_X1     g0152(.I(\in1[83] ), .ZN(new_n795_));
  INV_X1     g0153(.I(\in0[82] ), .ZN(new_n796_));
  INV_X1     g0154(.I(\in0[83] ), .ZN(new_n797_));
  AOI22_X1   g0155(.A1(new_n796_), .A2(\in1[82] ), .B1(new_n797_), .B2(\in1[83] ), .ZN(new_n798_));
  INV_X1     g0156(.I(\in1[81] ), .ZN(new_n799_));
  INV_X1     g0157(.I(\in1[82] ), .ZN(new_n800_));
  AOI22_X1   g0158(.A1(\in0[81] ), .A2(new_n799_), .B1(new_n800_), .B2(\in0[82] ), .ZN(new_n801_));
  NOR2_X1    g0159(.A1(new_n799_), .A2(\in0[81] ), .ZN(new_n802_));
  INV_X1     g0160(.I(\in1[80] ), .ZN(new_n803_));
  NAND2_X1   g0161(.A1(new_n803_), .A2(\in0[80] ), .ZN(new_n804_));
  OAI21_X1   g0162(.A1(new_n802_), .A2(new_n804_), .B(new_n801_), .ZN(new_n805_));
  AOI22_X1   g0163(.A1(new_n805_), .A2(new_n798_), .B1(\in0[83] ), .B2(new_n795_), .ZN(new_n806_));
  INV_X1     g0164(.I(new_n806_), .ZN(new_n807_));
  INV_X1     g0165(.I(\in1[79] ), .ZN(new_n808_));
  NOR2_X1    g0166(.A1(new_n808_), .A2(\in0[79] ), .ZN(new_n809_));
  INV_X1     g0167(.I(\in0[78] ), .ZN(new_n810_));
  AOI21_X1   g0168(.A1(new_n810_), .A2(\in1[78] ), .B(new_n809_), .ZN(new_n811_));
  INV_X1     g0169(.I(new_n811_), .ZN(new_n812_));
  INV_X1     g0170(.I(\in1[77] ), .ZN(new_n813_));
  NOR2_X1    g0171(.A1(new_n813_), .A2(\in0[77] ), .ZN(new_n814_));
  INV_X1     g0172(.I(\in1[76] ), .ZN(new_n815_));
  AOI22_X1   g0173(.A1(\in0[76] ), .A2(new_n815_), .B1(new_n813_), .B2(\in0[77] ), .ZN(new_n816_));
  NOR2_X1    g0174(.A1(new_n816_), .A2(new_n814_), .ZN(new_n817_));
  INV_X1     g0175(.I(new_n817_), .ZN(new_n818_));
  INV_X1     g0176(.I(\in1[78] ), .ZN(new_n819_));
  AOI22_X1   g0177(.A1(\in0[78] ), .A2(new_n819_), .B1(new_n808_), .B2(\in0[79] ), .ZN(new_n820_));
  OAI22_X1   g0178(.A1(new_n818_), .A2(new_n812_), .B1(new_n809_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1     g0179(.I(new_n821_), .ZN(new_n822_));
  NOR2_X1    g0180(.A1(new_n815_), .A2(\in0[76] ), .ZN(new_n823_));
  NOR3_X1    g0181(.A1(new_n812_), .A2(new_n814_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1     g0182(.I(new_n824_), .ZN(new_n825_));
  INV_X1     g0183(.I(\in1[73] ), .ZN(new_n826_));
  NOR2_X1    g0184(.A1(new_n826_), .A2(\in0[73] ), .ZN(new_n827_));
  INV_X1     g0185(.I(\in0[74] ), .ZN(new_n828_));
  INV_X1     g0186(.I(\in0[75] ), .ZN(new_n829_));
  AOI22_X1   g0187(.A1(new_n828_), .A2(\in1[74] ), .B1(new_n829_), .B2(\in1[75] ), .ZN(new_n830_));
  INV_X1     g0188(.I(new_n830_), .ZN(new_n831_));
  INV_X1     g0189(.I(\in1[72] ), .ZN(new_n832_));
  NOR2_X1    g0190(.A1(new_n832_), .A2(\in0[72] ), .ZN(new_n833_));
  NOR3_X1    g0191(.A1(new_n831_), .A2(new_n827_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1     g0192(.I(\in1[71] ), .ZN(new_n835_));
  NOR2_X1    g0193(.A1(new_n835_), .A2(\in0[71] ), .ZN(new_n836_));
  INV_X1     g0194(.I(\in0[70] ), .ZN(new_n837_));
  AOI21_X1   g0195(.A1(new_n837_), .A2(\in1[70] ), .B(new_n836_), .ZN(new_n838_));
  INV_X1     g0196(.I(new_n838_), .ZN(new_n839_));
  INV_X1     g0197(.I(\in1[69] ), .ZN(new_n840_));
  NOR2_X1    g0198(.A1(new_n840_), .A2(\in0[69] ), .ZN(new_n841_));
  INV_X1     g0199(.I(\in1[68] ), .ZN(new_n842_));
  AOI22_X1   g0200(.A1(\in0[68] ), .A2(new_n842_), .B1(new_n840_), .B2(\in0[69] ), .ZN(new_n843_));
  NOR2_X1    g0201(.A1(new_n843_), .A2(new_n841_), .ZN(new_n844_));
  INV_X1     g0202(.I(new_n844_), .ZN(new_n845_));
  INV_X1     g0203(.I(\in1[70] ), .ZN(new_n846_));
  AOI22_X1   g0204(.A1(\in0[70] ), .A2(new_n846_), .B1(new_n835_), .B2(\in0[71] ), .ZN(new_n847_));
  OAI22_X1   g0205(.A1(new_n845_), .A2(new_n839_), .B1(new_n836_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1     g0206(.I(new_n848_), .ZN(new_n849_));
  INV_X1     g0207(.I(\in1[67] ), .ZN(new_n850_));
  INV_X1     g0208(.I(\in0[66] ), .ZN(new_n851_));
  INV_X1     g0209(.I(\in0[67] ), .ZN(new_n852_));
  AOI22_X1   g0210(.A1(new_n851_), .A2(\in1[66] ), .B1(new_n852_), .B2(\in1[67] ), .ZN(new_n853_));
  INV_X1     g0211(.I(\in1[65] ), .ZN(new_n854_));
  INV_X1     g0212(.I(\in1[66] ), .ZN(new_n855_));
  AOI22_X1   g0213(.A1(\in0[65] ), .A2(new_n854_), .B1(new_n855_), .B2(\in0[66] ), .ZN(new_n856_));
  NOR2_X1    g0214(.A1(new_n854_), .A2(\in0[65] ), .ZN(new_n857_));
  INV_X1     g0215(.I(\in1[64] ), .ZN(new_n858_));
  NAND2_X1   g0216(.A1(new_n858_), .A2(\in0[64] ), .ZN(new_n859_));
  OAI21_X1   g0217(.A1(new_n857_), .A2(new_n859_), .B(new_n856_), .ZN(new_n860_));
  AOI22_X1   g0218(.A1(new_n860_), .A2(new_n853_), .B1(\in0[67] ), .B2(new_n850_), .ZN(new_n861_));
  INV_X1     g0219(.I(new_n861_), .ZN(new_n862_));
  INV_X1     g0220(.I(new_n853_), .ZN(new_n863_));
  NOR2_X1    g0221(.A1(new_n858_), .A2(\in0[64] ), .ZN(new_n864_));
  NOR3_X1    g0222(.A1(new_n863_), .A2(new_n857_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1     g0223(.I(\in0[56] ), .ZN(new_n866_));
  INV_X1     g0224(.I(\in0[57] ), .ZN(new_n867_));
  AOI22_X1   g0225(.A1(new_n866_), .A2(\in1[56] ), .B1(new_n867_), .B2(\in1[57] ), .ZN(new_n868_));
  INV_X1     g0226(.I(\in0[62] ), .ZN(new_n869_));
  INV_X1     g0227(.I(\in1[63] ), .ZN(new_n870_));
  NOR2_X1    g0228(.A1(new_n870_), .A2(\in0[63] ), .ZN(new_n871_));
  AOI21_X1   g0229(.A1(new_n869_), .A2(\in1[62] ), .B(new_n871_), .ZN(new_n872_));
  INV_X1     g0230(.I(\in0[60] ), .ZN(new_n873_));
  INV_X1     g0231(.I(\in0[61] ), .ZN(new_n874_));
  AOI22_X1   g0232(.A1(new_n873_), .A2(\in1[60] ), .B1(new_n874_), .B2(\in1[61] ), .ZN(new_n875_));
  NAND2_X1   g0233(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1     g0234(.I(new_n876_), .ZN(new_n877_));
  INV_X1     g0235(.I(\in0[58] ), .ZN(new_n878_));
  INV_X1     g0236(.I(\in0[59] ), .ZN(new_n879_));
  AOI22_X1   g0237(.A1(new_n878_), .A2(\in1[58] ), .B1(new_n879_), .B2(\in1[59] ), .ZN(new_n880_));
  NAND3_X1   g0238(.A1(new_n877_), .A2(new_n868_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1     g0239(.I(\in1[53] ), .ZN(new_n882_));
  NOR2_X1    g0240(.A1(new_n882_), .A2(\in0[53] ), .ZN(new_n883_));
  INV_X1     g0241(.I(\in0[54] ), .ZN(new_n884_));
  INV_X1     g0242(.I(\in0[55] ), .ZN(new_n885_));
  AOI22_X1   g0243(.A1(new_n884_), .A2(\in1[54] ), .B1(new_n885_), .B2(\in1[55] ), .ZN(new_n886_));
  INV_X1     g0244(.I(new_n886_), .ZN(new_n887_));
  INV_X1     g0245(.I(\in1[52] ), .ZN(new_n888_));
  NOR2_X1    g0246(.A1(new_n888_), .A2(\in0[52] ), .ZN(new_n889_));
  NOR3_X1    g0247(.A1(new_n887_), .A2(new_n883_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1     g0248(.I(\in0[50] ), .ZN(new_n891_));
  INV_X1     g0249(.I(\in0[51] ), .ZN(new_n892_));
  AOI22_X1   g0250(.A1(new_n891_), .A2(\in1[50] ), .B1(new_n892_), .B2(\in1[51] ), .ZN(new_n893_));
  INV_X1     g0251(.I(new_n893_), .ZN(new_n894_));
  INV_X1     g0252(.I(\in1[49] ), .ZN(new_n895_));
  INV_X1     g0253(.I(\in1[50] ), .ZN(new_n896_));
  AOI22_X1   g0254(.A1(\in0[49] ), .A2(new_n895_), .B1(new_n896_), .B2(\in0[50] ), .ZN(new_n897_));
  INV_X1     g0255(.I(\in0[48] ), .ZN(new_n898_));
  NOR2_X1    g0256(.A1(new_n895_), .A2(\in0[49] ), .ZN(new_n899_));
  NOR3_X1    g0257(.A1(new_n899_), .A2(new_n898_), .A3(\in1[48] ), .ZN(new_n900_));
  INV_X1     g0258(.I(new_n900_), .ZN(new_n901_));
  AOI21_X1   g0259(.A1(new_n901_), .A2(new_n897_), .B(new_n894_), .ZN(new_n902_));
  NOR2_X1    g0260(.A1(new_n892_), .A2(\in1[51] ), .ZN(new_n903_));
  OAI21_X1   g0261(.A1(new_n902_), .A2(new_n903_), .B(new_n890_), .ZN(new_n904_));
  INV_X1     g0262(.I(new_n904_), .ZN(new_n905_));
  INV_X1     g0263(.I(\in1[54] ), .ZN(new_n906_));
  AOI22_X1   g0264(.A1(\in0[53] ), .A2(new_n882_), .B1(new_n906_), .B2(\in0[54] ), .ZN(new_n907_));
  INV_X1     g0265(.I(new_n907_), .ZN(new_n908_));
  NOR2_X1    g0266(.A1(new_n883_), .A2(\in1[52] ), .ZN(new_n909_));
  AOI21_X1   g0267(.A1(\in0[52] ), .A2(new_n909_), .B(new_n908_), .ZN(new_n910_));
  OAI22_X1   g0268(.A1(new_n910_), .A2(new_n887_), .B1(new_n885_), .B2(\in1[55] ), .ZN(new_n911_));
  NOR2_X1    g0269(.A1(new_n905_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1     g0270(.I(new_n912_), .ZN(new_n913_));
  INV_X1     g0271(.I(\in0[46] ), .ZN(new_n914_));
  INV_X1     g0272(.I(\in1[47] ), .ZN(new_n915_));
  NOR2_X1    g0273(.A1(new_n915_), .A2(\in0[47] ), .ZN(new_n916_));
  AOI21_X1   g0274(.A1(new_n914_), .A2(\in1[46] ), .B(new_n916_), .ZN(new_n917_));
  INV_X1     g0275(.I(\in0[44] ), .ZN(new_n918_));
  INV_X1     g0276(.I(\in0[45] ), .ZN(new_n919_));
  AOI22_X1   g0277(.A1(new_n918_), .A2(\in1[44] ), .B1(new_n919_), .B2(\in1[45] ), .ZN(new_n920_));
  NAND2_X1   g0278(.A1(new_n917_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1     g0279(.I(new_n921_), .ZN(new_n922_));
  INV_X1     g0280(.I(\in0[43] ), .ZN(new_n923_));
  INV_X1     g0281(.I(\in0[42] ), .ZN(new_n924_));
  AOI22_X1   g0282(.A1(new_n924_), .A2(\in1[42] ), .B1(new_n923_), .B2(\in1[43] ), .ZN(new_n925_));
  INV_X1     g0283(.I(new_n925_), .ZN(new_n926_));
  INV_X1     g0284(.I(\in1[40] ), .ZN(new_n927_));
  INV_X1     g0285(.I(\in0[41] ), .ZN(new_n928_));
  OAI22_X1   g0286(.A1(new_n928_), .A2(\in1[41] ), .B1(new_n924_), .B2(\in1[42] ), .ZN(new_n929_));
  INV_X1     g0287(.I(\in0[40] ), .ZN(new_n930_));
  AOI21_X1   g0288(.A1(new_n928_), .A2(\in1[41] ), .B(new_n930_), .ZN(new_n931_));
  AOI21_X1   g0289(.A1(new_n927_), .A2(new_n931_), .B(new_n929_), .ZN(new_n932_));
  OAI22_X1   g0290(.A1(new_n932_), .A2(new_n926_), .B1(new_n923_), .B2(\in1[43] ), .ZN(new_n933_));
  NAND2_X1   g0291(.A1(new_n933_), .A2(new_n922_), .ZN(new_n934_));
  NOR2_X1    g0292(.A1(new_n918_), .A2(\in1[44] ), .ZN(new_n935_));
  NOR2_X1    g0293(.A1(new_n919_), .A2(\in1[45] ), .ZN(new_n936_));
  NOR2_X1    g0294(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1   g0295(.A1(new_n919_), .A2(\in1[45] ), .B(new_n937_), .ZN(new_n938_));
  INV_X1     g0296(.I(\in1[46] ), .ZN(new_n939_));
  AOI22_X1   g0297(.A1(\in0[46] ), .A2(new_n939_), .B1(new_n915_), .B2(\in0[47] ), .ZN(new_n940_));
  NOR2_X1    g0298(.A1(new_n940_), .A2(new_n916_), .ZN(new_n941_));
  AOI21_X1   g0299(.A1(new_n938_), .A2(new_n917_), .B(new_n941_), .ZN(new_n942_));
  AND2_X2    g0300(.A1(new_n934_), .A2(new_n942_), .Z(new_n943_));
  AOI22_X1   g0301(.A1(new_n930_), .A2(\in1[40] ), .B1(new_n928_), .B2(\in1[41] ), .ZN(new_n944_));
  NAND3_X1   g0302(.A1(new_n922_), .A2(new_n925_), .A3(new_n944_), .ZN(new_n945_));
  INV_X1     g0303(.I(\in0[32] ), .ZN(new_n946_));
  INV_X1     g0304(.I(\in0[33] ), .ZN(new_n947_));
  AOI22_X1   g0305(.A1(new_n946_), .A2(\in1[32] ), .B1(new_n947_), .B2(\in1[33] ), .ZN(new_n948_));
  INV_X1     g0306(.I(\in0[38] ), .ZN(new_n949_));
  INV_X1     g0307(.I(\in1[39] ), .ZN(new_n950_));
  NOR2_X1    g0308(.A1(new_n950_), .A2(\in0[39] ), .ZN(new_n951_));
  AOI21_X1   g0309(.A1(new_n949_), .A2(\in1[38] ), .B(new_n951_), .ZN(new_n952_));
  INV_X1     g0310(.I(\in0[36] ), .ZN(new_n953_));
  INV_X1     g0311(.I(\in0[37] ), .ZN(new_n954_));
  AOI22_X1   g0312(.A1(new_n953_), .A2(\in1[36] ), .B1(new_n954_), .B2(\in1[37] ), .ZN(new_n955_));
  NAND2_X1   g0313(.A1(new_n952_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1     g0314(.I(new_n956_), .ZN(new_n957_));
  INV_X1     g0315(.I(\in0[34] ), .ZN(new_n958_));
  INV_X1     g0316(.I(\in0[35] ), .ZN(new_n959_));
  AOI22_X1   g0317(.A1(new_n958_), .A2(\in1[34] ), .B1(new_n959_), .B2(\in1[35] ), .ZN(new_n960_));
  NAND3_X1   g0318(.A1(new_n957_), .A2(new_n948_), .A3(new_n960_), .ZN(new_n961_));
  INV_X1     g0319(.I(new_n961_), .ZN(new_n962_));
  INV_X1     g0320(.I(\in0[29] ), .ZN(new_n963_));
  NOR2_X1    g0321(.A1(new_n963_), .A2(\in1[29] ), .ZN(new_n964_));
  INV_X1     g0322(.I(new_n964_), .ZN(new_n965_));
  INV_X1     g0323(.I(\in1[29] ), .ZN(new_n966_));
  NOR2_X1    g0324(.A1(new_n966_), .A2(\in0[29] ), .ZN(new_n967_));
  INV_X1     g0325(.I(new_n967_), .ZN(new_n968_));
  INV_X1     g0326(.I(\in1[27] ), .ZN(new_n969_));
  INV_X1     g0327(.I(\in0[26] ), .ZN(new_n970_));
  NOR2_X1    g0328(.A1(new_n970_), .A2(\in1[26] ), .ZN(new_n971_));
  INV_X1     g0329(.I(new_n971_), .ZN(new_n972_));
  INV_X1     g0330(.I(\in1[26] ), .ZN(new_n973_));
  NOR2_X1    g0331(.A1(new_n973_), .A2(\in0[26] ), .ZN(new_n974_));
  INV_X1     g0332(.I(\in1[24] ), .ZN(new_n975_));
  NOR2_X1    g0333(.A1(new_n975_), .A2(\in0[24] ), .ZN(new_n976_));
  INV_X1     g0334(.I(\in1[23] ), .ZN(new_n977_));
  NOR2_X1    g0335(.A1(new_n977_), .A2(\in0[23] ), .ZN(new_n978_));
  INV_X1     g0336(.I(new_n978_), .ZN(new_n979_));
  INV_X1     g0337(.I(\in0[22] ), .ZN(new_n980_));
  INV_X1     g0338(.I(\in1[22] ), .ZN(new_n981_));
  INV_X1     g0339(.I(\in0[21] ), .ZN(new_n982_));
  NOR2_X1    g0340(.A1(new_n982_), .A2(\in1[21] ), .ZN(new_n983_));
  INV_X1     g0341(.I(\in1[21] ), .ZN(new_n984_));
  NOR2_X1    g0342(.A1(new_n984_), .A2(\in0[21] ), .ZN(new_n985_));
  INV_X1     g0343(.I(\in0[19] ), .ZN(new_n986_));
  INV_X1     g0344(.I(\in0[18] ), .ZN(new_n987_));
  NOR2_X1    g0345(.A1(new_n987_), .A2(\in1[18] ), .ZN(new_n988_));
  INV_X1     g0346(.I(\in1[18] ), .ZN(new_n989_));
  NOR2_X1    g0347(.A1(new_n989_), .A2(\in0[18] ), .ZN(new_n990_));
  INV_X1     g0348(.I(new_n990_), .ZN(new_n991_));
  INV_X1     g0349(.I(\in1[16] ), .ZN(new_n992_));
  NOR2_X1    g0350(.A1(new_n992_), .A2(\in0[16] ), .ZN(new_n993_));
  INV_X1     g0351(.I(new_n993_), .ZN(new_n994_));
  INV_X1     g0352(.I(\in1[15] ), .ZN(new_n995_));
  NOR2_X1    g0353(.A1(new_n995_), .A2(\in0[15] ), .ZN(new_n996_));
  INV_X1     g0354(.I(\in0[13] ), .ZN(new_n997_));
  NOR2_X1    g0355(.A1(new_n997_), .A2(\in1[13] ), .ZN(new_n998_));
  INV_X1     g0356(.I(new_n998_), .ZN(new_n999_));
  INV_X1     g0357(.I(\in1[13] ), .ZN(new_n1000_));
  NOR2_X1    g0358(.A1(new_n1000_), .A2(\in0[13] ), .ZN(new_n1001_));
  INV_X1     g0359(.I(new_n1001_), .ZN(new_n1002_));
  INV_X1     g0360(.I(\in1[11] ), .ZN(new_n1003_));
  INV_X1     g0361(.I(\in0[10] ), .ZN(new_n1004_));
  NOR2_X1    g0362(.A1(new_n1004_), .A2(\in1[10] ), .ZN(new_n1005_));
  INV_X1     g0363(.I(new_n1005_), .ZN(new_n1006_));
  INV_X1     g0364(.I(\in1[10] ), .ZN(new_n1007_));
  NOR2_X1    g0365(.A1(new_n1007_), .A2(\in0[10] ), .ZN(new_n1008_));
  INV_X1     g0366(.I(\in1[8] ), .ZN(new_n1009_));
  NOR2_X1    g0367(.A1(new_n1009_), .A2(\in0[8] ), .ZN(new_n1010_));
  INV_X1     g0368(.I(\in0[6] ), .ZN(new_n1011_));
  NOR2_X1    g0369(.A1(new_n1011_), .A2(\in1[6] ), .ZN(new_n1012_));
  INV_X1     g0370(.I(new_n1012_), .ZN(new_n1013_));
  INV_X1     g0371(.I(\in1[6] ), .ZN(new_n1014_));
  NOR2_X1    g0372(.A1(new_n1014_), .A2(\in0[6] ), .ZN(new_n1015_));
  INV_X1     g0373(.I(new_n1015_), .ZN(new_n1016_));
  INV_X1     g0374(.I(\in1[4] ), .ZN(new_n1017_));
  NOR2_X1    g0375(.A1(new_n1017_), .A2(\in0[4] ), .ZN(new_n1018_));
  INV_X1     g0376(.I(\in1[3] ), .ZN(new_n1019_));
  NOR2_X1    g0377(.A1(new_n1019_), .A2(\in0[3] ), .ZN(new_n1020_));
  INV_X1     g0378(.I(new_n1020_), .ZN(new_n1021_));
  INV_X1     g0379(.I(\in1[2] ), .ZN(new_n1022_));
  NAND2_X1   g0380(.A1(new_n643_), .A2(\in0[0] ), .ZN(new_n1023_));
  INV_X1     g0381(.I(\in1[1] ), .ZN(new_n1024_));
  NAND2_X1   g0382(.A1(new_n1024_), .A2(\in0[1] ), .ZN(new_n1025_));
  NOR2_X1    g0383(.A1(new_n1024_), .A2(\in0[1] ), .ZN(new_n1026_));
  AOI21_X1   g0384(.A1(new_n1023_), .A2(new_n1025_), .B(new_n1026_), .ZN(new_n1027_));
  OAI21_X1   g0385(.A1(new_n1027_), .A2(new_n1022_), .B(\in0[2] ), .ZN(new_n1028_));
  NAND2_X1   g0386(.A1(new_n1027_), .A2(new_n1022_), .ZN(new_n1029_));
  INV_X1     g0387(.I(\in0[3] ), .ZN(new_n1030_));
  NOR2_X1    g0388(.A1(new_n1030_), .A2(\in1[3] ), .ZN(new_n1031_));
  INV_X1     g0389(.I(new_n1031_), .ZN(new_n1032_));
  NAND3_X1   g0390(.A1(new_n1028_), .A2(new_n1029_), .A3(new_n1032_), .ZN(new_n1033_));
  INV_X1     g0391(.I(\in0[4] ), .ZN(new_n1034_));
  NOR2_X1    g0392(.A1(new_n1034_), .A2(\in1[4] ), .ZN(new_n1035_));
  AOI21_X1   g0393(.A1(new_n1033_), .A2(new_n1021_), .B(new_n1035_), .ZN(new_n1036_));
  INV_X1     g0394(.I(\in1[5] ), .ZN(new_n1037_));
  NOR2_X1    g0395(.A1(new_n1037_), .A2(\in0[5] ), .ZN(new_n1038_));
  NOR3_X1    g0396(.A1(new_n1036_), .A2(new_n1018_), .A3(new_n1038_), .ZN(new_n1039_));
  INV_X1     g0397(.I(\in0[5] ), .ZN(new_n1040_));
  NOR2_X1    g0398(.A1(new_n1040_), .A2(\in1[5] ), .ZN(new_n1041_));
  OAI21_X1   g0399(.A1(new_n1039_), .A2(new_n1041_), .B(new_n1016_), .ZN(new_n1042_));
  AOI21_X1   g0400(.A1(new_n1042_), .A2(new_n1013_), .B(\in1[7] ), .ZN(new_n1043_));
  NAND3_X1   g0401(.A1(new_n1042_), .A2(\in1[7] ), .A3(new_n1013_), .ZN(new_n1044_));
  OAI21_X1   g0402(.A1(\in0[7] ), .A2(new_n1043_), .B(new_n1044_), .ZN(new_n1045_));
  INV_X1     g0403(.I(\in0[8] ), .ZN(new_n1046_));
  NOR2_X1    g0404(.A1(new_n1046_), .A2(\in1[8] ), .ZN(new_n1047_));
  INV_X1     g0405(.I(new_n1047_), .ZN(new_n1048_));
  AOI21_X1   g0406(.A1(new_n1045_), .A2(new_n1048_), .B(new_n1010_), .ZN(new_n1049_));
  INV_X1     g0407(.I(\in1[9] ), .ZN(new_n1050_));
  NOR2_X1    g0408(.A1(new_n1050_), .A2(\in0[9] ), .ZN(new_n1051_));
  INV_X1     g0409(.I(new_n1051_), .ZN(new_n1052_));
  INV_X1     g0410(.I(\in0[9] ), .ZN(new_n1053_));
  NOR2_X1    g0411(.A1(new_n1053_), .A2(\in1[9] ), .ZN(new_n1054_));
  AOI21_X1   g0412(.A1(new_n1049_), .A2(new_n1052_), .B(new_n1054_), .ZN(new_n1055_));
  OAI21_X1   g0413(.A1(new_n1055_), .A2(new_n1008_), .B(new_n1006_), .ZN(new_n1056_));
  AOI21_X1   g0414(.A1(new_n1056_), .A2(new_n1003_), .B(\in0[11] ), .ZN(new_n1057_));
  NOR2_X1    g0415(.A1(new_n1056_), .A2(new_n1003_), .ZN(new_n1058_));
  INV_X1     g0416(.I(\in1[12] ), .ZN(new_n1059_));
  NOR2_X1    g0417(.A1(new_n1059_), .A2(\in0[12] ), .ZN(new_n1060_));
  NOR3_X1    g0418(.A1(new_n1057_), .A2(new_n1058_), .A3(new_n1060_), .ZN(new_n1061_));
  INV_X1     g0419(.I(\in0[12] ), .ZN(new_n1062_));
  NOR2_X1    g0420(.A1(new_n1062_), .A2(\in1[12] ), .ZN(new_n1063_));
  OAI21_X1   g0421(.A1(new_n1061_), .A2(new_n1063_), .B(new_n1002_), .ZN(new_n1064_));
  AOI21_X1   g0422(.A1(new_n1064_), .A2(new_n999_), .B(\in1[14] ), .ZN(new_n1065_));
  NAND3_X1   g0423(.A1(new_n1064_), .A2(\in1[14] ), .A3(new_n999_), .ZN(new_n1066_));
  OAI21_X1   g0424(.A1(\in0[14] ), .A2(new_n1065_), .B(new_n1066_), .ZN(new_n1067_));
  INV_X1     g0425(.I(\in0[15] ), .ZN(new_n1068_));
  NOR2_X1    g0426(.A1(new_n1068_), .A2(\in1[15] ), .ZN(new_n1069_));
  INV_X1     g0427(.I(new_n1069_), .ZN(new_n1070_));
  AOI21_X1   g0428(.A1(new_n1067_), .A2(new_n1070_), .B(new_n996_), .ZN(new_n1071_));
  INV_X1     g0429(.I(\in0[16] ), .ZN(new_n1072_));
  NOR2_X1    g0430(.A1(new_n1072_), .A2(\in1[16] ), .ZN(new_n1073_));
  OAI21_X1   g0431(.A1(new_n1071_), .A2(new_n1073_), .B(new_n994_), .ZN(new_n1074_));
  INV_X1     g0432(.I(\in1[17] ), .ZN(new_n1075_));
  NOR2_X1    g0433(.A1(new_n1075_), .A2(\in0[17] ), .ZN(new_n1076_));
  INV_X1     g0434(.I(\in0[17] ), .ZN(new_n1077_));
  NOR2_X1    g0435(.A1(new_n1077_), .A2(\in1[17] ), .ZN(new_n1078_));
  INV_X1     g0436(.I(new_n1078_), .ZN(new_n1079_));
  OAI21_X1   g0437(.A1(new_n1074_), .A2(new_n1076_), .B(new_n1079_), .ZN(new_n1080_));
  AOI21_X1   g0438(.A1(new_n1080_), .A2(new_n991_), .B(new_n988_), .ZN(new_n1081_));
  OAI21_X1   g0439(.A1(new_n1081_), .A2(\in1[19] ), .B(new_n986_), .ZN(new_n1082_));
  NAND2_X1   g0440(.A1(new_n1081_), .A2(\in1[19] ), .ZN(new_n1083_));
  INV_X1     g0441(.I(\in1[20] ), .ZN(new_n1084_));
  NOR2_X1    g0442(.A1(new_n1084_), .A2(\in0[20] ), .ZN(new_n1085_));
  INV_X1     g0443(.I(new_n1085_), .ZN(new_n1086_));
  NAND3_X1   g0444(.A1(new_n1082_), .A2(new_n1083_), .A3(new_n1086_), .ZN(new_n1087_));
  INV_X1     g0445(.I(\in0[20] ), .ZN(new_n1088_));
  NOR2_X1    g0446(.A1(new_n1088_), .A2(\in1[20] ), .ZN(new_n1089_));
  INV_X1     g0447(.I(new_n1089_), .ZN(new_n1090_));
  AOI21_X1   g0448(.A1(new_n1087_), .A2(new_n1090_), .B(new_n985_), .ZN(new_n1091_));
  OAI21_X1   g0449(.A1(new_n1091_), .A2(new_n983_), .B(new_n981_), .ZN(new_n1092_));
  NOR3_X1    g0450(.A1(new_n1091_), .A2(new_n981_), .A3(new_n983_), .ZN(new_n1093_));
  AOI21_X1   g0451(.A1(new_n980_), .A2(new_n1092_), .B(new_n1093_), .ZN(new_n1094_));
  INV_X1     g0452(.I(\in0[23] ), .ZN(new_n1095_));
  NOR2_X1    g0453(.A1(new_n1095_), .A2(\in1[23] ), .ZN(new_n1096_));
  OAI21_X1   g0454(.A1(new_n1094_), .A2(new_n1096_), .B(new_n979_), .ZN(new_n1097_));
  INV_X1     g0455(.I(\in0[24] ), .ZN(new_n1098_));
  NOR2_X1    g0456(.A1(new_n1098_), .A2(\in1[24] ), .ZN(new_n1099_));
  INV_X1     g0457(.I(new_n1099_), .ZN(new_n1100_));
  AOI21_X1   g0458(.A1(new_n1097_), .A2(new_n1100_), .B(new_n976_), .ZN(new_n1101_));
  INV_X1     g0459(.I(\in1[25] ), .ZN(new_n1102_));
  NOR2_X1    g0460(.A1(new_n1102_), .A2(\in0[25] ), .ZN(new_n1103_));
  INV_X1     g0461(.I(new_n1103_), .ZN(new_n1104_));
  INV_X1     g0462(.I(\in0[25] ), .ZN(new_n1105_));
  NOR2_X1    g0463(.A1(new_n1105_), .A2(\in1[25] ), .ZN(new_n1106_));
  AOI21_X1   g0464(.A1(new_n1101_), .A2(new_n1104_), .B(new_n1106_), .ZN(new_n1107_));
  OAI21_X1   g0465(.A1(new_n1107_), .A2(new_n974_), .B(new_n972_), .ZN(new_n1108_));
  AOI21_X1   g0466(.A1(new_n1108_), .A2(new_n969_), .B(\in0[27] ), .ZN(new_n1109_));
  NOR2_X1    g0467(.A1(new_n1108_), .A2(new_n969_), .ZN(new_n1110_));
  INV_X1     g0468(.I(\in1[28] ), .ZN(new_n1111_));
  NOR2_X1    g0469(.A1(new_n1111_), .A2(\in0[28] ), .ZN(new_n1112_));
  NOR3_X1    g0470(.A1(new_n1109_), .A2(new_n1110_), .A3(new_n1112_), .ZN(new_n1113_));
  INV_X1     g0471(.I(\in0[28] ), .ZN(new_n1114_));
  NOR2_X1    g0472(.A1(new_n1114_), .A2(\in1[28] ), .ZN(new_n1115_));
  OAI21_X1   g0473(.A1(new_n1113_), .A2(new_n1115_), .B(new_n968_), .ZN(new_n1116_));
  AOI21_X1   g0474(.A1(new_n1116_), .A2(new_n965_), .B(\in1[30] ), .ZN(new_n1117_));
  NAND3_X1   g0475(.A1(new_n1116_), .A2(\in1[30] ), .A3(new_n965_), .ZN(new_n1118_));
  OAI21_X1   g0476(.A1(\in0[30] ), .A2(new_n1117_), .B(new_n1118_), .ZN(new_n1119_));
  INV_X1     g0477(.I(\in1[31] ), .ZN(new_n1120_));
  NOR2_X1    g0478(.A1(new_n1120_), .A2(\in0[31] ), .ZN(new_n1121_));
  INV_X1     g0479(.I(\in0[31] ), .ZN(new_n1122_));
  NOR2_X1    g0480(.A1(new_n1122_), .A2(\in1[31] ), .ZN(new_n1123_));
  INV_X1     g0481(.I(new_n1123_), .ZN(new_n1124_));
  OAI21_X1   g0482(.A1(new_n1119_), .A2(new_n1121_), .B(new_n1124_), .ZN(new_n1125_));
  INV_X1     g0483(.I(new_n960_), .ZN(new_n1126_));
  INV_X1     g0484(.I(\in1[32] ), .ZN(new_n1127_));
  OAI22_X1   g0485(.A1(new_n947_), .A2(\in1[33] ), .B1(new_n958_), .B2(\in1[34] ), .ZN(new_n1128_));
  AOI21_X1   g0486(.A1(new_n947_), .A2(\in1[33] ), .B(new_n946_), .ZN(new_n1129_));
  AOI21_X1   g0487(.A1(new_n1127_), .A2(new_n1129_), .B(new_n1128_), .ZN(new_n1130_));
  OAI22_X1   g0488(.A1(new_n1130_), .A2(new_n1126_), .B1(new_n959_), .B2(\in1[35] ), .ZN(new_n1131_));
  NAND2_X1   g0489(.A1(new_n1131_), .A2(new_n957_), .ZN(new_n1132_));
  NOR2_X1    g0490(.A1(new_n953_), .A2(\in1[36] ), .ZN(new_n1133_));
  NOR2_X1    g0491(.A1(new_n954_), .A2(\in1[37] ), .ZN(new_n1134_));
  NOR2_X1    g0492(.A1(new_n1133_), .A2(new_n1134_), .ZN(new_n1135_));
  AOI21_X1   g0493(.A1(new_n954_), .A2(\in1[37] ), .B(new_n1135_), .ZN(new_n1136_));
  INV_X1     g0494(.I(\in1[38] ), .ZN(new_n1137_));
  AOI22_X1   g0495(.A1(\in0[38] ), .A2(new_n1137_), .B1(new_n950_), .B2(\in0[39] ), .ZN(new_n1138_));
  NOR2_X1    g0496(.A1(new_n1138_), .A2(new_n951_), .ZN(new_n1139_));
  AOI21_X1   g0497(.A1(new_n1136_), .A2(new_n952_), .B(new_n1139_), .ZN(new_n1140_));
  AND2_X2    g0498(.A1(new_n1132_), .A2(new_n1140_), .Z(new_n1141_));
  INV_X1     g0499(.I(new_n1141_), .ZN(new_n1142_));
  AOI21_X1   g0500(.A1(new_n1125_), .A2(new_n962_), .B(new_n1142_), .ZN(new_n1143_));
  OAI21_X1   g0501(.A1(new_n1143_), .A2(new_n945_), .B(new_n943_), .ZN(new_n1144_));
  AOI21_X1   g0502(.A1(new_n898_), .A2(\in1[48] ), .B(new_n899_), .ZN(new_n1145_));
  NAND3_X1   g0503(.A1(new_n890_), .A2(new_n893_), .A3(new_n1145_), .ZN(new_n1146_));
  INV_X1     g0504(.I(new_n1146_), .ZN(new_n1147_));
  AOI21_X1   g0505(.A1(new_n1144_), .A2(new_n1147_), .B(new_n913_), .ZN(new_n1148_));
  INV_X1     g0506(.I(new_n880_), .ZN(new_n1149_));
  INV_X1     g0507(.I(\in1[56] ), .ZN(new_n1150_));
  OAI22_X1   g0508(.A1(new_n867_), .A2(\in1[57] ), .B1(new_n878_), .B2(\in1[58] ), .ZN(new_n1151_));
  AOI21_X1   g0509(.A1(new_n867_), .A2(\in1[57] ), .B(new_n866_), .ZN(new_n1152_));
  AOI21_X1   g0510(.A1(new_n1150_), .A2(new_n1152_), .B(new_n1151_), .ZN(new_n1153_));
  OAI22_X1   g0511(.A1(new_n1153_), .A2(new_n1149_), .B1(new_n879_), .B2(\in1[59] ), .ZN(new_n1154_));
  NAND2_X1   g0512(.A1(new_n1154_), .A2(new_n877_), .ZN(new_n1155_));
  NOR2_X1    g0513(.A1(new_n873_), .A2(\in1[60] ), .ZN(new_n1156_));
  NOR2_X1    g0514(.A1(new_n874_), .A2(\in1[61] ), .ZN(new_n1157_));
  NOR2_X1    g0515(.A1(new_n1156_), .A2(new_n1157_), .ZN(new_n1158_));
  AOI21_X1   g0516(.A1(new_n874_), .A2(\in1[61] ), .B(new_n1158_), .ZN(new_n1159_));
  INV_X1     g0517(.I(\in1[62] ), .ZN(new_n1160_));
  AOI22_X1   g0518(.A1(\in0[62] ), .A2(new_n1160_), .B1(new_n870_), .B2(\in0[63] ), .ZN(new_n1161_));
  NOR2_X1    g0519(.A1(new_n1161_), .A2(new_n871_), .ZN(new_n1162_));
  AOI21_X1   g0520(.A1(new_n1159_), .A2(new_n872_), .B(new_n1162_), .ZN(new_n1163_));
  AND2_X2    g0521(.A1(new_n1155_), .A2(new_n1163_), .Z(new_n1164_));
  OAI21_X1   g0522(.A1(new_n1148_), .A2(new_n881_), .B(new_n1164_), .ZN(new_n1165_));
  AOI21_X1   g0523(.A1(new_n1165_), .A2(new_n865_), .B(new_n862_), .ZN(new_n1166_));
  NOR2_X1    g0524(.A1(new_n842_), .A2(\in0[68] ), .ZN(new_n1167_));
  NOR3_X1    g0525(.A1(new_n839_), .A2(new_n841_), .A3(new_n1167_), .ZN(new_n1168_));
  INV_X1     g0526(.I(new_n1168_), .ZN(new_n1169_));
  OAI21_X1   g0527(.A1(new_n1166_), .A2(new_n1169_), .B(new_n849_), .ZN(new_n1170_));
  INV_X1     g0528(.I(\in1[75] ), .ZN(new_n1171_));
  INV_X1     g0529(.I(\in1[74] ), .ZN(new_n1172_));
  AOI22_X1   g0530(.A1(\in0[73] ), .A2(new_n826_), .B1(new_n1172_), .B2(\in0[74] ), .ZN(new_n1173_));
  NAND2_X1   g0531(.A1(new_n832_), .A2(\in0[72] ), .ZN(new_n1174_));
  OAI21_X1   g0532(.A1(new_n827_), .A2(new_n1174_), .B(new_n1173_), .ZN(new_n1175_));
  AOI22_X1   g0533(.A1(new_n1175_), .A2(new_n830_), .B1(\in0[75] ), .B2(new_n1171_), .ZN(new_n1176_));
  INV_X1     g0534(.I(new_n1176_), .ZN(new_n1177_));
  AOI21_X1   g0535(.A1(new_n1170_), .A2(new_n834_), .B(new_n1177_), .ZN(new_n1178_));
  OAI21_X1   g0536(.A1(new_n1178_), .A2(new_n825_), .B(new_n822_), .ZN(new_n1179_));
  INV_X1     g0537(.I(new_n798_), .ZN(new_n1180_));
  NOR2_X1    g0538(.A1(new_n803_), .A2(\in0[80] ), .ZN(new_n1181_));
  NOR3_X1    g0539(.A1(new_n1180_), .A2(new_n802_), .A3(new_n1181_), .ZN(new_n1182_));
  AOI21_X1   g0540(.A1(new_n1179_), .A2(new_n1182_), .B(new_n807_), .ZN(new_n1183_));
  AOI22_X1   g0541(.A1(\in0[84] ), .A2(new_n789_), .B1(new_n791_), .B2(\in0[85] ), .ZN(new_n1184_));
  NOR2_X1    g0542(.A1(new_n1184_), .A2(new_n792_), .ZN(new_n1185_));
  INV_X1     g0543(.I(new_n1185_), .ZN(new_n1186_));
  INV_X1     g0544(.I(\in1[86] ), .ZN(new_n1187_));
  AOI22_X1   g0545(.A1(\in0[86] ), .A2(new_n1187_), .B1(new_n785_), .B2(\in0[87] ), .ZN(new_n1188_));
  OAI22_X1   g0546(.A1(new_n1186_), .A2(new_n788_), .B1(new_n786_), .B2(new_n1188_), .ZN(new_n1189_));
  INV_X1     g0547(.I(new_n1189_), .ZN(new_n1190_));
  OAI21_X1   g0548(.A1(new_n1183_), .A2(new_n794_), .B(new_n1190_), .ZN(new_n1191_));
  AOI21_X1   g0549(.A1(new_n1191_), .A2(new_n783_), .B(new_n780_), .ZN(new_n1192_));
  NOR2_X1    g0550(.A1(new_n760_), .A2(\in0[92] ), .ZN(new_n1193_));
  NOR3_X1    g0551(.A1(new_n757_), .A2(new_n759_), .A3(new_n1193_), .ZN(new_n1194_));
  INV_X1     g0552(.I(new_n1194_), .ZN(new_n1195_));
  OAI21_X1   g0553(.A1(new_n1192_), .A2(new_n1195_), .B(new_n767_), .ZN(new_n1196_));
  INV_X1     g0554(.I(\in1[99] ), .ZN(new_n1197_));
  INV_X1     g0555(.I(\in1[98] ), .ZN(new_n1198_));
  AOI22_X1   g0556(.A1(\in0[97] ), .A2(new_n744_), .B1(new_n1198_), .B2(\in0[98] ), .ZN(new_n1199_));
  NAND2_X1   g0557(.A1(new_n750_), .A2(\in0[96] ), .ZN(new_n1200_));
  OAI21_X1   g0558(.A1(new_n745_), .A2(new_n1200_), .B(new_n1199_), .ZN(new_n1201_));
  AOI22_X1   g0559(.A1(new_n1201_), .A2(new_n748_), .B1(\in0[99] ), .B2(new_n1197_), .ZN(new_n1202_));
  INV_X1     g0560(.I(new_n1202_), .ZN(new_n1203_));
  AOI21_X1   g0561(.A1(new_n1196_), .A2(new_n752_), .B(new_n1203_), .ZN(new_n1204_));
  OAI21_X1   g0562(.A1(new_n1204_), .A2(new_n743_), .B(new_n740_), .ZN(new_n1205_));
  INV_X1     g0563(.I(new_n716_), .ZN(new_n1206_));
  NOR2_X1    g0564(.A1(new_n721_), .A2(\in0[104] ), .ZN(new_n1207_));
  NOR3_X1    g0565(.A1(new_n1206_), .A2(new_n720_), .A3(new_n1207_), .ZN(new_n1208_));
  AOI21_X1   g0566(.A1(new_n1205_), .A2(new_n1208_), .B(new_n725_), .ZN(new_n1209_));
  AOI22_X1   g0567(.A1(\in0[108] ), .A2(new_n707_), .B1(new_n709_), .B2(\in0[109] ), .ZN(new_n1210_));
  NOR2_X1    g0568(.A1(new_n1210_), .A2(new_n710_), .ZN(new_n1211_));
  INV_X1     g0569(.I(new_n1211_), .ZN(new_n1212_));
  INV_X1     g0570(.I(\in1[110] ), .ZN(new_n1213_));
  AOI22_X1   g0571(.A1(\in0[110] ), .A2(new_n1213_), .B1(new_n703_), .B2(\in0[111] ), .ZN(new_n1214_));
  OAI22_X1   g0572(.A1(new_n1212_), .A2(new_n706_), .B1(new_n704_), .B2(new_n1214_), .ZN(new_n1215_));
  INV_X1     g0573(.I(new_n1215_), .ZN(new_n1216_));
  OAI21_X1   g0574(.A1(new_n1209_), .A2(new_n712_), .B(new_n1216_), .ZN(new_n1217_));
  AOI21_X1   g0575(.A1(new_n1217_), .A2(new_n701_), .B(new_n698_), .ZN(new_n1218_));
  NOR2_X1    g0576(.A1(new_n678_), .A2(\in0[116] ), .ZN(new_n1219_));
  NOR3_X1    g0577(.A1(new_n675_), .A2(new_n677_), .A3(new_n1219_), .ZN(new_n1220_));
  INV_X1     g0578(.I(new_n1220_), .ZN(new_n1221_));
  OAI21_X1   g0579(.A1(new_n1218_), .A2(new_n1221_), .B(new_n685_), .ZN(new_n1222_));
  INV_X1     g0580(.I(\in1[123] ), .ZN(new_n1223_));
  INV_X1     g0581(.I(\in1[122] ), .ZN(new_n1224_));
  AOI22_X1   g0582(.A1(\in0[121] ), .A2(new_n662_), .B1(new_n1224_), .B2(\in0[122] ), .ZN(new_n1225_));
  NAND2_X1   g0583(.A1(new_n668_), .A2(\in0[120] ), .ZN(new_n1226_));
  OAI21_X1   g0584(.A1(new_n663_), .A2(new_n1226_), .B(new_n1225_), .ZN(new_n1227_));
  AOI22_X1   g0585(.A1(new_n1227_), .A2(new_n666_), .B1(\in0[123] ), .B2(new_n1223_), .ZN(new_n1228_));
  INV_X1     g0586(.I(new_n1228_), .ZN(new_n1229_));
  AOI21_X1   g0587(.A1(new_n1222_), .A2(new_n670_), .B(new_n1229_), .ZN(new_n1230_));
  OAI21_X1   g0588(.A1(new_n1230_), .A2(new_n661_), .B(new_n657_), .ZN(new_n1231_));
  NAND2_X1   g0589(.A1(new_n644_), .A2(\in1[127] ), .ZN(new_n1232_));
  INV_X1     g0590(.I(new_n1232_), .ZN(new_n1233_));
  NOR3_X1    g0591(.A1(new_n1231_), .A2(new_n643_), .A3(new_n1233_), .ZN(new_n1234_));
  INV_X1     g0592(.I(\in0[0] ), .ZN(new_n1235_));
  INV_X1     g0593(.I(new_n670_), .ZN(new_n1236_));
  INV_X1     g0594(.I(new_n701_), .ZN(new_n1237_));
  INV_X1     g0595(.I(new_n752_), .ZN(new_n1238_));
  INV_X1     g0596(.I(new_n783_), .ZN(new_n1239_));
  INV_X1     g0597(.I(new_n834_), .ZN(new_n1240_));
  INV_X1     g0598(.I(new_n865_), .ZN(new_n1241_));
  INV_X1     g0599(.I(new_n881_), .ZN(new_n1242_));
  INV_X1     g0600(.I(new_n943_), .ZN(new_n1243_));
  INV_X1     g0601(.I(new_n945_), .ZN(new_n1244_));
  INV_X1     g0602(.I(\in0[30] ), .ZN(new_n1245_));
  INV_X1     g0603(.I(\in1[30] ), .ZN(new_n1246_));
  INV_X1     g0604(.I(\in0[27] ), .ZN(new_n1247_));
  INV_X1     g0605(.I(new_n974_), .ZN(new_n1248_));
  INV_X1     g0606(.I(new_n976_), .ZN(new_n1249_));
  INV_X1     g0607(.I(new_n983_), .ZN(new_n1250_));
  INV_X1     g0608(.I(new_n985_), .ZN(new_n1251_));
  INV_X1     g0609(.I(\in1[19] ), .ZN(new_n1252_));
  INV_X1     g0610(.I(new_n988_), .ZN(new_n1253_));
  INV_X1     g0611(.I(new_n996_), .ZN(new_n1254_));
  INV_X1     g0612(.I(\in0[14] ), .ZN(new_n1255_));
  INV_X1     g0613(.I(\in1[14] ), .ZN(new_n1256_));
  INV_X1     g0614(.I(\in0[11] ), .ZN(new_n1257_));
  INV_X1     g0615(.I(new_n1008_), .ZN(new_n1258_));
  INV_X1     g0616(.I(new_n1010_), .ZN(new_n1259_));
  INV_X1     g0617(.I(\in0[7] ), .ZN(new_n1260_));
  INV_X1     g0618(.I(\in1[7] ), .ZN(new_n1261_));
  INV_X1     g0619(.I(new_n1018_), .ZN(new_n1262_));
  INV_X1     g0620(.I(\in0[2] ), .ZN(new_n1263_));
  NOR2_X1    g0621(.A1(new_n1235_), .A2(\in1[0] ), .ZN(new_n1264_));
  INV_X1     g0622(.I(\in0[1] ), .ZN(new_n1265_));
  NOR2_X1    g0623(.A1(new_n1265_), .A2(\in1[1] ), .ZN(new_n1266_));
  NAND2_X1   g0624(.A1(new_n1265_), .A2(\in1[1] ), .ZN(new_n1267_));
  OAI21_X1   g0625(.A1(new_n1264_), .A2(new_n1266_), .B(new_n1267_), .ZN(new_n1268_));
  AOI21_X1   g0626(.A1(new_n1268_), .A2(\in1[2] ), .B(new_n1263_), .ZN(new_n1269_));
  NOR2_X1    g0627(.A1(new_n1268_), .A2(\in1[2] ), .ZN(new_n1270_));
  NOR3_X1    g0628(.A1(new_n1269_), .A2(new_n1270_), .A3(new_n1031_), .ZN(new_n1271_));
  OAI22_X1   g0629(.A1(new_n1271_), .A2(new_n1020_), .B1(new_n1034_), .B2(\in1[4] ), .ZN(new_n1272_));
  INV_X1     g0630(.I(new_n1038_), .ZN(new_n1273_));
  NAND3_X1   g0631(.A1(new_n1272_), .A2(new_n1262_), .A3(new_n1273_), .ZN(new_n1274_));
  INV_X1     g0632(.I(new_n1041_), .ZN(new_n1275_));
  AOI21_X1   g0633(.A1(new_n1274_), .A2(new_n1275_), .B(new_n1015_), .ZN(new_n1276_));
  OAI21_X1   g0634(.A1(new_n1276_), .A2(new_n1012_), .B(new_n1261_), .ZN(new_n1277_));
  NOR3_X1    g0635(.A1(new_n1276_), .A2(new_n1261_), .A3(new_n1012_), .ZN(new_n1278_));
  AOI21_X1   g0636(.A1(new_n1260_), .A2(new_n1277_), .B(new_n1278_), .ZN(new_n1279_));
  OAI21_X1   g0637(.A1(new_n1279_), .A2(new_n1047_), .B(new_n1259_), .ZN(new_n1280_));
  INV_X1     g0638(.I(new_n1054_), .ZN(new_n1281_));
  OAI21_X1   g0639(.A1(new_n1280_), .A2(new_n1051_), .B(new_n1281_), .ZN(new_n1282_));
  AOI21_X1   g0640(.A1(new_n1282_), .A2(new_n1258_), .B(new_n1005_), .ZN(new_n1283_));
  OAI21_X1   g0641(.A1(new_n1283_), .A2(\in1[11] ), .B(new_n1257_), .ZN(new_n1284_));
  NAND2_X1   g0642(.A1(new_n1277_), .A2(new_n1260_), .ZN(new_n1285_));
  AOI21_X1   g0643(.A1(new_n1285_), .A2(new_n1044_), .B(new_n1047_), .ZN(new_n1286_));
  NOR3_X1    g0644(.A1(new_n1286_), .A2(new_n1010_), .A3(new_n1051_), .ZN(new_n1287_));
  OAI21_X1   g0645(.A1(new_n1287_), .A2(new_n1054_), .B(new_n1258_), .ZN(new_n1288_));
  NAND3_X1   g0646(.A1(new_n1288_), .A2(\in1[11] ), .A3(new_n1006_), .ZN(new_n1289_));
  INV_X1     g0647(.I(new_n1060_), .ZN(new_n1290_));
  NAND3_X1   g0648(.A1(new_n1284_), .A2(new_n1289_), .A3(new_n1290_), .ZN(new_n1291_));
  INV_X1     g0649(.I(new_n1063_), .ZN(new_n1292_));
  AOI21_X1   g0650(.A1(new_n1291_), .A2(new_n1292_), .B(new_n1001_), .ZN(new_n1293_));
  OAI21_X1   g0651(.A1(new_n1293_), .A2(new_n998_), .B(new_n1256_), .ZN(new_n1294_));
  NOR3_X1    g0652(.A1(new_n1293_), .A2(new_n1256_), .A3(new_n998_), .ZN(new_n1295_));
  AOI21_X1   g0653(.A1(new_n1255_), .A2(new_n1294_), .B(new_n1295_), .ZN(new_n1296_));
  OAI21_X1   g0654(.A1(new_n1296_), .A2(new_n1069_), .B(new_n1254_), .ZN(new_n1297_));
  INV_X1     g0655(.I(new_n1073_), .ZN(new_n1298_));
  AOI21_X1   g0656(.A1(new_n1297_), .A2(new_n1298_), .B(new_n993_), .ZN(new_n1299_));
  INV_X1     g0657(.I(new_n1076_), .ZN(new_n1300_));
  AOI21_X1   g0658(.A1(new_n1299_), .A2(new_n1300_), .B(new_n1078_), .ZN(new_n1301_));
  OAI21_X1   g0659(.A1(new_n1301_), .A2(new_n990_), .B(new_n1253_), .ZN(new_n1302_));
  AOI21_X1   g0660(.A1(new_n1302_), .A2(new_n1252_), .B(\in0[19] ), .ZN(new_n1303_));
  NAND2_X1   g0661(.A1(new_n1294_), .A2(new_n1255_), .ZN(new_n1304_));
  AOI21_X1   g0662(.A1(new_n1304_), .A2(new_n1066_), .B(new_n1069_), .ZN(new_n1305_));
  OAI21_X1   g0663(.A1(new_n1305_), .A2(new_n996_), .B(new_n1298_), .ZN(new_n1306_));
  NAND3_X1   g0664(.A1(new_n1306_), .A2(new_n994_), .A3(new_n1300_), .ZN(new_n1307_));
  AOI21_X1   g0665(.A1(new_n1307_), .A2(new_n1079_), .B(new_n990_), .ZN(new_n1308_));
  NOR3_X1    g0666(.A1(new_n1308_), .A2(new_n1252_), .A3(new_n988_), .ZN(new_n1309_));
  NOR3_X1    g0667(.A1(new_n1303_), .A2(new_n1309_), .A3(new_n1085_), .ZN(new_n1310_));
  OAI21_X1   g0668(.A1(new_n1310_), .A2(new_n1089_), .B(new_n1251_), .ZN(new_n1311_));
  AOI21_X1   g0669(.A1(new_n1311_), .A2(new_n1250_), .B(\in1[22] ), .ZN(new_n1312_));
  NAND3_X1   g0670(.A1(new_n1311_), .A2(\in1[22] ), .A3(new_n1250_), .ZN(new_n1313_));
  OAI21_X1   g0671(.A1(\in0[22] ), .A2(new_n1312_), .B(new_n1313_), .ZN(new_n1314_));
  INV_X1     g0672(.I(new_n1096_), .ZN(new_n1315_));
  AOI21_X1   g0673(.A1(new_n1314_), .A2(new_n1315_), .B(new_n978_), .ZN(new_n1316_));
  OAI21_X1   g0674(.A1(new_n1316_), .A2(new_n1099_), .B(new_n1249_), .ZN(new_n1317_));
  INV_X1     g0675(.I(new_n1106_), .ZN(new_n1318_));
  OAI21_X1   g0676(.A1(new_n1317_), .A2(new_n1103_), .B(new_n1318_), .ZN(new_n1319_));
  AOI21_X1   g0677(.A1(new_n1319_), .A2(new_n1248_), .B(new_n971_), .ZN(new_n1320_));
  OAI21_X1   g0678(.A1(new_n1320_), .A2(\in1[27] ), .B(new_n1247_), .ZN(new_n1321_));
  OAI21_X1   g0679(.A1(new_n1308_), .A2(new_n988_), .B(new_n1252_), .ZN(new_n1322_));
  AOI21_X1   g0680(.A1(new_n986_), .A2(new_n1322_), .B(new_n1309_), .ZN(new_n1323_));
  AOI21_X1   g0681(.A1(new_n1323_), .A2(new_n1086_), .B(new_n1089_), .ZN(new_n1324_));
  OAI21_X1   g0682(.A1(new_n1324_), .A2(new_n985_), .B(new_n1250_), .ZN(new_n1325_));
  AOI21_X1   g0683(.A1(new_n1325_), .A2(new_n981_), .B(\in0[22] ), .ZN(new_n1326_));
  OAI21_X1   g0684(.A1(new_n1326_), .A2(new_n1093_), .B(new_n1315_), .ZN(new_n1327_));
  AOI21_X1   g0685(.A1(new_n1327_), .A2(new_n979_), .B(new_n1099_), .ZN(new_n1328_));
  NOR3_X1    g0686(.A1(new_n1328_), .A2(new_n976_), .A3(new_n1103_), .ZN(new_n1329_));
  OAI21_X1   g0687(.A1(new_n1329_), .A2(new_n1106_), .B(new_n1248_), .ZN(new_n1330_));
  NAND3_X1   g0688(.A1(new_n1330_), .A2(\in1[27] ), .A3(new_n972_), .ZN(new_n1331_));
  INV_X1     g0689(.I(new_n1112_), .ZN(new_n1332_));
  NAND3_X1   g0690(.A1(new_n1321_), .A2(new_n1331_), .A3(new_n1332_), .ZN(new_n1333_));
  INV_X1     g0691(.I(new_n1115_), .ZN(new_n1334_));
  AOI21_X1   g0692(.A1(new_n1333_), .A2(new_n1334_), .B(new_n967_), .ZN(new_n1335_));
  OAI21_X1   g0693(.A1(new_n1335_), .A2(new_n964_), .B(new_n1246_), .ZN(new_n1336_));
  NOR3_X1    g0694(.A1(new_n1335_), .A2(new_n1246_), .A3(new_n964_), .ZN(new_n1337_));
  AOI21_X1   g0695(.A1(new_n1245_), .A2(new_n1336_), .B(new_n1337_), .ZN(new_n1338_));
  INV_X1     g0696(.I(new_n1121_), .ZN(new_n1339_));
  AOI21_X1   g0697(.A1(new_n1338_), .A2(new_n1339_), .B(new_n1123_), .ZN(new_n1340_));
  OAI21_X1   g0698(.A1(new_n1340_), .A2(new_n961_), .B(new_n1141_), .ZN(new_n1341_));
  AOI21_X1   g0699(.A1(new_n1341_), .A2(new_n1244_), .B(new_n1243_), .ZN(new_n1342_));
  OAI21_X1   g0700(.A1(new_n1342_), .A2(new_n1146_), .B(new_n912_), .ZN(new_n1343_));
  INV_X1     g0701(.I(new_n1164_), .ZN(new_n1344_));
  AOI21_X1   g0702(.A1(new_n1343_), .A2(new_n1242_), .B(new_n1344_), .ZN(new_n1345_));
  OAI21_X1   g0703(.A1(new_n1345_), .A2(new_n1241_), .B(new_n861_), .ZN(new_n1346_));
  AOI21_X1   g0704(.A1(new_n1346_), .A2(new_n1168_), .B(new_n848_), .ZN(new_n1347_));
  OAI21_X1   g0705(.A1(new_n1347_), .A2(new_n1240_), .B(new_n1176_), .ZN(new_n1348_));
  AOI21_X1   g0706(.A1(new_n1348_), .A2(new_n824_), .B(new_n821_), .ZN(new_n1349_));
  INV_X1     g0707(.I(new_n1182_), .ZN(new_n1350_));
  OAI21_X1   g0708(.A1(new_n1349_), .A2(new_n1350_), .B(new_n806_), .ZN(new_n1351_));
  AOI21_X1   g0709(.A1(new_n1351_), .A2(new_n793_), .B(new_n1189_), .ZN(new_n1352_));
  OAI21_X1   g0710(.A1(new_n1352_), .A2(new_n1239_), .B(new_n779_), .ZN(new_n1353_));
  AOI21_X1   g0711(.A1(new_n1353_), .A2(new_n1194_), .B(new_n766_), .ZN(new_n1354_));
  OAI21_X1   g0712(.A1(new_n1354_), .A2(new_n1238_), .B(new_n1202_), .ZN(new_n1355_));
  AOI21_X1   g0713(.A1(new_n1355_), .A2(new_n742_), .B(new_n739_), .ZN(new_n1356_));
  INV_X1     g0714(.I(new_n1208_), .ZN(new_n1357_));
  OAI21_X1   g0715(.A1(new_n1356_), .A2(new_n1357_), .B(new_n724_), .ZN(new_n1358_));
  AOI21_X1   g0716(.A1(new_n1358_), .A2(new_n711_), .B(new_n1215_), .ZN(new_n1359_));
  OAI21_X1   g0717(.A1(new_n1359_), .A2(new_n1237_), .B(new_n697_), .ZN(new_n1360_));
  AOI21_X1   g0718(.A1(new_n1360_), .A2(new_n1220_), .B(new_n684_), .ZN(new_n1361_));
  OAI21_X1   g0719(.A1(new_n1361_), .A2(new_n1236_), .B(new_n1228_), .ZN(new_n1362_));
  AOI21_X1   g0720(.A1(new_n1362_), .A2(new_n660_), .B(new_n656_), .ZN(new_n1363_));
  AOI21_X1   g0721(.A1(new_n1363_), .A2(new_n1232_), .B(new_n1235_), .ZN(new_n1364_));
  NOR2_X1    g0722(.A1(new_n1364_), .A2(new_n1234_), .ZN(new_n1365_));
  OAI21_X1   g0723(.A1(new_n1231_), .A2(\in1[127] ), .B(\in0[127] ), .ZN(new_n1366_));
  INV_X1     g0724(.I(new_n1366_), .ZN(new_n1367_));
  INV_X1     g0725(.I(\in2[127] ), .ZN(new_n1368_));
  NOR2_X1    g0726(.A1(new_n1368_), .A2(\in3[127] ), .ZN(new_n1369_));
  INV_X1     g0727(.I(\in2[125] ), .ZN(new_n1370_));
  INV_X1     g0728(.I(\in2[126] ), .ZN(new_n1371_));
  AOI22_X1   g0729(.A1(new_n1370_), .A2(\in3[125] ), .B1(new_n1371_), .B2(\in3[126] ), .ZN(new_n1372_));
  INV_X1     g0730(.I(\in2[124] ), .ZN(new_n1373_));
  OAI22_X1   g0731(.A1(new_n1373_), .A2(\in3[124] ), .B1(new_n1370_), .B2(\in3[125] ), .ZN(new_n1374_));
  NAND2_X1   g0732(.A1(new_n1374_), .A2(new_n1372_), .ZN(new_n1375_));
  INV_X1     g0733(.I(\in3[126] ), .ZN(new_n1376_));
  NAND2_X1   g0734(.A1(new_n1376_), .A2(\in2[126] ), .ZN(new_n1377_));
  AOI21_X1   g0735(.A1(new_n1375_), .A2(new_n1377_), .B(new_n1369_), .ZN(new_n1378_));
  INV_X1     g0736(.I(new_n1378_), .ZN(new_n1379_));
  INV_X1     g0737(.I(new_n1372_), .ZN(new_n1380_));
  NAND2_X1   g0738(.A1(new_n1373_), .A2(\in3[124] ), .ZN(new_n1381_));
  INV_X1     g0739(.I(new_n1381_), .ZN(new_n1382_));
  NOR3_X1    g0740(.A1(new_n1380_), .A2(new_n1369_), .A3(new_n1382_), .ZN(new_n1383_));
  INV_X1     g0741(.I(new_n1383_), .ZN(new_n1384_));
  INV_X1     g0742(.I(\in3[121] ), .ZN(new_n1385_));
  NOR2_X1    g0743(.A1(new_n1385_), .A2(\in2[121] ), .ZN(new_n1386_));
  INV_X1     g0744(.I(\in2[122] ), .ZN(new_n1387_));
  INV_X1     g0745(.I(\in2[123] ), .ZN(new_n1388_));
  AOI22_X1   g0746(.A1(new_n1387_), .A2(\in3[122] ), .B1(new_n1388_), .B2(\in3[123] ), .ZN(new_n1389_));
  INV_X1     g0747(.I(new_n1389_), .ZN(new_n1390_));
  INV_X1     g0748(.I(\in3[120] ), .ZN(new_n1391_));
  NOR2_X1    g0749(.A1(new_n1391_), .A2(\in2[120] ), .ZN(new_n1392_));
  NOR3_X1    g0750(.A1(new_n1390_), .A2(new_n1386_), .A3(new_n1392_), .ZN(new_n1393_));
  INV_X1     g0751(.I(\in3[119] ), .ZN(new_n1394_));
  NOR2_X1    g0752(.A1(new_n1394_), .A2(\in2[119] ), .ZN(new_n1395_));
  INV_X1     g0753(.I(new_n1395_), .ZN(new_n1396_));
  INV_X1     g0754(.I(\in2[118] ), .ZN(new_n1397_));
  AOI21_X1   g0755(.A1(new_n1397_), .A2(\in3[118] ), .B(new_n1395_), .ZN(new_n1398_));
  INV_X1     g0756(.I(\in3[117] ), .ZN(new_n1399_));
  NOR2_X1    g0757(.A1(new_n1399_), .A2(\in2[117] ), .ZN(new_n1400_));
  INV_X1     g0758(.I(\in3[116] ), .ZN(new_n1401_));
  AOI22_X1   g0759(.A1(\in2[116] ), .A2(new_n1401_), .B1(new_n1399_), .B2(\in2[117] ), .ZN(new_n1402_));
  NOR2_X1    g0760(.A1(new_n1402_), .A2(new_n1400_), .ZN(new_n1403_));
  INV_X1     g0761(.I(\in2[119] ), .ZN(new_n1404_));
  OAI22_X1   g0762(.A1(new_n1397_), .A2(\in3[118] ), .B1(new_n1404_), .B2(\in3[119] ), .ZN(new_n1405_));
  AOI22_X1   g0763(.A1(new_n1403_), .A2(new_n1398_), .B1(new_n1396_), .B2(new_n1405_), .ZN(new_n1406_));
  INV_X1     g0764(.I(\in3[115] ), .ZN(new_n1407_));
  INV_X1     g0765(.I(\in2[114] ), .ZN(new_n1408_));
  INV_X1     g0766(.I(\in2[115] ), .ZN(new_n1409_));
  AOI22_X1   g0767(.A1(new_n1408_), .A2(\in3[114] ), .B1(new_n1409_), .B2(\in3[115] ), .ZN(new_n1410_));
  INV_X1     g0768(.I(\in2[113] ), .ZN(new_n1411_));
  OAI22_X1   g0769(.A1(new_n1411_), .A2(\in3[113] ), .B1(new_n1408_), .B2(\in3[114] ), .ZN(new_n1412_));
  INV_X1     g0770(.I(\in2[112] ), .ZN(new_n1413_));
  NAND2_X1   g0771(.A1(new_n1411_), .A2(\in3[113] ), .ZN(new_n1414_));
  INV_X1     g0772(.I(new_n1414_), .ZN(new_n1415_));
  NOR3_X1    g0773(.A1(new_n1415_), .A2(new_n1413_), .A3(\in3[112] ), .ZN(new_n1416_));
  OR2_X2     g0774(.A1(new_n1416_), .A2(new_n1412_), .Z(new_n1417_));
  AOI22_X1   g0775(.A1(new_n1417_), .A2(new_n1410_), .B1(\in2[115] ), .B2(new_n1407_), .ZN(new_n1418_));
  INV_X1     g0776(.I(new_n1418_), .ZN(new_n1419_));
  NAND2_X1   g0777(.A1(new_n1413_), .A2(\in3[112] ), .ZN(new_n1420_));
  NAND3_X1   g0778(.A1(new_n1410_), .A2(new_n1414_), .A3(new_n1420_), .ZN(new_n1421_));
  INV_X1     g0779(.I(new_n1421_), .ZN(new_n1422_));
  INV_X1     g0780(.I(\in2[110] ), .ZN(new_n1423_));
  INV_X1     g0781(.I(\in3[111] ), .ZN(new_n1424_));
  NOR2_X1    g0782(.A1(new_n1424_), .A2(\in2[111] ), .ZN(new_n1425_));
  AOI21_X1   g0783(.A1(new_n1423_), .A2(\in3[110] ), .B(new_n1425_), .ZN(new_n1426_));
  INV_X1     g0784(.I(new_n1426_), .ZN(new_n1427_));
  INV_X1     g0785(.I(\in3[108] ), .ZN(new_n1428_));
  NOR2_X1    g0786(.A1(new_n1428_), .A2(\in2[108] ), .ZN(new_n1429_));
  INV_X1     g0787(.I(\in3[109] ), .ZN(new_n1430_));
  NOR2_X1    g0788(.A1(new_n1430_), .A2(\in2[109] ), .ZN(new_n1431_));
  NOR3_X1    g0789(.A1(new_n1427_), .A2(new_n1429_), .A3(new_n1431_), .ZN(new_n1432_));
  INV_X1     g0790(.I(new_n1432_), .ZN(new_n1433_));
  INV_X1     g0791(.I(\in3[107] ), .ZN(new_n1434_));
  INV_X1     g0792(.I(\in2[106] ), .ZN(new_n1435_));
  INV_X1     g0793(.I(\in2[107] ), .ZN(new_n1436_));
  AOI22_X1   g0794(.A1(new_n1435_), .A2(\in3[106] ), .B1(new_n1436_), .B2(\in3[107] ), .ZN(new_n1437_));
  INV_X1     g0795(.I(\in2[105] ), .ZN(new_n1438_));
  OAI22_X1   g0796(.A1(new_n1438_), .A2(\in3[105] ), .B1(new_n1435_), .B2(\in3[106] ), .ZN(new_n1439_));
  INV_X1     g0797(.I(\in2[104] ), .ZN(new_n1440_));
  NAND2_X1   g0798(.A1(new_n1438_), .A2(\in3[105] ), .ZN(new_n1441_));
  INV_X1     g0799(.I(new_n1441_), .ZN(new_n1442_));
  NOR3_X1    g0800(.A1(new_n1442_), .A2(new_n1440_), .A3(\in3[104] ), .ZN(new_n1443_));
  OR2_X2     g0801(.A1(new_n1443_), .A2(new_n1439_), .Z(new_n1444_));
  AOI22_X1   g0802(.A1(new_n1444_), .A2(new_n1437_), .B1(\in2[107] ), .B2(new_n1434_), .ZN(new_n1445_));
  INV_X1     g0803(.I(new_n1445_), .ZN(new_n1446_));
  INV_X1     g0804(.I(\in3[103] ), .ZN(new_n1447_));
  NOR2_X1    g0805(.A1(new_n1447_), .A2(\in2[103] ), .ZN(new_n1448_));
  INV_X1     g0806(.I(new_n1448_), .ZN(new_n1449_));
  INV_X1     g0807(.I(\in2[102] ), .ZN(new_n1450_));
  AOI21_X1   g0808(.A1(new_n1450_), .A2(\in3[102] ), .B(new_n1448_), .ZN(new_n1451_));
  INV_X1     g0809(.I(\in3[101] ), .ZN(new_n1452_));
  NOR2_X1    g0810(.A1(new_n1452_), .A2(\in2[101] ), .ZN(new_n1453_));
  INV_X1     g0811(.I(\in3[100] ), .ZN(new_n1454_));
  AOI22_X1   g0812(.A1(\in2[100] ), .A2(new_n1454_), .B1(new_n1452_), .B2(\in2[101] ), .ZN(new_n1455_));
  NOR2_X1    g0813(.A1(new_n1455_), .A2(new_n1453_), .ZN(new_n1456_));
  INV_X1     g0814(.I(\in2[103] ), .ZN(new_n1457_));
  OAI22_X1   g0815(.A1(new_n1450_), .A2(\in3[102] ), .B1(new_n1457_), .B2(\in3[103] ), .ZN(new_n1458_));
  AOI22_X1   g0816(.A1(new_n1456_), .A2(new_n1451_), .B1(new_n1449_), .B2(new_n1458_), .ZN(new_n1459_));
  INV_X1     g0817(.I(new_n1451_), .ZN(new_n1460_));
  NOR2_X1    g0818(.A1(new_n1454_), .A2(\in2[100] ), .ZN(new_n1461_));
  NOR3_X1    g0819(.A1(new_n1460_), .A2(new_n1453_), .A3(new_n1461_), .ZN(new_n1462_));
  INV_X1     g0820(.I(new_n1462_), .ZN(new_n1463_));
  INV_X1     g0821(.I(\in3[97] ), .ZN(new_n1464_));
  NOR2_X1    g0822(.A1(new_n1464_), .A2(\in2[97] ), .ZN(new_n1465_));
  INV_X1     g0823(.I(\in2[98] ), .ZN(new_n1466_));
  INV_X1     g0824(.I(\in2[99] ), .ZN(new_n1467_));
  AOI22_X1   g0825(.A1(new_n1466_), .A2(\in3[98] ), .B1(new_n1467_), .B2(\in3[99] ), .ZN(new_n1468_));
  INV_X1     g0826(.I(new_n1468_), .ZN(new_n1469_));
  INV_X1     g0827(.I(\in3[96] ), .ZN(new_n1470_));
  NOR2_X1    g0828(.A1(new_n1470_), .A2(\in2[96] ), .ZN(new_n1471_));
  NOR3_X1    g0829(.A1(new_n1469_), .A2(new_n1465_), .A3(new_n1471_), .ZN(new_n1472_));
  INV_X1     g0830(.I(\in3[95] ), .ZN(new_n1473_));
  NOR2_X1    g0831(.A1(new_n1473_), .A2(\in2[95] ), .ZN(new_n1474_));
  INV_X1     g0832(.I(new_n1474_), .ZN(new_n1475_));
  INV_X1     g0833(.I(\in2[94] ), .ZN(new_n1476_));
  AOI21_X1   g0834(.A1(new_n1476_), .A2(\in3[94] ), .B(new_n1474_), .ZN(new_n1477_));
  INV_X1     g0835(.I(\in3[93] ), .ZN(new_n1478_));
  NOR2_X1    g0836(.A1(new_n1478_), .A2(\in2[93] ), .ZN(new_n1479_));
  INV_X1     g0837(.I(\in3[92] ), .ZN(new_n1480_));
  AOI22_X1   g0838(.A1(\in2[92] ), .A2(new_n1480_), .B1(new_n1478_), .B2(\in2[93] ), .ZN(new_n1481_));
  NOR2_X1    g0839(.A1(new_n1481_), .A2(new_n1479_), .ZN(new_n1482_));
  INV_X1     g0840(.I(\in2[95] ), .ZN(new_n1483_));
  OAI22_X1   g0841(.A1(new_n1476_), .A2(\in3[94] ), .B1(new_n1483_), .B2(\in3[95] ), .ZN(new_n1484_));
  AOI22_X1   g0842(.A1(new_n1482_), .A2(new_n1477_), .B1(new_n1475_), .B2(new_n1484_), .ZN(new_n1485_));
  INV_X1     g0843(.I(\in3[91] ), .ZN(new_n1486_));
  INV_X1     g0844(.I(\in2[90] ), .ZN(new_n1487_));
  INV_X1     g0845(.I(\in2[91] ), .ZN(new_n1488_));
  AOI22_X1   g0846(.A1(new_n1487_), .A2(\in3[90] ), .B1(new_n1488_), .B2(\in3[91] ), .ZN(new_n1489_));
  INV_X1     g0847(.I(\in2[89] ), .ZN(new_n1490_));
  OAI22_X1   g0848(.A1(new_n1490_), .A2(\in3[89] ), .B1(new_n1487_), .B2(\in3[90] ), .ZN(new_n1491_));
  INV_X1     g0849(.I(\in2[88] ), .ZN(new_n1492_));
  NAND2_X1   g0850(.A1(new_n1490_), .A2(\in3[89] ), .ZN(new_n1493_));
  INV_X1     g0851(.I(new_n1493_), .ZN(new_n1494_));
  NOR3_X1    g0852(.A1(new_n1494_), .A2(new_n1492_), .A3(\in3[88] ), .ZN(new_n1495_));
  OR2_X2     g0853(.A1(new_n1495_), .A2(new_n1491_), .Z(new_n1496_));
  AOI22_X1   g0854(.A1(new_n1496_), .A2(new_n1489_), .B1(\in2[91] ), .B2(new_n1486_), .ZN(new_n1497_));
  INV_X1     g0855(.I(new_n1497_), .ZN(new_n1498_));
  NAND2_X1   g0856(.A1(new_n1492_), .A2(\in3[88] ), .ZN(new_n1499_));
  NAND3_X1   g0857(.A1(new_n1489_), .A2(new_n1493_), .A3(new_n1499_), .ZN(new_n1500_));
  INV_X1     g0858(.I(new_n1500_), .ZN(new_n1501_));
  INV_X1     g0859(.I(\in2[86] ), .ZN(new_n1502_));
  INV_X1     g0860(.I(\in3[87] ), .ZN(new_n1503_));
  NOR2_X1    g0861(.A1(new_n1503_), .A2(\in2[87] ), .ZN(new_n1504_));
  AOI21_X1   g0862(.A1(new_n1502_), .A2(\in3[86] ), .B(new_n1504_), .ZN(new_n1505_));
  INV_X1     g0863(.I(new_n1505_), .ZN(new_n1506_));
  INV_X1     g0864(.I(\in3[84] ), .ZN(new_n1507_));
  NOR2_X1    g0865(.A1(new_n1507_), .A2(\in2[84] ), .ZN(new_n1508_));
  INV_X1     g0866(.I(\in3[85] ), .ZN(new_n1509_));
  NOR2_X1    g0867(.A1(new_n1509_), .A2(\in2[85] ), .ZN(new_n1510_));
  NOR3_X1    g0868(.A1(new_n1506_), .A2(new_n1508_), .A3(new_n1510_), .ZN(new_n1511_));
  INV_X1     g0869(.I(new_n1511_), .ZN(new_n1512_));
  INV_X1     g0870(.I(\in3[83] ), .ZN(new_n1513_));
  INV_X1     g0871(.I(\in2[82] ), .ZN(new_n1514_));
  INV_X1     g0872(.I(\in2[83] ), .ZN(new_n1515_));
  AOI22_X1   g0873(.A1(new_n1514_), .A2(\in3[82] ), .B1(new_n1515_), .B2(\in3[83] ), .ZN(new_n1516_));
  INV_X1     g0874(.I(\in2[81] ), .ZN(new_n1517_));
  OAI22_X1   g0875(.A1(new_n1517_), .A2(\in3[81] ), .B1(new_n1514_), .B2(\in3[82] ), .ZN(new_n1518_));
  INV_X1     g0876(.I(\in2[80] ), .ZN(new_n1519_));
  NAND2_X1   g0877(.A1(new_n1517_), .A2(\in3[81] ), .ZN(new_n1520_));
  INV_X1     g0878(.I(new_n1520_), .ZN(new_n1521_));
  NOR3_X1    g0879(.A1(new_n1521_), .A2(new_n1519_), .A3(\in3[80] ), .ZN(new_n1522_));
  OR2_X2     g0880(.A1(new_n1522_), .A2(new_n1518_), .Z(new_n1523_));
  AOI22_X1   g0881(.A1(new_n1523_), .A2(new_n1516_), .B1(\in2[83] ), .B2(new_n1513_), .ZN(new_n1524_));
  INV_X1     g0882(.I(new_n1524_), .ZN(new_n1525_));
  INV_X1     g0883(.I(\in3[79] ), .ZN(new_n1526_));
  NOR2_X1    g0884(.A1(new_n1526_), .A2(\in2[79] ), .ZN(new_n1527_));
  INV_X1     g0885(.I(new_n1527_), .ZN(new_n1528_));
  INV_X1     g0886(.I(\in2[78] ), .ZN(new_n1529_));
  AOI21_X1   g0887(.A1(new_n1529_), .A2(\in3[78] ), .B(new_n1527_), .ZN(new_n1530_));
  INV_X1     g0888(.I(\in3[77] ), .ZN(new_n1531_));
  NOR2_X1    g0889(.A1(new_n1531_), .A2(\in2[77] ), .ZN(new_n1532_));
  INV_X1     g0890(.I(\in3[76] ), .ZN(new_n1533_));
  AOI22_X1   g0891(.A1(\in2[76] ), .A2(new_n1533_), .B1(new_n1531_), .B2(\in2[77] ), .ZN(new_n1534_));
  NOR2_X1    g0892(.A1(new_n1534_), .A2(new_n1532_), .ZN(new_n1535_));
  INV_X1     g0893(.I(\in2[79] ), .ZN(new_n1536_));
  OAI22_X1   g0894(.A1(new_n1529_), .A2(\in3[78] ), .B1(new_n1536_), .B2(\in3[79] ), .ZN(new_n1537_));
  AOI22_X1   g0895(.A1(new_n1535_), .A2(new_n1530_), .B1(new_n1528_), .B2(new_n1537_), .ZN(new_n1538_));
  INV_X1     g0896(.I(new_n1530_), .ZN(new_n1539_));
  NOR2_X1    g0897(.A1(new_n1533_), .A2(\in2[76] ), .ZN(new_n1540_));
  NOR3_X1    g0898(.A1(new_n1539_), .A2(new_n1532_), .A3(new_n1540_), .ZN(new_n1541_));
  INV_X1     g0899(.I(new_n1541_), .ZN(new_n1542_));
  INV_X1     g0900(.I(\in3[73] ), .ZN(new_n1543_));
  NOR2_X1    g0901(.A1(new_n1543_), .A2(\in2[73] ), .ZN(new_n1544_));
  INV_X1     g0902(.I(\in2[74] ), .ZN(new_n1545_));
  INV_X1     g0903(.I(\in2[75] ), .ZN(new_n1546_));
  AOI22_X1   g0904(.A1(new_n1545_), .A2(\in3[74] ), .B1(new_n1546_), .B2(\in3[75] ), .ZN(new_n1547_));
  INV_X1     g0905(.I(new_n1547_), .ZN(new_n1548_));
  INV_X1     g0906(.I(\in3[72] ), .ZN(new_n1549_));
  NOR2_X1    g0907(.A1(new_n1549_), .A2(\in2[72] ), .ZN(new_n1550_));
  NOR3_X1    g0908(.A1(new_n1548_), .A2(new_n1544_), .A3(new_n1550_), .ZN(new_n1551_));
  INV_X1     g0909(.I(\in3[71] ), .ZN(new_n1552_));
  NOR2_X1    g0910(.A1(new_n1552_), .A2(\in2[71] ), .ZN(new_n1553_));
  INV_X1     g0911(.I(new_n1553_), .ZN(new_n1554_));
  INV_X1     g0912(.I(\in2[70] ), .ZN(new_n1555_));
  AOI21_X1   g0913(.A1(new_n1555_), .A2(\in3[70] ), .B(new_n1553_), .ZN(new_n1556_));
  INV_X1     g0914(.I(\in3[69] ), .ZN(new_n1557_));
  NOR2_X1    g0915(.A1(new_n1557_), .A2(\in2[69] ), .ZN(new_n1558_));
  INV_X1     g0916(.I(\in3[68] ), .ZN(new_n1559_));
  AOI22_X1   g0917(.A1(\in2[68] ), .A2(new_n1559_), .B1(new_n1557_), .B2(\in2[69] ), .ZN(new_n1560_));
  NOR2_X1    g0918(.A1(new_n1560_), .A2(new_n1558_), .ZN(new_n1561_));
  INV_X1     g0919(.I(\in2[71] ), .ZN(new_n1562_));
  OAI22_X1   g0920(.A1(new_n1555_), .A2(\in3[70] ), .B1(new_n1562_), .B2(\in3[71] ), .ZN(new_n1563_));
  AOI22_X1   g0921(.A1(new_n1561_), .A2(new_n1556_), .B1(new_n1554_), .B2(new_n1563_), .ZN(new_n1564_));
  INV_X1     g0922(.I(\in3[67] ), .ZN(new_n1565_));
  INV_X1     g0923(.I(\in2[66] ), .ZN(new_n1566_));
  INV_X1     g0924(.I(\in2[67] ), .ZN(new_n1567_));
  AOI22_X1   g0925(.A1(new_n1566_), .A2(\in3[66] ), .B1(new_n1567_), .B2(\in3[67] ), .ZN(new_n1568_));
  INV_X1     g0926(.I(\in2[65] ), .ZN(new_n1569_));
  OAI22_X1   g0927(.A1(new_n1569_), .A2(\in3[65] ), .B1(new_n1566_), .B2(\in3[66] ), .ZN(new_n1570_));
  INV_X1     g0928(.I(\in2[64] ), .ZN(new_n1571_));
  NAND2_X1   g0929(.A1(new_n1569_), .A2(\in3[65] ), .ZN(new_n1572_));
  INV_X1     g0930(.I(new_n1572_), .ZN(new_n1573_));
  NOR3_X1    g0931(.A1(new_n1573_), .A2(new_n1571_), .A3(\in3[64] ), .ZN(new_n1574_));
  OR2_X2     g0932(.A1(new_n1574_), .A2(new_n1570_), .Z(new_n1575_));
  AOI22_X1   g0933(.A1(new_n1575_), .A2(new_n1568_), .B1(\in2[67] ), .B2(new_n1565_), .ZN(new_n1576_));
  INV_X1     g0934(.I(new_n1576_), .ZN(new_n1577_));
  NAND2_X1   g0935(.A1(new_n1571_), .A2(\in3[64] ), .ZN(new_n1578_));
  NAND3_X1   g0936(.A1(new_n1568_), .A2(new_n1572_), .A3(new_n1578_), .ZN(new_n1579_));
  INV_X1     g0937(.I(new_n1579_), .ZN(new_n1580_));
  INV_X1     g0938(.I(\in2[56] ), .ZN(new_n1581_));
  INV_X1     g0939(.I(\in2[57] ), .ZN(new_n1582_));
  AOI22_X1   g0940(.A1(new_n1581_), .A2(\in3[56] ), .B1(new_n1582_), .B2(\in3[57] ), .ZN(new_n1583_));
  INV_X1     g0941(.I(\in2[62] ), .ZN(new_n1584_));
  INV_X1     g0942(.I(\in3[63] ), .ZN(new_n1585_));
  NOR2_X1    g0943(.A1(new_n1585_), .A2(\in2[63] ), .ZN(new_n1586_));
  AOI21_X1   g0944(.A1(new_n1584_), .A2(\in3[62] ), .B(new_n1586_), .ZN(new_n1587_));
  INV_X1     g0945(.I(\in2[60] ), .ZN(new_n1588_));
  NAND2_X1   g0946(.A1(new_n1588_), .A2(\in3[60] ), .ZN(new_n1589_));
  INV_X1     g0947(.I(\in2[61] ), .ZN(new_n1590_));
  NAND2_X1   g0948(.A1(new_n1590_), .A2(\in3[61] ), .ZN(new_n1591_));
  NAND3_X1   g0949(.A1(new_n1587_), .A2(new_n1589_), .A3(new_n1591_), .ZN(new_n1592_));
  INV_X1     g0950(.I(new_n1592_), .ZN(new_n1593_));
  INV_X1     g0951(.I(\in2[58] ), .ZN(new_n1594_));
  INV_X1     g0952(.I(\in2[59] ), .ZN(new_n1595_));
  AOI22_X1   g0953(.A1(new_n1594_), .A2(\in3[58] ), .B1(new_n1595_), .B2(\in3[59] ), .ZN(new_n1596_));
  NAND3_X1   g0954(.A1(new_n1593_), .A2(new_n1583_), .A3(new_n1596_), .ZN(new_n1597_));
  INV_X1     g0955(.I(\in3[53] ), .ZN(new_n1598_));
  NOR2_X1    g0956(.A1(new_n1598_), .A2(\in2[53] ), .ZN(new_n1599_));
  INV_X1     g0957(.I(\in2[54] ), .ZN(new_n1600_));
  INV_X1     g0958(.I(\in2[55] ), .ZN(new_n1601_));
  AOI22_X1   g0959(.A1(new_n1600_), .A2(\in3[54] ), .B1(new_n1601_), .B2(\in3[55] ), .ZN(new_n1602_));
  INV_X1     g0960(.I(new_n1602_), .ZN(new_n1603_));
  INV_X1     g0961(.I(\in3[52] ), .ZN(new_n1604_));
  NOR2_X1    g0962(.A1(new_n1604_), .A2(\in2[52] ), .ZN(new_n1605_));
  NOR3_X1    g0963(.A1(new_n1603_), .A2(new_n1599_), .A3(new_n1605_), .ZN(new_n1606_));
  INV_X1     g0964(.I(new_n1606_), .ZN(new_n1607_));
  INV_X1     g0965(.I(\in2[50] ), .ZN(new_n1608_));
  INV_X1     g0966(.I(\in2[51] ), .ZN(new_n1609_));
  AOI22_X1   g0967(.A1(new_n1608_), .A2(\in3[50] ), .B1(new_n1609_), .B2(\in3[51] ), .ZN(new_n1610_));
  INV_X1     g0968(.I(\in2[49] ), .ZN(new_n1611_));
  OAI22_X1   g0969(.A1(new_n1611_), .A2(\in3[49] ), .B1(new_n1608_), .B2(\in3[50] ), .ZN(new_n1612_));
  INV_X1     g0970(.I(\in2[48] ), .ZN(new_n1613_));
  INV_X1     g0971(.I(\in3[49] ), .ZN(new_n1614_));
  NOR2_X1    g0972(.A1(new_n1614_), .A2(\in2[49] ), .ZN(new_n1615_));
  NOR3_X1    g0973(.A1(new_n1615_), .A2(new_n1613_), .A3(\in3[48] ), .ZN(new_n1616_));
  OAI21_X1   g0974(.A1(new_n1616_), .A2(new_n1612_), .B(new_n1610_), .ZN(new_n1617_));
  NOR2_X1    g0975(.A1(new_n1609_), .A2(\in3[51] ), .ZN(new_n1618_));
  INV_X1     g0976(.I(new_n1618_), .ZN(new_n1619_));
  AOI21_X1   g0977(.A1(new_n1617_), .A2(new_n1619_), .B(new_n1607_), .ZN(new_n1620_));
  INV_X1     g0978(.I(\in2[53] ), .ZN(new_n1621_));
  OAI22_X1   g0979(.A1(new_n1621_), .A2(\in3[53] ), .B1(new_n1600_), .B2(\in3[54] ), .ZN(new_n1622_));
  NOR2_X1    g0980(.A1(new_n1599_), .A2(\in3[52] ), .ZN(new_n1623_));
  AOI21_X1   g0981(.A1(new_n1623_), .A2(\in2[52] ), .B(new_n1622_), .ZN(new_n1624_));
  OAI22_X1   g0982(.A1(new_n1624_), .A2(new_n1603_), .B1(new_n1601_), .B2(\in3[55] ), .ZN(new_n1625_));
  NOR2_X1    g0983(.A1(new_n1620_), .A2(new_n1625_), .ZN(new_n1626_));
  INV_X1     g0984(.I(new_n1626_), .ZN(new_n1627_));
  INV_X1     g0985(.I(\in2[46] ), .ZN(new_n1628_));
  INV_X1     g0986(.I(\in3[47] ), .ZN(new_n1629_));
  NOR2_X1    g0987(.A1(new_n1629_), .A2(\in2[47] ), .ZN(new_n1630_));
  AOI21_X1   g0988(.A1(new_n1628_), .A2(\in3[46] ), .B(new_n1630_), .ZN(new_n1631_));
  INV_X1     g0989(.I(\in2[44] ), .ZN(new_n1632_));
  NAND2_X1   g0990(.A1(new_n1632_), .A2(\in3[44] ), .ZN(new_n1633_));
  INV_X1     g0991(.I(\in2[45] ), .ZN(new_n1634_));
  NAND2_X1   g0992(.A1(new_n1634_), .A2(\in3[45] ), .ZN(new_n1635_));
  NAND3_X1   g0993(.A1(new_n1631_), .A2(new_n1633_), .A3(new_n1635_), .ZN(new_n1636_));
  INV_X1     g0994(.I(new_n1636_), .ZN(new_n1637_));
  INV_X1     g0995(.I(\in2[43] ), .ZN(new_n1638_));
  INV_X1     g0996(.I(\in2[42] ), .ZN(new_n1639_));
  AOI22_X1   g0997(.A1(new_n1639_), .A2(\in3[42] ), .B1(new_n1638_), .B2(\in3[43] ), .ZN(new_n1640_));
  INV_X1     g0998(.I(new_n1640_), .ZN(new_n1641_));
  INV_X1     g0999(.I(\in3[40] ), .ZN(new_n1642_));
  INV_X1     g1000(.I(\in2[41] ), .ZN(new_n1643_));
  OAI22_X1   g1001(.A1(new_n1643_), .A2(\in3[41] ), .B1(new_n1639_), .B2(\in3[42] ), .ZN(new_n1644_));
  INV_X1     g1002(.I(\in2[40] ), .ZN(new_n1645_));
  AOI21_X1   g1003(.A1(new_n1643_), .A2(\in3[41] ), .B(new_n1645_), .ZN(new_n1646_));
  AOI21_X1   g1004(.A1(new_n1642_), .A2(new_n1646_), .B(new_n1644_), .ZN(new_n1647_));
  OAI22_X1   g1005(.A1(new_n1647_), .A2(new_n1641_), .B1(new_n1638_), .B2(\in3[43] ), .ZN(new_n1648_));
  NAND2_X1   g1006(.A1(new_n1648_), .A2(new_n1637_), .ZN(new_n1649_));
  INV_X1     g1007(.I(new_n1630_), .ZN(new_n1650_));
  OAI22_X1   g1008(.A1(new_n1632_), .A2(\in3[44] ), .B1(new_n1634_), .B2(\in3[45] ), .ZN(new_n1651_));
  AND2_X2    g1009(.A1(new_n1651_), .A2(new_n1635_), .Z(new_n1652_));
  INV_X1     g1010(.I(\in2[47] ), .ZN(new_n1653_));
  OAI22_X1   g1011(.A1(new_n1628_), .A2(\in3[46] ), .B1(new_n1653_), .B2(\in3[47] ), .ZN(new_n1654_));
  AOI22_X1   g1012(.A1(new_n1652_), .A2(new_n1631_), .B1(new_n1650_), .B2(new_n1654_), .ZN(new_n1655_));
  AND2_X2    g1013(.A1(new_n1649_), .A2(new_n1655_), .Z(new_n1656_));
  AOI22_X1   g1014(.A1(new_n1645_), .A2(\in3[40] ), .B1(new_n1643_), .B2(\in3[41] ), .ZN(new_n1657_));
  NAND3_X1   g1015(.A1(new_n1637_), .A2(new_n1640_), .A3(new_n1657_), .ZN(new_n1658_));
  INV_X1     g1016(.I(\in2[32] ), .ZN(new_n1659_));
  INV_X1     g1017(.I(\in2[33] ), .ZN(new_n1660_));
  AOI22_X1   g1018(.A1(new_n1659_), .A2(\in3[32] ), .B1(new_n1660_), .B2(\in3[33] ), .ZN(new_n1661_));
  INV_X1     g1019(.I(\in2[38] ), .ZN(new_n1662_));
  INV_X1     g1020(.I(\in3[39] ), .ZN(new_n1663_));
  NOR2_X1    g1021(.A1(new_n1663_), .A2(\in2[39] ), .ZN(new_n1664_));
  AOI21_X1   g1022(.A1(new_n1662_), .A2(\in3[38] ), .B(new_n1664_), .ZN(new_n1665_));
  INV_X1     g1023(.I(\in2[36] ), .ZN(new_n1666_));
  NAND2_X1   g1024(.A1(new_n1666_), .A2(\in3[36] ), .ZN(new_n1667_));
  INV_X1     g1025(.I(\in2[37] ), .ZN(new_n1668_));
  NAND2_X1   g1026(.A1(new_n1668_), .A2(\in3[37] ), .ZN(new_n1669_));
  NAND3_X1   g1027(.A1(new_n1665_), .A2(new_n1667_), .A3(new_n1669_), .ZN(new_n1670_));
  INV_X1     g1028(.I(new_n1670_), .ZN(new_n1671_));
  INV_X1     g1029(.I(\in2[34] ), .ZN(new_n1672_));
  INV_X1     g1030(.I(\in2[35] ), .ZN(new_n1673_));
  AOI22_X1   g1031(.A1(new_n1672_), .A2(\in3[34] ), .B1(new_n1673_), .B2(\in3[35] ), .ZN(new_n1674_));
  NAND3_X1   g1032(.A1(new_n1671_), .A2(new_n1661_), .A3(new_n1674_), .ZN(new_n1675_));
  INV_X1     g1033(.I(new_n1675_), .ZN(new_n1676_));
  INV_X1     g1034(.I(\in2[29] ), .ZN(new_n1677_));
  NOR2_X1    g1035(.A1(new_n1677_), .A2(\in3[29] ), .ZN(new_n1678_));
  INV_X1     g1036(.I(new_n1678_), .ZN(new_n1679_));
  NAND2_X1   g1037(.A1(new_n1677_), .A2(\in3[29] ), .ZN(new_n1680_));
  INV_X1     g1038(.I(\in3[27] ), .ZN(new_n1681_));
  INV_X1     g1039(.I(\in2[26] ), .ZN(new_n1682_));
  NOR2_X1    g1040(.A1(new_n1682_), .A2(\in3[26] ), .ZN(new_n1683_));
  INV_X1     g1041(.I(new_n1683_), .ZN(new_n1684_));
  NAND2_X1   g1042(.A1(new_n1682_), .A2(\in3[26] ), .ZN(new_n1685_));
  INV_X1     g1043(.I(new_n1685_), .ZN(new_n1686_));
  INV_X1     g1044(.I(\in3[24] ), .ZN(new_n1687_));
  NOR2_X1    g1045(.A1(new_n1687_), .A2(\in2[24] ), .ZN(new_n1688_));
  INV_X1     g1046(.I(\in3[23] ), .ZN(new_n1689_));
  NOR2_X1    g1047(.A1(new_n1689_), .A2(\in2[23] ), .ZN(new_n1690_));
  INV_X1     g1048(.I(new_n1690_), .ZN(new_n1691_));
  INV_X1     g1049(.I(\in2[22] ), .ZN(new_n1692_));
  INV_X1     g1050(.I(\in3[22] ), .ZN(new_n1693_));
  INV_X1     g1051(.I(\in2[21] ), .ZN(new_n1694_));
  NOR2_X1    g1052(.A1(new_n1694_), .A2(\in3[21] ), .ZN(new_n1695_));
  NAND2_X1   g1053(.A1(new_n1694_), .A2(\in3[21] ), .ZN(new_n1696_));
  INV_X1     g1054(.I(new_n1696_), .ZN(new_n1697_));
  INV_X1     g1055(.I(\in2[19] ), .ZN(new_n1698_));
  INV_X1     g1056(.I(\in2[18] ), .ZN(new_n1699_));
  NOR2_X1    g1057(.A1(new_n1699_), .A2(\in3[18] ), .ZN(new_n1700_));
  NAND2_X1   g1058(.A1(new_n1699_), .A2(\in3[18] ), .ZN(new_n1701_));
  INV_X1     g1059(.I(\in3[16] ), .ZN(new_n1702_));
  NOR2_X1    g1060(.A1(new_n1702_), .A2(\in2[16] ), .ZN(new_n1703_));
  INV_X1     g1061(.I(new_n1703_), .ZN(new_n1704_));
  INV_X1     g1062(.I(\in3[15] ), .ZN(new_n1705_));
  NOR2_X1    g1063(.A1(new_n1705_), .A2(\in2[15] ), .ZN(new_n1706_));
  INV_X1     g1064(.I(\in2[13] ), .ZN(new_n1707_));
  NOR2_X1    g1065(.A1(new_n1707_), .A2(\in3[13] ), .ZN(new_n1708_));
  INV_X1     g1066(.I(new_n1708_), .ZN(new_n1709_));
  NAND2_X1   g1067(.A1(new_n1707_), .A2(\in3[13] ), .ZN(new_n1710_));
  INV_X1     g1068(.I(\in3[11] ), .ZN(new_n1711_));
  INV_X1     g1069(.I(\in2[10] ), .ZN(new_n1712_));
  NOR2_X1    g1070(.A1(new_n1712_), .A2(\in3[10] ), .ZN(new_n1713_));
  INV_X1     g1071(.I(new_n1713_), .ZN(new_n1714_));
  NAND2_X1   g1072(.A1(new_n1712_), .A2(\in3[10] ), .ZN(new_n1715_));
  INV_X1     g1073(.I(new_n1715_), .ZN(new_n1716_));
  INV_X1     g1074(.I(\in3[8] ), .ZN(new_n1717_));
  NOR2_X1    g1075(.A1(new_n1717_), .A2(\in2[8] ), .ZN(new_n1718_));
  INV_X1     g1076(.I(\in2[6] ), .ZN(new_n1719_));
  NOR2_X1    g1077(.A1(new_n1719_), .A2(\in3[6] ), .ZN(new_n1720_));
  INV_X1     g1078(.I(new_n1720_), .ZN(new_n1721_));
  NAND2_X1   g1079(.A1(new_n1719_), .A2(\in3[6] ), .ZN(new_n1722_));
  INV_X1     g1080(.I(\in3[4] ), .ZN(new_n1723_));
  NOR2_X1    g1081(.A1(new_n1723_), .A2(\in2[4] ), .ZN(new_n1724_));
  INV_X1     g1082(.I(\in3[3] ), .ZN(new_n1725_));
  NOR2_X1    g1083(.A1(new_n1725_), .A2(\in2[3] ), .ZN(new_n1726_));
  INV_X1     g1084(.I(new_n1726_), .ZN(new_n1727_));
  INV_X1     g1085(.I(\in3[2] ), .ZN(new_n1728_));
  INV_X1     g1086(.I(\in3[0] ), .ZN(new_n1729_));
  AOI21_X1   g1087(.A1(new_n1729_), .A2(\in2[0] ), .B(\in2[1] ), .ZN(new_n1730_));
  NAND3_X1   g1088(.A1(new_n1729_), .A2(\in2[0] ), .A3(\in2[1] ), .ZN(new_n1731_));
  AOI21_X1   g1089(.A1(\in3[1] ), .A2(new_n1731_), .B(new_n1730_), .ZN(new_n1732_));
  OAI21_X1   g1090(.A1(new_n1732_), .A2(new_n1728_), .B(\in2[2] ), .ZN(new_n1733_));
  NAND2_X1   g1091(.A1(new_n1732_), .A2(new_n1728_), .ZN(new_n1734_));
  INV_X1     g1092(.I(\in2[3] ), .ZN(new_n1735_));
  NOR2_X1    g1093(.A1(new_n1735_), .A2(\in3[3] ), .ZN(new_n1736_));
  INV_X1     g1094(.I(new_n1736_), .ZN(new_n1737_));
  NAND3_X1   g1095(.A1(new_n1733_), .A2(new_n1734_), .A3(new_n1737_), .ZN(new_n1738_));
  INV_X1     g1096(.I(\in2[4] ), .ZN(new_n1739_));
  NOR2_X1    g1097(.A1(new_n1739_), .A2(\in3[4] ), .ZN(new_n1740_));
  AOI21_X1   g1098(.A1(new_n1738_), .A2(new_n1727_), .B(new_n1740_), .ZN(new_n1741_));
  INV_X1     g1099(.I(\in3[5] ), .ZN(new_n1742_));
  NOR2_X1    g1100(.A1(new_n1742_), .A2(\in2[5] ), .ZN(new_n1743_));
  NOR3_X1    g1101(.A1(new_n1741_), .A2(new_n1724_), .A3(new_n1743_), .ZN(new_n1744_));
  INV_X1     g1102(.I(\in2[5] ), .ZN(new_n1745_));
  NOR2_X1    g1103(.A1(new_n1745_), .A2(\in3[5] ), .ZN(new_n1746_));
  OAI21_X1   g1104(.A1(new_n1744_), .A2(new_n1746_), .B(new_n1722_), .ZN(new_n1747_));
  AOI21_X1   g1105(.A1(new_n1747_), .A2(new_n1721_), .B(\in3[7] ), .ZN(new_n1748_));
  NAND3_X1   g1106(.A1(new_n1747_), .A2(\in3[7] ), .A3(new_n1721_), .ZN(new_n1749_));
  OAI21_X1   g1107(.A1(\in2[7] ), .A2(new_n1748_), .B(new_n1749_), .ZN(new_n1750_));
  INV_X1     g1108(.I(\in2[8] ), .ZN(new_n1751_));
  NOR2_X1    g1109(.A1(new_n1751_), .A2(\in3[8] ), .ZN(new_n1752_));
  INV_X1     g1110(.I(new_n1752_), .ZN(new_n1753_));
  AOI21_X1   g1111(.A1(new_n1750_), .A2(new_n1753_), .B(new_n1718_), .ZN(new_n1754_));
  INV_X1     g1112(.I(\in3[9] ), .ZN(new_n1755_));
  NOR2_X1    g1113(.A1(new_n1755_), .A2(\in2[9] ), .ZN(new_n1756_));
  INV_X1     g1114(.I(new_n1756_), .ZN(new_n1757_));
  INV_X1     g1115(.I(\in2[9] ), .ZN(new_n1758_));
  NOR2_X1    g1116(.A1(new_n1758_), .A2(\in3[9] ), .ZN(new_n1759_));
  AOI21_X1   g1117(.A1(new_n1754_), .A2(new_n1757_), .B(new_n1759_), .ZN(new_n1760_));
  OAI21_X1   g1118(.A1(new_n1760_), .A2(new_n1716_), .B(new_n1714_), .ZN(new_n1761_));
  AOI21_X1   g1119(.A1(new_n1761_), .A2(new_n1711_), .B(\in2[11] ), .ZN(new_n1762_));
  NOR2_X1    g1120(.A1(new_n1761_), .A2(new_n1711_), .ZN(new_n1763_));
  INV_X1     g1121(.I(\in3[12] ), .ZN(new_n1764_));
  NOR2_X1    g1122(.A1(new_n1764_), .A2(\in2[12] ), .ZN(new_n1765_));
  NOR3_X1    g1123(.A1(new_n1762_), .A2(new_n1763_), .A3(new_n1765_), .ZN(new_n1766_));
  INV_X1     g1124(.I(\in2[12] ), .ZN(new_n1767_));
  NOR2_X1    g1125(.A1(new_n1767_), .A2(\in3[12] ), .ZN(new_n1768_));
  OAI21_X1   g1126(.A1(new_n1766_), .A2(new_n1768_), .B(new_n1710_), .ZN(new_n1769_));
  AOI21_X1   g1127(.A1(new_n1769_), .A2(new_n1709_), .B(\in3[14] ), .ZN(new_n1770_));
  NAND3_X1   g1128(.A1(new_n1769_), .A2(\in3[14] ), .A3(new_n1709_), .ZN(new_n1771_));
  OAI21_X1   g1129(.A1(\in2[14] ), .A2(new_n1770_), .B(new_n1771_), .ZN(new_n1772_));
  INV_X1     g1130(.I(\in2[15] ), .ZN(new_n1773_));
  NOR2_X1    g1131(.A1(new_n1773_), .A2(\in3[15] ), .ZN(new_n1774_));
  INV_X1     g1132(.I(new_n1774_), .ZN(new_n1775_));
  AOI21_X1   g1133(.A1(new_n1772_), .A2(new_n1775_), .B(new_n1706_), .ZN(new_n1776_));
  INV_X1     g1134(.I(\in2[16] ), .ZN(new_n1777_));
  NOR2_X1    g1135(.A1(new_n1777_), .A2(\in3[16] ), .ZN(new_n1778_));
  OAI21_X1   g1136(.A1(new_n1776_), .A2(new_n1778_), .B(new_n1704_), .ZN(new_n1779_));
  INV_X1     g1137(.I(\in3[17] ), .ZN(new_n1780_));
  NOR2_X1    g1138(.A1(new_n1780_), .A2(\in2[17] ), .ZN(new_n1781_));
  INV_X1     g1139(.I(\in2[17] ), .ZN(new_n1782_));
  NOR2_X1    g1140(.A1(new_n1782_), .A2(\in3[17] ), .ZN(new_n1783_));
  INV_X1     g1141(.I(new_n1783_), .ZN(new_n1784_));
  OAI21_X1   g1142(.A1(new_n1779_), .A2(new_n1781_), .B(new_n1784_), .ZN(new_n1785_));
  AOI21_X1   g1143(.A1(new_n1785_), .A2(new_n1701_), .B(new_n1700_), .ZN(new_n1786_));
  OAI21_X1   g1144(.A1(new_n1786_), .A2(\in3[19] ), .B(new_n1698_), .ZN(new_n1787_));
  NAND2_X1   g1145(.A1(new_n1786_), .A2(\in3[19] ), .ZN(new_n1788_));
  INV_X1     g1146(.I(\in3[20] ), .ZN(new_n1789_));
  NOR2_X1    g1147(.A1(new_n1789_), .A2(\in2[20] ), .ZN(new_n1790_));
  INV_X1     g1148(.I(new_n1790_), .ZN(new_n1791_));
  NAND3_X1   g1149(.A1(new_n1787_), .A2(new_n1788_), .A3(new_n1791_), .ZN(new_n1792_));
  INV_X1     g1150(.I(\in2[20] ), .ZN(new_n1793_));
  NOR2_X1    g1151(.A1(new_n1793_), .A2(\in3[20] ), .ZN(new_n1794_));
  INV_X1     g1152(.I(new_n1794_), .ZN(new_n1795_));
  AOI21_X1   g1153(.A1(new_n1792_), .A2(new_n1795_), .B(new_n1697_), .ZN(new_n1796_));
  OAI21_X1   g1154(.A1(new_n1796_), .A2(new_n1695_), .B(new_n1693_), .ZN(new_n1797_));
  NOR3_X1    g1155(.A1(new_n1796_), .A2(new_n1693_), .A3(new_n1695_), .ZN(new_n1798_));
  AOI21_X1   g1156(.A1(new_n1692_), .A2(new_n1797_), .B(new_n1798_), .ZN(new_n1799_));
  INV_X1     g1157(.I(\in2[23] ), .ZN(new_n1800_));
  NOR2_X1    g1158(.A1(new_n1800_), .A2(\in3[23] ), .ZN(new_n1801_));
  OAI21_X1   g1159(.A1(new_n1799_), .A2(new_n1801_), .B(new_n1691_), .ZN(new_n1802_));
  INV_X1     g1160(.I(\in2[24] ), .ZN(new_n1803_));
  NOR2_X1    g1161(.A1(new_n1803_), .A2(\in3[24] ), .ZN(new_n1804_));
  INV_X1     g1162(.I(new_n1804_), .ZN(new_n1805_));
  AOI21_X1   g1163(.A1(new_n1802_), .A2(new_n1805_), .B(new_n1688_), .ZN(new_n1806_));
  INV_X1     g1164(.I(\in3[25] ), .ZN(new_n1807_));
  NOR2_X1    g1165(.A1(new_n1807_), .A2(\in2[25] ), .ZN(new_n1808_));
  INV_X1     g1166(.I(new_n1808_), .ZN(new_n1809_));
  INV_X1     g1167(.I(\in2[25] ), .ZN(new_n1810_));
  NOR2_X1    g1168(.A1(new_n1810_), .A2(\in3[25] ), .ZN(new_n1811_));
  AOI21_X1   g1169(.A1(new_n1806_), .A2(new_n1809_), .B(new_n1811_), .ZN(new_n1812_));
  OAI21_X1   g1170(.A1(new_n1812_), .A2(new_n1686_), .B(new_n1684_), .ZN(new_n1813_));
  AOI21_X1   g1171(.A1(new_n1813_), .A2(new_n1681_), .B(\in2[27] ), .ZN(new_n1814_));
  NOR2_X1    g1172(.A1(new_n1813_), .A2(new_n1681_), .ZN(new_n1815_));
  INV_X1     g1173(.I(\in3[28] ), .ZN(new_n1816_));
  NOR2_X1    g1174(.A1(new_n1816_), .A2(\in2[28] ), .ZN(new_n1817_));
  NOR3_X1    g1175(.A1(new_n1814_), .A2(new_n1815_), .A3(new_n1817_), .ZN(new_n1818_));
  INV_X1     g1176(.I(\in2[28] ), .ZN(new_n1819_));
  NOR2_X1    g1177(.A1(new_n1819_), .A2(\in3[28] ), .ZN(new_n1820_));
  OAI21_X1   g1178(.A1(new_n1818_), .A2(new_n1820_), .B(new_n1680_), .ZN(new_n1821_));
  AOI21_X1   g1179(.A1(new_n1821_), .A2(new_n1679_), .B(\in3[30] ), .ZN(new_n1822_));
  NAND3_X1   g1180(.A1(new_n1821_), .A2(\in3[30] ), .A3(new_n1679_), .ZN(new_n1823_));
  OAI21_X1   g1181(.A1(\in2[30] ), .A2(new_n1822_), .B(new_n1823_), .ZN(new_n1824_));
  INV_X1     g1182(.I(\in3[31] ), .ZN(new_n1825_));
  NOR2_X1    g1183(.A1(new_n1825_), .A2(\in2[31] ), .ZN(new_n1826_));
  INV_X1     g1184(.I(\in2[31] ), .ZN(new_n1827_));
  NOR2_X1    g1185(.A1(new_n1827_), .A2(\in3[31] ), .ZN(new_n1828_));
  INV_X1     g1186(.I(new_n1828_), .ZN(new_n1829_));
  OAI21_X1   g1187(.A1(new_n1824_), .A2(new_n1826_), .B(new_n1829_), .ZN(new_n1830_));
  INV_X1     g1188(.I(new_n1674_), .ZN(new_n1831_));
  INV_X1     g1189(.I(\in3[32] ), .ZN(new_n1832_));
  OAI22_X1   g1190(.A1(new_n1660_), .A2(\in3[33] ), .B1(new_n1672_), .B2(\in3[34] ), .ZN(new_n1833_));
  AOI21_X1   g1191(.A1(new_n1660_), .A2(\in3[33] ), .B(new_n1659_), .ZN(new_n1834_));
  AOI21_X1   g1192(.A1(new_n1832_), .A2(new_n1834_), .B(new_n1833_), .ZN(new_n1835_));
  OAI22_X1   g1193(.A1(new_n1835_), .A2(new_n1831_), .B1(new_n1673_), .B2(\in3[35] ), .ZN(new_n1836_));
  NAND2_X1   g1194(.A1(new_n1836_), .A2(new_n1671_), .ZN(new_n1837_));
  INV_X1     g1195(.I(new_n1664_), .ZN(new_n1838_));
  OAI22_X1   g1196(.A1(new_n1666_), .A2(\in3[36] ), .B1(new_n1668_), .B2(\in3[37] ), .ZN(new_n1839_));
  AND2_X2    g1197(.A1(new_n1839_), .A2(new_n1669_), .Z(new_n1840_));
  INV_X1     g1198(.I(\in2[39] ), .ZN(new_n1841_));
  OAI22_X1   g1199(.A1(new_n1662_), .A2(\in3[38] ), .B1(new_n1841_), .B2(\in3[39] ), .ZN(new_n1842_));
  AOI22_X1   g1200(.A1(new_n1840_), .A2(new_n1665_), .B1(new_n1838_), .B2(new_n1842_), .ZN(new_n1843_));
  AND2_X2    g1201(.A1(new_n1837_), .A2(new_n1843_), .Z(new_n1844_));
  INV_X1     g1202(.I(new_n1844_), .ZN(new_n1845_));
  AOI21_X1   g1203(.A1(new_n1830_), .A2(new_n1676_), .B(new_n1845_), .ZN(new_n1846_));
  OAI21_X1   g1204(.A1(new_n1846_), .A2(new_n1658_), .B(new_n1656_), .ZN(new_n1847_));
  AOI21_X1   g1205(.A1(new_n1613_), .A2(\in3[48] ), .B(new_n1615_), .ZN(new_n1848_));
  NAND3_X1   g1206(.A1(new_n1606_), .A2(new_n1610_), .A3(new_n1848_), .ZN(new_n1849_));
  INV_X1     g1207(.I(new_n1849_), .ZN(new_n1850_));
  AOI21_X1   g1208(.A1(new_n1847_), .A2(new_n1850_), .B(new_n1627_), .ZN(new_n1851_));
  INV_X1     g1209(.I(new_n1596_), .ZN(new_n1852_));
  INV_X1     g1210(.I(\in3[56] ), .ZN(new_n1853_));
  OAI22_X1   g1211(.A1(new_n1582_), .A2(\in3[57] ), .B1(new_n1594_), .B2(\in3[58] ), .ZN(new_n1854_));
  AOI21_X1   g1212(.A1(new_n1582_), .A2(\in3[57] ), .B(new_n1581_), .ZN(new_n1855_));
  AOI21_X1   g1213(.A1(new_n1853_), .A2(new_n1855_), .B(new_n1854_), .ZN(new_n1856_));
  OAI22_X1   g1214(.A1(new_n1856_), .A2(new_n1852_), .B1(new_n1595_), .B2(\in3[59] ), .ZN(new_n1857_));
  NAND2_X1   g1215(.A1(new_n1857_), .A2(new_n1593_), .ZN(new_n1858_));
  INV_X1     g1216(.I(new_n1586_), .ZN(new_n1859_));
  OAI22_X1   g1217(.A1(new_n1588_), .A2(\in3[60] ), .B1(new_n1590_), .B2(\in3[61] ), .ZN(new_n1860_));
  AND2_X2    g1218(.A1(new_n1860_), .A2(new_n1591_), .Z(new_n1861_));
  INV_X1     g1219(.I(\in2[63] ), .ZN(new_n1862_));
  OAI22_X1   g1220(.A1(new_n1584_), .A2(\in3[62] ), .B1(new_n1862_), .B2(\in3[63] ), .ZN(new_n1863_));
  AOI22_X1   g1221(.A1(new_n1861_), .A2(new_n1587_), .B1(new_n1859_), .B2(new_n1863_), .ZN(new_n1864_));
  AND2_X2    g1222(.A1(new_n1858_), .A2(new_n1864_), .Z(new_n1865_));
  OAI21_X1   g1223(.A1(new_n1851_), .A2(new_n1597_), .B(new_n1865_), .ZN(new_n1866_));
  AOI21_X1   g1224(.A1(new_n1866_), .A2(new_n1580_), .B(new_n1577_), .ZN(new_n1867_));
  INV_X1     g1225(.I(new_n1556_), .ZN(new_n1868_));
  NOR2_X1    g1226(.A1(new_n1559_), .A2(\in2[68] ), .ZN(new_n1869_));
  NOR3_X1    g1227(.A1(new_n1868_), .A2(new_n1558_), .A3(new_n1869_), .ZN(new_n1870_));
  INV_X1     g1228(.I(new_n1870_), .ZN(new_n1871_));
  OAI21_X1   g1229(.A1(new_n1867_), .A2(new_n1871_), .B(new_n1564_), .ZN(new_n1872_));
  INV_X1     g1230(.I(\in3[75] ), .ZN(new_n1873_));
  INV_X1     g1231(.I(\in2[73] ), .ZN(new_n1874_));
  OAI22_X1   g1232(.A1(new_n1874_), .A2(\in3[73] ), .B1(new_n1545_), .B2(\in3[74] ), .ZN(new_n1875_));
  INV_X1     g1233(.I(new_n1875_), .ZN(new_n1876_));
  NAND2_X1   g1234(.A1(new_n1549_), .A2(\in2[72] ), .ZN(new_n1877_));
  OAI21_X1   g1235(.A1(new_n1544_), .A2(new_n1877_), .B(new_n1876_), .ZN(new_n1878_));
  AOI22_X1   g1236(.A1(new_n1878_), .A2(new_n1547_), .B1(\in2[75] ), .B2(new_n1873_), .ZN(new_n1879_));
  INV_X1     g1237(.I(new_n1879_), .ZN(new_n1880_));
  AOI21_X1   g1238(.A1(new_n1872_), .A2(new_n1551_), .B(new_n1880_), .ZN(new_n1881_));
  OAI21_X1   g1239(.A1(new_n1881_), .A2(new_n1542_), .B(new_n1538_), .ZN(new_n1882_));
  NAND2_X1   g1240(.A1(new_n1519_), .A2(\in3[80] ), .ZN(new_n1883_));
  NAND3_X1   g1241(.A1(new_n1516_), .A2(new_n1520_), .A3(new_n1883_), .ZN(new_n1884_));
  INV_X1     g1242(.I(new_n1884_), .ZN(new_n1885_));
  AOI21_X1   g1243(.A1(new_n1882_), .A2(new_n1885_), .B(new_n1525_), .ZN(new_n1886_));
  INV_X1     g1244(.I(new_n1504_), .ZN(new_n1887_));
  AOI22_X1   g1245(.A1(\in2[84] ), .A2(new_n1507_), .B1(new_n1509_), .B2(\in2[85] ), .ZN(new_n1888_));
  NOR2_X1    g1246(.A1(new_n1888_), .A2(new_n1510_), .ZN(new_n1889_));
  INV_X1     g1247(.I(\in2[87] ), .ZN(new_n1890_));
  OAI22_X1   g1248(.A1(new_n1502_), .A2(\in3[86] ), .B1(new_n1890_), .B2(\in3[87] ), .ZN(new_n1891_));
  AOI22_X1   g1249(.A1(new_n1889_), .A2(new_n1505_), .B1(new_n1887_), .B2(new_n1891_), .ZN(new_n1892_));
  OAI21_X1   g1250(.A1(new_n1886_), .A2(new_n1512_), .B(new_n1892_), .ZN(new_n1893_));
  AOI21_X1   g1251(.A1(new_n1893_), .A2(new_n1501_), .B(new_n1498_), .ZN(new_n1894_));
  INV_X1     g1252(.I(new_n1477_), .ZN(new_n1895_));
  NOR2_X1    g1253(.A1(new_n1480_), .A2(\in2[92] ), .ZN(new_n1896_));
  NOR3_X1    g1254(.A1(new_n1895_), .A2(new_n1479_), .A3(new_n1896_), .ZN(new_n1897_));
  INV_X1     g1255(.I(new_n1897_), .ZN(new_n1898_));
  OAI21_X1   g1256(.A1(new_n1894_), .A2(new_n1898_), .B(new_n1485_), .ZN(new_n1899_));
  INV_X1     g1257(.I(\in3[99] ), .ZN(new_n1900_));
  INV_X1     g1258(.I(\in2[97] ), .ZN(new_n1901_));
  OAI22_X1   g1259(.A1(new_n1901_), .A2(\in3[97] ), .B1(new_n1466_), .B2(\in3[98] ), .ZN(new_n1902_));
  INV_X1     g1260(.I(new_n1902_), .ZN(new_n1903_));
  NAND2_X1   g1261(.A1(new_n1470_), .A2(\in2[96] ), .ZN(new_n1904_));
  OAI21_X1   g1262(.A1(new_n1465_), .A2(new_n1904_), .B(new_n1903_), .ZN(new_n1905_));
  AOI22_X1   g1263(.A1(new_n1905_), .A2(new_n1468_), .B1(\in2[99] ), .B2(new_n1900_), .ZN(new_n1906_));
  INV_X1     g1264(.I(new_n1906_), .ZN(new_n1907_));
  AOI21_X1   g1265(.A1(new_n1899_), .A2(new_n1472_), .B(new_n1907_), .ZN(new_n1908_));
  OAI21_X1   g1266(.A1(new_n1908_), .A2(new_n1463_), .B(new_n1459_), .ZN(new_n1909_));
  NAND2_X1   g1267(.A1(new_n1440_), .A2(\in3[104] ), .ZN(new_n1910_));
  NAND3_X1   g1268(.A1(new_n1437_), .A2(new_n1441_), .A3(new_n1910_), .ZN(new_n1911_));
  INV_X1     g1269(.I(new_n1911_), .ZN(new_n1912_));
  AOI21_X1   g1270(.A1(new_n1909_), .A2(new_n1912_), .B(new_n1446_), .ZN(new_n1913_));
  INV_X1     g1271(.I(new_n1425_), .ZN(new_n1914_));
  AOI22_X1   g1272(.A1(\in2[108] ), .A2(new_n1428_), .B1(new_n1430_), .B2(\in2[109] ), .ZN(new_n1915_));
  NOR2_X1    g1273(.A1(new_n1915_), .A2(new_n1431_), .ZN(new_n1916_));
  INV_X1     g1274(.I(\in2[111] ), .ZN(new_n1917_));
  OAI22_X1   g1275(.A1(new_n1423_), .A2(\in3[110] ), .B1(new_n1917_), .B2(\in3[111] ), .ZN(new_n1918_));
  AOI22_X1   g1276(.A1(new_n1916_), .A2(new_n1426_), .B1(new_n1914_), .B2(new_n1918_), .ZN(new_n1919_));
  OAI21_X1   g1277(.A1(new_n1913_), .A2(new_n1433_), .B(new_n1919_), .ZN(new_n1920_));
  AOI21_X1   g1278(.A1(new_n1920_), .A2(new_n1422_), .B(new_n1419_), .ZN(new_n1921_));
  INV_X1     g1279(.I(new_n1398_), .ZN(new_n1922_));
  NOR2_X1    g1280(.A1(new_n1401_), .A2(\in2[116] ), .ZN(new_n1923_));
  NOR3_X1    g1281(.A1(new_n1922_), .A2(new_n1400_), .A3(new_n1923_), .ZN(new_n1924_));
  INV_X1     g1282(.I(new_n1924_), .ZN(new_n1925_));
  OAI21_X1   g1283(.A1(new_n1921_), .A2(new_n1925_), .B(new_n1406_), .ZN(new_n1926_));
  INV_X1     g1284(.I(\in3[123] ), .ZN(new_n1927_));
  INV_X1     g1285(.I(\in2[121] ), .ZN(new_n1928_));
  OAI22_X1   g1286(.A1(new_n1928_), .A2(\in3[121] ), .B1(new_n1387_), .B2(\in3[122] ), .ZN(new_n1929_));
  INV_X1     g1287(.I(new_n1929_), .ZN(new_n1930_));
  NAND2_X1   g1288(.A1(new_n1391_), .A2(\in2[120] ), .ZN(new_n1931_));
  OAI21_X1   g1289(.A1(new_n1386_), .A2(new_n1931_), .B(new_n1930_), .ZN(new_n1932_));
  AOI22_X1   g1290(.A1(new_n1932_), .A2(new_n1389_), .B1(\in2[123] ), .B2(new_n1927_), .ZN(new_n1933_));
  INV_X1     g1291(.I(new_n1933_), .ZN(new_n1934_));
  AOI21_X1   g1292(.A1(new_n1926_), .A2(new_n1393_), .B(new_n1934_), .ZN(new_n1935_));
  OAI21_X1   g1293(.A1(new_n1935_), .A2(new_n1384_), .B(new_n1379_), .ZN(new_n1936_));
  OAI21_X1   g1294(.A1(new_n1936_), .A2(\in3[127] ), .B(\in2[127] ), .ZN(new_n1937_));
  NOR2_X1    g1295(.A1(new_n1367_), .A2(new_n1937_), .ZN(new_n1938_));
  NAND2_X1   g1296(.A1(new_n1367_), .A2(new_n1937_), .ZN(new_n1939_));
  INV_X1     g1297(.I(new_n1939_), .ZN(new_n1940_));
  INV_X1     g1298(.I(new_n1393_), .ZN(new_n1941_));
  INV_X1     g1299(.I(new_n1472_), .ZN(new_n1942_));
  INV_X1     g1300(.I(new_n1551_), .ZN(new_n1943_));
  INV_X1     g1301(.I(new_n1597_), .ZN(new_n1944_));
  INV_X1     g1302(.I(new_n1658_), .ZN(new_n1945_));
  INV_X1     g1303(.I(\in2[30] ), .ZN(new_n1946_));
  INV_X1     g1304(.I(new_n1695_), .ZN(new_n1947_));
  INV_X1     g1305(.I(\in3[19] ), .ZN(new_n1948_));
  INV_X1     g1306(.I(new_n1701_), .ZN(new_n1949_));
  INV_X1     g1307(.I(\in2[14] ), .ZN(new_n1950_));
  INV_X1     g1308(.I(\in2[7] ), .ZN(new_n1951_));
  INV_X1     g1309(.I(new_n1724_), .ZN(new_n1952_));
  INV_X1     g1310(.I(\in3[1] ), .ZN(new_n1953_));
  INV_X1     g1311(.I(\in2[0] ), .ZN(new_n1954_));
  NOR2_X1    g1312(.A1(new_n1954_), .A2(\in3[0] ), .ZN(new_n1955_));
  AOI21_X1   g1313(.A1(new_n1955_), .A2(\in2[1] ), .B(new_n1953_), .ZN(new_n1956_));
  OAI21_X1   g1314(.A1(new_n1956_), .A2(new_n1730_), .B(\in3[2] ), .ZN(new_n1957_));
  NOR3_X1    g1315(.A1(new_n1956_), .A2(\in3[2] ), .A3(new_n1730_), .ZN(new_n1958_));
  AOI21_X1   g1316(.A1(\in2[2] ), .A2(new_n1957_), .B(new_n1958_), .ZN(new_n1959_));
  AOI21_X1   g1317(.A1(new_n1959_), .A2(new_n1737_), .B(new_n1726_), .ZN(new_n1960_));
  OAI21_X1   g1318(.A1(new_n1960_), .A2(new_n1740_), .B(new_n1952_), .ZN(new_n1961_));
  INV_X1     g1319(.I(new_n1746_), .ZN(new_n1962_));
  OAI21_X1   g1320(.A1(new_n1961_), .A2(new_n1743_), .B(new_n1962_), .ZN(new_n1963_));
  AOI21_X1   g1321(.A1(new_n1963_), .A2(new_n1722_), .B(new_n1720_), .ZN(new_n1964_));
  OAI21_X1   g1322(.A1(new_n1964_), .A2(\in3[7] ), .B(new_n1951_), .ZN(new_n1965_));
  AOI21_X1   g1323(.A1(new_n1965_), .A2(new_n1749_), .B(new_n1752_), .ZN(new_n1966_));
  NOR3_X1    g1324(.A1(new_n1966_), .A2(new_n1718_), .A3(new_n1756_), .ZN(new_n1967_));
  OAI21_X1   g1325(.A1(new_n1967_), .A2(new_n1759_), .B(new_n1715_), .ZN(new_n1968_));
  AOI21_X1   g1326(.A1(new_n1968_), .A2(new_n1714_), .B(\in3[11] ), .ZN(new_n1969_));
  NAND3_X1   g1327(.A1(new_n1968_), .A2(\in3[11] ), .A3(new_n1714_), .ZN(new_n1970_));
  OAI21_X1   g1328(.A1(\in2[11] ), .A2(new_n1969_), .B(new_n1970_), .ZN(new_n1971_));
  INV_X1     g1329(.I(new_n1768_), .ZN(new_n1972_));
  OAI21_X1   g1330(.A1(new_n1971_), .A2(new_n1765_), .B(new_n1972_), .ZN(new_n1973_));
  AOI21_X1   g1331(.A1(new_n1973_), .A2(new_n1710_), .B(new_n1708_), .ZN(new_n1974_));
  OAI21_X1   g1332(.A1(new_n1974_), .A2(\in3[14] ), .B(new_n1950_), .ZN(new_n1975_));
  AOI21_X1   g1333(.A1(new_n1975_), .A2(new_n1771_), .B(new_n1774_), .ZN(new_n1976_));
  INV_X1     g1334(.I(new_n1778_), .ZN(new_n1977_));
  OAI21_X1   g1335(.A1(new_n1976_), .A2(new_n1706_), .B(new_n1977_), .ZN(new_n1978_));
  INV_X1     g1336(.I(new_n1781_), .ZN(new_n1979_));
  NAND3_X1   g1337(.A1(new_n1978_), .A2(new_n1704_), .A3(new_n1979_), .ZN(new_n1980_));
  AOI21_X1   g1338(.A1(new_n1980_), .A2(new_n1784_), .B(new_n1949_), .ZN(new_n1981_));
  OAI21_X1   g1339(.A1(new_n1981_), .A2(new_n1700_), .B(new_n1948_), .ZN(new_n1982_));
  NOR3_X1    g1340(.A1(new_n1981_), .A2(new_n1948_), .A3(new_n1700_), .ZN(new_n1983_));
  AOI21_X1   g1341(.A1(new_n1698_), .A2(new_n1982_), .B(new_n1983_), .ZN(new_n1984_));
  AOI21_X1   g1342(.A1(new_n1984_), .A2(new_n1791_), .B(new_n1794_), .ZN(new_n1985_));
  OAI21_X1   g1343(.A1(new_n1985_), .A2(new_n1697_), .B(new_n1947_), .ZN(new_n1986_));
  AOI21_X1   g1344(.A1(new_n1986_), .A2(new_n1693_), .B(\in2[22] ), .ZN(new_n1987_));
  INV_X1     g1345(.I(new_n1801_), .ZN(new_n1988_));
  OAI21_X1   g1346(.A1(new_n1987_), .A2(new_n1798_), .B(new_n1988_), .ZN(new_n1989_));
  AOI21_X1   g1347(.A1(new_n1989_), .A2(new_n1691_), .B(new_n1804_), .ZN(new_n1990_));
  NOR3_X1    g1348(.A1(new_n1990_), .A2(new_n1688_), .A3(new_n1808_), .ZN(new_n1991_));
  OAI21_X1   g1349(.A1(new_n1991_), .A2(new_n1811_), .B(new_n1685_), .ZN(new_n1992_));
  AOI21_X1   g1350(.A1(new_n1992_), .A2(new_n1684_), .B(\in3[27] ), .ZN(new_n1993_));
  NAND3_X1   g1351(.A1(new_n1992_), .A2(\in3[27] ), .A3(new_n1684_), .ZN(new_n1994_));
  OAI21_X1   g1352(.A1(\in2[27] ), .A2(new_n1993_), .B(new_n1994_), .ZN(new_n1995_));
  INV_X1     g1353(.I(new_n1820_), .ZN(new_n1996_));
  OAI21_X1   g1354(.A1(new_n1995_), .A2(new_n1817_), .B(new_n1996_), .ZN(new_n1997_));
  AOI21_X1   g1355(.A1(new_n1997_), .A2(new_n1680_), .B(new_n1678_), .ZN(new_n1998_));
  OAI21_X1   g1356(.A1(new_n1998_), .A2(\in3[30] ), .B(new_n1946_), .ZN(new_n1999_));
  INV_X1     g1357(.I(new_n1826_), .ZN(new_n2000_));
  NAND3_X1   g1358(.A1(new_n1999_), .A2(new_n1823_), .A3(new_n2000_), .ZN(new_n2001_));
  AOI21_X1   g1359(.A1(new_n2001_), .A2(new_n1829_), .B(new_n1675_), .ZN(new_n2002_));
  OAI21_X1   g1360(.A1(new_n2002_), .A2(new_n1845_), .B(new_n1945_), .ZN(new_n2003_));
  AOI21_X1   g1361(.A1(new_n2003_), .A2(new_n1656_), .B(new_n1849_), .ZN(new_n2004_));
  OAI21_X1   g1362(.A1(new_n2004_), .A2(new_n1627_), .B(new_n1944_), .ZN(new_n2005_));
  AOI21_X1   g1363(.A1(new_n2005_), .A2(new_n1865_), .B(new_n1579_), .ZN(new_n2006_));
  OAI21_X1   g1364(.A1(new_n2006_), .A2(new_n1577_), .B(new_n1870_), .ZN(new_n2007_));
  AOI21_X1   g1365(.A1(new_n2007_), .A2(new_n1564_), .B(new_n1943_), .ZN(new_n2008_));
  OAI21_X1   g1366(.A1(new_n2008_), .A2(new_n1880_), .B(new_n1541_), .ZN(new_n2009_));
  AOI21_X1   g1367(.A1(new_n2009_), .A2(new_n1538_), .B(new_n1884_), .ZN(new_n2010_));
  OAI21_X1   g1368(.A1(new_n2010_), .A2(new_n1525_), .B(new_n1511_), .ZN(new_n2011_));
  AOI21_X1   g1369(.A1(new_n2011_), .A2(new_n1892_), .B(new_n1500_), .ZN(new_n2012_));
  OAI21_X1   g1370(.A1(new_n2012_), .A2(new_n1498_), .B(new_n1897_), .ZN(new_n2013_));
  AOI21_X1   g1371(.A1(new_n2013_), .A2(new_n1485_), .B(new_n1942_), .ZN(new_n2014_));
  OAI21_X1   g1372(.A1(new_n2014_), .A2(new_n1907_), .B(new_n1462_), .ZN(new_n2015_));
  AOI21_X1   g1373(.A1(new_n2015_), .A2(new_n1459_), .B(new_n1911_), .ZN(new_n2016_));
  OAI21_X1   g1374(.A1(new_n2016_), .A2(new_n1446_), .B(new_n1432_), .ZN(new_n2017_));
  AOI21_X1   g1375(.A1(new_n2017_), .A2(new_n1919_), .B(new_n1421_), .ZN(new_n2018_));
  OAI21_X1   g1376(.A1(new_n2018_), .A2(new_n1419_), .B(new_n1924_), .ZN(new_n2019_));
  AOI21_X1   g1377(.A1(new_n2019_), .A2(new_n1406_), .B(new_n1941_), .ZN(new_n2020_));
  OAI21_X1   g1378(.A1(new_n2020_), .A2(new_n1934_), .B(new_n1383_), .ZN(new_n2021_));
  NAND2_X1   g1379(.A1(new_n1368_), .A2(\in3[127] ), .ZN(new_n2022_));
  NAND3_X1   g1380(.A1(new_n2021_), .A2(new_n1379_), .A3(new_n2022_), .ZN(new_n2023_));
  NOR2_X1    g1381(.A1(new_n2023_), .A2(\in3[126] ), .ZN(new_n2024_));
  AOI21_X1   g1382(.A1(new_n1371_), .A2(new_n2023_), .B(new_n2024_), .ZN(new_n2025_));
  INV_X1     g1383(.I(new_n2025_), .ZN(new_n2026_));
  NAND2_X1   g1384(.A1(new_n1336_), .A2(new_n1245_), .ZN(new_n2027_));
  NAND3_X1   g1385(.A1(new_n2027_), .A2(new_n1118_), .A3(new_n1339_), .ZN(new_n2028_));
  AOI21_X1   g1386(.A1(new_n2028_), .A2(new_n1124_), .B(new_n961_), .ZN(new_n2029_));
  OAI21_X1   g1387(.A1(new_n2029_), .A2(new_n1142_), .B(new_n1244_), .ZN(new_n2030_));
  AOI21_X1   g1388(.A1(new_n2030_), .A2(new_n943_), .B(new_n1146_), .ZN(new_n2031_));
  OAI21_X1   g1389(.A1(new_n2031_), .A2(new_n913_), .B(new_n1242_), .ZN(new_n2032_));
  AOI21_X1   g1390(.A1(new_n2032_), .A2(new_n1164_), .B(new_n1241_), .ZN(new_n2033_));
  OAI21_X1   g1391(.A1(new_n2033_), .A2(new_n862_), .B(new_n1168_), .ZN(new_n2034_));
  AOI21_X1   g1392(.A1(new_n2034_), .A2(new_n849_), .B(new_n1240_), .ZN(new_n2035_));
  OAI21_X1   g1393(.A1(new_n2035_), .A2(new_n1177_), .B(new_n824_), .ZN(new_n2036_));
  AOI21_X1   g1394(.A1(new_n2036_), .A2(new_n822_), .B(new_n1350_), .ZN(new_n2037_));
  OAI21_X1   g1395(.A1(new_n2037_), .A2(new_n807_), .B(new_n793_), .ZN(new_n2038_));
  AOI21_X1   g1396(.A1(new_n2038_), .A2(new_n1190_), .B(new_n1239_), .ZN(new_n2039_));
  OAI21_X1   g1397(.A1(new_n2039_), .A2(new_n780_), .B(new_n1194_), .ZN(new_n2040_));
  AOI21_X1   g1398(.A1(new_n2040_), .A2(new_n767_), .B(new_n1238_), .ZN(new_n2041_));
  OAI21_X1   g1399(.A1(new_n2041_), .A2(new_n1203_), .B(new_n742_), .ZN(new_n2042_));
  AOI21_X1   g1400(.A1(new_n2042_), .A2(new_n740_), .B(new_n1357_), .ZN(new_n2043_));
  OAI21_X1   g1401(.A1(new_n2043_), .A2(new_n725_), .B(new_n711_), .ZN(new_n2044_));
  AOI21_X1   g1402(.A1(new_n2044_), .A2(new_n1216_), .B(new_n1237_), .ZN(new_n2045_));
  OAI21_X1   g1403(.A1(new_n2045_), .A2(new_n698_), .B(new_n1220_), .ZN(new_n2046_));
  AOI21_X1   g1404(.A1(new_n2046_), .A2(new_n685_), .B(new_n1236_), .ZN(new_n2047_));
  OAI21_X1   g1405(.A1(new_n2047_), .A2(new_n1229_), .B(new_n660_), .ZN(new_n2048_));
  NAND3_X1   g1406(.A1(new_n2048_), .A2(new_n657_), .A3(new_n1232_), .ZN(new_n2049_));
  NOR2_X1    g1407(.A1(new_n2049_), .A2(\in1[126] ), .ZN(new_n2050_));
  AOI21_X1   g1408(.A1(new_n647_), .A2(new_n2049_), .B(new_n2050_), .ZN(new_n2051_));
  INV_X1     g1409(.I(new_n2051_), .ZN(new_n2052_));
  NOR2_X1    g1410(.A1(new_n2023_), .A2(\in3[125] ), .ZN(new_n2053_));
  AOI21_X1   g1411(.A1(new_n1370_), .A2(new_n2023_), .B(new_n2053_), .ZN(new_n2054_));
  NOR2_X1    g1412(.A1(new_n2049_), .A2(\in1[125] ), .ZN(new_n2055_));
  AOI21_X1   g1413(.A1(new_n646_), .A2(new_n2049_), .B(new_n2055_), .ZN(new_n2056_));
  INV_X1     g1414(.I(new_n2056_), .ZN(new_n2057_));
  AOI22_X1   g1415(.A1(new_n2025_), .A2(new_n2052_), .B1(new_n2057_), .B2(new_n2054_), .ZN(new_n2058_));
  NOR2_X1    g1416(.A1(new_n2023_), .A2(\in3[124] ), .ZN(new_n2059_));
  AOI21_X1   g1417(.A1(new_n1373_), .A2(new_n2023_), .B(new_n2059_), .ZN(new_n2060_));
  NOR2_X1    g1418(.A1(new_n2049_), .A2(\in1[124] ), .ZN(new_n2061_));
  INV_X1     g1419(.I(new_n2049_), .ZN(new_n2062_));
  NOR2_X1    g1420(.A1(new_n2062_), .A2(\in0[124] ), .ZN(new_n2063_));
  NOR2_X1    g1421(.A1(new_n2063_), .A2(new_n2061_), .ZN(new_n2064_));
  INV_X1     g1422(.I(new_n2064_), .ZN(new_n2065_));
  OAI22_X1   g1423(.A1(new_n2065_), .A2(new_n2060_), .B1(new_n2057_), .B2(new_n2054_), .ZN(new_n2066_));
  AOI22_X1   g1424(.A1(new_n2066_), .A2(new_n2058_), .B1(new_n2026_), .B2(new_n2051_), .ZN(new_n2067_));
  NOR2_X1    g1425(.A1(new_n2067_), .A2(new_n1940_), .ZN(new_n2068_));
  INV_X1     g1426(.I(new_n2058_), .ZN(new_n2069_));
  AOI21_X1   g1427(.A1(new_n2060_), .A2(new_n2065_), .B(new_n2069_), .ZN(new_n2070_));
  NAND2_X1   g1428(.A1(new_n2070_), .A2(new_n1939_), .ZN(new_n2071_));
  INV_X1     g1429(.I(\in2[120] ), .ZN(new_n2072_));
  NOR2_X1    g1430(.A1(new_n2023_), .A2(\in3[120] ), .ZN(new_n2073_));
  AOI21_X1   g1431(.A1(new_n2072_), .A2(new_n2023_), .B(new_n2073_), .ZN(new_n2074_));
  INV_X1     g1432(.I(new_n2074_), .ZN(new_n2075_));
  INV_X1     g1433(.I(\in0[120] ), .ZN(new_n2076_));
  NOR2_X1    g1434(.A1(new_n2049_), .A2(\in1[120] ), .ZN(new_n2077_));
  AOI21_X1   g1435(.A1(new_n2076_), .A2(new_n2049_), .B(new_n2077_), .ZN(new_n2078_));
  NOR2_X1    g1436(.A1(new_n2075_), .A2(new_n2078_), .ZN(new_n2079_));
  NOR2_X1    g1437(.A1(new_n2023_), .A2(\in3[123] ), .ZN(new_n2080_));
  AOI21_X1   g1438(.A1(new_n1388_), .A2(new_n2023_), .B(new_n2080_), .ZN(new_n2081_));
  NOR2_X1    g1439(.A1(new_n2049_), .A2(\in1[123] ), .ZN(new_n2082_));
  AOI21_X1   g1440(.A1(new_n665_), .A2(new_n2049_), .B(new_n2082_), .ZN(new_n2083_));
  INV_X1     g1441(.I(new_n2083_), .ZN(new_n2084_));
  NOR2_X1    g1442(.A1(new_n2023_), .A2(\in3[122] ), .ZN(new_n2085_));
  AOI21_X1   g1443(.A1(new_n1387_), .A2(new_n2023_), .B(new_n2085_), .ZN(new_n2086_));
  NOR2_X1    g1444(.A1(new_n2049_), .A2(\in1[122] ), .ZN(new_n2087_));
  AOI21_X1   g1445(.A1(new_n664_), .A2(new_n2049_), .B(new_n2087_), .ZN(new_n2088_));
  INV_X1     g1446(.I(new_n2088_), .ZN(new_n2089_));
  AOI22_X1   g1447(.A1(new_n2081_), .A2(new_n2084_), .B1(new_n2089_), .B2(new_n2086_), .ZN(new_n2090_));
  INV_X1     g1448(.I(new_n2090_), .ZN(new_n2091_));
  NOR2_X1    g1449(.A1(new_n2023_), .A2(\in3[121] ), .ZN(new_n2092_));
  AOI21_X1   g1450(.A1(new_n1928_), .A2(new_n2023_), .B(new_n2092_), .ZN(new_n2093_));
  INV_X1     g1451(.I(new_n2093_), .ZN(new_n2094_));
  NOR2_X1    g1452(.A1(new_n2049_), .A2(\in1[121] ), .ZN(new_n2095_));
  NOR2_X1    g1453(.A1(new_n2062_), .A2(\in0[121] ), .ZN(new_n2096_));
  NOR2_X1    g1454(.A1(new_n2096_), .A2(new_n2095_), .ZN(new_n2097_));
  NOR2_X1    g1455(.A1(new_n2094_), .A2(new_n2097_), .ZN(new_n2098_));
  NOR3_X1    g1456(.A1(new_n2091_), .A2(new_n2079_), .A3(new_n2098_), .ZN(new_n2099_));
  NOR2_X1    g1457(.A1(new_n2023_), .A2(\in3[119] ), .ZN(new_n2100_));
  AOI21_X1   g1458(.A1(new_n1404_), .A2(new_n2023_), .B(new_n2100_), .ZN(new_n2101_));
  INV_X1     g1459(.I(new_n2101_), .ZN(new_n2102_));
  NOR2_X1    g1460(.A1(new_n2049_), .A2(\in1[119] ), .ZN(new_n2103_));
  NOR2_X1    g1461(.A1(new_n2062_), .A2(\in0[119] ), .ZN(new_n2104_));
  NOR2_X1    g1462(.A1(new_n2104_), .A2(new_n2103_), .ZN(new_n2105_));
  NOR2_X1    g1463(.A1(new_n2102_), .A2(new_n2105_), .ZN(new_n2106_));
  NOR2_X1    g1464(.A1(new_n2023_), .A2(\in3[118] ), .ZN(new_n2107_));
  AOI21_X1   g1465(.A1(new_n1397_), .A2(new_n2023_), .B(new_n2107_), .ZN(new_n2108_));
  NOR2_X1    g1466(.A1(new_n2049_), .A2(\in1[118] ), .ZN(new_n2109_));
  AOI21_X1   g1467(.A1(new_n673_), .A2(new_n2049_), .B(new_n2109_), .ZN(new_n2110_));
  INV_X1     g1468(.I(new_n2110_), .ZN(new_n2111_));
  AOI21_X1   g1469(.A1(new_n2108_), .A2(new_n2111_), .B(new_n2106_), .ZN(new_n2112_));
  INV_X1     g1470(.I(new_n2112_), .ZN(new_n2113_));
  INV_X1     g1471(.I(\in2[117] ), .ZN(new_n2114_));
  NOR2_X1    g1472(.A1(new_n2023_), .A2(\in3[117] ), .ZN(new_n2115_));
  AOI21_X1   g1473(.A1(new_n2114_), .A2(new_n2023_), .B(new_n2115_), .ZN(new_n2116_));
  INV_X1     g1474(.I(new_n2116_), .ZN(new_n2117_));
  NOR2_X1    g1475(.A1(new_n2049_), .A2(\in1[117] ), .ZN(new_n2118_));
  NOR2_X1    g1476(.A1(new_n2062_), .A2(\in0[117] ), .ZN(new_n2119_));
  NOR2_X1    g1477(.A1(new_n2119_), .A2(new_n2118_), .ZN(new_n2120_));
  NOR2_X1    g1478(.A1(new_n2117_), .A2(new_n2120_), .ZN(new_n2121_));
  INV_X1     g1479(.I(new_n2121_), .ZN(new_n2122_));
  INV_X1     g1480(.I(new_n2120_), .ZN(new_n2123_));
  INV_X1     g1481(.I(new_n2022_), .ZN(new_n2124_));
  NOR2_X1    g1482(.A1(new_n1936_), .A2(new_n2124_), .ZN(new_n2125_));
  NOR2_X1    g1483(.A1(new_n2125_), .A2(\in2[116] ), .ZN(new_n2126_));
  AOI21_X1   g1484(.A1(new_n1401_), .A2(new_n2125_), .B(new_n2126_), .ZN(new_n2127_));
  NOR2_X1    g1485(.A1(new_n2062_), .A2(\in0[116] ), .ZN(new_n2128_));
  AOI21_X1   g1486(.A1(new_n678_), .A2(new_n2062_), .B(new_n2128_), .ZN(new_n2129_));
  INV_X1     g1487(.I(new_n2129_), .ZN(new_n2130_));
  OAI22_X1   g1488(.A1(new_n2116_), .A2(new_n2123_), .B1(new_n2130_), .B2(new_n2127_), .ZN(new_n2131_));
  NAND2_X1   g1489(.A1(new_n2131_), .A2(new_n2122_), .ZN(new_n2132_));
  INV_X1     g1490(.I(new_n2105_), .ZN(new_n2133_));
  OAI22_X1   g1491(.A1(new_n2133_), .A2(new_n2101_), .B1(new_n2111_), .B2(new_n2108_), .ZN(new_n2134_));
  INV_X1     g1492(.I(new_n2134_), .ZN(new_n2135_));
  OAI22_X1   g1493(.A1(new_n2132_), .A2(new_n2113_), .B1(new_n2106_), .B2(new_n2135_), .ZN(new_n2136_));
  NOR2_X1    g1494(.A1(new_n2023_), .A2(\in3[115] ), .ZN(new_n2137_));
  AOI21_X1   g1495(.A1(new_n1409_), .A2(new_n2023_), .B(new_n2137_), .ZN(new_n2138_));
  INV_X1     g1496(.I(new_n2138_), .ZN(new_n2139_));
  NOR2_X1    g1497(.A1(new_n2049_), .A2(\in1[115] ), .ZN(new_n2140_));
  AOI21_X1   g1498(.A1(new_n688_), .A2(new_n2049_), .B(new_n2140_), .ZN(new_n2141_));
  INV_X1     g1499(.I(new_n2141_), .ZN(new_n2142_));
  NOR2_X1    g1500(.A1(new_n2023_), .A2(\in3[114] ), .ZN(new_n2143_));
  AOI21_X1   g1501(.A1(new_n1408_), .A2(new_n2023_), .B(new_n2143_), .ZN(new_n2144_));
  NOR2_X1    g1502(.A1(new_n2049_), .A2(\in1[114] ), .ZN(new_n2145_));
  AOI21_X1   g1503(.A1(new_n687_), .A2(new_n2049_), .B(new_n2145_), .ZN(new_n2146_));
  INV_X1     g1504(.I(new_n2146_), .ZN(new_n2147_));
  AOI22_X1   g1505(.A1(new_n2138_), .A2(new_n2142_), .B1(new_n2147_), .B2(new_n2144_), .ZN(new_n2148_));
  NOR2_X1    g1506(.A1(new_n2023_), .A2(\in3[113] ), .ZN(new_n2149_));
  AOI21_X1   g1507(.A1(new_n1411_), .A2(new_n2023_), .B(new_n2149_), .ZN(new_n2150_));
  INV_X1     g1508(.I(new_n2150_), .ZN(new_n2151_));
  NOR2_X1    g1509(.A1(new_n2049_), .A2(\in1[113] ), .ZN(new_n2152_));
  NOR2_X1    g1510(.A1(new_n2062_), .A2(\in0[113] ), .ZN(new_n2153_));
  NOR2_X1    g1511(.A1(new_n2153_), .A2(new_n2152_), .ZN(new_n2154_));
  NOR2_X1    g1512(.A1(new_n2151_), .A2(new_n2154_), .ZN(new_n2155_));
  NOR2_X1    g1513(.A1(new_n2023_), .A2(\in3[112] ), .ZN(new_n2156_));
  AOI21_X1   g1514(.A1(new_n1413_), .A2(new_n2023_), .B(new_n2156_), .ZN(new_n2157_));
  INV_X1     g1515(.I(new_n2157_), .ZN(new_n2158_));
  INV_X1     g1516(.I(\in0[112] ), .ZN(new_n2159_));
  NOR2_X1    g1517(.A1(new_n2049_), .A2(\in1[112] ), .ZN(new_n2160_));
  AOI21_X1   g1518(.A1(new_n2159_), .A2(new_n2049_), .B(new_n2160_), .ZN(new_n2161_));
  AOI22_X1   g1519(.A1(new_n2151_), .A2(new_n2154_), .B1(new_n2158_), .B2(new_n2161_), .ZN(new_n2162_));
  OAI22_X1   g1520(.A1(new_n2162_), .A2(new_n2155_), .B1(new_n2144_), .B2(new_n2147_), .ZN(new_n2163_));
  AOI22_X1   g1521(.A1(new_n2163_), .A2(new_n2148_), .B1(new_n2139_), .B2(new_n2141_), .ZN(new_n2164_));
  INV_X1     g1522(.I(new_n2148_), .ZN(new_n2165_));
  NOR2_X1    g1523(.A1(new_n2158_), .A2(new_n2161_), .ZN(new_n2166_));
  NOR3_X1    g1524(.A1(new_n2165_), .A2(new_n2155_), .A3(new_n2166_), .ZN(new_n2167_));
  INV_X1     g1525(.I(\in2[109] ), .ZN(new_n2168_));
  NOR2_X1    g1526(.A1(new_n2023_), .A2(\in3[109] ), .ZN(new_n2169_));
  AOI21_X1   g1527(.A1(new_n2168_), .A2(new_n2023_), .B(new_n2169_), .ZN(new_n2170_));
  INV_X1     g1528(.I(new_n2170_), .ZN(new_n2171_));
  NOR2_X1    g1529(.A1(new_n2049_), .A2(\in1[109] ), .ZN(new_n2172_));
  NOR2_X1    g1530(.A1(new_n2062_), .A2(\in0[109] ), .ZN(new_n2173_));
  NOR2_X1    g1531(.A1(new_n2173_), .A2(new_n2172_), .ZN(new_n2174_));
  NOR2_X1    g1532(.A1(new_n2171_), .A2(new_n2174_), .ZN(new_n2175_));
  NOR2_X1    g1533(.A1(new_n2023_), .A2(\in3[111] ), .ZN(new_n2176_));
  AOI21_X1   g1534(.A1(new_n1917_), .A2(new_n2023_), .B(new_n2176_), .ZN(new_n2177_));
  INV_X1     g1535(.I(new_n2177_), .ZN(new_n2178_));
  NOR2_X1    g1536(.A1(new_n2049_), .A2(\in1[111] ), .ZN(new_n2179_));
  NOR2_X1    g1537(.A1(new_n2062_), .A2(\in0[111] ), .ZN(new_n2180_));
  NOR2_X1    g1538(.A1(new_n2180_), .A2(new_n2179_), .ZN(new_n2181_));
  NOR2_X1    g1539(.A1(new_n2178_), .A2(new_n2181_), .ZN(new_n2182_));
  NOR2_X1    g1540(.A1(new_n2023_), .A2(\in3[110] ), .ZN(new_n2183_));
  AOI21_X1   g1541(.A1(new_n1423_), .A2(new_n2023_), .B(new_n2183_), .ZN(new_n2184_));
  NOR2_X1    g1542(.A1(new_n2049_), .A2(\in1[110] ), .ZN(new_n2185_));
  AOI21_X1   g1543(.A1(new_n702_), .A2(new_n2049_), .B(new_n2185_), .ZN(new_n2186_));
  INV_X1     g1544(.I(new_n2186_), .ZN(new_n2187_));
  AOI21_X1   g1545(.A1(new_n2184_), .A2(new_n2187_), .B(new_n2182_), .ZN(new_n2188_));
  INV_X1     g1546(.I(new_n2188_), .ZN(new_n2189_));
  INV_X1     g1547(.I(\in2[108] ), .ZN(new_n2190_));
  NOR2_X1    g1548(.A1(new_n2023_), .A2(\in3[108] ), .ZN(new_n2191_));
  AOI21_X1   g1549(.A1(new_n2190_), .A2(new_n2023_), .B(new_n2191_), .ZN(new_n2192_));
  INV_X1     g1550(.I(new_n2192_), .ZN(new_n2193_));
  NOR2_X1    g1551(.A1(new_n2049_), .A2(\in1[108] ), .ZN(new_n2194_));
  NOR2_X1    g1552(.A1(new_n2062_), .A2(\in0[108] ), .ZN(new_n2195_));
  NOR2_X1    g1553(.A1(new_n2195_), .A2(new_n2194_), .ZN(new_n2196_));
  NOR2_X1    g1554(.A1(new_n2193_), .A2(new_n2196_), .ZN(new_n2197_));
  NOR3_X1    g1555(.A1(new_n2189_), .A2(new_n2175_), .A3(new_n2197_), .ZN(new_n2198_));
  INV_X1     g1556(.I(new_n2198_), .ZN(new_n2199_));
  NOR2_X1    g1557(.A1(new_n2023_), .A2(\in3[107] ), .ZN(new_n2200_));
  AOI21_X1   g1558(.A1(new_n1436_), .A2(new_n2023_), .B(new_n2200_), .ZN(new_n2201_));
  INV_X1     g1559(.I(new_n2201_), .ZN(new_n2202_));
  NOR2_X1    g1560(.A1(new_n2049_), .A2(\in1[107] ), .ZN(new_n2203_));
  AOI21_X1   g1561(.A1(new_n715_), .A2(new_n2049_), .B(new_n2203_), .ZN(new_n2204_));
  INV_X1     g1562(.I(new_n2204_), .ZN(new_n2205_));
  NOR2_X1    g1563(.A1(new_n2023_), .A2(\in3[106] ), .ZN(new_n2206_));
  AOI21_X1   g1564(.A1(new_n1435_), .A2(new_n2023_), .B(new_n2206_), .ZN(new_n2207_));
  NOR2_X1    g1565(.A1(new_n2049_), .A2(\in1[106] ), .ZN(new_n2208_));
  AOI21_X1   g1566(.A1(new_n714_), .A2(new_n2049_), .B(new_n2208_), .ZN(new_n2209_));
  INV_X1     g1567(.I(new_n2209_), .ZN(new_n2210_));
  AOI22_X1   g1568(.A1(new_n2201_), .A2(new_n2205_), .B1(new_n2210_), .B2(new_n2207_), .ZN(new_n2211_));
  NOR2_X1    g1569(.A1(new_n2023_), .A2(\in3[105] ), .ZN(new_n2212_));
  AOI21_X1   g1570(.A1(new_n1438_), .A2(new_n2023_), .B(new_n2212_), .ZN(new_n2213_));
  INV_X1     g1571(.I(new_n2213_), .ZN(new_n2214_));
  NOR2_X1    g1572(.A1(new_n2049_), .A2(\in1[105] ), .ZN(new_n2215_));
  NOR2_X1    g1573(.A1(new_n2062_), .A2(\in0[105] ), .ZN(new_n2216_));
  NOR2_X1    g1574(.A1(new_n2216_), .A2(new_n2215_), .ZN(new_n2217_));
  NOR2_X1    g1575(.A1(new_n2214_), .A2(new_n2217_), .ZN(new_n2218_));
  NOR2_X1    g1576(.A1(new_n2023_), .A2(\in3[104] ), .ZN(new_n2219_));
  AOI21_X1   g1577(.A1(new_n1440_), .A2(new_n2023_), .B(new_n2219_), .ZN(new_n2220_));
  INV_X1     g1578(.I(new_n2220_), .ZN(new_n2221_));
  INV_X1     g1579(.I(\in0[104] ), .ZN(new_n2222_));
  NOR2_X1    g1580(.A1(new_n2049_), .A2(\in1[104] ), .ZN(new_n2223_));
  AOI21_X1   g1581(.A1(new_n2222_), .A2(new_n2049_), .B(new_n2223_), .ZN(new_n2224_));
  AOI22_X1   g1582(.A1(new_n2214_), .A2(new_n2217_), .B1(new_n2221_), .B2(new_n2224_), .ZN(new_n2225_));
  OAI22_X1   g1583(.A1(new_n2225_), .A2(new_n2218_), .B1(new_n2207_), .B2(new_n2210_), .ZN(new_n2226_));
  AOI22_X1   g1584(.A1(new_n2226_), .A2(new_n2211_), .B1(new_n2202_), .B2(new_n2204_), .ZN(new_n2227_));
  NOR2_X1    g1585(.A1(new_n2023_), .A2(\in3[103] ), .ZN(new_n2228_));
  AOI21_X1   g1586(.A1(new_n1457_), .A2(new_n2023_), .B(new_n2228_), .ZN(new_n2229_));
  INV_X1     g1587(.I(new_n2229_), .ZN(new_n2230_));
  NOR2_X1    g1588(.A1(new_n2049_), .A2(\in1[103] ), .ZN(new_n2231_));
  NOR2_X1    g1589(.A1(new_n2062_), .A2(\in0[103] ), .ZN(new_n2232_));
  NOR2_X1    g1590(.A1(new_n2232_), .A2(new_n2231_), .ZN(new_n2233_));
  NOR2_X1    g1591(.A1(new_n2230_), .A2(new_n2233_), .ZN(new_n2234_));
  NOR2_X1    g1592(.A1(new_n2023_), .A2(\in3[102] ), .ZN(new_n2235_));
  AOI21_X1   g1593(.A1(new_n1450_), .A2(new_n2023_), .B(new_n2235_), .ZN(new_n2236_));
  NOR2_X1    g1594(.A1(new_n2049_), .A2(\in1[102] ), .ZN(new_n2237_));
  AOI21_X1   g1595(.A1(new_n728_), .A2(new_n2049_), .B(new_n2237_), .ZN(new_n2238_));
  INV_X1     g1596(.I(new_n2238_), .ZN(new_n2239_));
  AOI21_X1   g1597(.A1(new_n2236_), .A2(new_n2239_), .B(new_n2234_), .ZN(new_n2240_));
  INV_X1     g1598(.I(new_n2240_), .ZN(new_n2241_));
  INV_X1     g1599(.I(\in2[101] ), .ZN(new_n2242_));
  NOR2_X1    g1600(.A1(new_n2023_), .A2(\in3[101] ), .ZN(new_n2243_));
  AOI21_X1   g1601(.A1(new_n2242_), .A2(new_n2023_), .B(new_n2243_), .ZN(new_n2244_));
  INV_X1     g1602(.I(new_n2244_), .ZN(new_n2245_));
  NOR2_X1    g1603(.A1(new_n2049_), .A2(\in1[101] ), .ZN(new_n2246_));
  NOR2_X1    g1604(.A1(new_n2062_), .A2(\in0[101] ), .ZN(new_n2247_));
  NOR2_X1    g1605(.A1(new_n2247_), .A2(new_n2246_), .ZN(new_n2248_));
  NOR2_X1    g1606(.A1(new_n2245_), .A2(new_n2248_), .ZN(new_n2249_));
  INV_X1     g1607(.I(new_n2249_), .ZN(new_n2250_));
  INV_X1     g1608(.I(new_n2248_), .ZN(new_n2251_));
  NOR2_X1    g1609(.A1(new_n2125_), .A2(\in2[100] ), .ZN(new_n2252_));
  AOI21_X1   g1610(.A1(new_n1454_), .A2(new_n2125_), .B(new_n2252_), .ZN(new_n2253_));
  NOR2_X1    g1611(.A1(new_n2062_), .A2(\in0[100] ), .ZN(new_n2254_));
  AOI21_X1   g1612(.A1(new_n733_), .A2(new_n2062_), .B(new_n2254_), .ZN(new_n2255_));
  INV_X1     g1613(.I(new_n2255_), .ZN(new_n2256_));
  OAI22_X1   g1614(.A1(new_n2244_), .A2(new_n2251_), .B1(new_n2256_), .B2(new_n2253_), .ZN(new_n2257_));
  NAND2_X1   g1615(.A1(new_n2257_), .A2(new_n2250_), .ZN(new_n2258_));
  INV_X1     g1616(.I(new_n2233_), .ZN(new_n2259_));
  OAI22_X1   g1617(.A1(new_n2259_), .A2(new_n2229_), .B1(new_n2239_), .B2(new_n2236_), .ZN(new_n2260_));
  INV_X1     g1618(.I(new_n2260_), .ZN(new_n2261_));
  OAI22_X1   g1619(.A1(new_n2258_), .A2(new_n2241_), .B1(new_n2234_), .B2(new_n2261_), .ZN(new_n2262_));
  NAND2_X1   g1620(.A1(new_n2256_), .A2(new_n2253_), .ZN(new_n2263_));
  NAND3_X1   g1621(.A1(new_n2240_), .A2(new_n2250_), .A3(new_n2263_), .ZN(new_n2264_));
  INV_X1     g1622(.I(\in2[96] ), .ZN(new_n2265_));
  NOR2_X1    g1623(.A1(new_n2023_), .A2(\in3[96] ), .ZN(new_n2266_));
  AOI21_X1   g1624(.A1(new_n2265_), .A2(new_n2023_), .B(new_n2266_), .ZN(new_n2267_));
  INV_X1     g1625(.I(new_n2267_), .ZN(new_n2268_));
  INV_X1     g1626(.I(\in0[96] ), .ZN(new_n2269_));
  NOR2_X1    g1627(.A1(new_n2049_), .A2(\in1[96] ), .ZN(new_n2270_));
  AOI21_X1   g1628(.A1(new_n2269_), .A2(new_n2049_), .B(new_n2270_), .ZN(new_n2271_));
  NOR2_X1    g1629(.A1(new_n2268_), .A2(new_n2271_), .ZN(new_n2272_));
  NOR2_X1    g1630(.A1(new_n2023_), .A2(\in3[99] ), .ZN(new_n2273_));
  AOI21_X1   g1631(.A1(new_n1467_), .A2(new_n2023_), .B(new_n2273_), .ZN(new_n2274_));
  NOR2_X1    g1632(.A1(new_n2049_), .A2(\in1[99] ), .ZN(new_n2275_));
  AOI21_X1   g1633(.A1(new_n747_), .A2(new_n2049_), .B(new_n2275_), .ZN(new_n2276_));
  INV_X1     g1634(.I(new_n2276_), .ZN(new_n2277_));
  NOR2_X1    g1635(.A1(new_n2023_), .A2(\in3[98] ), .ZN(new_n2278_));
  AOI21_X1   g1636(.A1(new_n1466_), .A2(new_n2023_), .B(new_n2278_), .ZN(new_n2279_));
  NOR2_X1    g1637(.A1(new_n2049_), .A2(\in1[98] ), .ZN(new_n2280_));
  AOI21_X1   g1638(.A1(new_n746_), .A2(new_n2049_), .B(new_n2280_), .ZN(new_n2281_));
  INV_X1     g1639(.I(new_n2281_), .ZN(new_n2282_));
  AOI22_X1   g1640(.A1(new_n2274_), .A2(new_n2277_), .B1(new_n2282_), .B2(new_n2279_), .ZN(new_n2283_));
  INV_X1     g1641(.I(new_n2283_), .ZN(new_n2284_));
  NOR2_X1    g1642(.A1(new_n2023_), .A2(\in3[97] ), .ZN(new_n2285_));
  AOI21_X1   g1643(.A1(new_n1901_), .A2(new_n2023_), .B(new_n2285_), .ZN(new_n2286_));
  INV_X1     g1644(.I(new_n2286_), .ZN(new_n2287_));
  NOR2_X1    g1645(.A1(new_n2049_), .A2(\in1[97] ), .ZN(new_n2288_));
  NOR2_X1    g1646(.A1(new_n2062_), .A2(\in0[97] ), .ZN(new_n2289_));
  NOR2_X1    g1647(.A1(new_n2289_), .A2(new_n2288_), .ZN(new_n2290_));
  NOR2_X1    g1648(.A1(new_n2287_), .A2(new_n2290_), .ZN(new_n2291_));
  NOR3_X1    g1649(.A1(new_n2284_), .A2(new_n2272_), .A3(new_n2291_), .ZN(new_n2292_));
  NOR2_X1    g1650(.A1(new_n2023_), .A2(\in3[95] ), .ZN(new_n2293_));
  AOI21_X1   g1651(.A1(new_n1483_), .A2(new_n2023_), .B(new_n2293_), .ZN(new_n2294_));
  INV_X1     g1652(.I(new_n2294_), .ZN(new_n2295_));
  NOR2_X1    g1653(.A1(new_n2049_), .A2(\in1[95] ), .ZN(new_n2296_));
  NOR2_X1    g1654(.A1(new_n2062_), .A2(\in0[95] ), .ZN(new_n2297_));
  NOR2_X1    g1655(.A1(new_n2297_), .A2(new_n2296_), .ZN(new_n2298_));
  NOR2_X1    g1656(.A1(new_n2295_), .A2(new_n2298_), .ZN(new_n2299_));
  NOR2_X1    g1657(.A1(new_n2023_), .A2(\in3[94] ), .ZN(new_n2300_));
  AOI21_X1   g1658(.A1(new_n1476_), .A2(new_n2023_), .B(new_n2300_), .ZN(new_n2301_));
  NOR2_X1    g1659(.A1(new_n2049_), .A2(\in1[94] ), .ZN(new_n2302_));
  AOI21_X1   g1660(.A1(new_n755_), .A2(new_n2049_), .B(new_n2302_), .ZN(new_n2303_));
  INV_X1     g1661(.I(new_n2303_), .ZN(new_n2304_));
  AOI21_X1   g1662(.A1(new_n2301_), .A2(new_n2304_), .B(new_n2299_), .ZN(new_n2305_));
  INV_X1     g1663(.I(new_n2305_), .ZN(new_n2306_));
  INV_X1     g1664(.I(\in2[93] ), .ZN(new_n2307_));
  NOR2_X1    g1665(.A1(new_n2023_), .A2(\in3[93] ), .ZN(new_n2308_));
  AOI21_X1   g1666(.A1(new_n2307_), .A2(new_n2023_), .B(new_n2308_), .ZN(new_n2309_));
  INV_X1     g1667(.I(new_n2309_), .ZN(new_n2310_));
  NOR2_X1    g1668(.A1(new_n2049_), .A2(\in1[93] ), .ZN(new_n2311_));
  NOR2_X1    g1669(.A1(new_n2062_), .A2(\in0[93] ), .ZN(new_n2312_));
  NOR2_X1    g1670(.A1(new_n2312_), .A2(new_n2311_), .ZN(new_n2313_));
  NOR2_X1    g1671(.A1(new_n2310_), .A2(new_n2313_), .ZN(new_n2314_));
  INV_X1     g1672(.I(new_n2314_), .ZN(new_n2315_));
  INV_X1     g1673(.I(new_n2313_), .ZN(new_n2316_));
  NOR2_X1    g1674(.A1(new_n2125_), .A2(\in2[92] ), .ZN(new_n2317_));
  AOI21_X1   g1675(.A1(new_n1480_), .A2(new_n2125_), .B(new_n2317_), .ZN(new_n2318_));
  NOR2_X1    g1676(.A1(new_n2062_), .A2(\in0[92] ), .ZN(new_n2319_));
  AOI21_X1   g1677(.A1(new_n760_), .A2(new_n2062_), .B(new_n2319_), .ZN(new_n2320_));
  INV_X1     g1678(.I(new_n2320_), .ZN(new_n2321_));
  OAI22_X1   g1679(.A1(new_n2309_), .A2(new_n2316_), .B1(new_n2321_), .B2(new_n2318_), .ZN(new_n2322_));
  NAND2_X1   g1680(.A1(new_n2322_), .A2(new_n2315_), .ZN(new_n2323_));
  INV_X1     g1681(.I(new_n2298_), .ZN(new_n2324_));
  OAI22_X1   g1682(.A1(new_n2324_), .A2(new_n2294_), .B1(new_n2304_), .B2(new_n2301_), .ZN(new_n2325_));
  INV_X1     g1683(.I(new_n2325_), .ZN(new_n2326_));
  OAI22_X1   g1684(.A1(new_n2323_), .A2(new_n2306_), .B1(new_n2299_), .B2(new_n2326_), .ZN(new_n2327_));
  NOR2_X1    g1685(.A1(new_n2023_), .A2(\in3[91] ), .ZN(new_n2328_));
  AOI21_X1   g1686(.A1(new_n1488_), .A2(new_n2023_), .B(new_n2328_), .ZN(new_n2329_));
  INV_X1     g1687(.I(new_n2329_), .ZN(new_n2330_));
  NOR2_X1    g1688(.A1(new_n2049_), .A2(\in1[91] ), .ZN(new_n2331_));
  AOI21_X1   g1689(.A1(new_n770_), .A2(new_n2049_), .B(new_n2331_), .ZN(new_n2332_));
  INV_X1     g1690(.I(new_n2332_), .ZN(new_n2333_));
  NOR2_X1    g1691(.A1(new_n2023_), .A2(\in3[90] ), .ZN(new_n2334_));
  AOI21_X1   g1692(.A1(new_n1487_), .A2(new_n2023_), .B(new_n2334_), .ZN(new_n2335_));
  NOR2_X1    g1693(.A1(new_n2049_), .A2(\in1[90] ), .ZN(new_n2336_));
  AOI21_X1   g1694(.A1(new_n769_), .A2(new_n2049_), .B(new_n2336_), .ZN(new_n2337_));
  INV_X1     g1695(.I(new_n2337_), .ZN(new_n2338_));
  AOI22_X1   g1696(.A1(new_n2329_), .A2(new_n2333_), .B1(new_n2338_), .B2(new_n2335_), .ZN(new_n2339_));
  NOR2_X1    g1697(.A1(new_n2023_), .A2(\in3[89] ), .ZN(new_n2340_));
  AOI21_X1   g1698(.A1(new_n1490_), .A2(new_n2023_), .B(new_n2340_), .ZN(new_n2341_));
  INV_X1     g1699(.I(new_n2341_), .ZN(new_n2342_));
  NOR2_X1    g1700(.A1(new_n2049_), .A2(\in1[89] ), .ZN(new_n2343_));
  NOR2_X1    g1701(.A1(new_n2062_), .A2(\in0[89] ), .ZN(new_n2344_));
  NOR2_X1    g1702(.A1(new_n2344_), .A2(new_n2343_), .ZN(new_n2345_));
  NOR2_X1    g1703(.A1(new_n2342_), .A2(new_n2345_), .ZN(new_n2346_));
  NOR2_X1    g1704(.A1(new_n2023_), .A2(\in3[88] ), .ZN(new_n2347_));
  AOI21_X1   g1705(.A1(new_n1492_), .A2(new_n2023_), .B(new_n2347_), .ZN(new_n2348_));
  INV_X1     g1706(.I(new_n2348_), .ZN(new_n2349_));
  INV_X1     g1707(.I(\in0[88] ), .ZN(new_n2350_));
  NOR2_X1    g1708(.A1(new_n2049_), .A2(\in1[88] ), .ZN(new_n2351_));
  AOI21_X1   g1709(.A1(new_n2350_), .A2(new_n2049_), .B(new_n2351_), .ZN(new_n2352_));
  AOI22_X1   g1710(.A1(new_n2342_), .A2(new_n2345_), .B1(new_n2349_), .B2(new_n2352_), .ZN(new_n2353_));
  OAI22_X1   g1711(.A1(new_n2353_), .A2(new_n2346_), .B1(new_n2335_), .B2(new_n2338_), .ZN(new_n2354_));
  AOI22_X1   g1712(.A1(new_n2354_), .A2(new_n2339_), .B1(new_n2330_), .B2(new_n2332_), .ZN(new_n2355_));
  INV_X1     g1713(.I(new_n2339_), .ZN(new_n2356_));
  NOR2_X1    g1714(.A1(new_n2349_), .A2(new_n2352_), .ZN(new_n2357_));
  NOR3_X1    g1715(.A1(new_n2356_), .A2(new_n2346_), .A3(new_n2357_), .ZN(new_n2358_));
  INV_X1     g1716(.I(\in2[85] ), .ZN(new_n2359_));
  NOR2_X1    g1717(.A1(new_n2023_), .A2(\in3[85] ), .ZN(new_n2360_));
  AOI21_X1   g1718(.A1(new_n2359_), .A2(new_n2023_), .B(new_n2360_), .ZN(new_n2361_));
  INV_X1     g1719(.I(new_n2361_), .ZN(new_n2362_));
  NOR2_X1    g1720(.A1(new_n2049_), .A2(\in1[85] ), .ZN(new_n2363_));
  NOR2_X1    g1721(.A1(new_n2062_), .A2(\in0[85] ), .ZN(new_n2364_));
  NOR2_X1    g1722(.A1(new_n2364_), .A2(new_n2363_), .ZN(new_n2365_));
  NOR2_X1    g1723(.A1(new_n2362_), .A2(new_n2365_), .ZN(new_n2366_));
  NOR2_X1    g1724(.A1(new_n2023_), .A2(\in3[87] ), .ZN(new_n2367_));
  AOI21_X1   g1725(.A1(new_n1890_), .A2(new_n2023_), .B(new_n2367_), .ZN(new_n2368_));
  INV_X1     g1726(.I(new_n2368_), .ZN(new_n2369_));
  NOR2_X1    g1727(.A1(new_n2049_), .A2(\in1[87] ), .ZN(new_n2370_));
  NOR2_X1    g1728(.A1(new_n2062_), .A2(\in0[87] ), .ZN(new_n2371_));
  NOR2_X1    g1729(.A1(new_n2371_), .A2(new_n2370_), .ZN(new_n2372_));
  NOR2_X1    g1730(.A1(new_n2369_), .A2(new_n2372_), .ZN(new_n2373_));
  NOR2_X1    g1731(.A1(new_n2023_), .A2(\in3[86] ), .ZN(new_n2374_));
  AOI21_X1   g1732(.A1(new_n1502_), .A2(new_n2023_), .B(new_n2374_), .ZN(new_n2375_));
  NOR2_X1    g1733(.A1(new_n2049_), .A2(\in1[86] ), .ZN(new_n2376_));
  AOI21_X1   g1734(.A1(new_n784_), .A2(new_n2049_), .B(new_n2376_), .ZN(new_n2377_));
  INV_X1     g1735(.I(new_n2377_), .ZN(new_n2378_));
  AOI21_X1   g1736(.A1(new_n2375_), .A2(new_n2378_), .B(new_n2373_), .ZN(new_n2379_));
  INV_X1     g1737(.I(new_n2379_), .ZN(new_n2380_));
  INV_X1     g1738(.I(\in2[84] ), .ZN(new_n2381_));
  NOR2_X1    g1739(.A1(new_n2023_), .A2(\in3[84] ), .ZN(new_n2382_));
  AOI21_X1   g1740(.A1(new_n2381_), .A2(new_n2023_), .B(new_n2382_), .ZN(new_n2383_));
  INV_X1     g1741(.I(new_n2383_), .ZN(new_n2384_));
  NOR2_X1    g1742(.A1(new_n2049_), .A2(\in1[84] ), .ZN(new_n2385_));
  NOR2_X1    g1743(.A1(new_n2062_), .A2(\in0[84] ), .ZN(new_n2386_));
  NOR2_X1    g1744(.A1(new_n2386_), .A2(new_n2385_), .ZN(new_n2387_));
  NOR2_X1    g1745(.A1(new_n2384_), .A2(new_n2387_), .ZN(new_n2388_));
  NOR3_X1    g1746(.A1(new_n2380_), .A2(new_n2366_), .A3(new_n2388_), .ZN(new_n2389_));
  INV_X1     g1747(.I(new_n2389_), .ZN(new_n2390_));
  NOR2_X1    g1748(.A1(new_n2023_), .A2(\in3[83] ), .ZN(new_n2391_));
  AOI21_X1   g1749(.A1(new_n1515_), .A2(new_n2023_), .B(new_n2391_), .ZN(new_n2392_));
  INV_X1     g1750(.I(new_n2392_), .ZN(new_n2393_));
  NOR2_X1    g1751(.A1(new_n2049_), .A2(\in1[83] ), .ZN(new_n2394_));
  AOI21_X1   g1752(.A1(new_n797_), .A2(new_n2049_), .B(new_n2394_), .ZN(new_n2395_));
  INV_X1     g1753(.I(new_n2395_), .ZN(new_n2396_));
  NOR2_X1    g1754(.A1(new_n2023_), .A2(\in3[82] ), .ZN(new_n2397_));
  AOI21_X1   g1755(.A1(new_n1514_), .A2(new_n2023_), .B(new_n2397_), .ZN(new_n2398_));
  NOR2_X1    g1756(.A1(new_n2049_), .A2(\in1[82] ), .ZN(new_n2399_));
  AOI21_X1   g1757(.A1(new_n796_), .A2(new_n2049_), .B(new_n2399_), .ZN(new_n2400_));
  INV_X1     g1758(.I(new_n2400_), .ZN(new_n2401_));
  AOI22_X1   g1759(.A1(new_n2392_), .A2(new_n2396_), .B1(new_n2401_), .B2(new_n2398_), .ZN(new_n2402_));
  NOR2_X1    g1760(.A1(new_n2023_), .A2(\in3[81] ), .ZN(new_n2403_));
  AOI21_X1   g1761(.A1(new_n1517_), .A2(new_n2023_), .B(new_n2403_), .ZN(new_n2404_));
  INV_X1     g1762(.I(new_n2404_), .ZN(new_n2405_));
  NOR2_X1    g1763(.A1(new_n2049_), .A2(\in1[81] ), .ZN(new_n2406_));
  NOR2_X1    g1764(.A1(new_n2062_), .A2(\in0[81] ), .ZN(new_n2407_));
  NOR2_X1    g1765(.A1(new_n2407_), .A2(new_n2406_), .ZN(new_n2408_));
  NOR2_X1    g1766(.A1(new_n2405_), .A2(new_n2408_), .ZN(new_n2409_));
  NOR2_X1    g1767(.A1(new_n2023_), .A2(\in3[80] ), .ZN(new_n2410_));
  AOI21_X1   g1768(.A1(new_n1519_), .A2(new_n2023_), .B(new_n2410_), .ZN(new_n2411_));
  INV_X1     g1769(.I(new_n2411_), .ZN(new_n2412_));
  INV_X1     g1770(.I(\in0[80] ), .ZN(new_n2413_));
  NOR2_X1    g1771(.A1(new_n2049_), .A2(\in1[80] ), .ZN(new_n2414_));
  AOI21_X1   g1772(.A1(new_n2413_), .A2(new_n2049_), .B(new_n2414_), .ZN(new_n2415_));
  AOI22_X1   g1773(.A1(new_n2405_), .A2(new_n2408_), .B1(new_n2412_), .B2(new_n2415_), .ZN(new_n2416_));
  OAI22_X1   g1774(.A1(new_n2416_), .A2(new_n2409_), .B1(new_n2398_), .B2(new_n2401_), .ZN(new_n2417_));
  AOI22_X1   g1775(.A1(new_n2417_), .A2(new_n2402_), .B1(new_n2393_), .B2(new_n2395_), .ZN(new_n2418_));
  NOR2_X1    g1776(.A1(new_n2023_), .A2(\in3[79] ), .ZN(new_n2419_));
  AOI21_X1   g1777(.A1(new_n1536_), .A2(new_n2023_), .B(new_n2419_), .ZN(new_n2420_));
  INV_X1     g1778(.I(new_n2420_), .ZN(new_n2421_));
  NOR2_X1    g1779(.A1(new_n2049_), .A2(\in1[79] ), .ZN(new_n2422_));
  NOR2_X1    g1780(.A1(new_n2062_), .A2(\in0[79] ), .ZN(new_n2423_));
  NOR2_X1    g1781(.A1(new_n2423_), .A2(new_n2422_), .ZN(new_n2424_));
  NOR2_X1    g1782(.A1(new_n2421_), .A2(new_n2424_), .ZN(new_n2425_));
  NOR2_X1    g1783(.A1(new_n2023_), .A2(\in3[78] ), .ZN(new_n2426_));
  AOI21_X1   g1784(.A1(new_n1529_), .A2(new_n2023_), .B(new_n2426_), .ZN(new_n2427_));
  NOR2_X1    g1785(.A1(new_n2049_), .A2(\in1[78] ), .ZN(new_n2428_));
  AOI21_X1   g1786(.A1(new_n810_), .A2(new_n2049_), .B(new_n2428_), .ZN(new_n2429_));
  INV_X1     g1787(.I(new_n2429_), .ZN(new_n2430_));
  AOI21_X1   g1788(.A1(new_n2427_), .A2(new_n2430_), .B(new_n2425_), .ZN(new_n2431_));
  INV_X1     g1789(.I(new_n2431_), .ZN(new_n2432_));
  INV_X1     g1790(.I(\in2[77] ), .ZN(new_n2433_));
  NOR2_X1    g1791(.A1(new_n2023_), .A2(\in3[77] ), .ZN(new_n2434_));
  AOI21_X1   g1792(.A1(new_n2433_), .A2(new_n2023_), .B(new_n2434_), .ZN(new_n2435_));
  INV_X1     g1793(.I(new_n2435_), .ZN(new_n2436_));
  NOR2_X1    g1794(.A1(new_n2049_), .A2(\in1[77] ), .ZN(new_n2437_));
  NOR2_X1    g1795(.A1(new_n2062_), .A2(\in0[77] ), .ZN(new_n2438_));
  NOR2_X1    g1796(.A1(new_n2438_), .A2(new_n2437_), .ZN(new_n2439_));
  NOR2_X1    g1797(.A1(new_n2436_), .A2(new_n2439_), .ZN(new_n2440_));
  INV_X1     g1798(.I(new_n2440_), .ZN(new_n2441_));
  INV_X1     g1799(.I(new_n2439_), .ZN(new_n2442_));
  NOR2_X1    g1800(.A1(new_n2125_), .A2(\in2[76] ), .ZN(new_n2443_));
  AOI21_X1   g1801(.A1(new_n1533_), .A2(new_n2125_), .B(new_n2443_), .ZN(new_n2444_));
  NOR2_X1    g1802(.A1(new_n2062_), .A2(\in0[76] ), .ZN(new_n2445_));
  AOI21_X1   g1803(.A1(new_n815_), .A2(new_n2062_), .B(new_n2445_), .ZN(new_n2446_));
  INV_X1     g1804(.I(new_n2446_), .ZN(new_n2447_));
  OAI22_X1   g1805(.A1(new_n2435_), .A2(new_n2442_), .B1(new_n2447_), .B2(new_n2444_), .ZN(new_n2448_));
  NAND2_X1   g1806(.A1(new_n2448_), .A2(new_n2441_), .ZN(new_n2449_));
  INV_X1     g1807(.I(new_n2424_), .ZN(new_n2450_));
  OAI22_X1   g1808(.A1(new_n2450_), .A2(new_n2420_), .B1(new_n2430_), .B2(new_n2427_), .ZN(new_n2451_));
  INV_X1     g1809(.I(new_n2451_), .ZN(new_n2452_));
  OAI22_X1   g1810(.A1(new_n2449_), .A2(new_n2432_), .B1(new_n2425_), .B2(new_n2452_), .ZN(new_n2453_));
  NAND2_X1   g1811(.A1(new_n2447_), .A2(new_n2444_), .ZN(new_n2454_));
  NAND3_X1   g1812(.A1(new_n2431_), .A2(new_n2441_), .A3(new_n2454_), .ZN(new_n2455_));
  INV_X1     g1813(.I(\in2[72] ), .ZN(new_n2456_));
  NOR2_X1    g1814(.A1(new_n2023_), .A2(\in3[72] ), .ZN(new_n2457_));
  AOI21_X1   g1815(.A1(new_n2456_), .A2(new_n2023_), .B(new_n2457_), .ZN(new_n2458_));
  INV_X1     g1816(.I(new_n2458_), .ZN(new_n2459_));
  INV_X1     g1817(.I(\in0[72] ), .ZN(new_n2460_));
  NOR2_X1    g1818(.A1(new_n2049_), .A2(\in1[72] ), .ZN(new_n2461_));
  AOI21_X1   g1819(.A1(new_n2460_), .A2(new_n2049_), .B(new_n2461_), .ZN(new_n2462_));
  NOR2_X1    g1820(.A1(new_n2459_), .A2(new_n2462_), .ZN(new_n2463_));
  NOR2_X1    g1821(.A1(new_n2023_), .A2(\in3[75] ), .ZN(new_n2464_));
  AOI21_X1   g1822(.A1(new_n1546_), .A2(new_n2023_), .B(new_n2464_), .ZN(new_n2465_));
  NOR2_X1    g1823(.A1(new_n2049_), .A2(\in1[75] ), .ZN(new_n2466_));
  AOI21_X1   g1824(.A1(new_n829_), .A2(new_n2049_), .B(new_n2466_), .ZN(new_n2467_));
  INV_X1     g1825(.I(new_n2467_), .ZN(new_n2468_));
  NOR2_X1    g1826(.A1(new_n2023_), .A2(\in3[74] ), .ZN(new_n2469_));
  AOI21_X1   g1827(.A1(new_n1545_), .A2(new_n2023_), .B(new_n2469_), .ZN(new_n2470_));
  NOR2_X1    g1828(.A1(new_n2049_), .A2(\in1[74] ), .ZN(new_n2471_));
  AOI21_X1   g1829(.A1(new_n828_), .A2(new_n2049_), .B(new_n2471_), .ZN(new_n2472_));
  INV_X1     g1830(.I(new_n2472_), .ZN(new_n2473_));
  AOI22_X1   g1831(.A1(new_n2465_), .A2(new_n2468_), .B1(new_n2473_), .B2(new_n2470_), .ZN(new_n2474_));
  INV_X1     g1832(.I(new_n2474_), .ZN(new_n2475_));
  NOR2_X1    g1833(.A1(new_n2023_), .A2(\in3[73] ), .ZN(new_n2476_));
  AOI21_X1   g1834(.A1(new_n1874_), .A2(new_n2023_), .B(new_n2476_), .ZN(new_n2477_));
  INV_X1     g1835(.I(new_n2477_), .ZN(new_n2478_));
  NOR2_X1    g1836(.A1(new_n2049_), .A2(\in1[73] ), .ZN(new_n2479_));
  NOR2_X1    g1837(.A1(new_n2062_), .A2(\in0[73] ), .ZN(new_n2480_));
  NOR2_X1    g1838(.A1(new_n2480_), .A2(new_n2479_), .ZN(new_n2481_));
  NOR2_X1    g1839(.A1(new_n2478_), .A2(new_n2481_), .ZN(new_n2482_));
  NOR3_X1    g1840(.A1(new_n2475_), .A2(new_n2463_), .A3(new_n2482_), .ZN(new_n2483_));
  NOR2_X1    g1841(.A1(new_n2023_), .A2(\in3[71] ), .ZN(new_n2484_));
  AOI21_X1   g1842(.A1(new_n1562_), .A2(new_n2023_), .B(new_n2484_), .ZN(new_n2485_));
  INV_X1     g1843(.I(new_n2485_), .ZN(new_n2486_));
  NOR2_X1    g1844(.A1(new_n2049_), .A2(\in1[71] ), .ZN(new_n2487_));
  NOR2_X1    g1845(.A1(new_n2062_), .A2(\in0[71] ), .ZN(new_n2488_));
  NOR2_X1    g1846(.A1(new_n2488_), .A2(new_n2487_), .ZN(new_n2489_));
  NOR2_X1    g1847(.A1(new_n2486_), .A2(new_n2489_), .ZN(new_n2490_));
  NOR2_X1    g1848(.A1(new_n2023_), .A2(\in3[70] ), .ZN(new_n2491_));
  AOI21_X1   g1849(.A1(new_n1555_), .A2(new_n2023_), .B(new_n2491_), .ZN(new_n2492_));
  NOR2_X1    g1850(.A1(new_n2049_), .A2(\in1[70] ), .ZN(new_n2493_));
  AOI21_X1   g1851(.A1(new_n837_), .A2(new_n2049_), .B(new_n2493_), .ZN(new_n2494_));
  INV_X1     g1852(.I(new_n2494_), .ZN(new_n2495_));
  AOI21_X1   g1853(.A1(new_n2492_), .A2(new_n2495_), .B(new_n2490_), .ZN(new_n2496_));
  INV_X1     g1854(.I(new_n2496_), .ZN(new_n2497_));
  INV_X1     g1855(.I(\in2[69] ), .ZN(new_n2498_));
  NOR2_X1    g1856(.A1(new_n2023_), .A2(\in3[69] ), .ZN(new_n2499_));
  AOI21_X1   g1857(.A1(new_n2498_), .A2(new_n2023_), .B(new_n2499_), .ZN(new_n2500_));
  INV_X1     g1858(.I(new_n2500_), .ZN(new_n2501_));
  NOR2_X1    g1859(.A1(new_n2049_), .A2(\in1[69] ), .ZN(new_n2502_));
  NOR2_X1    g1860(.A1(new_n2062_), .A2(\in0[69] ), .ZN(new_n2503_));
  NOR2_X1    g1861(.A1(new_n2503_), .A2(new_n2502_), .ZN(new_n2504_));
  NOR2_X1    g1862(.A1(new_n2501_), .A2(new_n2504_), .ZN(new_n2505_));
  INV_X1     g1863(.I(new_n2505_), .ZN(new_n2506_));
  INV_X1     g1864(.I(new_n2504_), .ZN(new_n2507_));
  NOR2_X1    g1865(.A1(new_n2125_), .A2(\in2[68] ), .ZN(new_n2508_));
  AOI21_X1   g1866(.A1(new_n1559_), .A2(new_n2125_), .B(new_n2508_), .ZN(new_n2509_));
  NOR2_X1    g1867(.A1(new_n2062_), .A2(\in0[68] ), .ZN(new_n2510_));
  AOI21_X1   g1868(.A1(new_n842_), .A2(new_n2062_), .B(new_n2510_), .ZN(new_n2511_));
  INV_X1     g1869(.I(new_n2511_), .ZN(new_n2512_));
  OAI22_X1   g1870(.A1(new_n2500_), .A2(new_n2507_), .B1(new_n2512_), .B2(new_n2509_), .ZN(new_n2513_));
  NAND2_X1   g1871(.A1(new_n2513_), .A2(new_n2506_), .ZN(new_n2514_));
  INV_X1     g1872(.I(new_n2489_), .ZN(new_n2515_));
  OAI22_X1   g1873(.A1(new_n2515_), .A2(new_n2485_), .B1(new_n2495_), .B2(new_n2492_), .ZN(new_n2516_));
  INV_X1     g1874(.I(new_n2516_), .ZN(new_n2517_));
  OAI22_X1   g1875(.A1(new_n2514_), .A2(new_n2497_), .B1(new_n2490_), .B2(new_n2517_), .ZN(new_n2518_));
  NOR2_X1    g1876(.A1(new_n2023_), .A2(\in3[67] ), .ZN(new_n2519_));
  AOI21_X1   g1877(.A1(new_n1567_), .A2(new_n2023_), .B(new_n2519_), .ZN(new_n2520_));
  INV_X1     g1878(.I(new_n2520_), .ZN(new_n2521_));
  NOR2_X1    g1879(.A1(new_n2049_), .A2(\in1[67] ), .ZN(new_n2522_));
  AOI21_X1   g1880(.A1(new_n852_), .A2(new_n2049_), .B(new_n2522_), .ZN(new_n2523_));
  INV_X1     g1881(.I(new_n2523_), .ZN(new_n2524_));
  NOR2_X1    g1882(.A1(new_n2023_), .A2(\in3[66] ), .ZN(new_n2525_));
  AOI21_X1   g1883(.A1(new_n1566_), .A2(new_n2023_), .B(new_n2525_), .ZN(new_n2526_));
  NOR2_X1    g1884(.A1(new_n2049_), .A2(\in1[66] ), .ZN(new_n2527_));
  AOI21_X1   g1885(.A1(new_n851_), .A2(new_n2049_), .B(new_n2527_), .ZN(new_n2528_));
  INV_X1     g1886(.I(new_n2528_), .ZN(new_n2529_));
  AOI22_X1   g1887(.A1(new_n2520_), .A2(new_n2524_), .B1(new_n2529_), .B2(new_n2526_), .ZN(new_n2530_));
  NOR2_X1    g1888(.A1(new_n2023_), .A2(\in3[65] ), .ZN(new_n2531_));
  AOI21_X1   g1889(.A1(new_n1569_), .A2(new_n2023_), .B(new_n2531_), .ZN(new_n2532_));
  INV_X1     g1890(.I(new_n2532_), .ZN(new_n2533_));
  NOR2_X1    g1891(.A1(new_n2049_), .A2(\in1[65] ), .ZN(new_n2534_));
  NOR2_X1    g1892(.A1(new_n2062_), .A2(\in0[65] ), .ZN(new_n2535_));
  NOR2_X1    g1893(.A1(new_n2535_), .A2(new_n2534_), .ZN(new_n2536_));
  NOR2_X1    g1894(.A1(new_n2533_), .A2(new_n2536_), .ZN(new_n2537_));
  NOR2_X1    g1895(.A1(new_n2023_), .A2(\in3[64] ), .ZN(new_n2538_));
  AOI21_X1   g1896(.A1(new_n1571_), .A2(new_n2023_), .B(new_n2538_), .ZN(new_n2539_));
  INV_X1     g1897(.I(new_n2539_), .ZN(new_n2540_));
  INV_X1     g1898(.I(\in0[64] ), .ZN(new_n2541_));
  NOR2_X1    g1899(.A1(new_n2049_), .A2(\in1[64] ), .ZN(new_n2542_));
  AOI21_X1   g1900(.A1(new_n2541_), .A2(new_n2049_), .B(new_n2542_), .ZN(new_n2543_));
  AOI22_X1   g1901(.A1(new_n2533_), .A2(new_n2536_), .B1(new_n2540_), .B2(new_n2543_), .ZN(new_n2544_));
  OAI22_X1   g1902(.A1(new_n2544_), .A2(new_n2537_), .B1(new_n2526_), .B2(new_n2529_), .ZN(new_n2545_));
  AOI22_X1   g1903(.A1(new_n2545_), .A2(new_n2530_), .B1(new_n2521_), .B2(new_n2523_), .ZN(new_n2546_));
  INV_X1     g1904(.I(new_n2530_), .ZN(new_n2547_));
  NOR2_X1    g1905(.A1(new_n2540_), .A2(new_n2543_), .ZN(new_n2548_));
  NOR3_X1    g1906(.A1(new_n2547_), .A2(new_n2537_), .A3(new_n2548_), .ZN(new_n2549_));
  NOR2_X1    g1907(.A1(new_n2023_), .A2(\in3[57] ), .ZN(new_n2550_));
  AOI21_X1   g1908(.A1(new_n1582_), .A2(new_n2023_), .B(new_n2550_), .ZN(new_n2551_));
  INV_X1     g1909(.I(new_n2551_), .ZN(new_n2552_));
  NOR2_X1    g1910(.A1(new_n2049_), .A2(\in1[57] ), .ZN(new_n2553_));
  AOI21_X1   g1911(.A1(new_n867_), .A2(new_n2049_), .B(new_n2553_), .ZN(new_n2554_));
  NOR2_X1    g1912(.A1(new_n2552_), .A2(new_n2554_), .ZN(new_n2555_));
  NOR2_X1    g1913(.A1(new_n2023_), .A2(\in3[56] ), .ZN(new_n2556_));
  AOI21_X1   g1914(.A1(new_n1581_), .A2(new_n2023_), .B(new_n2556_), .ZN(new_n2557_));
  NOR2_X1    g1915(.A1(new_n2049_), .A2(\in1[56] ), .ZN(new_n2558_));
  AOI21_X1   g1916(.A1(new_n866_), .A2(new_n2049_), .B(new_n2558_), .ZN(new_n2559_));
  INV_X1     g1917(.I(new_n2559_), .ZN(new_n2560_));
  AOI21_X1   g1918(.A1(new_n2557_), .A2(new_n2560_), .B(new_n2555_), .ZN(new_n2561_));
  NOR2_X1    g1919(.A1(new_n2023_), .A2(\in3[61] ), .ZN(new_n2562_));
  AOI21_X1   g1920(.A1(new_n1590_), .A2(new_n2023_), .B(new_n2562_), .ZN(new_n2563_));
  INV_X1     g1921(.I(new_n2563_), .ZN(new_n2564_));
  NOR2_X1    g1922(.A1(new_n2049_), .A2(\in1[61] ), .ZN(new_n2565_));
  AOI21_X1   g1923(.A1(new_n874_), .A2(new_n2049_), .B(new_n2565_), .ZN(new_n2566_));
  NOR2_X1    g1924(.A1(new_n2564_), .A2(new_n2566_), .ZN(new_n2567_));
  NOR2_X1    g1925(.A1(new_n2023_), .A2(\in3[63] ), .ZN(new_n2568_));
  AOI21_X1   g1926(.A1(new_n1862_), .A2(new_n2023_), .B(new_n2568_), .ZN(new_n2569_));
  INV_X1     g1927(.I(new_n2569_), .ZN(new_n2570_));
  NOR2_X1    g1928(.A1(new_n2049_), .A2(\in1[63] ), .ZN(new_n2571_));
  NOR2_X1    g1929(.A1(new_n2062_), .A2(\in0[63] ), .ZN(new_n2572_));
  NOR2_X1    g1930(.A1(new_n2572_), .A2(new_n2571_), .ZN(new_n2573_));
  NOR2_X1    g1931(.A1(new_n2570_), .A2(new_n2573_), .ZN(new_n2574_));
  NOR2_X1    g1932(.A1(new_n2023_), .A2(\in3[62] ), .ZN(new_n2575_));
  AOI21_X1   g1933(.A1(new_n1584_), .A2(new_n2023_), .B(new_n2575_), .ZN(new_n2576_));
  NOR2_X1    g1934(.A1(new_n2049_), .A2(\in1[62] ), .ZN(new_n2577_));
  AOI21_X1   g1935(.A1(new_n869_), .A2(new_n2049_), .B(new_n2577_), .ZN(new_n2578_));
  INV_X1     g1936(.I(new_n2578_), .ZN(new_n2579_));
  AOI21_X1   g1937(.A1(new_n2576_), .A2(new_n2579_), .B(new_n2574_), .ZN(new_n2580_));
  INV_X1     g1938(.I(new_n2580_), .ZN(new_n2581_));
  NOR2_X1    g1939(.A1(new_n2023_), .A2(\in3[60] ), .ZN(new_n2582_));
  AOI21_X1   g1940(.A1(new_n1588_), .A2(new_n2023_), .B(new_n2582_), .ZN(new_n2583_));
  INV_X1     g1941(.I(new_n2583_), .ZN(new_n2584_));
  NOR2_X1    g1942(.A1(new_n2049_), .A2(\in1[60] ), .ZN(new_n2585_));
  AOI21_X1   g1943(.A1(new_n873_), .A2(new_n2049_), .B(new_n2585_), .ZN(new_n2586_));
  NOR2_X1    g1944(.A1(new_n2584_), .A2(new_n2586_), .ZN(new_n2587_));
  NOR3_X1    g1945(.A1(new_n2581_), .A2(new_n2567_), .A3(new_n2587_), .ZN(new_n2588_));
  NOR2_X1    g1946(.A1(new_n2023_), .A2(\in3[59] ), .ZN(new_n2589_));
  AOI21_X1   g1947(.A1(new_n1595_), .A2(new_n2023_), .B(new_n2589_), .ZN(new_n2590_));
  NOR2_X1    g1948(.A1(new_n2049_), .A2(\in1[59] ), .ZN(new_n2591_));
  AOI21_X1   g1949(.A1(new_n879_), .A2(new_n2049_), .B(new_n2591_), .ZN(new_n2592_));
  INV_X1     g1950(.I(new_n2592_), .ZN(new_n2593_));
  NOR2_X1    g1951(.A1(new_n2023_), .A2(\in3[58] ), .ZN(new_n2594_));
  AOI21_X1   g1952(.A1(new_n1594_), .A2(new_n2023_), .B(new_n2594_), .ZN(new_n2595_));
  NOR2_X1    g1953(.A1(new_n2049_), .A2(\in1[58] ), .ZN(new_n2596_));
  AOI21_X1   g1954(.A1(new_n878_), .A2(new_n2049_), .B(new_n2596_), .ZN(new_n2597_));
  INV_X1     g1955(.I(new_n2597_), .ZN(new_n2598_));
  AOI22_X1   g1956(.A1(new_n2590_), .A2(new_n2593_), .B1(new_n2598_), .B2(new_n2595_), .ZN(new_n2599_));
  NAND3_X1   g1957(.A1(new_n2588_), .A2(new_n2561_), .A3(new_n2599_), .ZN(new_n2600_));
  NOR2_X1    g1958(.A1(new_n2023_), .A2(\in3[55] ), .ZN(new_n2601_));
  AOI21_X1   g1959(.A1(new_n1601_), .A2(new_n2023_), .B(new_n2601_), .ZN(new_n2602_));
  INV_X1     g1960(.I(new_n2602_), .ZN(new_n2603_));
  NOR2_X1    g1961(.A1(new_n2049_), .A2(\in1[55] ), .ZN(new_n2604_));
  AOI21_X1   g1962(.A1(new_n885_), .A2(new_n2049_), .B(new_n2604_), .ZN(new_n2605_));
  INV_X1     g1963(.I(new_n2605_), .ZN(new_n2606_));
  NOR2_X1    g1964(.A1(new_n2023_), .A2(\in3[54] ), .ZN(new_n2607_));
  AOI21_X1   g1965(.A1(new_n1600_), .A2(new_n2023_), .B(new_n2607_), .ZN(new_n2608_));
  NOR2_X1    g1966(.A1(new_n2049_), .A2(\in1[54] ), .ZN(new_n2609_));
  AOI21_X1   g1967(.A1(new_n884_), .A2(new_n2049_), .B(new_n2609_), .ZN(new_n2610_));
  INV_X1     g1968(.I(new_n2610_), .ZN(new_n2611_));
  AOI22_X1   g1969(.A1(new_n2602_), .A2(new_n2606_), .B1(new_n2611_), .B2(new_n2608_), .ZN(new_n2612_));
  NOR2_X1    g1970(.A1(new_n2023_), .A2(\in3[53] ), .ZN(new_n2613_));
  AOI21_X1   g1971(.A1(new_n1621_), .A2(new_n2023_), .B(new_n2613_), .ZN(new_n2614_));
  INV_X1     g1972(.I(new_n2614_), .ZN(new_n2615_));
  NOR2_X1    g1973(.A1(new_n2049_), .A2(\in1[53] ), .ZN(new_n2616_));
  NOR2_X1    g1974(.A1(new_n2062_), .A2(\in0[53] ), .ZN(new_n2617_));
  NOR2_X1    g1975(.A1(new_n2617_), .A2(new_n2616_), .ZN(new_n2618_));
  NOR2_X1    g1976(.A1(new_n2615_), .A2(new_n2618_), .ZN(new_n2619_));
  INV_X1     g1977(.I(\in2[52] ), .ZN(new_n2620_));
  NOR2_X1    g1978(.A1(new_n2023_), .A2(\in3[52] ), .ZN(new_n2621_));
  AOI21_X1   g1979(.A1(new_n2620_), .A2(new_n2023_), .B(new_n2621_), .ZN(new_n2622_));
  INV_X1     g1980(.I(new_n2622_), .ZN(new_n2623_));
  NOR2_X1    g1981(.A1(new_n2049_), .A2(\in1[52] ), .ZN(new_n2624_));
  NOR2_X1    g1982(.A1(new_n2062_), .A2(\in0[52] ), .ZN(new_n2625_));
  NOR2_X1    g1983(.A1(new_n2625_), .A2(new_n2624_), .ZN(new_n2626_));
  AOI22_X1   g1984(.A1(new_n2615_), .A2(new_n2618_), .B1(new_n2623_), .B2(new_n2626_), .ZN(new_n2627_));
  OAI22_X1   g1985(.A1(new_n2627_), .A2(new_n2619_), .B1(new_n2608_), .B2(new_n2611_), .ZN(new_n2628_));
  AOI22_X1   g1986(.A1(new_n2628_), .A2(new_n2612_), .B1(new_n2603_), .B2(new_n2605_), .ZN(new_n2629_));
  INV_X1     g1987(.I(new_n2612_), .ZN(new_n2630_));
  NOR2_X1    g1988(.A1(new_n2623_), .A2(new_n2626_), .ZN(new_n2631_));
  NOR3_X1    g1989(.A1(new_n2630_), .A2(new_n2619_), .A3(new_n2631_), .ZN(new_n2632_));
  NOR2_X1    g1990(.A1(new_n2023_), .A2(\in3[49] ), .ZN(new_n2633_));
  AOI21_X1   g1991(.A1(new_n1611_), .A2(new_n2023_), .B(new_n2633_), .ZN(new_n2634_));
  INV_X1     g1992(.I(new_n2634_), .ZN(new_n2635_));
  NOR2_X1    g1993(.A1(new_n2049_), .A2(\in1[49] ), .ZN(new_n2636_));
  NOR2_X1    g1994(.A1(new_n2062_), .A2(\in0[49] ), .ZN(new_n2637_));
  NOR2_X1    g1995(.A1(new_n2637_), .A2(new_n2636_), .ZN(new_n2638_));
  NOR2_X1    g1996(.A1(new_n2023_), .A2(\in3[51] ), .ZN(new_n2639_));
  AOI21_X1   g1997(.A1(new_n1609_), .A2(new_n2023_), .B(new_n2639_), .ZN(new_n2640_));
  INV_X1     g1998(.I(new_n2640_), .ZN(new_n2641_));
  NOR2_X1    g1999(.A1(new_n2049_), .A2(\in1[51] ), .ZN(new_n2642_));
  AOI21_X1   g2000(.A1(new_n892_), .A2(new_n2049_), .B(new_n2642_), .ZN(new_n2643_));
  OAI22_X1   g2001(.A1(new_n2635_), .A2(new_n2638_), .B1(new_n2641_), .B2(new_n2643_), .ZN(new_n2644_));
  NOR2_X1    g2002(.A1(new_n2049_), .A2(\in1[50] ), .ZN(new_n2645_));
  AOI21_X1   g2003(.A1(new_n891_), .A2(new_n2049_), .B(new_n2645_), .ZN(new_n2646_));
  INV_X1     g2004(.I(new_n2646_), .ZN(new_n2647_));
  NOR2_X1    g2005(.A1(new_n2023_), .A2(\in3[50] ), .ZN(new_n2648_));
  AOI21_X1   g2006(.A1(new_n1608_), .A2(new_n2023_), .B(new_n2648_), .ZN(new_n2649_));
  AOI21_X1   g2007(.A1(new_n2647_), .A2(new_n2649_), .B(new_n2644_), .ZN(new_n2650_));
  INV_X1     g2008(.I(new_n2650_), .ZN(new_n2651_));
  NOR2_X1    g2009(.A1(new_n2049_), .A2(\in1[48] ), .ZN(new_n2652_));
  AOI21_X1   g2010(.A1(new_n898_), .A2(new_n2049_), .B(new_n2652_), .ZN(new_n2653_));
  NOR2_X1    g2011(.A1(new_n2023_), .A2(\in3[48] ), .ZN(new_n2654_));
  AOI21_X1   g2012(.A1(new_n1613_), .A2(new_n2023_), .B(new_n2654_), .ZN(new_n2655_));
  INV_X1     g2013(.I(new_n2655_), .ZN(new_n2656_));
  AOI22_X1   g2014(.A1(new_n2635_), .A2(new_n2638_), .B1(new_n2656_), .B2(new_n2653_), .ZN(new_n2657_));
  NOR2_X1    g2015(.A1(new_n2651_), .A2(new_n2657_), .ZN(new_n2658_));
  INV_X1     g2016(.I(new_n2643_), .ZN(new_n2659_));
  INV_X1     g2017(.I(new_n2649_), .ZN(new_n2660_));
  AOI22_X1   g2018(.A1(new_n2641_), .A2(new_n2643_), .B1(new_n2660_), .B2(new_n2646_), .ZN(new_n2661_));
  AOI21_X1   g2019(.A1(new_n2640_), .A2(new_n2659_), .B(new_n2661_), .ZN(new_n2662_));
  OAI21_X1   g2020(.A1(new_n2658_), .A2(new_n2662_), .B(new_n2632_), .ZN(new_n2663_));
  NAND2_X1   g2021(.A1(new_n2663_), .A2(new_n2629_), .ZN(new_n2664_));
  INV_X1     g2022(.I(new_n2664_), .ZN(new_n2665_));
  NOR2_X1    g2023(.A1(new_n2023_), .A2(\in3[47] ), .ZN(new_n2666_));
  AOI21_X1   g2024(.A1(new_n1653_), .A2(new_n2023_), .B(new_n2666_), .ZN(new_n2667_));
  INV_X1     g2025(.I(new_n2667_), .ZN(new_n2668_));
  NOR2_X1    g2026(.A1(new_n2049_), .A2(\in1[47] ), .ZN(new_n2669_));
  NOR2_X1    g2027(.A1(new_n2062_), .A2(\in0[47] ), .ZN(new_n2670_));
  NOR2_X1    g2028(.A1(new_n2670_), .A2(new_n2669_), .ZN(new_n2671_));
  NOR2_X1    g2029(.A1(new_n2668_), .A2(new_n2671_), .ZN(new_n2672_));
  NOR2_X1    g2030(.A1(new_n2023_), .A2(\in3[46] ), .ZN(new_n2673_));
  AOI21_X1   g2031(.A1(new_n1628_), .A2(new_n2023_), .B(new_n2673_), .ZN(new_n2674_));
  NOR2_X1    g2032(.A1(new_n2049_), .A2(\in1[46] ), .ZN(new_n2675_));
  AOI21_X1   g2033(.A1(new_n914_), .A2(new_n2049_), .B(new_n2675_), .ZN(new_n2676_));
  INV_X1     g2034(.I(new_n2676_), .ZN(new_n2677_));
  AOI21_X1   g2035(.A1(new_n2674_), .A2(new_n2677_), .B(new_n2672_), .ZN(new_n2678_));
  INV_X1     g2036(.I(new_n2678_), .ZN(new_n2679_));
  NOR2_X1    g2037(.A1(new_n2023_), .A2(\in3[45] ), .ZN(new_n2680_));
  AOI21_X1   g2038(.A1(new_n1634_), .A2(new_n2023_), .B(new_n2680_), .ZN(new_n2681_));
  INV_X1     g2039(.I(new_n2681_), .ZN(new_n2682_));
  NOR2_X1    g2040(.A1(new_n2049_), .A2(\in1[45] ), .ZN(new_n2683_));
  AOI21_X1   g2041(.A1(new_n919_), .A2(new_n2049_), .B(new_n2683_), .ZN(new_n2684_));
  NAND2_X1   g2042(.A1(new_n2682_), .A2(new_n2684_), .ZN(new_n2685_));
  NOR2_X1    g2043(.A1(new_n2682_), .A2(new_n2684_), .ZN(new_n2686_));
  NOR2_X1    g2044(.A1(new_n2023_), .A2(\in3[44] ), .ZN(new_n2687_));
  AOI21_X1   g2045(.A1(new_n1632_), .A2(new_n2023_), .B(new_n2687_), .ZN(new_n2688_));
  NOR2_X1    g2046(.A1(new_n2049_), .A2(\in1[44] ), .ZN(new_n2689_));
  AOI21_X1   g2047(.A1(new_n918_), .A2(new_n2049_), .B(new_n2689_), .ZN(new_n2690_));
  INV_X1     g2048(.I(new_n2690_), .ZN(new_n2691_));
  OR3_X2     g2049(.A1(new_n2686_), .A2(new_n2688_), .A3(new_n2691_), .Z(new_n2692_));
  AOI21_X1   g2050(.A1(new_n2685_), .A2(new_n2692_), .B(new_n2679_), .ZN(new_n2693_));
  INV_X1     g2051(.I(new_n2688_), .ZN(new_n2694_));
  NOR2_X1    g2052(.A1(new_n2694_), .A2(new_n2690_), .ZN(new_n2695_));
  NOR2_X1    g2053(.A1(new_n2023_), .A2(\in3[43] ), .ZN(new_n2696_));
  AOI21_X1   g2054(.A1(new_n1638_), .A2(new_n2023_), .B(new_n2696_), .ZN(new_n2697_));
  INV_X1     g2055(.I(new_n2697_), .ZN(new_n2698_));
  NOR2_X1    g2056(.A1(new_n2049_), .A2(\in1[43] ), .ZN(new_n2699_));
  AOI21_X1   g2057(.A1(new_n923_), .A2(new_n2049_), .B(new_n2699_), .ZN(new_n2700_));
  INV_X1     g2058(.I(new_n2700_), .ZN(new_n2701_));
  NOR2_X1    g2059(.A1(new_n2023_), .A2(\in3[42] ), .ZN(new_n2702_));
  AOI21_X1   g2060(.A1(new_n1639_), .A2(new_n2023_), .B(new_n2702_), .ZN(new_n2703_));
  NOR2_X1    g2061(.A1(new_n2049_), .A2(\in1[42] ), .ZN(new_n2704_));
  AOI21_X1   g2062(.A1(new_n924_), .A2(new_n2049_), .B(new_n2704_), .ZN(new_n2705_));
  INV_X1     g2063(.I(new_n2705_), .ZN(new_n2706_));
  AOI22_X1   g2064(.A1(new_n2697_), .A2(new_n2701_), .B1(new_n2706_), .B2(new_n2703_), .ZN(new_n2707_));
  NOR2_X1    g2065(.A1(new_n2023_), .A2(\in3[41] ), .ZN(new_n2708_));
  AOI21_X1   g2066(.A1(new_n1643_), .A2(new_n2023_), .B(new_n2708_), .ZN(new_n2709_));
  INV_X1     g2067(.I(new_n2709_), .ZN(new_n2710_));
  NOR2_X1    g2068(.A1(new_n2049_), .A2(\in1[41] ), .ZN(new_n2711_));
  AOI21_X1   g2069(.A1(new_n928_), .A2(new_n2049_), .B(new_n2711_), .ZN(new_n2712_));
  NOR2_X1    g2070(.A1(new_n2710_), .A2(new_n2712_), .ZN(new_n2713_));
  NOR2_X1    g2071(.A1(new_n2023_), .A2(\in3[40] ), .ZN(new_n2714_));
  AOI21_X1   g2072(.A1(new_n1645_), .A2(new_n2023_), .B(new_n2714_), .ZN(new_n2715_));
  INV_X1     g2073(.I(new_n2715_), .ZN(new_n2716_));
  NOR2_X1    g2074(.A1(new_n2049_), .A2(\in1[40] ), .ZN(new_n2717_));
  AOI21_X1   g2075(.A1(new_n930_), .A2(new_n2049_), .B(new_n2717_), .ZN(new_n2718_));
  AOI22_X1   g2076(.A1(new_n2710_), .A2(new_n2712_), .B1(new_n2716_), .B2(new_n2718_), .ZN(new_n2719_));
  OAI22_X1   g2077(.A1(new_n2719_), .A2(new_n2713_), .B1(new_n2703_), .B2(new_n2706_), .ZN(new_n2720_));
  AOI22_X1   g2078(.A1(new_n2720_), .A2(new_n2707_), .B1(new_n2698_), .B2(new_n2700_), .ZN(new_n2721_));
  NOR4_X1    g2079(.A1(new_n2721_), .A2(new_n2679_), .A3(new_n2686_), .A4(new_n2695_), .ZN(new_n2722_));
  INV_X1     g2080(.I(new_n2674_), .ZN(new_n2723_));
  AOI22_X1   g2081(.A1(new_n2668_), .A2(new_n2671_), .B1(new_n2723_), .B2(new_n2676_), .ZN(new_n2724_));
  NOR2_X1    g2082(.A1(new_n2724_), .A2(new_n2672_), .ZN(new_n2725_));
  NOR3_X1    g2083(.A1(new_n2722_), .A2(new_n2693_), .A3(new_n2725_), .ZN(new_n2726_));
  INV_X1     g2084(.I(new_n2726_), .ZN(new_n2727_));
  NOR3_X1    g2085(.A1(new_n2679_), .A2(new_n2686_), .A3(new_n2695_), .ZN(new_n2728_));
  INV_X1     g2086(.I(new_n2718_), .ZN(new_n2729_));
  AOI21_X1   g2087(.A1(new_n2715_), .A2(new_n2729_), .B(new_n2713_), .ZN(new_n2730_));
  NAND3_X1   g2088(.A1(new_n2728_), .A2(new_n2707_), .A3(new_n2730_), .ZN(new_n2731_));
  NOR2_X1    g2089(.A1(new_n2023_), .A2(\in3[33] ), .ZN(new_n2732_));
  AOI21_X1   g2090(.A1(new_n1660_), .A2(new_n2023_), .B(new_n2732_), .ZN(new_n2733_));
  INV_X1     g2091(.I(new_n2733_), .ZN(new_n2734_));
  NOR2_X1    g2092(.A1(new_n2049_), .A2(\in1[33] ), .ZN(new_n2735_));
  AOI21_X1   g2093(.A1(new_n947_), .A2(new_n2049_), .B(new_n2735_), .ZN(new_n2736_));
  NOR2_X1    g2094(.A1(new_n2023_), .A2(\in3[35] ), .ZN(new_n2737_));
  AOI21_X1   g2095(.A1(new_n1673_), .A2(new_n2023_), .B(new_n2737_), .ZN(new_n2738_));
  INV_X1     g2096(.I(new_n2738_), .ZN(new_n2739_));
  NOR2_X1    g2097(.A1(new_n2049_), .A2(\in1[35] ), .ZN(new_n2740_));
  AOI21_X1   g2098(.A1(new_n959_), .A2(new_n2049_), .B(new_n2740_), .ZN(new_n2741_));
  OAI22_X1   g2099(.A1(new_n2734_), .A2(new_n2736_), .B1(new_n2739_), .B2(new_n2741_), .ZN(new_n2742_));
  NOR2_X1    g2100(.A1(new_n2049_), .A2(\in1[34] ), .ZN(new_n2743_));
  AOI21_X1   g2101(.A1(new_n958_), .A2(new_n2049_), .B(new_n2743_), .ZN(new_n2744_));
  INV_X1     g2102(.I(new_n2744_), .ZN(new_n2745_));
  NOR2_X1    g2103(.A1(new_n2023_), .A2(\in3[34] ), .ZN(new_n2746_));
  AOI21_X1   g2104(.A1(new_n1672_), .A2(new_n2023_), .B(new_n2746_), .ZN(new_n2747_));
  AOI21_X1   g2105(.A1(new_n2745_), .A2(new_n2747_), .B(new_n2742_), .ZN(new_n2748_));
  INV_X1     g2106(.I(new_n2748_), .ZN(new_n2749_));
  NOR2_X1    g2107(.A1(new_n2023_), .A2(\in3[37] ), .ZN(new_n2750_));
  AOI21_X1   g2108(.A1(new_n1668_), .A2(new_n2023_), .B(new_n2750_), .ZN(new_n2751_));
  INV_X1     g2109(.I(new_n2751_), .ZN(new_n2752_));
  NOR2_X1    g2110(.A1(new_n2049_), .A2(\in1[37] ), .ZN(new_n2753_));
  AOI21_X1   g2111(.A1(new_n954_), .A2(new_n2049_), .B(new_n2753_), .ZN(new_n2754_));
  NOR2_X1    g2112(.A1(new_n2752_), .A2(new_n2754_), .ZN(new_n2755_));
  NOR2_X1    g2113(.A1(new_n2023_), .A2(\in3[39] ), .ZN(new_n2756_));
  AOI21_X1   g2114(.A1(new_n1841_), .A2(new_n2023_), .B(new_n2756_), .ZN(new_n2757_));
  NOR2_X1    g2115(.A1(new_n2062_), .A2(\in0[39] ), .ZN(new_n2758_));
  AOI21_X1   g2116(.A1(new_n950_), .A2(new_n2062_), .B(new_n2758_), .ZN(new_n2759_));
  INV_X1     g2117(.I(new_n2759_), .ZN(new_n2760_));
  NOR2_X1    g2118(.A1(new_n2023_), .A2(\in3[38] ), .ZN(new_n2761_));
  AOI21_X1   g2119(.A1(new_n1662_), .A2(new_n2023_), .B(new_n2761_), .ZN(new_n2762_));
  NOR2_X1    g2120(.A1(new_n2049_), .A2(\in1[38] ), .ZN(new_n2763_));
  AOI21_X1   g2121(.A1(new_n949_), .A2(new_n2049_), .B(new_n2763_), .ZN(new_n2764_));
  INV_X1     g2122(.I(new_n2764_), .ZN(new_n2765_));
  AOI22_X1   g2123(.A1(new_n2760_), .A2(new_n2757_), .B1(new_n2762_), .B2(new_n2765_), .ZN(new_n2766_));
  INV_X1     g2124(.I(new_n2766_), .ZN(new_n2767_));
  NOR2_X1    g2125(.A1(new_n2023_), .A2(\in3[36] ), .ZN(new_n2768_));
  AOI21_X1   g2126(.A1(new_n1666_), .A2(new_n2023_), .B(new_n2768_), .ZN(new_n2769_));
  INV_X1     g2127(.I(new_n2769_), .ZN(new_n2770_));
  NOR2_X1    g2128(.A1(new_n2049_), .A2(\in1[36] ), .ZN(new_n2771_));
  AOI21_X1   g2129(.A1(new_n953_), .A2(new_n2049_), .B(new_n2771_), .ZN(new_n2772_));
  NOR2_X1    g2130(.A1(new_n2770_), .A2(new_n2772_), .ZN(new_n2773_));
  NOR3_X1    g2131(.A1(new_n2767_), .A2(new_n2755_), .A3(new_n2773_), .ZN(new_n2774_));
  INV_X1     g2132(.I(new_n2774_), .ZN(new_n2775_));
  NOR2_X1    g2133(.A1(new_n2049_), .A2(\in1[32] ), .ZN(new_n2776_));
  AOI21_X1   g2134(.A1(new_n946_), .A2(new_n2049_), .B(new_n2776_), .ZN(new_n2777_));
  NOR2_X1    g2135(.A1(new_n2023_), .A2(\in3[32] ), .ZN(new_n2778_));
  AOI21_X1   g2136(.A1(new_n1659_), .A2(new_n2023_), .B(new_n2778_), .ZN(new_n2779_));
  INV_X1     g2137(.I(new_n2779_), .ZN(new_n2780_));
  NOR2_X1    g2138(.A1(new_n2780_), .A2(new_n2777_), .ZN(new_n2781_));
  NOR3_X1    g2139(.A1(new_n2775_), .A2(new_n2749_), .A3(new_n2781_), .ZN(new_n2782_));
  NOR2_X1    g2140(.A1(new_n2049_), .A2(\in1[30] ), .ZN(new_n2783_));
  AOI21_X1   g2141(.A1(new_n1245_), .A2(new_n2049_), .B(new_n2783_), .ZN(new_n2784_));
  NOR2_X1    g2142(.A1(new_n2023_), .A2(\in3[30] ), .ZN(new_n2785_));
  AOI21_X1   g2143(.A1(new_n1946_), .A2(new_n2023_), .B(new_n2785_), .ZN(new_n2786_));
  INV_X1     g2144(.I(new_n2786_), .ZN(new_n2787_));
  NOR2_X1    g2145(.A1(new_n2023_), .A2(\in3[29] ), .ZN(new_n2788_));
  AOI21_X1   g2146(.A1(new_n1677_), .A2(new_n2023_), .B(new_n2788_), .ZN(new_n2789_));
  INV_X1     g2147(.I(new_n2789_), .ZN(new_n2790_));
  NOR2_X1    g2148(.A1(new_n2049_), .A2(\in1[29] ), .ZN(new_n2791_));
  AOI21_X1   g2149(.A1(new_n963_), .A2(new_n2049_), .B(new_n2791_), .ZN(new_n2792_));
  NOR2_X1    g2150(.A1(new_n2790_), .A2(new_n2792_), .ZN(new_n2793_));
  NOR2_X1    g2151(.A1(new_n2049_), .A2(\in1[27] ), .ZN(new_n2794_));
  AOI21_X1   g2152(.A1(new_n1247_), .A2(new_n2049_), .B(new_n2794_), .ZN(new_n2795_));
  INV_X1     g2153(.I(new_n2795_), .ZN(new_n2796_));
  INV_X1     g2154(.I(\in2[27] ), .ZN(new_n2797_));
  NOR2_X1    g2155(.A1(new_n2023_), .A2(\in3[27] ), .ZN(new_n2798_));
  AOI21_X1   g2156(.A1(new_n2797_), .A2(new_n2023_), .B(new_n2798_), .ZN(new_n2799_));
  INV_X1     g2157(.I(new_n2799_), .ZN(new_n2800_));
  NOR2_X1    g2158(.A1(new_n2023_), .A2(\in3[26] ), .ZN(new_n2801_));
  AOI21_X1   g2159(.A1(new_n1682_), .A2(new_n2023_), .B(new_n2801_), .ZN(new_n2802_));
  INV_X1     g2160(.I(new_n2802_), .ZN(new_n2803_));
  NOR2_X1    g2161(.A1(new_n2049_), .A2(\in1[26] ), .ZN(new_n2804_));
  AOI21_X1   g2162(.A1(new_n970_), .A2(new_n2049_), .B(new_n2804_), .ZN(new_n2805_));
  NOR2_X1    g2163(.A1(new_n2803_), .A2(new_n2805_), .ZN(new_n2806_));
  NOR2_X1    g2164(.A1(new_n2023_), .A2(\in3[24] ), .ZN(new_n2807_));
  AOI21_X1   g2165(.A1(new_n1803_), .A2(new_n2023_), .B(new_n2807_), .ZN(new_n2808_));
  INV_X1     g2166(.I(new_n2808_), .ZN(new_n2809_));
  NOR2_X1    g2167(.A1(new_n2049_), .A2(\in1[24] ), .ZN(new_n2810_));
  AOI21_X1   g2168(.A1(new_n1098_), .A2(new_n2049_), .B(new_n2810_), .ZN(new_n2811_));
  NOR2_X1    g2169(.A1(new_n2809_), .A2(new_n2811_), .ZN(new_n2812_));
  INV_X1     g2170(.I(new_n2812_), .ZN(new_n2813_));
  NOR2_X1    g2171(.A1(new_n2023_), .A2(\in3[23] ), .ZN(new_n2814_));
  AOI21_X1   g2172(.A1(new_n1800_), .A2(new_n2023_), .B(new_n2814_), .ZN(new_n2815_));
  INV_X1     g2173(.I(new_n2815_), .ZN(new_n2816_));
  NOR2_X1    g2174(.A1(new_n2049_), .A2(\in1[23] ), .ZN(new_n2817_));
  AOI21_X1   g2175(.A1(new_n1095_), .A2(new_n2049_), .B(new_n2817_), .ZN(new_n2818_));
  NOR2_X1    g2176(.A1(new_n2816_), .A2(new_n2818_), .ZN(new_n2819_));
  NOR2_X1    g2177(.A1(new_n2049_), .A2(\in1[22] ), .ZN(new_n2820_));
  AOI21_X1   g2178(.A1(new_n980_), .A2(new_n2049_), .B(new_n2820_), .ZN(new_n2821_));
  INV_X1     g2179(.I(new_n2821_), .ZN(new_n2822_));
  NOR2_X1    g2180(.A1(new_n2023_), .A2(\in3[22] ), .ZN(new_n2823_));
  AOI21_X1   g2181(.A1(new_n1692_), .A2(new_n2023_), .B(new_n2823_), .ZN(new_n2824_));
  NOR2_X1    g2182(.A1(new_n2023_), .A2(\in3[21] ), .ZN(new_n2825_));
  AOI21_X1   g2183(.A1(new_n1694_), .A2(new_n2023_), .B(new_n2825_), .ZN(new_n2826_));
  INV_X1     g2184(.I(new_n2826_), .ZN(new_n2827_));
  NOR2_X1    g2185(.A1(new_n2049_), .A2(\in1[21] ), .ZN(new_n2828_));
  AOI21_X1   g2186(.A1(new_n982_), .A2(new_n2049_), .B(new_n2828_), .ZN(new_n2829_));
  NOR2_X1    g2187(.A1(new_n2827_), .A2(new_n2829_), .ZN(new_n2830_));
  INV_X1     g2188(.I(new_n2830_), .ZN(new_n2831_));
  NOR2_X1    g2189(.A1(new_n2049_), .A2(\in1[19] ), .ZN(new_n2832_));
  AOI21_X1   g2190(.A1(new_n986_), .A2(new_n2049_), .B(new_n2832_), .ZN(new_n2833_));
  NOR2_X1    g2191(.A1(new_n2023_), .A2(\in3[19] ), .ZN(new_n2834_));
  AOI21_X1   g2192(.A1(new_n1698_), .A2(new_n2023_), .B(new_n2834_), .ZN(new_n2835_));
  NOR2_X1    g2193(.A1(new_n2023_), .A2(\in3[18] ), .ZN(new_n2836_));
  AOI21_X1   g2194(.A1(new_n1699_), .A2(new_n2023_), .B(new_n2836_), .ZN(new_n2837_));
  INV_X1     g2195(.I(new_n2837_), .ZN(new_n2838_));
  NOR2_X1    g2196(.A1(new_n2049_), .A2(\in1[18] ), .ZN(new_n2839_));
  AOI21_X1   g2197(.A1(new_n987_), .A2(new_n2049_), .B(new_n2839_), .ZN(new_n2840_));
  NOR2_X1    g2198(.A1(new_n2838_), .A2(new_n2840_), .ZN(new_n2841_));
  INV_X1     g2199(.I(new_n2841_), .ZN(new_n2842_));
  NOR2_X1    g2200(.A1(new_n2023_), .A2(\in3[16] ), .ZN(new_n2843_));
  AOI21_X1   g2201(.A1(new_n1777_), .A2(new_n2023_), .B(new_n2843_), .ZN(new_n2844_));
  INV_X1     g2202(.I(new_n2844_), .ZN(new_n2845_));
  NOR2_X1    g2203(.A1(new_n2049_), .A2(\in1[16] ), .ZN(new_n2846_));
  AOI21_X1   g2204(.A1(new_n1072_), .A2(new_n2049_), .B(new_n2846_), .ZN(new_n2847_));
  NOR2_X1    g2205(.A1(new_n2845_), .A2(new_n2847_), .ZN(new_n2848_));
  NOR2_X1    g2206(.A1(new_n2023_), .A2(\in3[15] ), .ZN(new_n2849_));
  AOI21_X1   g2207(.A1(new_n1773_), .A2(new_n2023_), .B(new_n2849_), .ZN(new_n2850_));
  INV_X1     g2208(.I(new_n2850_), .ZN(new_n2851_));
  NOR2_X1    g2209(.A1(new_n2049_), .A2(\in1[15] ), .ZN(new_n2852_));
  AOI21_X1   g2210(.A1(new_n1068_), .A2(new_n2049_), .B(new_n2852_), .ZN(new_n2853_));
  NOR2_X1    g2211(.A1(new_n2851_), .A2(new_n2853_), .ZN(new_n2854_));
  INV_X1     g2212(.I(new_n2854_), .ZN(new_n2855_));
  NOR2_X1    g2213(.A1(new_n2049_), .A2(\in1[14] ), .ZN(new_n2856_));
  AOI21_X1   g2214(.A1(new_n1255_), .A2(new_n2049_), .B(new_n2856_), .ZN(new_n2857_));
  NOR2_X1    g2215(.A1(new_n2023_), .A2(\in3[14] ), .ZN(new_n2858_));
  AOI21_X1   g2216(.A1(new_n1950_), .A2(new_n2023_), .B(new_n2858_), .ZN(new_n2859_));
  INV_X1     g2217(.I(new_n2859_), .ZN(new_n2860_));
  NOR2_X1    g2218(.A1(new_n2023_), .A2(\in3[13] ), .ZN(new_n2861_));
  AOI21_X1   g2219(.A1(new_n1707_), .A2(new_n2023_), .B(new_n2861_), .ZN(new_n2862_));
  INV_X1     g2220(.I(new_n2862_), .ZN(new_n2863_));
  NOR2_X1    g2221(.A1(new_n2049_), .A2(\in1[13] ), .ZN(new_n2864_));
  AOI21_X1   g2222(.A1(new_n997_), .A2(new_n2049_), .B(new_n2864_), .ZN(new_n2865_));
  NOR2_X1    g2223(.A1(new_n2863_), .A2(new_n2865_), .ZN(new_n2866_));
  NOR2_X1    g2224(.A1(new_n2049_), .A2(\in1[11] ), .ZN(new_n2867_));
  AOI21_X1   g2225(.A1(new_n1257_), .A2(new_n2049_), .B(new_n2867_), .ZN(new_n2868_));
  INV_X1     g2226(.I(new_n2868_), .ZN(new_n2869_));
  INV_X1     g2227(.I(\in2[11] ), .ZN(new_n2870_));
  NOR2_X1    g2228(.A1(new_n2023_), .A2(\in3[11] ), .ZN(new_n2871_));
  AOI21_X1   g2229(.A1(new_n2870_), .A2(new_n2023_), .B(new_n2871_), .ZN(new_n2872_));
  INV_X1     g2230(.I(new_n2872_), .ZN(new_n2873_));
  NOR2_X1    g2231(.A1(new_n2023_), .A2(\in3[10] ), .ZN(new_n2874_));
  AOI21_X1   g2232(.A1(new_n1712_), .A2(new_n2023_), .B(new_n2874_), .ZN(new_n2875_));
  INV_X1     g2233(.I(new_n2875_), .ZN(new_n2876_));
  NOR2_X1    g2234(.A1(new_n2049_), .A2(\in1[10] ), .ZN(new_n2877_));
  AOI21_X1   g2235(.A1(new_n1004_), .A2(new_n2049_), .B(new_n2877_), .ZN(new_n2878_));
  NOR2_X1    g2236(.A1(new_n2876_), .A2(new_n2878_), .ZN(new_n2879_));
  NOR2_X1    g2237(.A1(new_n2023_), .A2(\in3[8] ), .ZN(new_n2880_));
  AOI21_X1   g2238(.A1(new_n1751_), .A2(new_n2023_), .B(new_n2880_), .ZN(new_n2881_));
  NOR2_X1    g2239(.A1(new_n2049_), .A2(\in1[8] ), .ZN(new_n2882_));
  AOI21_X1   g2240(.A1(new_n1046_), .A2(new_n2049_), .B(new_n2882_), .ZN(new_n2883_));
  INV_X1     g2241(.I(new_n2883_), .ZN(new_n2884_));
  NOR2_X1    g2242(.A1(new_n2049_), .A2(\in1[7] ), .ZN(new_n2885_));
  AOI21_X1   g2243(.A1(new_n1260_), .A2(new_n2049_), .B(new_n2885_), .ZN(new_n2886_));
  INV_X1     g2244(.I(new_n2886_), .ZN(new_n2887_));
  NOR2_X1    g2245(.A1(new_n2023_), .A2(\in3[7] ), .ZN(new_n2888_));
  AOI21_X1   g2246(.A1(new_n1951_), .A2(new_n2023_), .B(new_n2888_), .ZN(new_n2889_));
  NOR2_X1    g2247(.A1(new_n2887_), .A2(new_n2889_), .ZN(new_n2890_));
  NAND2_X1   g2248(.A1(new_n2887_), .A2(new_n2889_), .ZN(new_n2891_));
  NOR2_X1    g2249(.A1(new_n2023_), .A2(\in3[5] ), .ZN(new_n2892_));
  AOI21_X1   g2250(.A1(new_n1745_), .A2(new_n2023_), .B(new_n2892_), .ZN(new_n2893_));
  INV_X1     g2251(.I(new_n2893_), .ZN(new_n2894_));
  NOR2_X1    g2252(.A1(new_n2049_), .A2(\in1[5] ), .ZN(new_n2895_));
  AOI21_X1   g2253(.A1(new_n1040_), .A2(new_n2049_), .B(new_n2895_), .ZN(new_n2896_));
  NOR2_X1    g2254(.A1(new_n2894_), .A2(new_n2896_), .ZN(new_n2897_));
  INV_X1     g2255(.I(new_n2897_), .ZN(new_n2898_));
  NOR2_X1    g2256(.A1(new_n2023_), .A2(\in3[4] ), .ZN(new_n2899_));
  AOI21_X1   g2257(.A1(new_n1739_), .A2(new_n2023_), .B(new_n2899_), .ZN(new_n2900_));
  INV_X1     g2258(.I(new_n2900_), .ZN(new_n2901_));
  NOR2_X1    g2259(.A1(new_n2049_), .A2(\in1[4] ), .ZN(new_n2902_));
  AOI21_X1   g2260(.A1(new_n1034_), .A2(new_n2049_), .B(new_n2902_), .ZN(new_n2903_));
  NOR2_X1    g2261(.A1(new_n2901_), .A2(new_n2903_), .ZN(new_n2904_));
  NOR2_X1    g2262(.A1(new_n2049_), .A2(\in1[3] ), .ZN(new_n2905_));
  AOI21_X1   g2263(.A1(new_n1030_), .A2(new_n2049_), .B(new_n2905_), .ZN(new_n2906_));
  NOR2_X1    g2264(.A1(new_n2023_), .A2(\in3[3] ), .ZN(new_n2907_));
  AOI21_X1   g2265(.A1(new_n1735_), .A2(new_n2023_), .B(new_n2907_), .ZN(new_n2908_));
  NOR2_X1    g2266(.A1(new_n2125_), .A2(\in2[2] ), .ZN(new_n2909_));
  NOR2_X1    g2267(.A1(new_n2023_), .A2(\in3[2] ), .ZN(new_n2910_));
  NOR2_X1    g2268(.A1(new_n2909_), .A2(new_n2910_), .ZN(new_n2911_));
  NAND3_X1   g2269(.A1(new_n1363_), .A2(new_n1022_), .A3(new_n1232_), .ZN(new_n2912_));
  OAI21_X1   g2270(.A1(new_n2062_), .A2(\in0[2] ), .B(new_n2912_), .ZN(new_n2913_));
  NAND2_X1   g2271(.A1(new_n2911_), .A2(new_n2913_), .ZN(new_n2914_));
  NAND3_X1   g2272(.A1(new_n1363_), .A2(new_n1024_), .A3(new_n1232_), .ZN(new_n2915_));
  OAI21_X1   g2273(.A1(new_n2062_), .A2(\in0[1] ), .B(new_n2915_), .ZN(new_n2916_));
  INV_X1     g2274(.I(new_n1406_), .ZN(new_n2917_));
  INV_X1     g2275(.I(new_n1459_), .ZN(new_n2918_));
  INV_X1     g2276(.I(new_n1485_), .ZN(new_n2919_));
  INV_X1     g2277(.I(new_n1538_), .ZN(new_n2920_));
  INV_X1     g2278(.I(new_n1564_), .ZN(new_n2921_));
  INV_X1     g2279(.I(new_n1656_), .ZN(new_n2922_));
  INV_X1     g2280(.I(\in3[30] ), .ZN(new_n2923_));
  INV_X1     g2281(.I(new_n1680_), .ZN(new_n2924_));
  INV_X1     g2282(.I(new_n1688_), .ZN(new_n2925_));
  INV_X1     g2283(.I(new_n1700_), .ZN(new_n2926_));
  INV_X1     g2284(.I(new_n1706_), .ZN(new_n2927_));
  INV_X1     g2285(.I(\in3[14] ), .ZN(new_n2928_));
  INV_X1     g2286(.I(new_n1710_), .ZN(new_n2929_));
  INV_X1     g2287(.I(new_n1718_), .ZN(new_n2930_));
  INV_X1     g2288(.I(\in3[7] ), .ZN(new_n2931_));
  INV_X1     g2289(.I(new_n1722_), .ZN(new_n2932_));
  INV_X1     g2290(.I(\in2[2] ), .ZN(new_n2933_));
  INV_X1     g2291(.I(\in2[1] ), .ZN(new_n2934_));
  OAI21_X1   g2292(.A1(new_n1954_), .A2(\in3[0] ), .B(new_n2934_), .ZN(new_n2935_));
  NOR3_X1    g2293(.A1(new_n1954_), .A2(new_n2934_), .A3(\in3[0] ), .ZN(new_n2936_));
  OAI21_X1   g2294(.A1(new_n1953_), .A2(new_n2936_), .B(new_n2935_), .ZN(new_n2937_));
  AOI21_X1   g2295(.A1(new_n2937_), .A2(\in3[2] ), .B(new_n2933_), .ZN(new_n2938_));
  NOR3_X1    g2296(.A1(new_n2938_), .A2(new_n1958_), .A3(new_n1736_), .ZN(new_n2939_));
  INV_X1     g2297(.I(new_n1740_), .ZN(new_n2940_));
  OAI21_X1   g2298(.A1(new_n2939_), .A2(new_n1726_), .B(new_n2940_), .ZN(new_n2941_));
  INV_X1     g2299(.I(new_n1743_), .ZN(new_n2942_));
  NAND3_X1   g2300(.A1(new_n2941_), .A2(new_n1952_), .A3(new_n2942_), .ZN(new_n2943_));
  AOI21_X1   g2301(.A1(new_n2943_), .A2(new_n1962_), .B(new_n2932_), .ZN(new_n2944_));
  OAI21_X1   g2302(.A1(new_n2944_), .A2(new_n1720_), .B(new_n2931_), .ZN(new_n2945_));
  NOR3_X1    g2303(.A1(new_n2944_), .A2(new_n2931_), .A3(new_n1720_), .ZN(new_n2946_));
  AOI21_X1   g2304(.A1(new_n1951_), .A2(new_n2945_), .B(new_n2946_), .ZN(new_n2947_));
  OAI21_X1   g2305(.A1(new_n2947_), .A2(new_n1752_), .B(new_n2930_), .ZN(new_n2948_));
  INV_X1     g2306(.I(new_n1759_), .ZN(new_n2949_));
  OAI21_X1   g2307(.A1(new_n2948_), .A2(new_n1756_), .B(new_n2949_), .ZN(new_n2950_));
  AOI21_X1   g2308(.A1(new_n2950_), .A2(new_n1715_), .B(new_n1713_), .ZN(new_n2951_));
  OAI21_X1   g2309(.A1(new_n2951_), .A2(\in3[11] ), .B(new_n2870_), .ZN(new_n2952_));
  INV_X1     g2310(.I(new_n1765_), .ZN(new_n2953_));
  NAND3_X1   g2311(.A1(new_n2952_), .A2(new_n1970_), .A3(new_n2953_), .ZN(new_n2954_));
  AOI21_X1   g2312(.A1(new_n2954_), .A2(new_n1972_), .B(new_n2929_), .ZN(new_n2955_));
  OAI21_X1   g2313(.A1(new_n2955_), .A2(new_n1708_), .B(new_n2928_), .ZN(new_n2956_));
  NOR3_X1    g2314(.A1(new_n2955_), .A2(new_n2928_), .A3(new_n1708_), .ZN(new_n2957_));
  AOI21_X1   g2315(.A1(new_n1950_), .A2(new_n2956_), .B(new_n2957_), .ZN(new_n2958_));
  OAI21_X1   g2316(.A1(new_n2958_), .A2(new_n1774_), .B(new_n2927_), .ZN(new_n2959_));
  AOI21_X1   g2317(.A1(new_n2959_), .A2(new_n1977_), .B(new_n1703_), .ZN(new_n2960_));
  AOI21_X1   g2318(.A1(new_n2960_), .A2(new_n1979_), .B(new_n1783_), .ZN(new_n2961_));
  OAI21_X1   g2319(.A1(new_n2961_), .A2(new_n1949_), .B(new_n2926_), .ZN(new_n2962_));
  AOI21_X1   g2320(.A1(new_n2962_), .A2(new_n1948_), .B(\in2[19] ), .ZN(new_n2963_));
  NOR3_X1    g2321(.A1(new_n2963_), .A2(new_n1983_), .A3(new_n1790_), .ZN(new_n2964_));
  OAI21_X1   g2322(.A1(new_n2964_), .A2(new_n1794_), .B(new_n1696_), .ZN(new_n2965_));
  AOI21_X1   g2323(.A1(new_n2965_), .A2(new_n1947_), .B(\in3[22] ), .ZN(new_n2966_));
  NAND3_X1   g2324(.A1(new_n2965_), .A2(\in3[22] ), .A3(new_n1947_), .ZN(new_n2967_));
  OAI21_X1   g2325(.A1(\in2[22] ), .A2(new_n2966_), .B(new_n2967_), .ZN(new_n2968_));
  AOI21_X1   g2326(.A1(new_n2968_), .A2(new_n1988_), .B(new_n1690_), .ZN(new_n2969_));
  OAI21_X1   g2327(.A1(new_n2969_), .A2(new_n1804_), .B(new_n2925_), .ZN(new_n2970_));
  INV_X1     g2328(.I(new_n1811_), .ZN(new_n2971_));
  OAI21_X1   g2329(.A1(new_n2970_), .A2(new_n1808_), .B(new_n2971_), .ZN(new_n2972_));
  AOI21_X1   g2330(.A1(new_n2972_), .A2(new_n1685_), .B(new_n1683_), .ZN(new_n2973_));
  OAI21_X1   g2331(.A1(new_n2973_), .A2(\in3[27] ), .B(new_n2797_), .ZN(new_n2974_));
  INV_X1     g2332(.I(new_n1817_), .ZN(new_n2975_));
  NAND3_X1   g2333(.A1(new_n2974_), .A2(new_n1994_), .A3(new_n2975_), .ZN(new_n2976_));
  AOI21_X1   g2334(.A1(new_n2976_), .A2(new_n1996_), .B(new_n2924_), .ZN(new_n2977_));
  OAI21_X1   g2335(.A1(new_n2977_), .A2(new_n1678_), .B(new_n2923_), .ZN(new_n2978_));
  NOR3_X1    g2336(.A1(new_n2977_), .A2(new_n2923_), .A3(new_n1678_), .ZN(new_n2979_));
  AOI21_X1   g2337(.A1(new_n1946_), .A2(new_n2978_), .B(new_n2979_), .ZN(new_n2980_));
  AOI21_X1   g2338(.A1(new_n2980_), .A2(new_n2000_), .B(new_n1828_), .ZN(new_n2981_));
  OAI21_X1   g2339(.A1(new_n2981_), .A2(new_n1675_), .B(new_n1844_), .ZN(new_n2982_));
  AOI21_X1   g2340(.A1(new_n2982_), .A2(new_n1945_), .B(new_n2922_), .ZN(new_n2983_));
  OAI21_X1   g2341(.A1(new_n2983_), .A2(new_n1849_), .B(new_n1626_), .ZN(new_n2984_));
  INV_X1     g2342(.I(new_n1865_), .ZN(new_n2985_));
  AOI21_X1   g2343(.A1(new_n2984_), .A2(new_n1944_), .B(new_n2985_), .ZN(new_n2986_));
  OAI21_X1   g2344(.A1(new_n2986_), .A2(new_n1579_), .B(new_n1576_), .ZN(new_n2987_));
  AOI21_X1   g2345(.A1(new_n2987_), .A2(new_n1870_), .B(new_n2921_), .ZN(new_n2988_));
  OAI21_X1   g2346(.A1(new_n2988_), .A2(new_n1943_), .B(new_n1879_), .ZN(new_n2989_));
  AOI21_X1   g2347(.A1(new_n2989_), .A2(new_n1541_), .B(new_n2920_), .ZN(new_n2990_));
  OAI21_X1   g2348(.A1(new_n2990_), .A2(new_n1884_), .B(new_n1524_), .ZN(new_n2991_));
  INV_X1     g2349(.I(new_n1892_), .ZN(new_n2992_));
  AOI21_X1   g2350(.A1(new_n2991_), .A2(new_n1511_), .B(new_n2992_), .ZN(new_n2993_));
  OAI21_X1   g2351(.A1(new_n2993_), .A2(new_n1500_), .B(new_n1497_), .ZN(new_n2994_));
  AOI21_X1   g2352(.A1(new_n2994_), .A2(new_n1897_), .B(new_n2919_), .ZN(new_n2995_));
  OAI21_X1   g2353(.A1(new_n2995_), .A2(new_n1942_), .B(new_n1906_), .ZN(new_n2996_));
  AOI21_X1   g2354(.A1(new_n2996_), .A2(new_n1462_), .B(new_n2918_), .ZN(new_n2997_));
  OAI21_X1   g2355(.A1(new_n2997_), .A2(new_n1911_), .B(new_n1445_), .ZN(new_n2998_));
  INV_X1     g2356(.I(new_n1919_), .ZN(new_n2999_));
  AOI21_X1   g2357(.A1(new_n2998_), .A2(new_n1432_), .B(new_n2999_), .ZN(new_n3000_));
  OAI21_X1   g2358(.A1(new_n3000_), .A2(new_n1421_), .B(new_n1418_), .ZN(new_n3001_));
  AOI21_X1   g2359(.A1(new_n3001_), .A2(new_n1924_), .B(new_n2917_), .ZN(new_n3002_));
  OAI21_X1   g2360(.A1(new_n3002_), .A2(new_n1941_), .B(new_n1933_), .ZN(new_n3003_));
  AOI21_X1   g2361(.A1(new_n3003_), .A2(new_n1383_), .B(new_n1378_), .ZN(new_n3004_));
  AOI21_X1   g2362(.A1(new_n3004_), .A2(new_n2022_), .B(\in2[0] ), .ZN(new_n3005_));
  NOR3_X1    g2363(.A1(new_n1936_), .A2(\in3[0] ), .A3(new_n2124_), .ZN(new_n3006_));
  OAI22_X1   g2364(.A1(new_n3005_), .A2(new_n3006_), .B1(new_n1364_), .B2(new_n1234_), .ZN(new_n3007_));
  NOR2_X1    g2365(.A1(new_n3007_), .A2(new_n2916_), .ZN(new_n3008_));
  NOR3_X1    g2366(.A1(new_n1936_), .A2(\in3[1] ), .A3(new_n2124_), .ZN(new_n3009_));
  AOI21_X1   g2367(.A1(new_n2934_), .A2(new_n2023_), .B(new_n3009_), .ZN(new_n3010_));
  AOI21_X1   g2368(.A1(new_n3007_), .A2(new_n2916_), .B(new_n3010_), .ZN(new_n3011_));
  OAI21_X1   g2369(.A1(new_n3011_), .A2(new_n3008_), .B(new_n2914_), .ZN(new_n3012_));
  NOR2_X1    g2370(.A1(new_n2911_), .A2(new_n2913_), .ZN(new_n3013_));
  INV_X1     g2371(.I(new_n3013_), .ZN(new_n3014_));
  AOI21_X1   g2372(.A1(new_n3012_), .A2(new_n3014_), .B(new_n2908_), .ZN(new_n3015_));
  NAND3_X1   g2373(.A1(new_n3012_), .A2(new_n2908_), .A3(new_n3014_), .ZN(new_n3016_));
  OAI21_X1   g2374(.A1(new_n2906_), .A2(new_n3015_), .B(new_n3016_), .ZN(new_n3017_));
  INV_X1     g2375(.I(new_n2903_), .ZN(new_n3018_));
  NOR2_X1    g2376(.A1(new_n3018_), .A2(new_n2900_), .ZN(new_n3019_));
  INV_X1     g2377(.I(new_n3019_), .ZN(new_n3020_));
  AOI21_X1   g2378(.A1(new_n3017_), .A2(new_n3020_), .B(new_n2904_), .ZN(new_n3021_));
  INV_X1     g2379(.I(new_n2896_), .ZN(new_n3022_));
  NOR2_X1    g2380(.A1(new_n3022_), .A2(new_n2893_), .ZN(new_n3023_));
  OAI21_X1   g2381(.A1(new_n3021_), .A2(new_n3023_), .B(new_n2898_), .ZN(new_n3024_));
  NOR2_X1    g2382(.A1(new_n2049_), .A2(\in1[6] ), .ZN(new_n3025_));
  AOI21_X1   g2383(.A1(new_n1011_), .A2(new_n2049_), .B(new_n3025_), .ZN(new_n3026_));
  NOR2_X1    g2384(.A1(new_n2023_), .A2(\in3[6] ), .ZN(new_n3027_));
  AOI21_X1   g2385(.A1(new_n1719_), .A2(new_n2023_), .B(new_n3027_), .ZN(new_n3028_));
  INV_X1     g2386(.I(new_n3028_), .ZN(new_n3029_));
  NOR2_X1    g2387(.A1(new_n3029_), .A2(new_n3026_), .ZN(new_n3030_));
  INV_X1     g2388(.I(new_n3026_), .ZN(new_n3031_));
  NOR2_X1    g2389(.A1(new_n3031_), .A2(new_n3028_), .ZN(new_n3032_));
  INV_X1     g2390(.I(new_n3032_), .ZN(new_n3033_));
  OAI21_X1   g2391(.A1(new_n3024_), .A2(new_n3030_), .B(new_n3033_), .ZN(new_n3034_));
  AOI21_X1   g2392(.A1(new_n3034_), .A2(new_n2891_), .B(new_n2890_), .ZN(new_n3035_));
  OAI21_X1   g2393(.A1(new_n3035_), .A2(new_n2884_), .B(new_n2881_), .ZN(new_n3036_));
  NAND2_X1   g2394(.A1(new_n3035_), .A2(new_n2884_), .ZN(new_n3037_));
  NOR2_X1    g2395(.A1(new_n2049_), .A2(\in1[9] ), .ZN(new_n3038_));
  AOI21_X1   g2396(.A1(new_n1053_), .A2(new_n2049_), .B(new_n3038_), .ZN(new_n3039_));
  NOR2_X1    g2397(.A1(new_n2023_), .A2(\in3[9] ), .ZN(new_n3040_));
  AOI21_X1   g2398(.A1(new_n1758_), .A2(new_n2023_), .B(new_n3040_), .ZN(new_n3041_));
  INV_X1     g2399(.I(new_n3041_), .ZN(new_n3042_));
  NOR2_X1    g2400(.A1(new_n3042_), .A2(new_n3039_), .ZN(new_n3043_));
  INV_X1     g2401(.I(new_n3043_), .ZN(new_n3044_));
  NAND3_X1   g2402(.A1(new_n3036_), .A2(new_n3037_), .A3(new_n3044_), .ZN(new_n3045_));
  INV_X1     g2403(.I(new_n3039_), .ZN(new_n3046_));
  NOR2_X1    g2404(.A1(new_n3046_), .A2(new_n3041_), .ZN(new_n3047_));
  INV_X1     g2405(.I(new_n3047_), .ZN(new_n3048_));
  AOI21_X1   g2406(.A1(new_n3045_), .A2(new_n3048_), .B(new_n2879_), .ZN(new_n3049_));
  INV_X1     g2407(.I(new_n2878_), .ZN(new_n3050_));
  NOR2_X1    g2408(.A1(new_n3050_), .A2(new_n2875_), .ZN(new_n3051_));
  OAI21_X1   g2409(.A1(new_n3049_), .A2(new_n3051_), .B(new_n2873_), .ZN(new_n3052_));
  NOR3_X1    g2410(.A1(new_n3049_), .A2(new_n2873_), .A3(new_n3051_), .ZN(new_n3053_));
  AOI21_X1   g2411(.A1(new_n2869_), .A2(new_n3052_), .B(new_n3053_), .ZN(new_n3054_));
  NOR2_X1    g2412(.A1(new_n2049_), .A2(\in1[12] ), .ZN(new_n3055_));
  AOI21_X1   g2413(.A1(new_n1062_), .A2(new_n2049_), .B(new_n3055_), .ZN(new_n3056_));
  NOR2_X1    g2414(.A1(new_n2023_), .A2(\in3[12] ), .ZN(new_n3057_));
  AOI21_X1   g2415(.A1(new_n1767_), .A2(new_n2023_), .B(new_n3057_), .ZN(new_n3058_));
  INV_X1     g2416(.I(new_n3058_), .ZN(new_n3059_));
  NOR2_X1    g2417(.A1(new_n3059_), .A2(new_n3056_), .ZN(new_n3060_));
  INV_X1     g2418(.I(new_n3060_), .ZN(new_n3061_));
  INV_X1     g2419(.I(new_n3056_), .ZN(new_n3062_));
  NOR2_X1    g2420(.A1(new_n3062_), .A2(new_n3058_), .ZN(new_n3063_));
  AOI21_X1   g2421(.A1(new_n3054_), .A2(new_n3061_), .B(new_n3063_), .ZN(new_n3064_));
  INV_X1     g2422(.I(new_n2865_), .ZN(new_n3065_));
  NOR2_X1    g2423(.A1(new_n3065_), .A2(new_n2862_), .ZN(new_n3066_));
  INV_X1     g2424(.I(new_n3066_), .ZN(new_n3067_));
  OAI21_X1   g2425(.A1(new_n3064_), .A2(new_n2866_), .B(new_n3067_), .ZN(new_n3068_));
  AOI21_X1   g2426(.A1(new_n3068_), .A2(new_n2860_), .B(new_n2857_), .ZN(new_n3069_));
  NOR2_X1    g2427(.A1(new_n3068_), .A2(new_n2860_), .ZN(new_n3070_));
  INV_X1     g2428(.I(new_n2853_), .ZN(new_n3071_));
  NOR2_X1    g2429(.A1(new_n3071_), .A2(new_n2850_), .ZN(new_n3072_));
  INV_X1     g2430(.I(new_n3072_), .ZN(new_n3073_));
  OAI21_X1   g2431(.A1(new_n3069_), .A2(new_n3070_), .B(new_n3073_), .ZN(new_n3074_));
  INV_X1     g2432(.I(new_n2847_), .ZN(new_n3075_));
  NOR2_X1    g2433(.A1(new_n3075_), .A2(new_n2844_), .ZN(new_n3076_));
  AOI21_X1   g2434(.A1(new_n3074_), .A2(new_n2855_), .B(new_n3076_), .ZN(new_n3077_));
  NOR2_X1    g2435(.A1(new_n2049_), .A2(\in1[17] ), .ZN(new_n3078_));
  AOI21_X1   g2436(.A1(new_n1077_), .A2(new_n2049_), .B(new_n3078_), .ZN(new_n3079_));
  NOR2_X1    g2437(.A1(new_n2023_), .A2(\in3[17] ), .ZN(new_n3080_));
  AOI21_X1   g2438(.A1(new_n1782_), .A2(new_n2023_), .B(new_n3080_), .ZN(new_n3081_));
  INV_X1     g2439(.I(new_n3081_), .ZN(new_n3082_));
  NOR2_X1    g2440(.A1(new_n3082_), .A2(new_n3079_), .ZN(new_n3083_));
  NOR3_X1    g2441(.A1(new_n3077_), .A2(new_n2848_), .A3(new_n3083_), .ZN(new_n3084_));
  INV_X1     g2442(.I(new_n3079_), .ZN(new_n3085_));
  NOR2_X1    g2443(.A1(new_n3085_), .A2(new_n3081_), .ZN(new_n3086_));
  OAI21_X1   g2444(.A1(new_n3084_), .A2(new_n3086_), .B(new_n2842_), .ZN(new_n3087_));
  INV_X1     g2445(.I(new_n2840_), .ZN(new_n3088_));
  NOR2_X1    g2446(.A1(new_n3088_), .A2(new_n2837_), .ZN(new_n3089_));
  INV_X1     g2447(.I(new_n3089_), .ZN(new_n3090_));
  AOI21_X1   g2448(.A1(new_n3087_), .A2(new_n3090_), .B(new_n2835_), .ZN(new_n3091_));
  NAND3_X1   g2449(.A1(new_n3087_), .A2(new_n2835_), .A3(new_n3090_), .ZN(new_n3092_));
  OAI21_X1   g2450(.A1(new_n2833_), .A2(new_n3091_), .B(new_n3092_), .ZN(new_n3093_));
  NOR2_X1    g2451(.A1(new_n2049_), .A2(\in1[20] ), .ZN(new_n3094_));
  AOI21_X1   g2452(.A1(new_n1088_), .A2(new_n2049_), .B(new_n3094_), .ZN(new_n3095_));
  NOR2_X1    g2453(.A1(new_n2023_), .A2(\in3[20] ), .ZN(new_n3096_));
  AOI21_X1   g2454(.A1(new_n1793_), .A2(new_n2023_), .B(new_n3096_), .ZN(new_n3097_));
  INV_X1     g2455(.I(new_n3097_), .ZN(new_n3098_));
  NOR2_X1    g2456(.A1(new_n3098_), .A2(new_n3095_), .ZN(new_n3099_));
  INV_X1     g2457(.I(new_n3095_), .ZN(new_n3100_));
  NOR2_X1    g2458(.A1(new_n3100_), .A2(new_n3097_), .ZN(new_n3101_));
  INV_X1     g2459(.I(new_n3101_), .ZN(new_n3102_));
  OAI21_X1   g2460(.A1(new_n3093_), .A2(new_n3099_), .B(new_n3102_), .ZN(new_n3103_));
  INV_X1     g2461(.I(new_n2829_), .ZN(new_n3104_));
  NOR2_X1    g2462(.A1(new_n3104_), .A2(new_n2826_), .ZN(new_n3105_));
  AOI21_X1   g2463(.A1(new_n3103_), .A2(new_n2831_), .B(new_n3105_), .ZN(new_n3106_));
  OAI21_X1   g2464(.A1(new_n3106_), .A2(new_n2824_), .B(new_n2822_), .ZN(new_n3107_));
  NAND2_X1   g2465(.A1(new_n3106_), .A2(new_n2824_), .ZN(new_n3108_));
  INV_X1     g2466(.I(new_n2818_), .ZN(new_n3109_));
  NOR2_X1    g2467(.A1(new_n3109_), .A2(new_n2815_), .ZN(new_n3110_));
  AOI21_X1   g2468(.A1(new_n3107_), .A2(new_n3108_), .B(new_n3110_), .ZN(new_n3111_));
  INV_X1     g2469(.I(new_n2811_), .ZN(new_n3112_));
  NOR2_X1    g2470(.A1(new_n3112_), .A2(new_n2808_), .ZN(new_n3113_));
  INV_X1     g2471(.I(new_n3113_), .ZN(new_n3114_));
  OAI21_X1   g2472(.A1(new_n3111_), .A2(new_n2819_), .B(new_n3114_), .ZN(new_n3115_));
  NOR2_X1    g2473(.A1(new_n2049_), .A2(\in1[25] ), .ZN(new_n3116_));
  AOI21_X1   g2474(.A1(new_n1105_), .A2(new_n2049_), .B(new_n3116_), .ZN(new_n3117_));
  NOR2_X1    g2475(.A1(new_n2023_), .A2(\in3[25] ), .ZN(new_n3118_));
  AOI21_X1   g2476(.A1(new_n1810_), .A2(new_n2023_), .B(new_n3118_), .ZN(new_n3119_));
  INV_X1     g2477(.I(new_n3119_), .ZN(new_n3120_));
  NOR2_X1    g2478(.A1(new_n3120_), .A2(new_n3117_), .ZN(new_n3121_));
  INV_X1     g2479(.I(new_n3121_), .ZN(new_n3122_));
  NAND3_X1   g2480(.A1(new_n3115_), .A2(new_n2813_), .A3(new_n3122_), .ZN(new_n3123_));
  INV_X1     g2481(.I(new_n3117_), .ZN(new_n3124_));
  NOR2_X1    g2482(.A1(new_n3124_), .A2(new_n3119_), .ZN(new_n3125_));
  INV_X1     g2483(.I(new_n3125_), .ZN(new_n3126_));
  AOI21_X1   g2484(.A1(new_n3123_), .A2(new_n3126_), .B(new_n2806_), .ZN(new_n3127_));
  INV_X1     g2485(.I(new_n2805_), .ZN(new_n3128_));
  NOR2_X1    g2486(.A1(new_n3128_), .A2(new_n2802_), .ZN(new_n3129_));
  OAI21_X1   g2487(.A1(new_n3127_), .A2(new_n3129_), .B(new_n2800_), .ZN(new_n3130_));
  NOR3_X1    g2488(.A1(new_n3127_), .A2(new_n2800_), .A3(new_n3129_), .ZN(new_n3131_));
  AOI21_X1   g2489(.A1(new_n2796_), .A2(new_n3130_), .B(new_n3131_), .ZN(new_n3132_));
  NOR2_X1    g2490(.A1(new_n2049_), .A2(\in1[28] ), .ZN(new_n3133_));
  AOI21_X1   g2491(.A1(new_n1114_), .A2(new_n2049_), .B(new_n3133_), .ZN(new_n3134_));
  NOR2_X1    g2492(.A1(new_n2023_), .A2(\in3[28] ), .ZN(new_n3135_));
  AOI21_X1   g2493(.A1(new_n1819_), .A2(new_n2023_), .B(new_n3135_), .ZN(new_n3136_));
  INV_X1     g2494(.I(new_n3136_), .ZN(new_n3137_));
  NOR2_X1    g2495(.A1(new_n3137_), .A2(new_n3134_), .ZN(new_n3138_));
  INV_X1     g2496(.I(new_n3138_), .ZN(new_n3139_));
  INV_X1     g2497(.I(new_n3134_), .ZN(new_n3140_));
  NOR2_X1    g2498(.A1(new_n3140_), .A2(new_n3136_), .ZN(new_n3141_));
  AOI21_X1   g2499(.A1(new_n3132_), .A2(new_n3139_), .B(new_n3141_), .ZN(new_n3142_));
  INV_X1     g2500(.I(new_n2792_), .ZN(new_n3143_));
  NOR2_X1    g2501(.A1(new_n3143_), .A2(new_n2789_), .ZN(new_n3144_));
  INV_X1     g2502(.I(new_n3144_), .ZN(new_n3145_));
  OAI21_X1   g2503(.A1(new_n3142_), .A2(new_n2793_), .B(new_n3145_), .ZN(new_n3146_));
  AOI21_X1   g2504(.A1(new_n3146_), .A2(new_n2787_), .B(new_n2784_), .ZN(new_n3147_));
  NOR2_X1    g2505(.A1(new_n3146_), .A2(new_n2787_), .ZN(new_n3148_));
  NOR2_X1    g2506(.A1(new_n2049_), .A2(\in1[31] ), .ZN(new_n3149_));
  AOI21_X1   g2507(.A1(new_n1122_), .A2(new_n2049_), .B(new_n3149_), .ZN(new_n3150_));
  NOR2_X1    g2508(.A1(new_n2023_), .A2(\in3[31] ), .ZN(new_n3151_));
  AOI21_X1   g2509(.A1(new_n1827_), .A2(new_n2023_), .B(new_n3151_), .ZN(new_n3152_));
  INV_X1     g2510(.I(new_n3152_), .ZN(new_n3153_));
  NOR2_X1    g2511(.A1(new_n3153_), .A2(new_n3150_), .ZN(new_n3154_));
  NOR3_X1    g2512(.A1(new_n3147_), .A2(new_n3148_), .A3(new_n3154_), .ZN(new_n3155_));
  INV_X1     g2513(.I(new_n3150_), .ZN(new_n3156_));
  NOR2_X1    g2514(.A1(new_n3156_), .A2(new_n3152_), .ZN(new_n3157_));
  OAI21_X1   g2515(.A1(new_n3155_), .A2(new_n3157_), .B(new_n2782_), .ZN(new_n3158_));
  NOR2_X1    g2516(.A1(new_n2739_), .A2(new_n2741_), .ZN(new_n3159_));
  AOI22_X1   g2517(.A1(new_n2734_), .A2(new_n2736_), .B1(new_n2780_), .B2(new_n2777_), .ZN(new_n3160_));
  INV_X1     g2518(.I(new_n2747_), .ZN(new_n3161_));
  AOI22_X1   g2519(.A1(new_n2739_), .A2(new_n2741_), .B1(new_n3161_), .B2(new_n2744_), .ZN(new_n3162_));
  OAI22_X1   g2520(.A1(new_n2749_), .A2(new_n3160_), .B1(new_n3159_), .B2(new_n3162_), .ZN(new_n3163_));
  NAND2_X1   g2521(.A1(new_n3163_), .A2(new_n2774_), .ZN(new_n3164_));
  NAND2_X1   g2522(.A1(new_n2760_), .A2(new_n2757_), .ZN(new_n3165_));
  AOI22_X1   g2523(.A1(new_n2752_), .A2(new_n2754_), .B1(new_n2770_), .B2(new_n2772_), .ZN(new_n3166_));
  NOR2_X1    g2524(.A1(new_n3166_), .A2(new_n2755_), .ZN(new_n3167_));
  OAI22_X1   g2525(.A1(new_n2760_), .A2(new_n2757_), .B1(new_n2762_), .B2(new_n2765_), .ZN(new_n3168_));
  AOI22_X1   g2526(.A1(new_n3167_), .A2(new_n2766_), .B1(new_n3165_), .B2(new_n3168_), .ZN(new_n3169_));
  NAND2_X1   g2527(.A1(new_n3164_), .A2(new_n3169_), .ZN(new_n3170_));
  INV_X1     g2528(.I(new_n3170_), .ZN(new_n3171_));
  AOI21_X1   g2529(.A1(new_n3158_), .A2(new_n3171_), .B(new_n2731_), .ZN(new_n3172_));
  INV_X1     g2530(.I(new_n2632_), .ZN(new_n3173_));
  NOR2_X1    g2531(.A1(new_n2656_), .A2(new_n2653_), .ZN(new_n3174_));
  NOR3_X1    g2532(.A1(new_n3173_), .A2(new_n2651_), .A3(new_n3174_), .ZN(new_n3175_));
  OAI21_X1   g2533(.A1(new_n3172_), .A2(new_n2727_), .B(new_n3175_), .ZN(new_n3176_));
  AOI21_X1   g2534(.A1(new_n3176_), .A2(new_n2665_), .B(new_n2600_), .ZN(new_n3177_));
  NAND2_X1   g2535(.A1(new_n2564_), .A2(new_n2566_), .ZN(new_n3178_));
  INV_X1     g2536(.I(new_n2586_), .ZN(new_n3179_));
  OR3_X2     g2537(.A1(new_n2567_), .A2(new_n2583_), .A3(new_n3179_), .Z(new_n3180_));
  AOI21_X1   g2538(.A1(new_n3178_), .A2(new_n3180_), .B(new_n2581_), .ZN(new_n3181_));
  INV_X1     g2539(.I(new_n2590_), .ZN(new_n3182_));
  INV_X1     g2540(.I(new_n2557_), .ZN(new_n3183_));
  AOI22_X1   g2541(.A1(new_n2552_), .A2(new_n2554_), .B1(new_n3183_), .B2(new_n2559_), .ZN(new_n3184_));
  OAI22_X1   g2542(.A1(new_n3184_), .A2(new_n2555_), .B1(new_n2595_), .B2(new_n2598_), .ZN(new_n3185_));
  AOI22_X1   g2543(.A1(new_n3185_), .A2(new_n2599_), .B1(new_n3182_), .B2(new_n2592_), .ZN(new_n3186_));
  NOR4_X1    g2544(.A1(new_n3186_), .A2(new_n2567_), .A3(new_n2581_), .A4(new_n2587_), .ZN(new_n3187_));
  INV_X1     g2545(.I(new_n2576_), .ZN(new_n3188_));
  AOI22_X1   g2546(.A1(new_n2570_), .A2(new_n2573_), .B1(new_n3188_), .B2(new_n2578_), .ZN(new_n3189_));
  NOR2_X1    g2547(.A1(new_n3189_), .A2(new_n2574_), .ZN(new_n3190_));
  NOR3_X1    g2548(.A1(new_n3187_), .A2(new_n3181_), .A3(new_n3190_), .ZN(new_n3191_));
  INV_X1     g2549(.I(new_n3191_), .ZN(new_n3192_));
  OAI21_X1   g2550(.A1(new_n3177_), .A2(new_n3192_), .B(new_n2549_), .ZN(new_n3193_));
  NAND2_X1   g2551(.A1(new_n2512_), .A2(new_n2509_), .ZN(new_n3194_));
  NAND3_X1   g2552(.A1(new_n2496_), .A2(new_n2506_), .A3(new_n3194_), .ZN(new_n3195_));
  AOI21_X1   g2553(.A1(new_n3193_), .A2(new_n2546_), .B(new_n3195_), .ZN(new_n3196_));
  OAI21_X1   g2554(.A1(new_n3196_), .A2(new_n2518_), .B(new_n2483_), .ZN(new_n3197_));
  INV_X1     g2555(.I(new_n2465_), .ZN(new_n3198_));
  AOI22_X1   g2556(.A1(new_n2459_), .A2(new_n2462_), .B1(new_n2478_), .B2(new_n2481_), .ZN(new_n3199_));
  OAI22_X1   g2557(.A1(new_n3199_), .A2(new_n2482_), .B1(new_n2470_), .B2(new_n2473_), .ZN(new_n3200_));
  AOI22_X1   g2558(.A1(new_n3200_), .A2(new_n2474_), .B1(new_n3198_), .B2(new_n2467_), .ZN(new_n3201_));
  AOI21_X1   g2559(.A1(new_n3197_), .A2(new_n3201_), .B(new_n2455_), .ZN(new_n3202_));
  INV_X1     g2560(.I(new_n2402_), .ZN(new_n3203_));
  NOR2_X1    g2561(.A1(new_n2412_), .A2(new_n2415_), .ZN(new_n3204_));
  NOR3_X1    g2562(.A1(new_n3203_), .A2(new_n2409_), .A3(new_n3204_), .ZN(new_n3205_));
  OAI21_X1   g2563(.A1(new_n3202_), .A2(new_n2453_), .B(new_n3205_), .ZN(new_n3206_));
  AOI21_X1   g2564(.A1(new_n3206_), .A2(new_n2418_), .B(new_n2390_), .ZN(new_n3207_));
  INV_X1     g2565(.I(new_n2373_), .ZN(new_n3208_));
  AOI22_X1   g2566(.A1(new_n2362_), .A2(new_n2365_), .B1(new_n2384_), .B2(new_n2387_), .ZN(new_n3209_));
  NOR2_X1    g2567(.A1(new_n3209_), .A2(new_n2366_), .ZN(new_n3210_));
  INV_X1     g2568(.I(new_n2372_), .ZN(new_n3211_));
  OAI22_X1   g2569(.A1(new_n3211_), .A2(new_n2368_), .B1(new_n2378_), .B2(new_n2375_), .ZN(new_n3212_));
  AOI22_X1   g2570(.A1(new_n3210_), .A2(new_n2379_), .B1(new_n3208_), .B2(new_n3212_), .ZN(new_n3213_));
  INV_X1     g2571(.I(new_n3213_), .ZN(new_n3214_));
  OAI21_X1   g2572(.A1(new_n3207_), .A2(new_n3214_), .B(new_n2358_), .ZN(new_n3215_));
  NAND2_X1   g2573(.A1(new_n2321_), .A2(new_n2318_), .ZN(new_n3216_));
  NAND3_X1   g2574(.A1(new_n2305_), .A2(new_n2315_), .A3(new_n3216_), .ZN(new_n3217_));
  AOI21_X1   g2575(.A1(new_n3215_), .A2(new_n2355_), .B(new_n3217_), .ZN(new_n3218_));
  OAI21_X1   g2576(.A1(new_n3218_), .A2(new_n2327_), .B(new_n2292_), .ZN(new_n3219_));
  INV_X1     g2577(.I(new_n2274_), .ZN(new_n3220_));
  AOI22_X1   g2578(.A1(new_n2268_), .A2(new_n2271_), .B1(new_n2287_), .B2(new_n2290_), .ZN(new_n3221_));
  OAI22_X1   g2579(.A1(new_n3221_), .A2(new_n2291_), .B1(new_n2279_), .B2(new_n2282_), .ZN(new_n3222_));
  AOI22_X1   g2580(.A1(new_n3222_), .A2(new_n2283_), .B1(new_n3220_), .B2(new_n2276_), .ZN(new_n3223_));
  AOI21_X1   g2581(.A1(new_n3219_), .A2(new_n3223_), .B(new_n2264_), .ZN(new_n3224_));
  INV_X1     g2582(.I(new_n2211_), .ZN(new_n3225_));
  NOR2_X1    g2583(.A1(new_n2221_), .A2(new_n2224_), .ZN(new_n3226_));
  NOR3_X1    g2584(.A1(new_n3225_), .A2(new_n2218_), .A3(new_n3226_), .ZN(new_n3227_));
  OAI21_X1   g2585(.A1(new_n3224_), .A2(new_n2262_), .B(new_n3227_), .ZN(new_n3228_));
  AOI21_X1   g2586(.A1(new_n3228_), .A2(new_n2227_), .B(new_n2199_), .ZN(new_n3229_));
  INV_X1     g2587(.I(new_n2182_), .ZN(new_n3230_));
  AOI22_X1   g2588(.A1(new_n2171_), .A2(new_n2174_), .B1(new_n2193_), .B2(new_n2196_), .ZN(new_n3231_));
  NOR2_X1    g2589(.A1(new_n3231_), .A2(new_n2175_), .ZN(new_n3232_));
  INV_X1     g2590(.I(new_n2181_), .ZN(new_n3233_));
  OAI22_X1   g2591(.A1(new_n3233_), .A2(new_n2177_), .B1(new_n2187_), .B2(new_n2184_), .ZN(new_n3234_));
  AOI22_X1   g2592(.A1(new_n3232_), .A2(new_n2188_), .B1(new_n3230_), .B2(new_n3234_), .ZN(new_n3235_));
  INV_X1     g2593(.I(new_n3235_), .ZN(new_n3236_));
  OAI21_X1   g2594(.A1(new_n3229_), .A2(new_n3236_), .B(new_n2167_), .ZN(new_n3237_));
  NAND2_X1   g2595(.A1(new_n2130_), .A2(new_n2127_), .ZN(new_n3238_));
  NAND3_X1   g2596(.A1(new_n2112_), .A2(new_n2122_), .A3(new_n3238_), .ZN(new_n3239_));
  AOI21_X1   g2597(.A1(new_n3237_), .A2(new_n2164_), .B(new_n3239_), .ZN(new_n3240_));
  OAI21_X1   g2598(.A1(new_n3240_), .A2(new_n2136_), .B(new_n2099_), .ZN(new_n3241_));
  INV_X1     g2599(.I(new_n2081_), .ZN(new_n3242_));
  AOI22_X1   g2600(.A1(new_n2075_), .A2(new_n2078_), .B1(new_n2094_), .B2(new_n2097_), .ZN(new_n3243_));
  OAI22_X1   g2601(.A1(new_n3243_), .A2(new_n2098_), .B1(new_n2086_), .B2(new_n2089_), .ZN(new_n3244_));
  AOI22_X1   g2602(.A1(new_n3244_), .A2(new_n2090_), .B1(new_n3242_), .B2(new_n2083_), .ZN(new_n3245_));
  AOI21_X1   g2603(.A1(new_n3241_), .A2(new_n3245_), .B(new_n2071_), .ZN(new_n3246_));
  NOR3_X1    g2604(.A1(new_n3246_), .A2(new_n1938_), .A3(new_n2068_), .ZN(\address[1] ));
  INV_X1     g2605(.I(new_n1938_), .ZN(new_n3248_));
  INV_X1     g2606(.I(new_n2068_), .ZN(new_n3249_));
  NOR2_X1    g2607(.A1(new_n3005_), .A2(new_n3006_), .ZN(new_n3250_));
  INV_X1     g2608(.I(new_n2071_), .ZN(new_n3251_));
  INV_X1     g2609(.I(new_n2099_), .ZN(new_n3252_));
  INV_X1     g2610(.I(new_n2136_), .ZN(new_n3253_));
  INV_X1     g2611(.I(new_n2164_), .ZN(new_n3254_));
  INV_X1     g2612(.I(new_n2167_), .ZN(new_n3255_));
  INV_X1     g2613(.I(new_n2227_), .ZN(new_n3256_));
  INV_X1     g2614(.I(new_n2262_), .ZN(new_n3257_));
  INV_X1     g2615(.I(new_n2264_), .ZN(new_n3258_));
  INV_X1     g2616(.I(new_n2292_), .ZN(new_n3259_));
  INV_X1     g2617(.I(new_n2327_), .ZN(new_n3260_));
  INV_X1     g2618(.I(new_n2355_), .ZN(new_n3261_));
  INV_X1     g2619(.I(new_n2358_), .ZN(new_n3262_));
  INV_X1     g2620(.I(new_n2418_), .ZN(new_n3263_));
  INV_X1     g2621(.I(new_n2453_), .ZN(new_n3264_));
  INV_X1     g2622(.I(new_n2455_), .ZN(new_n3265_));
  INV_X1     g2623(.I(new_n2483_), .ZN(new_n3266_));
  INV_X1     g2624(.I(new_n2518_), .ZN(new_n3267_));
  INV_X1     g2625(.I(new_n2546_), .ZN(new_n3268_));
  INV_X1     g2626(.I(new_n2549_), .ZN(new_n3269_));
  INV_X1     g2627(.I(new_n2600_), .ZN(new_n3270_));
  INV_X1     g2628(.I(new_n2731_), .ZN(new_n3271_));
  INV_X1     g2629(.I(new_n2782_), .ZN(new_n3272_));
  INV_X1     g2630(.I(new_n2784_), .ZN(new_n3273_));
  INV_X1     g2631(.I(new_n2793_), .ZN(new_n3274_));
  INV_X1     g2632(.I(new_n2806_), .ZN(new_n3275_));
  INV_X1     g2633(.I(new_n2819_), .ZN(new_n3276_));
  INV_X1     g2634(.I(new_n2824_), .ZN(new_n3277_));
  INV_X1     g2635(.I(new_n2833_), .ZN(new_n3278_));
  INV_X1     g2636(.I(new_n2835_), .ZN(new_n3279_));
  INV_X1     g2637(.I(new_n2848_), .ZN(new_n3280_));
  INV_X1     g2638(.I(new_n2857_), .ZN(new_n3281_));
  INV_X1     g2639(.I(new_n2866_), .ZN(new_n3282_));
  INV_X1     g2640(.I(new_n2879_), .ZN(new_n3283_));
  INV_X1     g2641(.I(new_n2881_), .ZN(new_n3284_));
  INV_X1     g2642(.I(new_n2890_), .ZN(new_n3285_));
  INV_X1     g2643(.I(new_n2891_), .ZN(new_n3286_));
  INV_X1     g2644(.I(new_n2904_), .ZN(new_n3287_));
  INV_X1     g2645(.I(new_n2906_), .ZN(new_n3288_));
  INV_X1     g2646(.I(new_n2908_), .ZN(new_n3289_));
  NOR2_X1    g2647(.A1(new_n1117_), .A2(\in0[30] ), .ZN(new_n3290_));
  NOR3_X1    g2648(.A1(new_n3290_), .A2(new_n1337_), .A3(new_n1121_), .ZN(new_n3291_));
  OAI21_X1   g2649(.A1(new_n3291_), .A2(new_n1123_), .B(new_n962_), .ZN(new_n3292_));
  AOI21_X1   g2650(.A1(new_n3292_), .A2(new_n1141_), .B(new_n945_), .ZN(new_n3293_));
  OAI21_X1   g2651(.A1(new_n3293_), .A2(new_n1243_), .B(new_n1147_), .ZN(new_n3294_));
  AOI21_X1   g2652(.A1(new_n3294_), .A2(new_n912_), .B(new_n881_), .ZN(new_n3295_));
  OAI21_X1   g2653(.A1(new_n3295_), .A2(new_n1344_), .B(new_n865_), .ZN(new_n3296_));
  AOI21_X1   g2654(.A1(new_n3296_), .A2(new_n861_), .B(new_n1169_), .ZN(new_n3297_));
  OAI21_X1   g2655(.A1(new_n3297_), .A2(new_n848_), .B(new_n834_), .ZN(new_n3298_));
  AOI21_X1   g2656(.A1(new_n3298_), .A2(new_n1176_), .B(new_n825_), .ZN(new_n3299_));
  OAI21_X1   g2657(.A1(new_n3299_), .A2(new_n821_), .B(new_n1182_), .ZN(new_n3300_));
  AOI21_X1   g2658(.A1(new_n3300_), .A2(new_n806_), .B(new_n794_), .ZN(new_n3301_));
  OAI21_X1   g2659(.A1(new_n3301_), .A2(new_n1189_), .B(new_n783_), .ZN(new_n3302_));
  AOI21_X1   g2660(.A1(new_n3302_), .A2(new_n779_), .B(new_n1195_), .ZN(new_n3303_));
  OAI21_X1   g2661(.A1(new_n3303_), .A2(new_n766_), .B(new_n752_), .ZN(new_n3304_));
  AOI21_X1   g2662(.A1(new_n3304_), .A2(new_n1202_), .B(new_n743_), .ZN(new_n3305_));
  OAI21_X1   g2663(.A1(new_n3305_), .A2(new_n739_), .B(new_n1208_), .ZN(new_n3306_));
  AOI21_X1   g2664(.A1(new_n3306_), .A2(new_n724_), .B(new_n712_), .ZN(new_n3307_));
  OAI21_X1   g2665(.A1(new_n3307_), .A2(new_n1215_), .B(new_n701_), .ZN(new_n3308_));
  AOI21_X1   g2666(.A1(new_n3308_), .A2(new_n697_), .B(new_n1221_), .ZN(new_n3309_));
  OAI21_X1   g2667(.A1(new_n3309_), .A2(new_n684_), .B(new_n670_), .ZN(new_n3310_));
  AOI21_X1   g2668(.A1(new_n3310_), .A2(new_n1228_), .B(new_n661_), .ZN(new_n3311_));
  NOR4_X1    g2669(.A1(new_n3311_), .A2(\in1[2] ), .A3(new_n656_), .A4(new_n1233_), .ZN(new_n3312_));
  AOI21_X1   g2670(.A1(new_n1263_), .A2(new_n2049_), .B(new_n3312_), .ZN(new_n3313_));
  NOR3_X1    g2671(.A1(new_n3313_), .A2(new_n2909_), .A3(new_n2910_), .ZN(new_n3314_));
  NOR3_X1    g2672(.A1(new_n1231_), .A2(\in1[1] ), .A3(new_n1233_), .ZN(new_n3315_));
  AOI21_X1   g2673(.A1(new_n1265_), .A2(new_n2049_), .B(new_n3315_), .ZN(new_n3316_));
  NAND4_X1   g2674(.A1(new_n2048_), .A2(\in1[0] ), .A3(new_n657_), .A4(new_n1232_), .ZN(new_n3317_));
  OAI21_X1   g2675(.A1(new_n1231_), .A2(new_n1233_), .B(\in0[0] ), .ZN(new_n3318_));
  OAI21_X1   g2676(.A1(new_n1936_), .A2(new_n2124_), .B(new_n1954_), .ZN(new_n3319_));
  NAND4_X1   g2677(.A1(new_n2021_), .A2(new_n1729_), .A3(new_n1379_), .A4(new_n2022_), .ZN(new_n3320_));
  AOI22_X1   g2678(.A1(new_n3319_), .A2(new_n3320_), .B1(new_n3318_), .B2(new_n3317_), .ZN(new_n3321_));
  NAND2_X1   g2679(.A1(new_n3321_), .A2(new_n3316_), .ZN(new_n3322_));
  NAND4_X1   g2680(.A1(new_n2021_), .A2(new_n1953_), .A3(new_n1379_), .A4(new_n2022_), .ZN(new_n3323_));
  OAI21_X1   g2681(.A1(\in2[1] ), .A2(new_n2125_), .B(new_n3323_), .ZN(new_n3324_));
  OAI21_X1   g2682(.A1(new_n3321_), .A2(new_n3316_), .B(new_n3324_), .ZN(new_n3325_));
  AOI21_X1   g2683(.A1(new_n3325_), .A2(new_n3322_), .B(new_n3314_), .ZN(new_n3326_));
  OAI21_X1   g2684(.A1(new_n3326_), .A2(new_n3013_), .B(new_n3289_), .ZN(new_n3327_));
  NOR3_X1    g2685(.A1(new_n3326_), .A2(new_n3289_), .A3(new_n3013_), .ZN(new_n3328_));
  AOI21_X1   g2686(.A1(new_n3288_), .A2(new_n3327_), .B(new_n3328_), .ZN(new_n3329_));
  OAI21_X1   g2687(.A1(new_n3329_), .A2(new_n3019_), .B(new_n3287_), .ZN(new_n3330_));
  INV_X1     g2688(.I(new_n3023_), .ZN(new_n3331_));
  AOI21_X1   g2689(.A1(new_n3330_), .A2(new_n3331_), .B(new_n2897_), .ZN(new_n3332_));
  INV_X1     g2690(.I(new_n3030_), .ZN(new_n3333_));
  AOI21_X1   g2691(.A1(new_n3332_), .A2(new_n3333_), .B(new_n3032_), .ZN(new_n3334_));
  OAI21_X1   g2692(.A1(new_n3334_), .A2(new_n3286_), .B(new_n3285_), .ZN(new_n3335_));
  AOI21_X1   g2693(.A1(new_n3335_), .A2(new_n2883_), .B(new_n3284_), .ZN(new_n3336_));
  NOR2_X1    g2694(.A1(new_n3335_), .A2(new_n2883_), .ZN(new_n3337_));
  NOR3_X1    g2695(.A1(new_n3336_), .A2(new_n3337_), .A3(new_n3043_), .ZN(new_n3338_));
  OAI21_X1   g2696(.A1(new_n3338_), .A2(new_n3047_), .B(new_n3283_), .ZN(new_n3339_));
  INV_X1     g2697(.I(new_n3051_), .ZN(new_n3340_));
  AOI21_X1   g2698(.A1(new_n3339_), .A2(new_n3340_), .B(new_n2872_), .ZN(new_n3341_));
  NAND3_X1   g2699(.A1(new_n3339_), .A2(new_n2872_), .A3(new_n3340_), .ZN(new_n3342_));
  OAI21_X1   g2700(.A1(new_n2868_), .A2(new_n3341_), .B(new_n3342_), .ZN(new_n3343_));
  INV_X1     g2701(.I(new_n3063_), .ZN(new_n3344_));
  OAI21_X1   g2702(.A1(new_n3343_), .A2(new_n3060_), .B(new_n3344_), .ZN(new_n3345_));
  AOI21_X1   g2703(.A1(new_n3345_), .A2(new_n3282_), .B(new_n3066_), .ZN(new_n3346_));
  OAI21_X1   g2704(.A1(new_n3346_), .A2(new_n2859_), .B(new_n3281_), .ZN(new_n3347_));
  NAND2_X1   g2705(.A1(new_n3346_), .A2(new_n2859_), .ZN(new_n3348_));
  AOI21_X1   g2706(.A1(new_n3347_), .A2(new_n3348_), .B(new_n3072_), .ZN(new_n3349_));
  INV_X1     g2707(.I(new_n3076_), .ZN(new_n3350_));
  OAI21_X1   g2708(.A1(new_n3349_), .A2(new_n2854_), .B(new_n3350_), .ZN(new_n3351_));
  INV_X1     g2709(.I(new_n3083_), .ZN(new_n3352_));
  NAND3_X1   g2710(.A1(new_n3351_), .A2(new_n3280_), .A3(new_n3352_), .ZN(new_n3353_));
  INV_X1     g2711(.I(new_n3086_), .ZN(new_n3354_));
  AOI21_X1   g2712(.A1(new_n3353_), .A2(new_n3354_), .B(new_n2841_), .ZN(new_n3355_));
  OAI21_X1   g2713(.A1(new_n3355_), .A2(new_n3089_), .B(new_n3279_), .ZN(new_n3356_));
  NOR3_X1    g2714(.A1(new_n3355_), .A2(new_n3279_), .A3(new_n3089_), .ZN(new_n3357_));
  AOI21_X1   g2715(.A1(new_n3278_), .A2(new_n3356_), .B(new_n3357_), .ZN(new_n3358_));
  INV_X1     g2716(.I(new_n3099_), .ZN(new_n3359_));
  AOI21_X1   g2717(.A1(new_n3358_), .A2(new_n3359_), .B(new_n3101_), .ZN(new_n3360_));
  INV_X1     g2718(.I(new_n3105_), .ZN(new_n3361_));
  OAI21_X1   g2719(.A1(new_n3360_), .A2(new_n2830_), .B(new_n3361_), .ZN(new_n3362_));
  AOI21_X1   g2720(.A1(new_n3362_), .A2(new_n3277_), .B(new_n2821_), .ZN(new_n3363_));
  NOR2_X1    g2721(.A1(new_n3362_), .A2(new_n3277_), .ZN(new_n3364_));
  INV_X1     g2722(.I(new_n3110_), .ZN(new_n3365_));
  OAI21_X1   g2723(.A1(new_n3363_), .A2(new_n3364_), .B(new_n3365_), .ZN(new_n3366_));
  AOI21_X1   g2724(.A1(new_n3366_), .A2(new_n3276_), .B(new_n3113_), .ZN(new_n3367_));
  NOR3_X1    g2725(.A1(new_n3367_), .A2(new_n2812_), .A3(new_n3121_), .ZN(new_n3368_));
  OAI21_X1   g2726(.A1(new_n3368_), .A2(new_n3125_), .B(new_n3275_), .ZN(new_n3369_));
  INV_X1     g2727(.I(new_n3129_), .ZN(new_n3370_));
  AOI21_X1   g2728(.A1(new_n3369_), .A2(new_n3370_), .B(new_n2799_), .ZN(new_n3371_));
  NAND3_X1   g2729(.A1(new_n3369_), .A2(new_n2799_), .A3(new_n3370_), .ZN(new_n3372_));
  OAI21_X1   g2730(.A1(new_n2795_), .A2(new_n3371_), .B(new_n3372_), .ZN(new_n3373_));
  INV_X1     g2731(.I(new_n3141_), .ZN(new_n3374_));
  OAI21_X1   g2732(.A1(new_n3373_), .A2(new_n3138_), .B(new_n3374_), .ZN(new_n3375_));
  AOI21_X1   g2733(.A1(new_n3375_), .A2(new_n3274_), .B(new_n3144_), .ZN(new_n3376_));
  OAI21_X1   g2734(.A1(new_n3376_), .A2(new_n2786_), .B(new_n3273_), .ZN(new_n3377_));
  NAND2_X1   g2735(.A1(new_n3376_), .A2(new_n2786_), .ZN(new_n3378_));
  INV_X1     g2736(.I(new_n3154_), .ZN(new_n3379_));
  NAND3_X1   g2737(.A1(new_n3377_), .A2(new_n3378_), .A3(new_n3379_), .ZN(new_n3380_));
  INV_X1     g2738(.I(new_n3157_), .ZN(new_n3381_));
  AOI21_X1   g2739(.A1(new_n3380_), .A2(new_n3381_), .B(new_n3272_), .ZN(new_n3382_));
  OAI21_X1   g2740(.A1(new_n3382_), .A2(new_n3170_), .B(new_n3271_), .ZN(new_n3383_));
  INV_X1     g2741(.I(new_n3175_), .ZN(new_n3384_));
  AOI21_X1   g2742(.A1(new_n3383_), .A2(new_n2726_), .B(new_n3384_), .ZN(new_n3385_));
  OAI21_X1   g2743(.A1(new_n3385_), .A2(new_n2664_), .B(new_n3270_), .ZN(new_n3386_));
  AOI21_X1   g2744(.A1(new_n3386_), .A2(new_n3191_), .B(new_n3269_), .ZN(new_n3387_));
  INV_X1     g2745(.I(new_n3195_), .ZN(new_n3388_));
  OAI21_X1   g2746(.A1(new_n3387_), .A2(new_n3268_), .B(new_n3388_), .ZN(new_n3389_));
  AOI21_X1   g2747(.A1(new_n3389_), .A2(new_n3267_), .B(new_n3266_), .ZN(new_n3390_));
  INV_X1     g2748(.I(new_n3201_), .ZN(new_n3391_));
  OAI21_X1   g2749(.A1(new_n3390_), .A2(new_n3391_), .B(new_n3265_), .ZN(new_n3392_));
  INV_X1     g2750(.I(new_n3205_), .ZN(new_n3393_));
  AOI21_X1   g2751(.A1(new_n3392_), .A2(new_n3264_), .B(new_n3393_), .ZN(new_n3394_));
  OAI21_X1   g2752(.A1(new_n3394_), .A2(new_n3263_), .B(new_n2389_), .ZN(new_n3395_));
  AOI21_X1   g2753(.A1(new_n3395_), .A2(new_n3213_), .B(new_n3262_), .ZN(new_n3396_));
  INV_X1     g2754(.I(new_n3217_), .ZN(new_n3397_));
  OAI21_X1   g2755(.A1(new_n3396_), .A2(new_n3261_), .B(new_n3397_), .ZN(new_n3398_));
  AOI21_X1   g2756(.A1(new_n3398_), .A2(new_n3260_), .B(new_n3259_), .ZN(new_n3399_));
  INV_X1     g2757(.I(new_n3223_), .ZN(new_n3400_));
  OAI21_X1   g2758(.A1(new_n3399_), .A2(new_n3400_), .B(new_n3258_), .ZN(new_n3401_));
  INV_X1     g2759(.I(new_n3227_), .ZN(new_n3402_));
  AOI21_X1   g2760(.A1(new_n3401_), .A2(new_n3257_), .B(new_n3402_), .ZN(new_n3403_));
  OAI21_X1   g2761(.A1(new_n3403_), .A2(new_n3256_), .B(new_n2198_), .ZN(new_n3404_));
  AOI21_X1   g2762(.A1(new_n3404_), .A2(new_n3235_), .B(new_n3255_), .ZN(new_n3405_));
  INV_X1     g2763(.I(new_n3239_), .ZN(new_n3406_));
  OAI21_X1   g2764(.A1(new_n3405_), .A2(new_n3254_), .B(new_n3406_), .ZN(new_n3407_));
  AOI21_X1   g2765(.A1(new_n3407_), .A2(new_n3253_), .B(new_n3252_), .ZN(new_n3408_));
  INV_X1     g2766(.I(new_n3245_), .ZN(new_n3409_));
  OAI21_X1   g2767(.A1(new_n3408_), .A2(new_n3409_), .B(new_n3251_), .ZN(new_n3410_));
  NAND4_X1   g2768(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3250_), .ZN(new_n3411_));
  OAI21_X1   g2769(.A1(\address[1] ), .A2(new_n1365_), .B(new_n3411_), .ZN(\result[0] ));
  NAND4_X1   g2770(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3010_), .ZN(new_n3413_));
  OAI21_X1   g2771(.A1(\address[1] ), .A2(new_n2916_), .B(new_n3413_), .ZN(\result[1] ));
  NAND4_X1   g2772(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2911_), .ZN(new_n3415_));
  OAI21_X1   g2773(.A1(\address[1] ), .A2(new_n2913_), .B(new_n3415_), .ZN(\result[2] ));
  NAND4_X1   g2774(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2908_), .ZN(new_n3417_));
  OAI21_X1   g2775(.A1(\address[1] ), .A2(new_n3288_), .B(new_n3417_), .ZN(\result[3] ));
  NAND4_X1   g2776(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2900_), .ZN(new_n3419_));
  OAI21_X1   g2777(.A1(\address[1] ), .A2(new_n3018_), .B(new_n3419_), .ZN(\result[4] ));
  NAND4_X1   g2778(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2893_), .ZN(new_n3421_));
  OAI21_X1   g2779(.A1(\address[1] ), .A2(new_n3022_), .B(new_n3421_), .ZN(\result[5] ));
  NAND4_X1   g2780(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3028_), .ZN(new_n3423_));
  OAI21_X1   g2781(.A1(\address[1] ), .A2(new_n3031_), .B(new_n3423_), .ZN(\result[6] ));
  NAND4_X1   g2782(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2889_), .ZN(new_n3425_));
  OAI21_X1   g2783(.A1(\address[1] ), .A2(new_n2887_), .B(new_n3425_), .ZN(\result[7] ));
  NAND4_X1   g2784(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2881_), .ZN(new_n3427_));
  OAI21_X1   g2785(.A1(\address[1] ), .A2(new_n2884_), .B(new_n3427_), .ZN(\result[8] ));
  NAND4_X1   g2786(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3041_), .ZN(new_n3429_));
  OAI21_X1   g2787(.A1(\address[1] ), .A2(new_n3046_), .B(new_n3429_), .ZN(\result[9] ));
  NAND4_X1   g2788(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2875_), .ZN(new_n3431_));
  OAI21_X1   g2789(.A1(\address[1] ), .A2(new_n3050_), .B(new_n3431_), .ZN(\result[10] ));
  NAND4_X1   g2790(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2872_), .ZN(new_n3433_));
  OAI21_X1   g2791(.A1(\address[1] ), .A2(new_n2869_), .B(new_n3433_), .ZN(\result[11] ));
  NAND4_X1   g2792(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3058_), .ZN(new_n3435_));
  OAI21_X1   g2793(.A1(\address[1] ), .A2(new_n3062_), .B(new_n3435_), .ZN(\result[12] ));
  NAND4_X1   g2794(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2862_), .ZN(new_n3437_));
  OAI21_X1   g2795(.A1(\address[1] ), .A2(new_n3065_), .B(new_n3437_), .ZN(\result[13] ));
  NAND4_X1   g2796(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2859_), .ZN(new_n3439_));
  OAI21_X1   g2797(.A1(\address[1] ), .A2(new_n3281_), .B(new_n3439_), .ZN(\result[14] ));
  NAND4_X1   g2798(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2850_), .ZN(new_n3441_));
  OAI21_X1   g2799(.A1(\address[1] ), .A2(new_n3071_), .B(new_n3441_), .ZN(\result[15] ));
  NAND4_X1   g2800(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2844_), .ZN(new_n3443_));
  OAI21_X1   g2801(.A1(\address[1] ), .A2(new_n3075_), .B(new_n3443_), .ZN(\result[16] ));
  NAND4_X1   g2802(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3081_), .ZN(new_n3445_));
  OAI21_X1   g2803(.A1(\address[1] ), .A2(new_n3085_), .B(new_n3445_), .ZN(\result[17] ));
  NAND4_X1   g2804(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2837_), .ZN(new_n3447_));
  OAI21_X1   g2805(.A1(\address[1] ), .A2(new_n3088_), .B(new_n3447_), .ZN(\result[18] ));
  NAND4_X1   g2806(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2835_), .ZN(new_n3449_));
  OAI21_X1   g2807(.A1(\address[1] ), .A2(new_n3278_), .B(new_n3449_), .ZN(\result[19] ));
  NAND4_X1   g2808(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3097_), .ZN(new_n3451_));
  OAI21_X1   g2809(.A1(\address[1] ), .A2(new_n3100_), .B(new_n3451_), .ZN(\result[20] ));
  NAND4_X1   g2810(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2826_), .ZN(new_n3453_));
  OAI21_X1   g2811(.A1(\address[1] ), .A2(new_n3104_), .B(new_n3453_), .ZN(\result[21] ));
  NAND4_X1   g2812(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2824_), .ZN(new_n3455_));
  OAI21_X1   g2813(.A1(\address[1] ), .A2(new_n2822_), .B(new_n3455_), .ZN(\result[22] ));
  NAND4_X1   g2814(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2815_), .ZN(new_n3457_));
  OAI21_X1   g2815(.A1(\address[1] ), .A2(new_n3109_), .B(new_n3457_), .ZN(\result[23] ));
  NAND4_X1   g2816(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2808_), .ZN(new_n3459_));
  OAI21_X1   g2817(.A1(\address[1] ), .A2(new_n3112_), .B(new_n3459_), .ZN(\result[24] ));
  NAND4_X1   g2818(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3119_), .ZN(new_n3461_));
  OAI21_X1   g2819(.A1(\address[1] ), .A2(new_n3124_), .B(new_n3461_), .ZN(\result[25] ));
  NAND4_X1   g2820(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2802_), .ZN(new_n3463_));
  OAI21_X1   g2821(.A1(\address[1] ), .A2(new_n3128_), .B(new_n3463_), .ZN(\result[26] ));
  NAND4_X1   g2822(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2799_), .ZN(new_n3465_));
  OAI21_X1   g2823(.A1(\address[1] ), .A2(new_n2796_), .B(new_n3465_), .ZN(\result[27] ));
  NAND4_X1   g2824(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3136_), .ZN(new_n3467_));
  OAI21_X1   g2825(.A1(\address[1] ), .A2(new_n3140_), .B(new_n3467_), .ZN(\result[28] ));
  NAND4_X1   g2826(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2789_), .ZN(new_n3469_));
  OAI21_X1   g2827(.A1(\address[1] ), .A2(new_n3143_), .B(new_n3469_), .ZN(\result[29] ));
  NAND4_X1   g2828(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2786_), .ZN(new_n3471_));
  OAI21_X1   g2829(.A1(\address[1] ), .A2(new_n3273_), .B(new_n3471_), .ZN(\result[30] ));
  NAND4_X1   g2830(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n3152_), .ZN(new_n3473_));
  OAI21_X1   g2831(.A1(\address[1] ), .A2(new_n3156_), .B(new_n3473_), .ZN(\result[31] ));
  INV_X1     g2832(.I(new_n2777_), .ZN(new_n3475_));
  NAND4_X1   g2833(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2779_), .ZN(new_n3476_));
  OAI21_X1   g2834(.A1(\address[1] ), .A2(new_n3475_), .B(new_n3476_), .ZN(\result[32] ));
  INV_X1     g2835(.I(new_n2736_), .ZN(new_n3478_));
  NAND4_X1   g2836(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2733_), .ZN(new_n3479_));
  OAI21_X1   g2837(.A1(\address[1] ), .A2(new_n3478_), .B(new_n3479_), .ZN(\result[33] ));
  NAND4_X1   g2838(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2747_), .ZN(new_n3481_));
  OAI21_X1   g2839(.A1(\address[1] ), .A2(new_n2745_), .B(new_n3481_), .ZN(\result[34] ));
  INV_X1     g2840(.I(new_n2741_), .ZN(new_n3483_));
  NAND4_X1   g2841(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2738_), .ZN(new_n3484_));
  OAI21_X1   g2842(.A1(\address[1] ), .A2(new_n3483_), .B(new_n3484_), .ZN(\result[35] ));
  INV_X1     g2843(.I(new_n2772_), .ZN(new_n3486_));
  NAND4_X1   g2844(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2769_), .ZN(new_n3487_));
  OAI21_X1   g2845(.A1(\address[1] ), .A2(new_n3486_), .B(new_n3487_), .ZN(\result[36] ));
  INV_X1     g2846(.I(new_n2754_), .ZN(new_n3489_));
  NAND4_X1   g2847(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2751_), .ZN(new_n3490_));
  OAI21_X1   g2848(.A1(\address[1] ), .A2(new_n3489_), .B(new_n3490_), .ZN(\result[37] ));
  NAND4_X1   g2849(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2762_), .ZN(new_n3492_));
  OAI21_X1   g2850(.A1(\address[1] ), .A2(new_n2765_), .B(new_n3492_), .ZN(\result[38] ));
  NAND4_X1   g2851(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2757_), .ZN(new_n3494_));
  OAI21_X1   g2852(.A1(\address[1] ), .A2(new_n2760_), .B(new_n3494_), .ZN(\result[39] ));
  NAND4_X1   g2853(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2715_), .ZN(new_n3496_));
  OAI21_X1   g2854(.A1(\address[1] ), .A2(new_n2729_), .B(new_n3496_), .ZN(\result[40] ));
  INV_X1     g2855(.I(new_n2712_), .ZN(new_n3498_));
  NAND4_X1   g2856(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2709_), .ZN(new_n3499_));
  OAI21_X1   g2857(.A1(\address[1] ), .A2(new_n3498_), .B(new_n3499_), .ZN(\result[41] ));
  NAND4_X1   g2858(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2703_), .ZN(new_n3501_));
  OAI21_X1   g2859(.A1(\address[1] ), .A2(new_n2706_), .B(new_n3501_), .ZN(\result[42] ));
  NAND4_X1   g2860(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2697_), .ZN(new_n3503_));
  OAI21_X1   g2861(.A1(\address[1] ), .A2(new_n2701_), .B(new_n3503_), .ZN(\result[43] ));
  NAND4_X1   g2862(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2688_), .ZN(new_n3505_));
  OAI21_X1   g2863(.A1(\address[1] ), .A2(new_n2691_), .B(new_n3505_), .ZN(\result[44] ));
  INV_X1     g2864(.I(new_n2684_), .ZN(new_n3507_));
  NAND4_X1   g2865(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2681_), .ZN(new_n3508_));
  OAI21_X1   g2866(.A1(\address[1] ), .A2(new_n3507_), .B(new_n3508_), .ZN(\result[45] ));
  NAND4_X1   g2867(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2674_), .ZN(new_n3510_));
  OAI21_X1   g2868(.A1(\address[1] ), .A2(new_n2677_), .B(new_n3510_), .ZN(\result[46] ));
  INV_X1     g2869(.I(new_n2671_), .ZN(new_n3512_));
  NAND4_X1   g2870(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2667_), .ZN(new_n3513_));
  OAI21_X1   g2871(.A1(\address[1] ), .A2(new_n3512_), .B(new_n3513_), .ZN(\result[47] ));
  INV_X1     g2872(.I(new_n2653_), .ZN(new_n3515_));
  NAND4_X1   g2873(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2655_), .ZN(new_n3516_));
  OAI21_X1   g2874(.A1(\address[1] ), .A2(new_n3515_), .B(new_n3516_), .ZN(\result[48] ));
  INV_X1     g2875(.I(new_n2638_), .ZN(new_n3518_));
  NAND4_X1   g2876(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2634_), .ZN(new_n3519_));
  OAI21_X1   g2877(.A1(\address[1] ), .A2(new_n3518_), .B(new_n3519_), .ZN(\result[49] ));
  NAND4_X1   g2878(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2649_), .ZN(new_n3521_));
  OAI21_X1   g2879(.A1(\address[1] ), .A2(new_n2647_), .B(new_n3521_), .ZN(\result[50] ));
  NAND4_X1   g2880(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2640_), .ZN(new_n3523_));
  OAI21_X1   g2881(.A1(\address[1] ), .A2(new_n2659_), .B(new_n3523_), .ZN(\result[51] ));
  INV_X1     g2882(.I(new_n2626_), .ZN(new_n3525_));
  NAND4_X1   g2883(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2622_), .ZN(new_n3526_));
  OAI21_X1   g2884(.A1(\address[1] ), .A2(new_n3525_), .B(new_n3526_), .ZN(\result[52] ));
  INV_X1     g2885(.I(new_n2618_), .ZN(new_n3528_));
  NAND4_X1   g2886(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2614_), .ZN(new_n3529_));
  OAI21_X1   g2887(.A1(\address[1] ), .A2(new_n3528_), .B(new_n3529_), .ZN(\result[53] ));
  NAND4_X1   g2888(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2608_), .ZN(new_n3531_));
  OAI21_X1   g2889(.A1(\address[1] ), .A2(new_n2611_), .B(new_n3531_), .ZN(\result[54] ));
  NAND4_X1   g2890(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2602_), .ZN(new_n3533_));
  OAI21_X1   g2891(.A1(\address[1] ), .A2(new_n2606_), .B(new_n3533_), .ZN(\result[55] ));
  NAND4_X1   g2892(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2557_), .ZN(new_n3535_));
  OAI21_X1   g2893(.A1(\address[1] ), .A2(new_n2560_), .B(new_n3535_), .ZN(\result[56] ));
  INV_X1     g2894(.I(new_n2554_), .ZN(new_n3537_));
  NAND4_X1   g2895(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2551_), .ZN(new_n3538_));
  OAI21_X1   g2896(.A1(\address[1] ), .A2(new_n3537_), .B(new_n3538_), .ZN(\result[57] ));
  NAND4_X1   g2897(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2595_), .ZN(new_n3540_));
  OAI21_X1   g2898(.A1(\address[1] ), .A2(new_n2598_), .B(new_n3540_), .ZN(\result[58] ));
  NAND4_X1   g2899(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2590_), .ZN(new_n3542_));
  OAI21_X1   g2900(.A1(\address[1] ), .A2(new_n2593_), .B(new_n3542_), .ZN(\result[59] ));
  NAND4_X1   g2901(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2583_), .ZN(new_n3544_));
  OAI21_X1   g2902(.A1(\address[1] ), .A2(new_n3179_), .B(new_n3544_), .ZN(\result[60] ));
  INV_X1     g2903(.I(new_n2566_), .ZN(new_n3546_));
  NAND4_X1   g2904(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2563_), .ZN(new_n3547_));
  OAI21_X1   g2905(.A1(\address[1] ), .A2(new_n3546_), .B(new_n3547_), .ZN(\result[61] ));
  NAND4_X1   g2906(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2576_), .ZN(new_n3549_));
  OAI21_X1   g2907(.A1(\address[1] ), .A2(new_n2579_), .B(new_n3549_), .ZN(\result[62] ));
  INV_X1     g2908(.I(new_n2573_), .ZN(new_n3551_));
  NAND4_X1   g2909(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2569_), .ZN(new_n3552_));
  OAI21_X1   g2910(.A1(\address[1] ), .A2(new_n3551_), .B(new_n3552_), .ZN(\result[63] ));
  INV_X1     g2911(.I(new_n2543_), .ZN(new_n3554_));
  NAND4_X1   g2912(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2539_), .ZN(new_n3555_));
  OAI21_X1   g2913(.A1(\address[1] ), .A2(new_n3554_), .B(new_n3555_), .ZN(\result[64] ));
  INV_X1     g2914(.I(new_n2536_), .ZN(new_n3557_));
  NAND4_X1   g2915(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2532_), .ZN(new_n3558_));
  OAI21_X1   g2916(.A1(\address[1] ), .A2(new_n3557_), .B(new_n3558_), .ZN(\result[65] ));
  NAND4_X1   g2917(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2526_), .ZN(new_n3560_));
  OAI21_X1   g2918(.A1(\address[1] ), .A2(new_n2529_), .B(new_n3560_), .ZN(\result[66] ));
  NAND4_X1   g2919(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2520_), .ZN(new_n3562_));
  OAI21_X1   g2920(.A1(\address[1] ), .A2(new_n2524_), .B(new_n3562_), .ZN(\result[67] ));
  NAND4_X1   g2921(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2509_), .ZN(new_n3564_));
  OAI21_X1   g2922(.A1(\address[1] ), .A2(new_n2512_), .B(new_n3564_), .ZN(\result[68] ));
  NAND4_X1   g2923(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2500_), .ZN(new_n3566_));
  OAI21_X1   g2924(.A1(\address[1] ), .A2(new_n2507_), .B(new_n3566_), .ZN(\result[69] ));
  NAND4_X1   g2925(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2492_), .ZN(new_n3568_));
  OAI21_X1   g2926(.A1(\address[1] ), .A2(new_n2495_), .B(new_n3568_), .ZN(\result[70] ));
  NAND4_X1   g2927(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2485_), .ZN(new_n3570_));
  OAI21_X1   g2928(.A1(\address[1] ), .A2(new_n2515_), .B(new_n3570_), .ZN(\result[71] ));
  INV_X1     g2929(.I(new_n2462_), .ZN(new_n3572_));
  NAND4_X1   g2930(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2458_), .ZN(new_n3573_));
  OAI21_X1   g2931(.A1(\address[1] ), .A2(new_n3572_), .B(new_n3573_), .ZN(\result[72] ));
  INV_X1     g2932(.I(new_n2481_), .ZN(new_n3575_));
  NAND4_X1   g2933(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2477_), .ZN(new_n3576_));
  OAI21_X1   g2934(.A1(\address[1] ), .A2(new_n3575_), .B(new_n3576_), .ZN(\result[73] ));
  NAND4_X1   g2935(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2470_), .ZN(new_n3578_));
  OAI21_X1   g2936(.A1(\address[1] ), .A2(new_n2473_), .B(new_n3578_), .ZN(\result[74] ));
  NAND4_X1   g2937(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2465_), .ZN(new_n3580_));
  OAI21_X1   g2938(.A1(\address[1] ), .A2(new_n2468_), .B(new_n3580_), .ZN(\result[75] ));
  NAND4_X1   g2939(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2444_), .ZN(new_n3582_));
  OAI21_X1   g2940(.A1(\address[1] ), .A2(new_n2447_), .B(new_n3582_), .ZN(\result[76] ));
  NAND4_X1   g2941(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2435_), .ZN(new_n3584_));
  OAI21_X1   g2942(.A1(\address[1] ), .A2(new_n2442_), .B(new_n3584_), .ZN(\result[77] ));
  NAND4_X1   g2943(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2427_), .ZN(new_n3586_));
  OAI21_X1   g2944(.A1(\address[1] ), .A2(new_n2430_), .B(new_n3586_), .ZN(\result[78] ));
  NAND4_X1   g2945(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2420_), .ZN(new_n3588_));
  OAI21_X1   g2946(.A1(\address[1] ), .A2(new_n2450_), .B(new_n3588_), .ZN(\result[79] ));
  INV_X1     g2947(.I(new_n2415_), .ZN(new_n3590_));
  NAND4_X1   g2948(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2411_), .ZN(new_n3591_));
  OAI21_X1   g2949(.A1(\address[1] ), .A2(new_n3590_), .B(new_n3591_), .ZN(\result[80] ));
  INV_X1     g2950(.I(new_n2408_), .ZN(new_n3593_));
  NAND4_X1   g2951(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2404_), .ZN(new_n3594_));
  OAI21_X1   g2952(.A1(\address[1] ), .A2(new_n3593_), .B(new_n3594_), .ZN(\result[81] ));
  NAND4_X1   g2953(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2398_), .ZN(new_n3596_));
  OAI21_X1   g2954(.A1(\address[1] ), .A2(new_n2401_), .B(new_n3596_), .ZN(\result[82] ));
  NAND4_X1   g2955(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2392_), .ZN(new_n3598_));
  OAI21_X1   g2956(.A1(\address[1] ), .A2(new_n2396_), .B(new_n3598_), .ZN(\result[83] ));
  INV_X1     g2957(.I(new_n2387_), .ZN(new_n3600_));
  NAND4_X1   g2958(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2383_), .ZN(new_n3601_));
  OAI21_X1   g2959(.A1(\address[1] ), .A2(new_n3600_), .B(new_n3601_), .ZN(\result[84] ));
  INV_X1     g2960(.I(new_n2365_), .ZN(new_n3603_));
  NAND4_X1   g2961(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2361_), .ZN(new_n3604_));
  OAI21_X1   g2962(.A1(\address[1] ), .A2(new_n3603_), .B(new_n3604_), .ZN(\result[85] ));
  NAND4_X1   g2963(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2375_), .ZN(new_n3606_));
  OAI21_X1   g2964(.A1(\address[1] ), .A2(new_n2378_), .B(new_n3606_), .ZN(\result[86] ));
  NAND4_X1   g2965(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2368_), .ZN(new_n3608_));
  OAI21_X1   g2966(.A1(\address[1] ), .A2(new_n3211_), .B(new_n3608_), .ZN(\result[87] ));
  INV_X1     g2967(.I(new_n2352_), .ZN(new_n3610_));
  NAND4_X1   g2968(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2348_), .ZN(new_n3611_));
  OAI21_X1   g2969(.A1(\address[1] ), .A2(new_n3610_), .B(new_n3611_), .ZN(\result[88] ));
  INV_X1     g2970(.I(new_n2345_), .ZN(new_n3613_));
  NAND4_X1   g2971(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2341_), .ZN(new_n3614_));
  OAI21_X1   g2972(.A1(\address[1] ), .A2(new_n3613_), .B(new_n3614_), .ZN(\result[89] ));
  NAND4_X1   g2973(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2335_), .ZN(new_n3616_));
  OAI21_X1   g2974(.A1(\address[1] ), .A2(new_n2338_), .B(new_n3616_), .ZN(\result[90] ));
  NAND4_X1   g2975(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2329_), .ZN(new_n3618_));
  OAI21_X1   g2976(.A1(\address[1] ), .A2(new_n2333_), .B(new_n3618_), .ZN(\result[91] ));
  NAND4_X1   g2977(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2318_), .ZN(new_n3620_));
  OAI21_X1   g2978(.A1(\address[1] ), .A2(new_n2321_), .B(new_n3620_), .ZN(\result[92] ));
  NAND4_X1   g2979(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2309_), .ZN(new_n3622_));
  OAI21_X1   g2980(.A1(\address[1] ), .A2(new_n2316_), .B(new_n3622_), .ZN(\result[93] ));
  NAND4_X1   g2981(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2301_), .ZN(new_n3624_));
  OAI21_X1   g2982(.A1(\address[1] ), .A2(new_n2304_), .B(new_n3624_), .ZN(\result[94] ));
  NAND4_X1   g2983(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2294_), .ZN(new_n3626_));
  OAI21_X1   g2984(.A1(\address[1] ), .A2(new_n2324_), .B(new_n3626_), .ZN(\result[95] ));
  INV_X1     g2985(.I(new_n2271_), .ZN(new_n3628_));
  NAND4_X1   g2986(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2267_), .ZN(new_n3629_));
  OAI21_X1   g2987(.A1(\address[1] ), .A2(new_n3628_), .B(new_n3629_), .ZN(\result[96] ));
  INV_X1     g2988(.I(new_n2290_), .ZN(new_n3631_));
  NAND4_X1   g2989(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2286_), .ZN(new_n3632_));
  OAI21_X1   g2990(.A1(\address[1] ), .A2(new_n3631_), .B(new_n3632_), .ZN(\result[97] ));
  NAND4_X1   g2991(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2279_), .ZN(new_n3634_));
  OAI21_X1   g2992(.A1(\address[1] ), .A2(new_n2282_), .B(new_n3634_), .ZN(\result[98] ));
  NAND4_X1   g2993(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2274_), .ZN(new_n3636_));
  OAI21_X1   g2994(.A1(\address[1] ), .A2(new_n2277_), .B(new_n3636_), .ZN(\result[99] ));
  NAND4_X1   g2995(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2253_), .ZN(new_n3638_));
  OAI21_X1   g2996(.A1(\address[1] ), .A2(new_n2256_), .B(new_n3638_), .ZN(\result[100] ));
  NAND4_X1   g2997(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2244_), .ZN(new_n3640_));
  OAI21_X1   g2998(.A1(\address[1] ), .A2(new_n2251_), .B(new_n3640_), .ZN(\result[101] ));
  NAND4_X1   g2999(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2236_), .ZN(new_n3642_));
  OAI21_X1   g3000(.A1(\address[1] ), .A2(new_n2239_), .B(new_n3642_), .ZN(\result[102] ));
  NAND4_X1   g3001(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2229_), .ZN(new_n3644_));
  OAI21_X1   g3002(.A1(\address[1] ), .A2(new_n2259_), .B(new_n3644_), .ZN(\result[103] ));
  INV_X1     g3003(.I(new_n2224_), .ZN(new_n3646_));
  NAND4_X1   g3004(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2220_), .ZN(new_n3647_));
  OAI21_X1   g3005(.A1(\address[1] ), .A2(new_n3646_), .B(new_n3647_), .ZN(\result[104] ));
  INV_X1     g3006(.I(new_n2217_), .ZN(new_n3649_));
  NAND4_X1   g3007(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2213_), .ZN(new_n3650_));
  OAI21_X1   g3008(.A1(\address[1] ), .A2(new_n3649_), .B(new_n3650_), .ZN(\result[105] ));
  NAND4_X1   g3009(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2207_), .ZN(new_n3652_));
  OAI21_X1   g3010(.A1(\address[1] ), .A2(new_n2210_), .B(new_n3652_), .ZN(\result[106] ));
  NAND4_X1   g3011(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2201_), .ZN(new_n3654_));
  OAI21_X1   g3012(.A1(\address[1] ), .A2(new_n2205_), .B(new_n3654_), .ZN(\result[107] ));
  INV_X1     g3013(.I(new_n2196_), .ZN(new_n3656_));
  NAND4_X1   g3014(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2192_), .ZN(new_n3657_));
  OAI21_X1   g3015(.A1(\address[1] ), .A2(new_n3656_), .B(new_n3657_), .ZN(\result[108] ));
  INV_X1     g3016(.I(new_n2174_), .ZN(new_n3659_));
  NAND4_X1   g3017(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2170_), .ZN(new_n3660_));
  OAI21_X1   g3018(.A1(\address[1] ), .A2(new_n3659_), .B(new_n3660_), .ZN(\result[109] ));
  NAND4_X1   g3019(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2184_), .ZN(new_n3662_));
  OAI21_X1   g3020(.A1(\address[1] ), .A2(new_n2187_), .B(new_n3662_), .ZN(\result[110] ));
  NAND4_X1   g3021(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2177_), .ZN(new_n3664_));
  OAI21_X1   g3022(.A1(\address[1] ), .A2(new_n3233_), .B(new_n3664_), .ZN(\result[111] ));
  INV_X1     g3023(.I(new_n2161_), .ZN(new_n3666_));
  NAND4_X1   g3024(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2157_), .ZN(new_n3667_));
  OAI21_X1   g3025(.A1(\address[1] ), .A2(new_n3666_), .B(new_n3667_), .ZN(\result[112] ));
  INV_X1     g3026(.I(new_n2154_), .ZN(new_n3669_));
  NAND4_X1   g3027(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2150_), .ZN(new_n3670_));
  OAI21_X1   g3028(.A1(\address[1] ), .A2(new_n3669_), .B(new_n3670_), .ZN(\result[113] ));
  NAND4_X1   g3029(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2144_), .ZN(new_n3672_));
  OAI21_X1   g3030(.A1(\address[1] ), .A2(new_n2147_), .B(new_n3672_), .ZN(\result[114] ));
  NAND4_X1   g3031(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2138_), .ZN(new_n3674_));
  OAI21_X1   g3032(.A1(\address[1] ), .A2(new_n2142_), .B(new_n3674_), .ZN(\result[115] ));
  NAND4_X1   g3033(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2127_), .ZN(new_n3676_));
  OAI21_X1   g3034(.A1(\address[1] ), .A2(new_n2130_), .B(new_n3676_), .ZN(\result[116] ));
  NAND4_X1   g3035(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2116_), .ZN(new_n3678_));
  OAI21_X1   g3036(.A1(\address[1] ), .A2(new_n2123_), .B(new_n3678_), .ZN(\result[117] ));
  NAND4_X1   g3037(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2108_), .ZN(new_n3680_));
  OAI21_X1   g3038(.A1(\address[1] ), .A2(new_n2111_), .B(new_n3680_), .ZN(\result[118] ));
  NAND4_X1   g3039(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2101_), .ZN(new_n3682_));
  OAI21_X1   g3040(.A1(\address[1] ), .A2(new_n2133_), .B(new_n3682_), .ZN(\result[119] ));
  INV_X1     g3041(.I(new_n2078_), .ZN(new_n3684_));
  NAND4_X1   g3042(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2074_), .ZN(new_n3685_));
  OAI21_X1   g3043(.A1(\address[1] ), .A2(new_n3684_), .B(new_n3685_), .ZN(\result[120] ));
  INV_X1     g3044(.I(new_n2097_), .ZN(new_n3687_));
  NAND4_X1   g3045(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2093_), .ZN(new_n3688_));
  OAI21_X1   g3046(.A1(\address[1] ), .A2(new_n3687_), .B(new_n3688_), .ZN(\result[121] ));
  NAND4_X1   g3047(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2086_), .ZN(new_n3690_));
  OAI21_X1   g3048(.A1(\address[1] ), .A2(new_n2089_), .B(new_n3690_), .ZN(\result[122] ));
  NAND4_X1   g3049(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n3249_), .A4(new_n2081_), .ZN(new_n3692_));
  OAI21_X1   g3050(.A1(\address[1] ), .A2(new_n2084_), .B(new_n3692_), .ZN(\result[123] ));
  NAND4_X1   g3051(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n2060_), .A4(new_n3249_), .ZN(new_n3694_));
  OAI21_X1   g3052(.A1(\address[1] ), .A2(new_n2065_), .B(new_n3694_), .ZN(\result[124] ));
  NAND4_X1   g3053(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n2054_), .A4(new_n3249_), .ZN(new_n3696_));
  OAI21_X1   g3054(.A1(\address[1] ), .A2(new_n2057_), .B(new_n3696_), .ZN(\result[125] ));
  NAND4_X1   g3055(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n2025_), .A4(new_n3249_), .ZN(new_n3698_));
  OAI21_X1   g3056(.A1(\address[1] ), .A2(new_n2052_), .B(new_n3698_), .ZN(\result[126] ));
  NOR2_X1    g3057(.A1(new_n1937_), .A2(new_n1366_), .ZN(\result[127] ));
  NAND4_X1   g3058(.A1(new_n3410_), .A2(new_n3248_), .A3(new_n2125_), .A4(new_n3249_), .ZN(new_n3702_));
  OAI21_X1   g3059(.A1(\address[1] ), .A2(new_n2049_), .B(new_n3702_), .ZN(\address[0] ));
endmodule


