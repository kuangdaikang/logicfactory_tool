// Benchmark "max" written by ABC on Thu Sep 14 20:19:42 2023

module max ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2865_, new_n2866_, new_n2867_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2879_,
    new_n2880_, new_n2881_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2888_, new_n2889_, new_n2891_, new_n2892_, new_n2893_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2905_, new_n2906_, new_n2908_, new_n2909_, new_n2910_,
    new_n2912_, new_n2913_, new_n2915_, new_n2916_, new_n2918_, new_n2919_,
    new_n2921_, new_n2922_, new_n2924_, new_n2925_, new_n2926_, new_n2928_,
    new_n2929_, new_n2931_, new_n2932_, new_n2934_, new_n2935_, new_n2936_,
    new_n2938_, new_n2939_, new_n2941_, new_n2942_, new_n2944_, new_n2945_,
    new_n2947_, new_n2948_, new_n2950_, new_n2951_, new_n2952_, new_n2954_,
    new_n2955_, new_n2957_, new_n2958_, new_n2960_, new_n2961_, new_n2962_,
    new_n2964_, new_n2965_, new_n2967_, new_n2968_, new_n2970_, new_n2971_,
    new_n2973_, new_n2974_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2981_, new_n2982_, new_n2983_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2990_, new_n2991_, new_n2992_, new_n2994_, new_n2995_,
    new_n2997_, new_n2998_, new_n3000_, new_n3001_, new_n3003_, new_n3004_,
    new_n3005_, new_n3007_, new_n3008_, new_n3010_, new_n3011_, new_n3013_,
    new_n3014_, new_n3016_, new_n3017_, new_n3019_, new_n3020_, new_n3021_,
    new_n3023_, new_n3024_, new_n3026_, new_n3027_, new_n3029_, new_n3030_,
    new_n3032_, new_n3033_, new_n3034_, new_n3036_, new_n3037_, new_n3038_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3045_, new_n3046_,
    new_n3048_, new_n3049_, new_n3050_, new_n3052_, new_n3053_, new_n3054_,
    new_n3056_, new_n3057_, new_n3058_, new_n3060_, new_n3061_, new_n3062_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3069_, new_n3070_,
    new_n3071_, new_n3073_, new_n3074_, new_n3076_, new_n3077_, new_n3079_,
    new_n3080_, new_n3082_, new_n3083_, new_n3085_, new_n3086_, new_n3088_,
    new_n3089_, new_n3090_, new_n3092_, new_n3093_, new_n3095_, new_n3096_,
    new_n3098_, new_n3099_, new_n3101_, new_n3102_, new_n3104_, new_n3105_,
    new_n3106_, new_n3108_, new_n3109_, new_n3111_, new_n3112_, new_n3114_,
    new_n3115_, new_n3116_, new_n3118_, new_n3119_, new_n3121_, new_n3122_,
    new_n3124_, new_n3125_, new_n3127_, new_n3128_, new_n3130_, new_n3131_,
    new_n3133_, new_n3134_, new_n3136_, new_n3137_, new_n3139_, new_n3140_,
    new_n3141_, new_n3143_, new_n3144_, new_n3146_, new_n3147_, new_n3148_,
    new_n3150_, new_n3151_, new_n3152_, new_n3154_, new_n3155_, new_n3156_,
    new_n3158_, new_n3159_, new_n3161_, new_n3162_, new_n3163_, new_n3165_,
    new_n3166_, new_n3167_, new_n3169_, new_n3170_, new_n3172_, new_n3173_,
    new_n3174_, new_n3176_, new_n3177_, new_n3178_, new_n3180_, new_n3181_,
    new_n3182_, new_n3184_, new_n3185_, new_n3187_, new_n3188_, new_n3190_,
    new_n3191_, new_n3193_, new_n3194_, new_n3196_, new_n3197_, new_n3199_,
    new_n3200_, new_n3202_, new_n3203_, new_n3205_, new_n3206_, new_n3208_,
    new_n3209_, new_n3211_, new_n3212_, new_n3214_, new_n3215_, new_n3217_,
    new_n3218_, new_n3220_, new_n3221_, new_n3222_, new_n3224_, new_n3225_,
    new_n3227_, new_n3228_, new_n3229_, new_n3231_, new_n3232_, new_n3233_,
    new_n3235_, new_n3236_, new_n3237_, new_n3239_, new_n3240_, new_n3242_,
    new_n3243_, new_n3244_, new_n3246_, new_n3247_, new_n3248_, new_n3250_,
    new_n3251_, new_n3253_, new_n3254_, new_n3255_, new_n3257_, new_n3258_,
    new_n3259_, new_n3261_, new_n3262_, new_n3263_, new_n3265_, new_n3266_,
    new_n3268_, new_n3269_, new_n3271_, new_n3272_, new_n3274_, new_n3275_,
    new_n3277_, new_n3278_, new_n3280_, new_n3281_, new_n3283_, new_n3284_,
    new_n3286_, new_n3287_, new_n3289_, new_n3290_, new_n3292_, new_n3293_,
    new_n3295_, new_n3296_, new_n3297_, new_n3300_, new_n3301_, new_n3302_,
    new_n3304_;
  INV_X1     g0000(.I(\in3[127] ), .ZN(new_n643_));
  NOR2_X1    g0001(.A1(new_n643_), .A2(\in2[127] ), .ZN(new_n644_));
  INV_X1     g0002(.I(\in2[29] ), .ZN(new_n645_));
  INV_X1     g0003(.I(\in2[30] ), .ZN(new_n646_));
  NOR3_X1    g0004(.A1(new_n645_), .A2(new_n646_), .A3(\in3[29] ), .ZN(new_n647_));
  INV_X1     g0005(.I(new_n647_), .ZN(new_n648_));
  INV_X1     g0006(.I(\in2[26] ), .ZN(new_n649_));
  INV_X1     g0007(.I(\in2[27] ), .ZN(new_n650_));
  NOR3_X1    g0008(.A1(new_n649_), .A2(new_n650_), .A3(\in3[26] ), .ZN(new_n651_));
  INV_X1     g0009(.I(\in3[24] ), .ZN(new_n652_));
  NOR2_X1    g0010(.A1(new_n652_), .A2(\in2[24] ), .ZN(new_n653_));
  INV_X1     g0011(.I(new_n653_), .ZN(new_n654_));
  INV_X1     g0012(.I(\in3[23] ), .ZN(new_n655_));
  NOR2_X1    g0013(.A1(new_n655_), .A2(\in2[23] ), .ZN(new_n656_));
  INV_X1     g0014(.I(\in2[21] ), .ZN(new_n657_));
  INV_X1     g0015(.I(\in2[22] ), .ZN(new_n658_));
  NOR3_X1    g0016(.A1(new_n657_), .A2(new_n658_), .A3(\in3[21] ), .ZN(new_n659_));
  INV_X1     g0017(.I(new_n659_), .ZN(new_n660_));
  INV_X1     g0018(.I(\in2[18] ), .ZN(new_n661_));
  INV_X1     g0019(.I(\in2[19] ), .ZN(new_n662_));
  NOR3_X1    g0020(.A1(new_n661_), .A2(new_n662_), .A3(\in3[18] ), .ZN(new_n663_));
  INV_X1     g0021(.I(\in3[16] ), .ZN(new_n664_));
  NOR2_X1    g0022(.A1(new_n664_), .A2(\in2[16] ), .ZN(new_n665_));
  INV_X1     g0023(.I(new_n665_), .ZN(new_n666_));
  INV_X1     g0024(.I(\in3[15] ), .ZN(new_n667_));
  NOR2_X1    g0025(.A1(new_n667_), .A2(\in2[15] ), .ZN(new_n668_));
  INV_X1     g0026(.I(\in2[13] ), .ZN(new_n669_));
  INV_X1     g0027(.I(\in2[14] ), .ZN(new_n670_));
  NOR3_X1    g0028(.A1(new_n669_), .A2(new_n670_), .A3(\in3[13] ), .ZN(new_n671_));
  INV_X1     g0029(.I(new_n671_), .ZN(new_n672_));
  INV_X1     g0030(.I(\in2[10] ), .ZN(new_n673_));
  INV_X1     g0031(.I(\in2[11] ), .ZN(new_n674_));
  NOR3_X1    g0032(.A1(new_n673_), .A2(new_n674_), .A3(\in3[10] ), .ZN(new_n675_));
  INV_X1     g0033(.I(\in3[8] ), .ZN(new_n676_));
  NOR2_X1    g0034(.A1(new_n676_), .A2(\in2[8] ), .ZN(new_n677_));
  INV_X1     g0035(.I(new_n677_), .ZN(new_n678_));
  INV_X1     g0036(.I(\in2[6] ), .ZN(new_n679_));
  INV_X1     g0037(.I(\in2[7] ), .ZN(new_n680_));
  NOR3_X1    g0038(.A1(new_n679_), .A2(new_n680_), .A3(\in3[6] ), .ZN(new_n681_));
  INV_X1     g0039(.I(\in3[4] ), .ZN(new_n682_));
  NOR2_X1    g0040(.A1(new_n682_), .A2(\in2[4] ), .ZN(new_n683_));
  INV_X1     g0041(.I(new_n683_), .ZN(new_n684_));
  INV_X1     g0042(.I(\in2[3] ), .ZN(new_n685_));
  NAND2_X1   g0043(.A1(new_n685_), .A2(\in3[3] ), .ZN(new_n686_));
  INV_X1     g0044(.I(new_n686_), .ZN(new_n687_));
  INV_X1     g0045(.I(\in2[2] ), .ZN(new_n688_));
  INV_X1     g0046(.I(\in3[2] ), .ZN(new_n689_));
  NOR2_X1    g0047(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1     g0048(.I(new_n690_), .ZN(new_n691_));
  OR3_X2     g0049(.A1(\in2[0] ), .A2(\in2[1] ), .A3(\in3[1] ), .Z(new_n692_));
  NOR2_X1    g0050(.A1(\in2[2] ), .A2(\in3[2] ), .ZN(new_n693_));
  INV_X1     g0051(.I(new_n693_), .ZN(new_n694_));
  INV_X1     g0052(.I(\in3[0] ), .ZN(new_n695_));
  NAND2_X1   g0053(.A1(new_n695_), .A2(\in2[0] ), .ZN(new_n696_));
  NOR2_X1    g0054(.A1(new_n695_), .A2(\in2[1] ), .ZN(new_n697_));
  NAND4_X1   g0055(.A1(new_n692_), .A2(new_n694_), .A3(new_n697_), .A4(new_n696_), .ZN(new_n698_));
  NOR2_X1    g0056(.A1(new_n685_), .A2(\in3[3] ), .ZN(new_n699_));
  AOI21_X1   g0057(.A1(new_n698_), .A2(new_n691_), .B(new_n699_), .ZN(new_n700_));
  NAND2_X1   g0058(.A1(new_n682_), .A2(\in2[4] ), .ZN(new_n701_));
  OAI21_X1   g0059(.A1(new_n700_), .A2(new_n687_), .B(new_n701_), .ZN(new_n702_));
  INV_X1     g0060(.I(\in3[6] ), .ZN(new_n703_));
  NOR2_X1    g0061(.A1(new_n703_), .A2(\in2[6] ), .ZN(new_n704_));
  AOI21_X1   g0062(.A1(new_n704_), .A2(\in2[5] ), .B(\in3[5] ), .ZN(new_n705_));
  AOI21_X1   g0063(.A1(new_n703_), .A2(\in2[6] ), .B(\in2[7] ), .ZN(new_n706_));
  OAI21_X1   g0064(.A1(new_n704_), .A2(\in2[5] ), .B(\in3[7] ), .ZN(new_n707_));
  NOR3_X1    g0065(.A1(new_n705_), .A2(new_n707_), .A3(new_n706_), .ZN(new_n708_));
  INV_X1     g0066(.I(new_n708_), .ZN(new_n709_));
  AOI21_X1   g0067(.A1(new_n702_), .A2(new_n684_), .B(new_n709_), .ZN(new_n710_));
  NAND2_X1   g0068(.A1(new_n676_), .A2(\in2[8] ), .ZN(new_n711_));
  OAI21_X1   g0069(.A1(new_n710_), .A2(new_n681_), .B(new_n711_), .ZN(new_n712_));
  INV_X1     g0070(.I(\in3[10] ), .ZN(new_n713_));
  NOR2_X1    g0071(.A1(new_n713_), .A2(\in2[10] ), .ZN(new_n714_));
  AOI21_X1   g0072(.A1(new_n714_), .A2(\in2[9] ), .B(\in3[9] ), .ZN(new_n715_));
  AOI21_X1   g0073(.A1(new_n713_), .A2(\in2[10] ), .B(\in2[11] ), .ZN(new_n716_));
  OAI21_X1   g0074(.A1(new_n714_), .A2(\in2[9] ), .B(\in3[11] ), .ZN(new_n717_));
  NOR3_X1    g0075(.A1(new_n715_), .A2(new_n717_), .A3(new_n716_), .ZN(new_n718_));
  INV_X1     g0076(.I(new_n718_), .ZN(new_n719_));
  AOI21_X1   g0077(.A1(new_n712_), .A2(new_n678_), .B(new_n719_), .ZN(new_n720_));
  INV_X1     g0078(.I(\in3[13] ), .ZN(new_n721_));
  NOR2_X1    g0079(.A1(new_n721_), .A2(\in2[13] ), .ZN(new_n722_));
  AOI21_X1   g0080(.A1(new_n722_), .A2(\in2[12] ), .B(\in3[12] ), .ZN(new_n723_));
  AOI21_X1   g0081(.A1(new_n721_), .A2(\in2[13] ), .B(\in2[14] ), .ZN(new_n724_));
  OAI21_X1   g0082(.A1(new_n722_), .A2(\in2[12] ), .B(\in3[14] ), .ZN(new_n725_));
  NOR3_X1    g0083(.A1(new_n723_), .A2(new_n725_), .A3(new_n724_), .ZN(new_n726_));
  OAI21_X1   g0084(.A1(new_n720_), .A2(new_n675_), .B(new_n726_), .ZN(new_n727_));
  NAND2_X1   g0085(.A1(new_n667_), .A2(\in2[15] ), .ZN(new_n728_));
  INV_X1     g0086(.I(new_n728_), .ZN(new_n729_));
  AOI21_X1   g0087(.A1(new_n727_), .A2(new_n672_), .B(new_n729_), .ZN(new_n730_));
  NAND2_X1   g0088(.A1(new_n664_), .A2(\in2[16] ), .ZN(new_n731_));
  OAI21_X1   g0089(.A1(new_n730_), .A2(new_n668_), .B(new_n731_), .ZN(new_n732_));
  INV_X1     g0090(.I(\in3[18] ), .ZN(new_n733_));
  NOR2_X1    g0091(.A1(new_n733_), .A2(\in2[18] ), .ZN(new_n734_));
  AOI21_X1   g0092(.A1(new_n734_), .A2(\in2[17] ), .B(\in3[17] ), .ZN(new_n735_));
  AOI21_X1   g0093(.A1(new_n733_), .A2(\in2[18] ), .B(\in2[19] ), .ZN(new_n736_));
  OAI21_X1   g0094(.A1(new_n734_), .A2(\in2[17] ), .B(\in3[19] ), .ZN(new_n737_));
  NOR3_X1    g0095(.A1(new_n735_), .A2(new_n737_), .A3(new_n736_), .ZN(new_n738_));
  INV_X1     g0096(.I(new_n738_), .ZN(new_n739_));
  AOI21_X1   g0097(.A1(new_n732_), .A2(new_n666_), .B(new_n739_), .ZN(new_n740_));
  INV_X1     g0098(.I(\in3[21] ), .ZN(new_n741_));
  NOR2_X1    g0099(.A1(new_n741_), .A2(\in2[21] ), .ZN(new_n742_));
  AOI21_X1   g0100(.A1(new_n742_), .A2(\in2[20] ), .B(\in3[20] ), .ZN(new_n743_));
  AOI21_X1   g0101(.A1(new_n741_), .A2(\in2[21] ), .B(\in2[22] ), .ZN(new_n744_));
  OAI21_X1   g0102(.A1(new_n742_), .A2(\in2[20] ), .B(\in3[22] ), .ZN(new_n745_));
  NOR3_X1    g0103(.A1(new_n743_), .A2(new_n745_), .A3(new_n744_), .ZN(new_n746_));
  OAI21_X1   g0104(.A1(new_n740_), .A2(new_n663_), .B(new_n746_), .ZN(new_n747_));
  NAND2_X1   g0105(.A1(new_n655_), .A2(\in2[23] ), .ZN(new_n748_));
  INV_X1     g0106(.I(new_n748_), .ZN(new_n749_));
  AOI21_X1   g0107(.A1(new_n747_), .A2(new_n660_), .B(new_n749_), .ZN(new_n750_));
  NAND2_X1   g0108(.A1(new_n652_), .A2(\in2[24] ), .ZN(new_n751_));
  OAI21_X1   g0109(.A1(new_n750_), .A2(new_n656_), .B(new_n751_), .ZN(new_n752_));
  INV_X1     g0110(.I(\in3[26] ), .ZN(new_n753_));
  NOR2_X1    g0111(.A1(new_n753_), .A2(\in2[26] ), .ZN(new_n754_));
  AOI21_X1   g0112(.A1(new_n754_), .A2(\in2[25] ), .B(\in3[25] ), .ZN(new_n755_));
  AOI21_X1   g0113(.A1(new_n753_), .A2(\in2[26] ), .B(\in2[27] ), .ZN(new_n756_));
  OAI21_X1   g0114(.A1(new_n754_), .A2(\in2[25] ), .B(\in3[27] ), .ZN(new_n757_));
  NOR3_X1    g0115(.A1(new_n755_), .A2(new_n757_), .A3(new_n756_), .ZN(new_n758_));
  INV_X1     g0116(.I(new_n758_), .ZN(new_n759_));
  AOI21_X1   g0117(.A1(new_n752_), .A2(new_n654_), .B(new_n759_), .ZN(new_n760_));
  INV_X1     g0118(.I(\in3[29] ), .ZN(new_n761_));
  NOR2_X1    g0119(.A1(new_n761_), .A2(\in2[29] ), .ZN(new_n762_));
  AOI21_X1   g0120(.A1(new_n762_), .A2(\in2[28] ), .B(\in3[28] ), .ZN(new_n763_));
  AOI21_X1   g0121(.A1(new_n761_), .A2(\in2[29] ), .B(\in2[30] ), .ZN(new_n764_));
  OAI21_X1   g0122(.A1(new_n762_), .A2(\in2[28] ), .B(\in3[30] ), .ZN(new_n765_));
  NOR3_X1    g0123(.A1(new_n763_), .A2(new_n765_), .A3(new_n764_), .ZN(new_n766_));
  OAI21_X1   g0124(.A1(new_n760_), .A2(new_n651_), .B(new_n766_), .ZN(new_n767_));
  AOI22_X1   g0125(.A1(\in2[94] ), .A2(\in3[95] ), .B1(\in2[95] ), .B2(\in3[94] ), .ZN(new_n768_));
  AOI22_X1   g0126(.A1(\in2[92] ), .A2(\in3[93] ), .B1(\in2[93] ), .B2(\in3[92] ), .ZN(new_n769_));
  INV_X1     g0127(.I(\in2[93] ), .ZN(new_n770_));
  INV_X1     g0128(.I(\in3[93] ), .ZN(new_n771_));
  NAND2_X1   g0129(.A1(\in2[92] ), .A2(\in3[92] ), .ZN(new_n772_));
  AOI21_X1   g0130(.A1(new_n770_), .A2(new_n771_), .B(new_n772_), .ZN(new_n773_));
  NOR2_X1    g0131(.A1(new_n770_), .A2(new_n771_), .ZN(new_n774_));
  NOR3_X1    g0132(.A1(new_n773_), .A2(new_n768_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1     g0133(.I(\in3[97] ), .ZN(new_n776_));
  AOI22_X1   g0134(.A1(\in2[98] ), .A2(\in3[99] ), .B1(\in2[99] ), .B2(\in3[98] ), .ZN(new_n777_));
  OAI21_X1   g0135(.A1(\in2[97] ), .A2(new_n776_), .B(new_n777_), .ZN(new_n778_));
  NAND2_X1   g0136(.A1(\in2[95] ), .A2(\in3[95] ), .ZN(new_n779_));
  NOR2_X1    g0137(.A1(\in2[95] ), .A2(\in3[95] ), .ZN(new_n780_));
  NAND2_X1   g0138(.A1(\in2[94] ), .A2(\in3[94] ), .ZN(new_n781_));
  OAI21_X1   g0139(.A1(new_n780_), .A2(new_n781_), .B(new_n779_), .ZN(new_n782_));
  NAND4_X1   g0140(.A1(new_n778_), .A2(\in2[96] ), .A3(\in3[96] ), .A4(new_n782_), .ZN(new_n783_));
  OAI22_X1   g0141(.A1(new_n783_), .A2(new_n775_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n784_));
  INV_X1     g0142(.I(\in3[105] ), .ZN(new_n785_));
  NOR2_X1    g0143(.A1(new_n785_), .A2(\in2[105] ), .ZN(new_n786_));
  INV_X1     g0144(.I(\in2[106] ), .ZN(new_n787_));
  INV_X1     g0145(.I(\in2[107] ), .ZN(new_n788_));
  INV_X1     g0146(.I(\in3[106] ), .ZN(new_n789_));
  INV_X1     g0147(.I(\in3[107] ), .ZN(new_n790_));
  OAI22_X1   g0148(.A1(new_n787_), .A2(new_n790_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n791_));
  NOR2_X1    g0149(.A1(new_n791_), .A2(new_n786_), .ZN(new_n792_));
  NAND2_X1   g0150(.A1(\in2[104] ), .A2(\in3[104] ), .ZN(new_n793_));
  INV_X1     g0151(.I(\in2[104] ), .ZN(new_n794_));
  INV_X1     g0152(.I(\in3[104] ), .ZN(new_n795_));
  NAND2_X1   g0153(.A1(\in2[106] ), .A2(\in3[105] ), .ZN(new_n796_));
  NAND2_X1   g0154(.A1(\in2[105] ), .A2(\in3[106] ), .ZN(new_n797_));
  NAND4_X1   g0155(.A1(new_n796_), .A2(new_n797_), .A3(new_n794_), .A4(new_n795_), .ZN(new_n798_));
  NOR3_X1    g0156(.A1(new_n788_), .A2(new_n785_), .A3(\in2[105] ), .ZN(new_n799_));
  AOI22_X1   g0157(.A1(new_n798_), .A2(new_n799_), .B1(new_n791_), .B2(\in3[107] ), .ZN(new_n800_));
  AOI22_X1   g0158(.A1(\in2[110] ), .A2(\in3[111] ), .B1(\in2[111] ), .B2(\in3[110] ), .ZN(new_n801_));
  AOI22_X1   g0159(.A1(\in2[108] ), .A2(\in3[109] ), .B1(\in2[109] ), .B2(\in3[108] ), .ZN(new_n802_));
  OR2_X2     g0160(.A1(new_n801_), .A2(new_n802_), .Z(new_n803_));
  OAI22_X1   g0161(.A1(new_n800_), .A2(new_n803_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n804_));
  INV_X1     g0162(.I(\in2[111] ), .ZN(new_n805_));
  INV_X1     g0163(.I(\in3[111] ), .ZN(new_n806_));
  NOR2_X1    g0164(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1   g0165(.A1(new_n805_), .A2(new_n806_), .ZN(new_n808_));
  AND2_X2    g0166(.A1(\in2[110] ), .A2(\in3[110] ), .Z(new_n809_));
  AOI21_X1   g0167(.A1(new_n808_), .A2(new_n809_), .B(new_n807_), .ZN(new_n810_));
  INV_X1     g0168(.I(\in2[109] ), .ZN(new_n811_));
  INV_X1     g0169(.I(\in3[109] ), .ZN(new_n812_));
  NAND2_X1   g0170(.A1(\in2[108] ), .A2(\in3[108] ), .ZN(new_n813_));
  AOI21_X1   g0171(.A1(new_n811_), .A2(new_n812_), .B(new_n813_), .ZN(new_n814_));
  NOR2_X1    g0172(.A1(new_n811_), .A2(new_n812_), .ZN(new_n815_));
  NOR3_X1    g0173(.A1(new_n814_), .A2(new_n801_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1     g0174(.I(\in2[114] ), .ZN(new_n817_));
  INV_X1     g0175(.I(\in2[115] ), .ZN(new_n818_));
  INV_X1     g0176(.I(\in3[114] ), .ZN(new_n819_));
  INV_X1     g0177(.I(\in3[115] ), .ZN(new_n820_));
  OAI22_X1   g0178(.A1(new_n817_), .A2(new_n820_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n821_));
  INV_X1     g0179(.I(\in2[112] ), .ZN(new_n822_));
  INV_X1     g0180(.I(\in3[112] ), .ZN(new_n823_));
  NAND2_X1   g0181(.A1(\in2[114] ), .A2(\in3[113] ), .ZN(new_n824_));
  NAND2_X1   g0182(.A1(\in2[113] ), .A2(\in3[114] ), .ZN(new_n825_));
  NAND4_X1   g0183(.A1(new_n824_), .A2(new_n825_), .A3(new_n822_), .A4(new_n823_), .ZN(new_n826_));
  INV_X1     g0184(.I(\in3[113] ), .ZN(new_n827_));
  NOR3_X1    g0185(.A1(new_n818_), .A2(new_n827_), .A3(\in2[113] ), .ZN(new_n828_));
  AOI22_X1   g0186(.A1(new_n826_), .A2(new_n828_), .B1(new_n821_), .B2(\in3[115] ), .ZN(new_n829_));
  NOR2_X1    g0187(.A1(new_n827_), .A2(\in2[113] ), .ZN(new_n830_));
  NOR2_X1    g0188(.A1(new_n822_), .A2(new_n823_), .ZN(new_n831_));
  OAI21_X1   g0189(.A1(new_n821_), .A2(new_n830_), .B(new_n831_), .ZN(new_n832_));
  OAI22_X1   g0190(.A1(new_n829_), .A2(new_n832_), .B1(new_n810_), .B2(new_n816_), .ZN(new_n833_));
  AOI22_X1   g0191(.A1(\in2[118] ), .A2(\in3[119] ), .B1(\in2[119] ), .B2(\in3[118] ), .ZN(new_n834_));
  AOI22_X1   g0192(.A1(\in2[116] ), .A2(\in3[117] ), .B1(\in2[117] ), .B2(\in3[116] ), .ZN(new_n835_));
  INV_X1     g0193(.I(\in2[117] ), .ZN(new_n836_));
  INV_X1     g0194(.I(\in3[117] ), .ZN(new_n837_));
  NAND2_X1   g0195(.A1(\in2[116] ), .A2(\in3[116] ), .ZN(new_n838_));
  AOI21_X1   g0196(.A1(new_n836_), .A2(new_n837_), .B(new_n838_), .ZN(new_n839_));
  NOR2_X1    g0197(.A1(new_n836_), .A2(new_n837_), .ZN(new_n840_));
  NOR3_X1    g0198(.A1(new_n839_), .A2(new_n834_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1     g0199(.I(\in3[121] ), .ZN(new_n842_));
  AOI22_X1   g0200(.A1(\in2[122] ), .A2(\in3[123] ), .B1(\in2[123] ), .B2(\in3[122] ), .ZN(new_n843_));
  OAI21_X1   g0201(.A1(\in2[121] ), .A2(new_n842_), .B(new_n843_), .ZN(new_n844_));
  NAND2_X1   g0202(.A1(\in2[119] ), .A2(\in3[119] ), .ZN(new_n845_));
  NOR2_X1    g0203(.A1(\in2[119] ), .A2(\in3[119] ), .ZN(new_n846_));
  NAND2_X1   g0204(.A1(\in2[118] ), .A2(\in3[118] ), .ZN(new_n847_));
  OAI21_X1   g0205(.A1(new_n846_), .A2(new_n847_), .B(new_n845_), .ZN(new_n848_));
  NAND4_X1   g0206(.A1(new_n844_), .A2(\in2[120] ), .A3(\in3[120] ), .A4(new_n848_), .ZN(new_n849_));
  OAI22_X1   g0207(.A1(new_n849_), .A2(new_n841_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n850_));
  NAND4_X1   g0208(.A1(new_n784_), .A2(new_n850_), .A3(new_n804_), .A4(new_n833_), .ZN(new_n851_));
  AOI22_X1   g0209(.A1(\in2[124] ), .A2(\in2[127] ), .B1(\in3[124] ), .B2(\in3[127] ), .ZN(new_n852_));
  AOI22_X1   g0210(.A1(\in2[125] ), .A2(\in3[126] ), .B1(\in2[126] ), .B2(\in3[125] ), .ZN(new_n853_));
  INV_X1     g0211(.I(\in2[127] ), .ZN(new_n854_));
  NOR2_X1    g0212(.A1(new_n854_), .A2(\in3[127] ), .ZN(new_n855_));
  OR3_X2     g0213(.A1(new_n852_), .A2(new_n853_), .A3(new_n855_), .Z(new_n856_));
  INV_X1     g0214(.I(\in2[126] ), .ZN(new_n857_));
  INV_X1     g0215(.I(\in3[126] ), .ZN(new_n858_));
  AOI22_X1   g0216(.A1(\in2[124] ), .A2(\in3[125] ), .B1(\in2[125] ), .B2(\in3[124] ), .ZN(new_n859_));
  OAI22_X1   g0217(.A1(new_n857_), .A2(new_n859_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n860_));
  INV_X1     g0218(.I(new_n843_), .ZN(new_n861_));
  INV_X1     g0219(.I(\in2[120] ), .ZN(new_n862_));
  INV_X1     g0220(.I(\in3[120] ), .ZN(new_n863_));
  NAND2_X1   g0221(.A1(\in2[122] ), .A2(\in3[121] ), .ZN(new_n864_));
  NAND2_X1   g0222(.A1(\in2[121] ), .A2(\in3[122] ), .ZN(new_n865_));
  NAND4_X1   g0223(.A1(new_n864_), .A2(new_n865_), .A3(new_n862_), .A4(new_n863_), .ZN(new_n866_));
  INV_X1     g0224(.I(\in2[123] ), .ZN(new_n867_));
  NOR3_X1    g0225(.A1(new_n867_), .A2(new_n842_), .A3(\in2[121] ), .ZN(new_n868_));
  AOI22_X1   g0226(.A1(new_n866_), .A2(new_n868_), .B1(new_n861_), .B2(\in3[123] ), .ZN(new_n869_));
  OAI21_X1   g0227(.A1(new_n856_), .A2(new_n860_), .B(new_n869_), .ZN(new_n870_));
  INV_X1     g0228(.I(\in2[77] ), .ZN(new_n871_));
  INV_X1     g0229(.I(\in3[77] ), .ZN(new_n872_));
  NAND2_X1   g0230(.A1(\in2[76] ), .A2(\in3[76] ), .ZN(new_n873_));
  AOI21_X1   g0231(.A1(new_n871_), .A2(new_n872_), .B(new_n873_), .ZN(new_n874_));
  AOI22_X1   g0232(.A1(\in2[78] ), .A2(\in3[79] ), .B1(\in2[79] ), .B2(\in3[78] ), .ZN(new_n875_));
  NOR2_X1    g0233(.A1(new_n871_), .A2(new_n872_), .ZN(new_n876_));
  NOR3_X1    g0234(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  NOR2_X1    g0235(.A1(\in2[79] ), .A2(\in3[79] ), .ZN(new_n878_));
  NAND2_X1   g0236(.A1(\in2[78] ), .A2(\in3[78] ), .ZN(new_n879_));
  NOR2_X1    g0237(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1   g0238(.A1(\in2[79] ), .A2(\in3[79] ), .B(new_n880_), .ZN(new_n881_));
  AOI22_X1   g0239(.A1(\in2[76] ), .A2(\in3[77] ), .B1(\in2[77] ), .B2(\in3[76] ), .ZN(new_n882_));
  OR3_X2     g0240(.A1(new_n881_), .A2(new_n875_), .A3(new_n882_), .Z(new_n883_));
  AOI22_X1   g0241(.A1(\in2[74] ), .A2(\in3[75] ), .B1(\in2[75] ), .B2(\in3[74] ), .ZN(new_n884_));
  INV_X1     g0242(.I(new_n884_), .ZN(new_n885_));
  INV_X1     g0243(.I(\in2[72] ), .ZN(new_n886_));
  INV_X1     g0244(.I(\in3[72] ), .ZN(new_n887_));
  NAND2_X1   g0245(.A1(\in2[74] ), .A2(\in3[73] ), .ZN(new_n888_));
  NAND2_X1   g0246(.A1(\in2[73] ), .A2(\in3[74] ), .ZN(new_n889_));
  NAND4_X1   g0247(.A1(new_n888_), .A2(new_n889_), .A3(new_n886_), .A4(new_n887_), .ZN(new_n890_));
  INV_X1     g0248(.I(\in2[75] ), .ZN(new_n891_));
  INV_X1     g0249(.I(\in3[73] ), .ZN(new_n892_));
  NOR3_X1    g0250(.A1(new_n891_), .A2(new_n892_), .A3(\in2[73] ), .ZN(new_n893_));
  AOI22_X1   g0251(.A1(new_n890_), .A2(new_n893_), .B1(new_n885_), .B2(\in3[75] ), .ZN(new_n894_));
  OAI21_X1   g0252(.A1(new_n883_), .A2(new_n877_), .B(new_n894_), .ZN(new_n895_));
  INV_X1     g0253(.I(\in2[101] ), .ZN(new_n896_));
  INV_X1     g0254(.I(\in3[101] ), .ZN(new_n897_));
  NAND2_X1   g0255(.A1(\in2[100] ), .A2(\in3[100] ), .ZN(new_n898_));
  AOI21_X1   g0256(.A1(new_n896_), .A2(new_n897_), .B(new_n898_), .ZN(new_n899_));
  AOI22_X1   g0257(.A1(\in2[102] ), .A2(\in3[103] ), .B1(\in2[103] ), .B2(\in3[102] ), .ZN(new_n900_));
  NOR2_X1    g0258(.A1(new_n896_), .A2(new_n897_), .ZN(new_n901_));
  NOR3_X1    g0259(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  NOR2_X1    g0260(.A1(\in2[103] ), .A2(\in3[103] ), .ZN(new_n903_));
  NAND2_X1   g0261(.A1(\in2[102] ), .A2(\in3[102] ), .ZN(new_n904_));
  NOR2_X1    g0262(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1   g0263(.A1(\in2[103] ), .A2(\in3[103] ), .B(new_n905_), .ZN(new_n906_));
  AOI22_X1   g0264(.A1(\in2[100] ), .A2(\in3[101] ), .B1(\in2[101] ), .B2(\in3[100] ), .ZN(new_n907_));
  OR3_X2     g0265(.A1(new_n906_), .A2(new_n900_), .A3(new_n907_), .Z(new_n908_));
  INV_X1     g0266(.I(new_n777_), .ZN(new_n909_));
  INV_X1     g0267(.I(\in2[96] ), .ZN(new_n910_));
  INV_X1     g0268(.I(\in3[96] ), .ZN(new_n911_));
  NAND2_X1   g0269(.A1(\in2[98] ), .A2(\in3[97] ), .ZN(new_n912_));
  NAND2_X1   g0270(.A1(\in2[97] ), .A2(\in3[98] ), .ZN(new_n913_));
  NAND4_X1   g0271(.A1(new_n912_), .A2(new_n913_), .A3(new_n910_), .A4(new_n911_), .ZN(new_n914_));
  INV_X1     g0272(.I(\in2[99] ), .ZN(new_n915_));
  NOR3_X1    g0273(.A1(new_n915_), .A2(new_n776_), .A3(\in2[97] ), .ZN(new_n916_));
  AOI22_X1   g0274(.A1(new_n914_), .A2(new_n916_), .B1(new_n909_), .B2(\in3[99] ), .ZN(new_n917_));
  OAI21_X1   g0275(.A1(new_n908_), .A2(new_n902_), .B(new_n917_), .ZN(new_n918_));
  NAND3_X1   g0276(.A1(new_n895_), .A2(new_n918_), .A3(new_n870_), .ZN(new_n919_));
  AOI22_X1   g0277(.A1(\in2[70] ), .A2(\in3[71] ), .B1(\in2[71] ), .B2(\in3[70] ), .ZN(new_n920_));
  AOI22_X1   g0278(.A1(\in2[68] ), .A2(\in3[69] ), .B1(\in2[69] ), .B2(\in3[68] ), .ZN(new_n921_));
  INV_X1     g0279(.I(\in2[69] ), .ZN(new_n922_));
  INV_X1     g0280(.I(\in3[69] ), .ZN(new_n923_));
  NAND2_X1   g0281(.A1(\in2[68] ), .A2(\in3[68] ), .ZN(new_n924_));
  AOI21_X1   g0282(.A1(new_n922_), .A2(new_n923_), .B(new_n924_), .ZN(new_n925_));
  NOR2_X1    g0283(.A1(new_n922_), .A2(new_n923_), .ZN(new_n926_));
  NOR3_X1    g0284(.A1(new_n925_), .A2(new_n920_), .A3(new_n926_), .ZN(new_n927_));
  OAI21_X1   g0285(.A1(\in2[73] ), .A2(new_n892_), .B(new_n884_), .ZN(new_n928_));
  NAND2_X1   g0286(.A1(\in2[71] ), .A2(\in3[71] ), .ZN(new_n929_));
  NOR2_X1    g0287(.A1(\in2[71] ), .A2(\in3[71] ), .ZN(new_n930_));
  NAND2_X1   g0288(.A1(\in2[70] ), .A2(\in3[70] ), .ZN(new_n931_));
  OAI21_X1   g0289(.A1(new_n930_), .A2(new_n931_), .B(new_n929_), .ZN(new_n932_));
  NAND4_X1   g0290(.A1(new_n928_), .A2(\in2[72] ), .A3(\in3[72] ), .A4(new_n932_), .ZN(new_n933_));
  OAI22_X1   g0291(.A1(new_n933_), .A2(new_n927_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n934_));
  INV_X1     g0292(.I(\in2[31] ), .ZN(new_n935_));
  AOI22_X1   g0293(.A1(\in2[38] ), .A2(\in3[39] ), .B1(\in2[39] ), .B2(\in3[38] ), .ZN(new_n936_));
  NAND2_X1   g0294(.A1(\in2[37] ), .A2(\in3[36] ), .ZN(new_n937_));
  NAND2_X1   g0295(.A1(\in2[36] ), .A2(\in3[37] ), .ZN(new_n938_));
  AOI21_X1   g0296(.A1(new_n937_), .A2(new_n938_), .B(new_n936_), .ZN(new_n939_));
  INV_X1     g0297(.I(\in2[32] ), .ZN(new_n940_));
  INV_X1     g0298(.I(\in2[33] ), .ZN(new_n941_));
  INV_X1     g0299(.I(\in3[32] ), .ZN(new_n942_));
  INV_X1     g0300(.I(\in3[33] ), .ZN(new_n943_));
  OAI22_X1   g0301(.A1(new_n940_), .A2(new_n943_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n944_));
  INV_X1     g0302(.I(\in2[34] ), .ZN(new_n945_));
  INV_X1     g0303(.I(\in2[35] ), .ZN(new_n946_));
  INV_X1     g0304(.I(\in3[34] ), .ZN(new_n947_));
  INV_X1     g0305(.I(\in3[35] ), .ZN(new_n948_));
  OAI22_X1   g0306(.A1(new_n945_), .A2(new_n948_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n949_));
  NAND3_X1   g0307(.A1(new_n939_), .A2(new_n944_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1   g0308(.A1(new_n950_), .A2(new_n935_), .ZN(new_n951_));
  INV_X1     g0309(.I(\in3[31] ), .ZN(new_n952_));
  OAI21_X1   g0310(.A1(new_n950_), .A2(new_n935_), .B(new_n952_), .ZN(new_n953_));
  NAND3_X1   g0311(.A1(new_n934_), .A2(new_n951_), .A3(new_n953_), .ZN(new_n954_));
  INV_X1     g0312(.I(\in3[81] ), .ZN(new_n955_));
  NOR2_X1    g0313(.A1(new_n955_), .A2(\in2[81] ), .ZN(new_n956_));
  INV_X1     g0314(.I(\in2[82] ), .ZN(new_n957_));
  INV_X1     g0315(.I(\in2[83] ), .ZN(new_n958_));
  INV_X1     g0316(.I(\in3[82] ), .ZN(new_n959_));
  INV_X1     g0317(.I(\in3[83] ), .ZN(new_n960_));
  OAI22_X1   g0318(.A1(new_n957_), .A2(new_n960_), .B1(new_n958_), .B2(new_n959_), .ZN(new_n961_));
  NOR2_X1    g0319(.A1(new_n961_), .A2(new_n956_), .ZN(new_n962_));
  NAND2_X1   g0320(.A1(\in2[80] ), .A2(\in3[80] ), .ZN(new_n963_));
  INV_X1     g0321(.I(\in2[80] ), .ZN(new_n964_));
  INV_X1     g0322(.I(\in3[80] ), .ZN(new_n965_));
  NAND2_X1   g0323(.A1(\in2[82] ), .A2(\in3[81] ), .ZN(new_n966_));
  NAND2_X1   g0324(.A1(\in2[81] ), .A2(\in3[82] ), .ZN(new_n967_));
  NAND4_X1   g0325(.A1(new_n966_), .A2(new_n967_), .A3(new_n964_), .A4(new_n965_), .ZN(new_n968_));
  NOR3_X1    g0326(.A1(new_n958_), .A2(new_n955_), .A3(\in2[81] ), .ZN(new_n969_));
  AOI22_X1   g0327(.A1(new_n968_), .A2(new_n969_), .B1(new_n961_), .B2(\in3[83] ), .ZN(new_n970_));
  AOI22_X1   g0328(.A1(\in2[86] ), .A2(\in3[87] ), .B1(\in2[87] ), .B2(\in3[86] ), .ZN(new_n971_));
  AOI22_X1   g0329(.A1(\in2[84] ), .A2(\in3[85] ), .B1(\in2[85] ), .B2(\in3[84] ), .ZN(new_n972_));
  OR2_X2     g0330(.A1(new_n971_), .A2(new_n972_), .Z(new_n973_));
  OAI22_X1   g0331(.A1(new_n970_), .A2(new_n973_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n974_));
  INV_X1     g0332(.I(\in2[87] ), .ZN(new_n975_));
  INV_X1     g0333(.I(\in3[87] ), .ZN(new_n976_));
  NOR2_X1    g0334(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  NAND2_X1   g0335(.A1(new_n975_), .A2(new_n976_), .ZN(new_n978_));
  AND2_X2    g0336(.A1(\in2[86] ), .A2(\in3[86] ), .Z(new_n979_));
  AOI21_X1   g0337(.A1(new_n978_), .A2(new_n979_), .B(new_n977_), .ZN(new_n980_));
  INV_X1     g0338(.I(\in2[85] ), .ZN(new_n981_));
  INV_X1     g0339(.I(\in3[85] ), .ZN(new_n982_));
  NAND2_X1   g0340(.A1(\in2[84] ), .A2(\in3[84] ), .ZN(new_n983_));
  AOI21_X1   g0341(.A1(new_n981_), .A2(new_n982_), .B(new_n983_), .ZN(new_n984_));
  NOR2_X1    g0342(.A1(new_n981_), .A2(new_n982_), .ZN(new_n985_));
  NOR3_X1    g0343(.A1(new_n984_), .A2(new_n971_), .A3(new_n985_), .ZN(new_n986_));
  INV_X1     g0344(.I(\in2[90] ), .ZN(new_n987_));
  INV_X1     g0345(.I(\in2[91] ), .ZN(new_n988_));
  INV_X1     g0346(.I(\in3[90] ), .ZN(new_n989_));
  INV_X1     g0347(.I(\in3[91] ), .ZN(new_n990_));
  OAI22_X1   g0348(.A1(new_n987_), .A2(new_n990_), .B1(new_n988_), .B2(new_n989_), .ZN(new_n991_));
  INV_X1     g0349(.I(\in2[88] ), .ZN(new_n992_));
  INV_X1     g0350(.I(\in3[88] ), .ZN(new_n993_));
  NAND2_X1   g0351(.A1(\in2[90] ), .A2(\in3[89] ), .ZN(new_n994_));
  NAND2_X1   g0352(.A1(\in2[89] ), .A2(\in3[90] ), .ZN(new_n995_));
  NAND4_X1   g0353(.A1(new_n994_), .A2(new_n995_), .A3(new_n992_), .A4(new_n993_), .ZN(new_n996_));
  INV_X1     g0354(.I(\in3[89] ), .ZN(new_n997_));
  NOR3_X1    g0355(.A1(new_n988_), .A2(new_n997_), .A3(\in2[89] ), .ZN(new_n998_));
  AOI22_X1   g0356(.A1(new_n996_), .A2(new_n998_), .B1(new_n991_), .B2(\in3[91] ), .ZN(new_n999_));
  NOR2_X1    g0357(.A1(new_n997_), .A2(\in2[89] ), .ZN(new_n1000_));
  NOR2_X1    g0358(.A1(new_n992_), .A2(new_n993_), .ZN(new_n1001_));
  OAI21_X1   g0359(.A1(new_n991_), .A2(new_n1000_), .B(new_n1001_), .ZN(new_n1002_));
  OAI22_X1   g0360(.A1(new_n999_), .A2(new_n1002_), .B1(new_n980_), .B2(new_n986_), .ZN(new_n1003_));
  NAND2_X1   g0361(.A1(new_n1003_), .A2(new_n974_), .ZN(new_n1004_));
  NOR4_X1    g0362(.A1(new_n919_), .A2(new_n851_), .A3(new_n954_), .A4(new_n1004_), .ZN(new_n1005_));
  INV_X1     g0363(.I(\in2[59] ), .ZN(new_n1006_));
  AOI22_X1   g0364(.A1(\in2[57] ), .A2(\in3[58] ), .B1(\in2[58] ), .B2(\in3[57] ), .ZN(new_n1007_));
  OR2_X2     g0365(.A1(\in2[56] ), .A2(\in3[56] ), .Z(new_n1008_));
  AND2_X2    g0366(.A1(\in2[57] ), .A2(\in3[57] ), .Z(new_n1009_));
  AOI21_X1   g0367(.A1(new_n1009_), .A2(new_n1008_), .B(new_n1007_), .ZN(new_n1010_));
  NAND2_X1   g0368(.A1(\in2[63] ), .A2(\in3[62] ), .ZN(new_n1011_));
  NAND2_X1   g0369(.A1(\in2[62] ), .A2(\in3[63] ), .ZN(new_n1012_));
  NAND2_X1   g0370(.A1(new_n1011_), .A2(new_n1012_), .ZN(new_n1013_));
  NAND2_X1   g0371(.A1(\in2[61] ), .A2(\in3[60] ), .ZN(new_n1014_));
  NAND2_X1   g0372(.A1(\in2[60] ), .A2(\in3[61] ), .ZN(new_n1015_));
  NAND2_X1   g0373(.A1(new_n1014_), .A2(new_n1015_), .ZN(new_n1016_));
  INV_X1     g0374(.I(\in2[58] ), .ZN(new_n1017_));
  INV_X1     g0375(.I(\in3[58] ), .ZN(new_n1018_));
  INV_X1     g0376(.I(\in3[59] ), .ZN(new_n1019_));
  OAI22_X1   g0377(.A1(new_n1017_), .A2(new_n1019_), .B1(new_n1006_), .B2(new_n1018_), .ZN(new_n1020_));
  NAND3_X1   g0378(.A1(new_n1020_), .A2(new_n1013_), .A3(new_n1016_), .ZN(new_n1021_));
  OAI21_X1   g0379(.A1(new_n1021_), .A2(new_n1010_), .B(new_n1006_), .ZN(new_n1022_));
  NAND2_X1   g0380(.A1(\in2[63] ), .A2(\in3[63] ), .ZN(new_n1023_));
  NOR2_X1    g0381(.A1(\in2[63] ), .A2(\in3[63] ), .ZN(new_n1024_));
  NAND2_X1   g0382(.A1(\in2[62] ), .A2(\in3[62] ), .ZN(new_n1025_));
  OAI21_X1   g0383(.A1(new_n1024_), .A2(new_n1025_), .B(new_n1023_), .ZN(new_n1026_));
  AOI21_X1   g0384(.A1(new_n1022_), .A2(\in3[59] ), .B(new_n1026_), .ZN(new_n1027_));
  NAND2_X1   g0385(.A1(\in2[61] ), .A2(\in3[61] ), .ZN(new_n1028_));
  NOR2_X1    g0386(.A1(\in2[61] ), .A2(\in3[61] ), .ZN(new_n1029_));
  NAND2_X1   g0387(.A1(\in2[60] ), .A2(\in3[60] ), .ZN(new_n1030_));
  OAI21_X1   g0388(.A1(new_n1029_), .A2(new_n1030_), .B(new_n1028_), .ZN(new_n1031_));
  NAND2_X1   g0389(.A1(new_n1031_), .A2(new_n1013_), .ZN(new_n1032_));
  INV_X1     g0390(.I(\in3[67] ), .ZN(new_n1033_));
  AOI22_X1   g0391(.A1(\in2[66] ), .A2(\in3[67] ), .B1(\in2[67] ), .B2(\in3[66] ), .ZN(new_n1034_));
  NOR2_X1    g0392(.A1(new_n1034_), .A2(new_n1033_), .ZN(new_n1035_));
  NAND2_X1   g0393(.A1(\in2[66] ), .A2(\in3[65] ), .ZN(new_n1036_));
  INV_X1     g0394(.I(\in2[65] ), .ZN(new_n1037_));
  INV_X1     g0395(.I(\in3[66] ), .ZN(new_n1038_));
  NOR2_X1    g0396(.A1(new_n1037_), .A2(new_n1038_), .ZN(new_n1039_));
  NOR3_X1    g0397(.A1(new_n1039_), .A2(\in2[64] ), .A3(\in3[64] ), .ZN(new_n1040_));
  NAND3_X1   g0398(.A1(new_n1037_), .A2(\in2[67] ), .A3(\in3[65] ), .ZN(new_n1041_));
  AOI21_X1   g0399(.A1(new_n1040_), .A2(new_n1036_), .B(new_n1041_), .ZN(new_n1042_));
  NOR2_X1    g0400(.A1(new_n1042_), .A2(new_n1035_), .ZN(new_n1043_));
  INV_X1     g0401(.I(\in3[65] ), .ZN(new_n1044_));
  OAI21_X1   g0402(.A1(\in2[65] ), .A2(new_n1044_), .B(new_n1034_), .ZN(new_n1045_));
  NAND3_X1   g0403(.A1(new_n1045_), .A2(\in2[64] ), .A3(\in3[64] ), .ZN(new_n1046_));
  OAI22_X1   g0404(.A1(new_n1027_), .A2(new_n1032_), .B1(new_n1043_), .B2(new_n1046_), .ZN(new_n1047_));
  AOI22_X1   g0405(.A1(\in2[33] ), .A2(\in3[34] ), .B1(\in2[34] ), .B2(\in3[33] ), .ZN(new_n1048_));
  NAND2_X1   g0406(.A1(new_n940_), .A2(new_n942_), .ZN(new_n1049_));
  NOR2_X1    g0407(.A1(new_n941_), .A2(new_n943_), .ZN(new_n1050_));
  AOI21_X1   g0408(.A1(new_n1050_), .A2(new_n1049_), .B(new_n1048_), .ZN(new_n1051_));
  NAND2_X1   g0409(.A1(new_n939_), .A2(new_n949_), .ZN(new_n1052_));
  OAI21_X1   g0410(.A1(new_n1052_), .A2(new_n1051_), .B(new_n946_), .ZN(new_n1053_));
  NAND2_X1   g0411(.A1(\in2[39] ), .A2(\in3[39] ), .ZN(new_n1054_));
  NOR2_X1    g0412(.A1(\in2[39] ), .A2(\in3[39] ), .ZN(new_n1055_));
  NAND2_X1   g0413(.A1(\in2[38] ), .A2(\in3[38] ), .ZN(new_n1056_));
  OAI21_X1   g0414(.A1(new_n1055_), .A2(new_n1056_), .B(new_n1054_), .ZN(new_n1057_));
  AOI21_X1   g0415(.A1(new_n1053_), .A2(\in3[35] ), .B(new_n1057_), .ZN(new_n1058_));
  INV_X1     g0416(.I(new_n936_), .ZN(new_n1059_));
  NAND2_X1   g0417(.A1(\in2[37] ), .A2(\in3[37] ), .ZN(new_n1060_));
  NOR2_X1    g0418(.A1(\in2[37] ), .A2(\in3[37] ), .ZN(new_n1061_));
  NAND2_X1   g0419(.A1(\in2[36] ), .A2(\in3[36] ), .ZN(new_n1062_));
  OAI21_X1   g0420(.A1(new_n1061_), .A2(new_n1062_), .B(new_n1060_), .ZN(new_n1063_));
  NAND2_X1   g0421(.A1(new_n1063_), .A2(new_n1059_), .ZN(new_n1064_));
  INV_X1     g0422(.I(\in2[43] ), .ZN(new_n1065_));
  AOI22_X1   g0423(.A1(\in2[41] ), .A2(\in3[42] ), .B1(\in2[42] ), .B2(\in3[41] ), .ZN(new_n1066_));
  INV_X1     g0424(.I(\in2[40] ), .ZN(new_n1067_));
  INV_X1     g0425(.I(\in3[40] ), .ZN(new_n1068_));
  NAND2_X1   g0426(.A1(new_n1067_), .A2(new_n1068_), .ZN(new_n1069_));
  INV_X1     g0427(.I(\in2[41] ), .ZN(new_n1070_));
  INV_X1     g0428(.I(\in3[41] ), .ZN(new_n1071_));
  NOR2_X1    g0429(.A1(new_n1070_), .A2(new_n1071_), .ZN(new_n1072_));
  AOI21_X1   g0430(.A1(new_n1072_), .A2(new_n1069_), .B(new_n1066_), .ZN(new_n1073_));
  AOI22_X1   g0431(.A1(\in2[46] ), .A2(\in3[47] ), .B1(\in2[47] ), .B2(\in3[46] ), .ZN(new_n1074_));
  AOI22_X1   g0432(.A1(\in2[44] ), .A2(\in3[45] ), .B1(\in2[45] ), .B2(\in3[44] ), .ZN(new_n1075_));
  AOI22_X1   g0433(.A1(\in2[42] ), .A2(\in3[43] ), .B1(\in2[43] ), .B2(\in3[42] ), .ZN(new_n1076_));
  NOR3_X1    g0434(.A1(new_n1074_), .A2(new_n1075_), .A3(new_n1076_), .ZN(new_n1077_));
  INV_X1     g0435(.I(new_n1077_), .ZN(new_n1078_));
  OAI21_X1   g0436(.A1(new_n1078_), .A2(new_n1073_), .B(new_n1065_), .ZN(new_n1079_));
  NAND2_X1   g0437(.A1(\in2[47] ), .A2(\in3[47] ), .ZN(new_n1080_));
  NOR2_X1    g0438(.A1(\in2[47] ), .A2(\in3[47] ), .ZN(new_n1081_));
  NAND2_X1   g0439(.A1(\in2[46] ), .A2(\in3[46] ), .ZN(new_n1082_));
  OAI21_X1   g0440(.A1(new_n1081_), .A2(new_n1082_), .B(new_n1080_), .ZN(new_n1083_));
  AOI21_X1   g0441(.A1(new_n1079_), .A2(\in3[43] ), .B(new_n1083_), .ZN(new_n1084_));
  INV_X1     g0442(.I(new_n1074_), .ZN(new_n1085_));
  NAND2_X1   g0443(.A1(\in2[45] ), .A2(\in3[45] ), .ZN(new_n1086_));
  NOR2_X1    g0444(.A1(\in2[45] ), .A2(\in3[45] ), .ZN(new_n1087_));
  NAND2_X1   g0445(.A1(\in2[44] ), .A2(\in3[44] ), .ZN(new_n1088_));
  OAI21_X1   g0446(.A1(new_n1087_), .A2(new_n1088_), .B(new_n1086_), .ZN(new_n1089_));
  OAI22_X1   g0447(.A1(new_n1067_), .A2(new_n1071_), .B1(new_n1070_), .B2(new_n1068_), .ZN(new_n1090_));
  NAND4_X1   g0448(.A1(new_n1077_), .A2(new_n1085_), .A3(new_n1089_), .A4(new_n1090_), .ZN(new_n1091_));
  OAI22_X1   g0449(.A1(new_n1058_), .A2(new_n1064_), .B1(new_n1084_), .B2(new_n1091_), .ZN(new_n1092_));
  INV_X1     g0450(.I(\in3[53] ), .ZN(new_n1093_));
  NOR2_X1    g0451(.A1(new_n1093_), .A2(\in2[53] ), .ZN(new_n1094_));
  INV_X1     g0452(.I(new_n1094_), .ZN(new_n1095_));
  AOI22_X1   g0453(.A1(\in2[54] ), .A2(\in3[55] ), .B1(\in2[55] ), .B2(\in3[54] ), .ZN(new_n1096_));
  NAND2_X1   g0454(.A1(\in2[52] ), .A2(\in3[52] ), .ZN(new_n1097_));
  AOI21_X1   g0455(.A1(new_n1095_), .A2(new_n1096_), .B(new_n1097_), .ZN(new_n1098_));
  INV_X1     g0456(.I(new_n1098_), .ZN(new_n1099_));
  INV_X1     g0457(.I(\in2[48] ), .ZN(new_n1100_));
  INV_X1     g0458(.I(\in2[49] ), .ZN(new_n1101_));
  INV_X1     g0459(.I(\in3[48] ), .ZN(new_n1102_));
  INV_X1     g0460(.I(\in3[49] ), .ZN(new_n1103_));
  OAI22_X1   g0461(.A1(new_n1100_), .A2(new_n1103_), .B1(new_n1101_), .B2(new_n1102_), .ZN(new_n1104_));
  INV_X1     g0462(.I(\in2[50] ), .ZN(new_n1105_));
  INV_X1     g0463(.I(\in2[51] ), .ZN(new_n1106_));
  INV_X1     g0464(.I(\in3[50] ), .ZN(new_n1107_));
  INV_X1     g0465(.I(\in3[51] ), .ZN(new_n1108_));
  OAI22_X1   g0466(.A1(new_n1105_), .A2(new_n1108_), .B1(new_n1106_), .B2(new_n1107_), .ZN(new_n1109_));
  NAND2_X1   g0467(.A1(new_n1104_), .A2(new_n1109_), .ZN(new_n1110_));
  AOI22_X1   g0468(.A1(\in2[49] ), .A2(\in3[50] ), .B1(\in2[50] ), .B2(\in3[49] ), .ZN(new_n1111_));
  NOR2_X1    g0469(.A1(\in2[48] ), .A2(\in3[48] ), .ZN(new_n1112_));
  NOR3_X1    g0470(.A1(new_n1112_), .A2(new_n1101_), .A3(new_n1103_), .ZN(new_n1113_));
  OAI21_X1   g0471(.A1(new_n1111_), .A2(new_n1113_), .B(new_n1109_), .ZN(new_n1114_));
  OAI21_X1   g0472(.A1(new_n1099_), .A2(new_n1114_), .B(new_n1106_), .ZN(new_n1115_));
  NAND2_X1   g0473(.A1(\in2[53] ), .A2(\in3[54] ), .ZN(new_n1116_));
  NAND2_X1   g0474(.A1(\in2[54] ), .A2(\in3[53] ), .ZN(new_n1117_));
  NAND2_X1   g0475(.A1(new_n1116_), .A2(new_n1117_), .ZN(new_n1118_));
  INV_X1     g0476(.I(\in3[52] ), .ZN(new_n1119_));
  NAND3_X1   g0477(.A1(new_n1095_), .A2(\in2[52] ), .A3(new_n1119_), .ZN(new_n1120_));
  AOI21_X1   g0478(.A1(new_n1120_), .A2(new_n1118_), .B(new_n1096_), .ZN(new_n1121_));
  AOI21_X1   g0479(.A1(new_n1115_), .A2(\in3[51] ), .B(new_n1121_), .ZN(new_n1122_));
  AOI22_X1   g0480(.A1(\in2[56] ), .A2(\in3[57] ), .B1(\in2[57] ), .B2(\in3[56] ), .ZN(new_n1123_));
  NAND2_X1   g0481(.A1(\in2[55] ), .A2(\in3[55] ), .ZN(new_n1124_));
  NOR2_X1    g0482(.A1(new_n1123_), .A2(new_n1124_), .ZN(new_n1125_));
  NAND4_X1   g0483(.A1(new_n1125_), .A2(new_n1020_), .A3(new_n1013_), .A4(new_n1016_), .ZN(new_n1126_));
  OAI22_X1   g0484(.A1(new_n1122_), .A2(new_n1126_), .B1(new_n1099_), .B2(new_n1110_), .ZN(new_n1127_));
  NAND4_X1   g0485(.A1(new_n1005_), .A2(new_n1047_), .A3(new_n1092_), .A4(new_n1127_), .ZN(new_n1128_));
  AOI21_X1   g0486(.A1(new_n767_), .A2(new_n648_), .B(new_n1128_), .ZN(new_n1129_));
  NAND4_X1   g0487(.A1(new_n1129_), .A2(\in2[0] ), .A3(\in3[0] ), .A4(new_n644_), .ZN(new_n1130_));
  INV_X1     g0488(.I(\in2[0] ), .ZN(new_n1131_));
  NAND4_X1   g0489(.A1(new_n1129_), .A2(new_n1131_), .A3(new_n695_), .A4(new_n644_), .ZN(new_n1132_));
  NAND2_X1   g0490(.A1(new_n1130_), .A2(new_n1132_), .ZN(new_n1133_));
  INV_X1     g0491(.I(\in0[127] ), .ZN(new_n1134_));
  INV_X1     g0492(.I(\in1[127] ), .ZN(new_n1135_));
  INV_X1     g0493(.I(\in0[29] ), .ZN(new_n1136_));
  INV_X1     g0494(.I(\in0[30] ), .ZN(new_n1137_));
  NOR3_X1    g0495(.A1(new_n1136_), .A2(new_n1137_), .A3(\in1[29] ), .ZN(new_n1138_));
  INV_X1     g0496(.I(new_n1138_), .ZN(new_n1139_));
  INV_X1     g0497(.I(\in0[26] ), .ZN(new_n1140_));
  INV_X1     g0498(.I(\in0[27] ), .ZN(new_n1141_));
  NOR3_X1    g0499(.A1(new_n1140_), .A2(new_n1141_), .A3(\in1[26] ), .ZN(new_n1142_));
  INV_X1     g0500(.I(\in1[24] ), .ZN(new_n1143_));
  NOR2_X1    g0501(.A1(new_n1143_), .A2(\in0[24] ), .ZN(new_n1144_));
  INV_X1     g0502(.I(new_n1144_), .ZN(new_n1145_));
  INV_X1     g0503(.I(\in0[23] ), .ZN(new_n1146_));
  NAND2_X1   g0504(.A1(new_n1146_), .A2(\in1[23] ), .ZN(new_n1147_));
  INV_X1     g0505(.I(new_n1147_), .ZN(new_n1148_));
  INV_X1     g0506(.I(\in0[21] ), .ZN(new_n1149_));
  INV_X1     g0507(.I(\in0[22] ), .ZN(new_n1150_));
  NOR3_X1    g0508(.A1(new_n1149_), .A2(new_n1150_), .A3(\in1[21] ), .ZN(new_n1151_));
  INV_X1     g0509(.I(new_n1151_), .ZN(new_n1152_));
  INV_X1     g0510(.I(\in0[18] ), .ZN(new_n1153_));
  INV_X1     g0511(.I(\in0[19] ), .ZN(new_n1154_));
  NOR3_X1    g0512(.A1(new_n1153_), .A2(new_n1154_), .A3(\in1[18] ), .ZN(new_n1155_));
  INV_X1     g0513(.I(\in1[16] ), .ZN(new_n1156_));
  NOR2_X1    g0514(.A1(new_n1156_), .A2(\in0[16] ), .ZN(new_n1157_));
  INV_X1     g0515(.I(new_n1157_), .ZN(new_n1158_));
  INV_X1     g0516(.I(\in0[15] ), .ZN(new_n1159_));
  NAND2_X1   g0517(.A1(new_n1159_), .A2(\in1[15] ), .ZN(new_n1160_));
  INV_X1     g0518(.I(new_n1160_), .ZN(new_n1161_));
  INV_X1     g0519(.I(\in0[13] ), .ZN(new_n1162_));
  INV_X1     g0520(.I(\in0[14] ), .ZN(new_n1163_));
  NOR3_X1    g0521(.A1(new_n1162_), .A2(new_n1163_), .A3(\in1[13] ), .ZN(new_n1164_));
  INV_X1     g0522(.I(new_n1164_), .ZN(new_n1165_));
  INV_X1     g0523(.I(\in0[10] ), .ZN(new_n1166_));
  INV_X1     g0524(.I(\in0[11] ), .ZN(new_n1167_));
  NOR3_X1    g0525(.A1(new_n1166_), .A2(new_n1167_), .A3(\in1[10] ), .ZN(new_n1168_));
  INV_X1     g0526(.I(\in1[8] ), .ZN(new_n1169_));
  NOR2_X1    g0527(.A1(new_n1169_), .A2(\in0[8] ), .ZN(new_n1170_));
  INV_X1     g0528(.I(new_n1170_), .ZN(new_n1171_));
  INV_X1     g0529(.I(\in0[6] ), .ZN(new_n1172_));
  INV_X1     g0530(.I(\in0[7] ), .ZN(new_n1173_));
  NOR3_X1    g0531(.A1(new_n1172_), .A2(new_n1173_), .A3(\in1[6] ), .ZN(new_n1174_));
  INV_X1     g0532(.I(\in1[4] ), .ZN(new_n1175_));
  NOR2_X1    g0533(.A1(new_n1175_), .A2(\in0[4] ), .ZN(new_n1176_));
  INV_X1     g0534(.I(new_n1176_), .ZN(new_n1177_));
  INV_X1     g0535(.I(\in0[3] ), .ZN(new_n1178_));
  NAND2_X1   g0536(.A1(new_n1178_), .A2(\in1[3] ), .ZN(new_n1179_));
  INV_X1     g0537(.I(\in0[2] ), .ZN(new_n1180_));
  INV_X1     g0538(.I(\in1[2] ), .ZN(new_n1181_));
  NOR2_X1    g0539(.A1(new_n1180_), .A2(new_n1181_), .ZN(new_n1182_));
  INV_X1     g0540(.I(\in1[1] ), .ZN(new_n1183_));
  AOI22_X1   g0541(.A1(\in0[0] ), .A2(\in1[1] ), .B1(\in0[1] ), .B2(\in1[0] ), .ZN(new_n1184_));
  NOR2_X1    g0542(.A1(\in0[2] ), .A2(\in1[2] ), .ZN(new_n1185_));
  NOR4_X1    g0543(.A1(new_n1184_), .A2(\in0[1] ), .A3(new_n1183_), .A4(new_n1185_), .ZN(new_n1186_));
  OAI22_X1   g0544(.A1(new_n1186_), .A2(new_n1182_), .B1(new_n1178_), .B2(\in1[3] ), .ZN(new_n1187_));
  NAND2_X1   g0545(.A1(new_n1187_), .A2(new_n1179_), .ZN(new_n1188_));
  NAND2_X1   g0546(.A1(new_n1175_), .A2(\in0[4] ), .ZN(new_n1189_));
  NAND2_X1   g0547(.A1(new_n1188_), .A2(new_n1189_), .ZN(new_n1190_));
  INV_X1     g0548(.I(\in1[6] ), .ZN(new_n1191_));
  NOR2_X1    g0549(.A1(new_n1191_), .A2(\in0[6] ), .ZN(new_n1192_));
  AOI21_X1   g0550(.A1(new_n1192_), .A2(\in0[5] ), .B(\in1[5] ), .ZN(new_n1193_));
  AOI21_X1   g0551(.A1(new_n1191_), .A2(\in0[6] ), .B(\in0[7] ), .ZN(new_n1194_));
  OAI21_X1   g0552(.A1(new_n1192_), .A2(\in0[5] ), .B(\in1[7] ), .ZN(new_n1195_));
  NOR3_X1    g0553(.A1(new_n1193_), .A2(new_n1195_), .A3(new_n1194_), .ZN(new_n1196_));
  INV_X1     g0554(.I(new_n1196_), .ZN(new_n1197_));
  AOI21_X1   g0555(.A1(new_n1190_), .A2(new_n1177_), .B(new_n1197_), .ZN(new_n1198_));
  NAND2_X1   g0556(.A1(new_n1169_), .A2(\in0[8] ), .ZN(new_n1199_));
  OAI21_X1   g0557(.A1(new_n1198_), .A2(new_n1174_), .B(new_n1199_), .ZN(new_n1200_));
  INV_X1     g0558(.I(\in1[10] ), .ZN(new_n1201_));
  NOR2_X1    g0559(.A1(new_n1201_), .A2(\in0[10] ), .ZN(new_n1202_));
  AOI21_X1   g0560(.A1(new_n1202_), .A2(\in0[9] ), .B(\in1[9] ), .ZN(new_n1203_));
  AOI21_X1   g0561(.A1(new_n1201_), .A2(\in0[10] ), .B(\in0[11] ), .ZN(new_n1204_));
  OAI21_X1   g0562(.A1(new_n1202_), .A2(\in0[9] ), .B(\in1[11] ), .ZN(new_n1205_));
  NOR3_X1    g0563(.A1(new_n1203_), .A2(new_n1205_), .A3(new_n1204_), .ZN(new_n1206_));
  INV_X1     g0564(.I(new_n1206_), .ZN(new_n1207_));
  AOI21_X1   g0565(.A1(new_n1200_), .A2(new_n1171_), .B(new_n1207_), .ZN(new_n1208_));
  INV_X1     g0566(.I(\in1[13] ), .ZN(new_n1209_));
  NOR2_X1    g0567(.A1(new_n1209_), .A2(\in0[13] ), .ZN(new_n1210_));
  AOI21_X1   g0568(.A1(new_n1210_), .A2(\in0[12] ), .B(\in1[12] ), .ZN(new_n1211_));
  AOI21_X1   g0569(.A1(new_n1209_), .A2(\in0[13] ), .B(\in0[14] ), .ZN(new_n1212_));
  OAI21_X1   g0570(.A1(new_n1210_), .A2(\in0[12] ), .B(\in1[14] ), .ZN(new_n1213_));
  NOR3_X1    g0571(.A1(new_n1211_), .A2(new_n1213_), .A3(new_n1212_), .ZN(new_n1214_));
  OAI21_X1   g0572(.A1(new_n1208_), .A2(new_n1168_), .B(new_n1214_), .ZN(new_n1215_));
  NOR2_X1    g0573(.A1(new_n1159_), .A2(\in1[15] ), .ZN(new_n1216_));
  AOI21_X1   g0574(.A1(new_n1215_), .A2(new_n1165_), .B(new_n1216_), .ZN(new_n1217_));
  INV_X1     g0575(.I(\in0[16] ), .ZN(new_n1218_));
  NOR2_X1    g0576(.A1(new_n1218_), .A2(\in1[16] ), .ZN(new_n1219_));
  INV_X1     g0577(.I(new_n1219_), .ZN(new_n1220_));
  OAI21_X1   g0578(.A1(new_n1217_), .A2(new_n1161_), .B(new_n1220_), .ZN(new_n1221_));
  INV_X1     g0579(.I(\in1[18] ), .ZN(new_n1222_));
  NOR2_X1    g0580(.A1(new_n1222_), .A2(\in0[18] ), .ZN(new_n1223_));
  AOI21_X1   g0581(.A1(new_n1223_), .A2(\in0[17] ), .B(\in1[17] ), .ZN(new_n1224_));
  AOI21_X1   g0582(.A1(new_n1222_), .A2(\in0[18] ), .B(\in0[19] ), .ZN(new_n1225_));
  OAI21_X1   g0583(.A1(new_n1223_), .A2(\in0[17] ), .B(\in1[19] ), .ZN(new_n1226_));
  NOR3_X1    g0584(.A1(new_n1224_), .A2(new_n1226_), .A3(new_n1225_), .ZN(new_n1227_));
  INV_X1     g0585(.I(new_n1227_), .ZN(new_n1228_));
  AOI21_X1   g0586(.A1(new_n1221_), .A2(new_n1158_), .B(new_n1228_), .ZN(new_n1229_));
  INV_X1     g0587(.I(\in1[21] ), .ZN(new_n1230_));
  NOR2_X1    g0588(.A1(new_n1230_), .A2(\in0[21] ), .ZN(new_n1231_));
  AOI21_X1   g0589(.A1(new_n1231_), .A2(\in0[20] ), .B(\in1[20] ), .ZN(new_n1232_));
  AOI21_X1   g0590(.A1(new_n1230_), .A2(\in0[21] ), .B(\in0[22] ), .ZN(new_n1233_));
  OAI21_X1   g0591(.A1(new_n1231_), .A2(\in0[20] ), .B(\in1[22] ), .ZN(new_n1234_));
  NOR3_X1    g0592(.A1(new_n1232_), .A2(new_n1234_), .A3(new_n1233_), .ZN(new_n1235_));
  OAI21_X1   g0593(.A1(new_n1229_), .A2(new_n1155_), .B(new_n1235_), .ZN(new_n1236_));
  NOR2_X1    g0594(.A1(new_n1146_), .A2(\in1[23] ), .ZN(new_n1237_));
  AOI21_X1   g0595(.A1(new_n1236_), .A2(new_n1152_), .B(new_n1237_), .ZN(new_n1238_));
  INV_X1     g0596(.I(\in0[24] ), .ZN(new_n1239_));
  NOR2_X1    g0597(.A1(new_n1239_), .A2(\in1[24] ), .ZN(new_n1240_));
  INV_X1     g0598(.I(new_n1240_), .ZN(new_n1241_));
  OAI21_X1   g0599(.A1(new_n1238_), .A2(new_n1148_), .B(new_n1241_), .ZN(new_n1242_));
  INV_X1     g0600(.I(\in1[26] ), .ZN(new_n1243_));
  NOR2_X1    g0601(.A1(new_n1243_), .A2(\in0[26] ), .ZN(new_n1244_));
  AOI21_X1   g0602(.A1(new_n1244_), .A2(\in0[25] ), .B(\in1[25] ), .ZN(new_n1245_));
  AOI21_X1   g0603(.A1(new_n1243_), .A2(\in0[26] ), .B(\in0[27] ), .ZN(new_n1246_));
  OAI21_X1   g0604(.A1(new_n1244_), .A2(\in0[25] ), .B(\in1[27] ), .ZN(new_n1247_));
  NOR3_X1    g0605(.A1(new_n1245_), .A2(new_n1247_), .A3(new_n1246_), .ZN(new_n1248_));
  INV_X1     g0606(.I(new_n1248_), .ZN(new_n1249_));
  AOI21_X1   g0607(.A1(new_n1242_), .A2(new_n1145_), .B(new_n1249_), .ZN(new_n1250_));
  INV_X1     g0608(.I(\in1[29] ), .ZN(new_n1251_));
  NOR2_X1    g0609(.A1(new_n1251_), .A2(\in0[29] ), .ZN(new_n1252_));
  AOI21_X1   g0610(.A1(new_n1252_), .A2(\in0[28] ), .B(\in1[28] ), .ZN(new_n1253_));
  AOI21_X1   g0611(.A1(new_n1251_), .A2(\in0[29] ), .B(\in0[30] ), .ZN(new_n1254_));
  OAI21_X1   g0612(.A1(new_n1252_), .A2(\in0[28] ), .B(\in1[30] ), .ZN(new_n1255_));
  NOR3_X1    g0613(.A1(new_n1253_), .A2(new_n1255_), .A3(new_n1254_), .ZN(new_n1256_));
  OAI21_X1   g0614(.A1(new_n1250_), .A2(new_n1142_), .B(new_n1256_), .ZN(new_n1257_));
  AOI22_X1   g0615(.A1(\in0[94] ), .A2(\in1[95] ), .B1(\in0[95] ), .B2(\in1[94] ), .ZN(new_n1258_));
  AOI22_X1   g0616(.A1(\in0[92] ), .A2(\in1[93] ), .B1(\in0[93] ), .B2(\in1[92] ), .ZN(new_n1259_));
  INV_X1     g0617(.I(\in0[93] ), .ZN(new_n1260_));
  INV_X1     g0618(.I(\in1[93] ), .ZN(new_n1261_));
  NAND2_X1   g0619(.A1(\in0[92] ), .A2(\in1[92] ), .ZN(new_n1262_));
  AOI21_X1   g0620(.A1(new_n1260_), .A2(new_n1261_), .B(new_n1262_), .ZN(new_n1263_));
  NOR2_X1    g0621(.A1(new_n1260_), .A2(new_n1261_), .ZN(new_n1264_));
  NOR3_X1    g0622(.A1(new_n1263_), .A2(new_n1258_), .A3(new_n1264_), .ZN(new_n1265_));
  INV_X1     g0623(.I(\in1[97] ), .ZN(new_n1266_));
  AOI22_X1   g0624(.A1(\in0[98] ), .A2(\in1[99] ), .B1(\in0[99] ), .B2(\in1[98] ), .ZN(new_n1267_));
  OAI21_X1   g0625(.A1(\in0[97] ), .A2(new_n1266_), .B(new_n1267_), .ZN(new_n1268_));
  NAND2_X1   g0626(.A1(\in0[95] ), .A2(\in1[95] ), .ZN(new_n1269_));
  NOR2_X1    g0627(.A1(\in0[95] ), .A2(\in1[95] ), .ZN(new_n1270_));
  NAND2_X1   g0628(.A1(\in0[94] ), .A2(\in1[94] ), .ZN(new_n1271_));
  OAI21_X1   g0629(.A1(new_n1270_), .A2(new_n1271_), .B(new_n1269_), .ZN(new_n1272_));
  NAND4_X1   g0630(.A1(new_n1268_), .A2(\in0[96] ), .A3(\in1[96] ), .A4(new_n1272_), .ZN(new_n1273_));
  OAI22_X1   g0631(.A1(new_n1273_), .A2(new_n1265_), .B1(new_n1258_), .B2(new_n1259_), .ZN(new_n1274_));
  INV_X1     g0632(.I(\in0[105] ), .ZN(new_n1275_));
  NAND2_X1   g0633(.A1(\in0[107] ), .A2(\in1[106] ), .ZN(new_n1276_));
  NAND2_X1   g0634(.A1(\in0[106] ), .A2(\in1[107] ), .ZN(new_n1277_));
  NAND2_X1   g0635(.A1(new_n1276_), .A2(new_n1277_), .ZN(new_n1278_));
  AOI21_X1   g0636(.A1(new_n1275_), .A2(\in1[105] ), .B(new_n1278_), .ZN(new_n1279_));
  NAND2_X1   g0637(.A1(\in0[104] ), .A2(\in1[104] ), .ZN(new_n1280_));
  INV_X1     g0638(.I(\in0[104] ), .ZN(new_n1281_));
  INV_X1     g0639(.I(\in1[104] ), .ZN(new_n1282_));
  NAND2_X1   g0640(.A1(\in0[106] ), .A2(\in1[105] ), .ZN(new_n1283_));
  NAND2_X1   g0641(.A1(\in0[105] ), .A2(\in1[106] ), .ZN(new_n1284_));
  NAND4_X1   g0642(.A1(new_n1283_), .A2(new_n1284_), .A3(new_n1281_), .A4(new_n1282_), .ZN(new_n1285_));
  AND3_X2    g0643(.A1(new_n1275_), .A2(\in0[107] ), .A3(\in1[105] ), .Z(new_n1286_));
  AOI22_X1   g0644(.A1(new_n1286_), .A2(new_n1285_), .B1(\in1[107] ), .B2(new_n1278_), .ZN(new_n1287_));
  AOI22_X1   g0645(.A1(\in0[110] ), .A2(\in1[111] ), .B1(\in0[111] ), .B2(\in1[110] ), .ZN(new_n1288_));
  AOI22_X1   g0646(.A1(\in0[108] ), .A2(\in1[109] ), .B1(\in0[109] ), .B2(\in1[108] ), .ZN(new_n1289_));
  OR2_X2     g0647(.A1(new_n1288_), .A2(new_n1289_), .Z(new_n1290_));
  OAI22_X1   g0648(.A1(new_n1287_), .A2(new_n1290_), .B1(new_n1279_), .B2(new_n1280_), .ZN(new_n1291_));
  INV_X1     g0649(.I(\in0[111] ), .ZN(new_n1292_));
  INV_X1     g0650(.I(\in1[111] ), .ZN(new_n1293_));
  NOR2_X1    g0651(.A1(new_n1292_), .A2(new_n1293_), .ZN(new_n1294_));
  NAND2_X1   g0652(.A1(new_n1292_), .A2(new_n1293_), .ZN(new_n1295_));
  AND2_X2    g0653(.A1(\in0[110] ), .A2(\in1[110] ), .Z(new_n1296_));
  AOI21_X1   g0654(.A1(new_n1295_), .A2(new_n1296_), .B(new_n1294_), .ZN(new_n1297_));
  INV_X1     g0655(.I(\in0[109] ), .ZN(new_n1298_));
  INV_X1     g0656(.I(\in1[109] ), .ZN(new_n1299_));
  NAND2_X1   g0657(.A1(\in0[108] ), .A2(\in1[108] ), .ZN(new_n1300_));
  AOI21_X1   g0658(.A1(new_n1298_), .A2(new_n1299_), .B(new_n1300_), .ZN(new_n1301_));
  NOR2_X1    g0659(.A1(new_n1298_), .A2(new_n1299_), .ZN(new_n1302_));
  NOR3_X1    g0660(.A1(new_n1301_), .A2(new_n1288_), .A3(new_n1302_), .ZN(new_n1303_));
  NAND2_X1   g0661(.A1(\in0[115] ), .A2(\in1[114] ), .ZN(new_n1304_));
  NAND2_X1   g0662(.A1(\in0[114] ), .A2(\in1[115] ), .ZN(new_n1305_));
  NAND2_X1   g0663(.A1(new_n1304_), .A2(new_n1305_), .ZN(new_n1306_));
  INV_X1     g0664(.I(\in0[112] ), .ZN(new_n1307_));
  INV_X1     g0665(.I(\in1[112] ), .ZN(new_n1308_));
  NAND2_X1   g0666(.A1(\in0[114] ), .A2(\in1[113] ), .ZN(new_n1309_));
  NAND2_X1   g0667(.A1(\in0[113] ), .A2(\in1[114] ), .ZN(new_n1310_));
  NAND4_X1   g0668(.A1(new_n1309_), .A2(new_n1310_), .A3(new_n1307_), .A4(new_n1308_), .ZN(new_n1311_));
  INV_X1     g0669(.I(\in0[115] ), .ZN(new_n1312_));
  INV_X1     g0670(.I(\in1[113] ), .ZN(new_n1313_));
  NOR3_X1    g0671(.A1(new_n1312_), .A2(new_n1313_), .A3(\in0[113] ), .ZN(new_n1314_));
  AOI22_X1   g0672(.A1(new_n1311_), .A2(new_n1314_), .B1(new_n1306_), .B2(\in1[115] ), .ZN(new_n1315_));
  NOR2_X1    g0673(.A1(new_n1313_), .A2(\in0[113] ), .ZN(new_n1316_));
  NOR2_X1    g0674(.A1(new_n1307_), .A2(new_n1308_), .ZN(new_n1317_));
  OAI21_X1   g0675(.A1(new_n1306_), .A2(new_n1316_), .B(new_n1317_), .ZN(new_n1318_));
  OAI22_X1   g0676(.A1(new_n1315_), .A2(new_n1318_), .B1(new_n1303_), .B2(new_n1297_), .ZN(new_n1319_));
  AOI22_X1   g0677(.A1(\in0[118] ), .A2(\in1[119] ), .B1(\in0[119] ), .B2(\in1[118] ), .ZN(new_n1320_));
  AOI22_X1   g0678(.A1(\in0[116] ), .A2(\in1[117] ), .B1(\in0[117] ), .B2(\in1[116] ), .ZN(new_n1321_));
  INV_X1     g0679(.I(\in0[117] ), .ZN(new_n1322_));
  INV_X1     g0680(.I(\in1[117] ), .ZN(new_n1323_));
  NAND2_X1   g0681(.A1(\in0[116] ), .A2(\in1[116] ), .ZN(new_n1324_));
  AOI21_X1   g0682(.A1(new_n1322_), .A2(new_n1323_), .B(new_n1324_), .ZN(new_n1325_));
  NOR2_X1    g0683(.A1(new_n1322_), .A2(new_n1323_), .ZN(new_n1326_));
  NOR3_X1    g0684(.A1(new_n1325_), .A2(new_n1320_), .A3(new_n1326_), .ZN(new_n1327_));
  INV_X1     g0685(.I(\in1[121] ), .ZN(new_n1328_));
  AOI22_X1   g0686(.A1(\in0[122] ), .A2(\in1[123] ), .B1(\in0[123] ), .B2(\in1[122] ), .ZN(new_n1329_));
  OAI21_X1   g0687(.A1(\in0[121] ), .A2(new_n1328_), .B(new_n1329_), .ZN(new_n1330_));
  NAND2_X1   g0688(.A1(\in0[119] ), .A2(\in1[119] ), .ZN(new_n1331_));
  NOR2_X1    g0689(.A1(\in0[119] ), .A2(\in1[119] ), .ZN(new_n1332_));
  NAND2_X1   g0690(.A1(\in0[118] ), .A2(\in1[118] ), .ZN(new_n1333_));
  OAI21_X1   g0691(.A1(new_n1332_), .A2(new_n1333_), .B(new_n1331_), .ZN(new_n1334_));
  NAND4_X1   g0692(.A1(new_n1330_), .A2(\in0[120] ), .A3(\in1[120] ), .A4(new_n1334_), .ZN(new_n1335_));
  OAI22_X1   g0693(.A1(new_n1335_), .A2(new_n1327_), .B1(new_n1320_), .B2(new_n1321_), .ZN(new_n1336_));
  NAND4_X1   g0694(.A1(new_n1274_), .A2(new_n1336_), .A3(new_n1291_), .A4(new_n1319_), .ZN(new_n1337_));
  AOI22_X1   g0695(.A1(\in0[124] ), .A2(\in0[127] ), .B1(\in1[124] ), .B2(\in1[127] ), .ZN(new_n1338_));
  AOI22_X1   g0696(.A1(\in0[125] ), .A2(\in1[126] ), .B1(\in0[126] ), .B2(\in1[125] ), .ZN(new_n1339_));
  NOR2_X1    g0697(.A1(new_n1134_), .A2(\in1[127] ), .ZN(new_n1340_));
  OR3_X2     g0698(.A1(new_n1338_), .A2(new_n1339_), .A3(new_n1340_), .Z(new_n1341_));
  INV_X1     g0699(.I(\in0[126] ), .ZN(new_n1342_));
  INV_X1     g0700(.I(\in1[126] ), .ZN(new_n1343_));
  AOI22_X1   g0701(.A1(\in0[124] ), .A2(\in1[125] ), .B1(\in0[125] ), .B2(\in1[124] ), .ZN(new_n1344_));
  OAI22_X1   g0702(.A1(new_n1342_), .A2(new_n1344_), .B1(new_n1339_), .B2(new_n1343_), .ZN(new_n1345_));
  INV_X1     g0703(.I(new_n1329_), .ZN(new_n1346_));
  INV_X1     g0704(.I(\in0[120] ), .ZN(new_n1347_));
  INV_X1     g0705(.I(\in1[120] ), .ZN(new_n1348_));
  NAND2_X1   g0706(.A1(\in0[122] ), .A2(\in1[121] ), .ZN(new_n1349_));
  NAND2_X1   g0707(.A1(\in0[121] ), .A2(\in1[122] ), .ZN(new_n1350_));
  NAND4_X1   g0708(.A1(new_n1349_), .A2(new_n1350_), .A3(new_n1347_), .A4(new_n1348_), .ZN(new_n1351_));
  INV_X1     g0709(.I(\in0[123] ), .ZN(new_n1352_));
  NOR3_X1    g0710(.A1(new_n1352_), .A2(new_n1328_), .A3(\in0[121] ), .ZN(new_n1353_));
  AOI22_X1   g0711(.A1(new_n1351_), .A2(new_n1353_), .B1(new_n1346_), .B2(\in1[123] ), .ZN(new_n1354_));
  OAI21_X1   g0712(.A1(new_n1341_), .A2(new_n1345_), .B(new_n1354_), .ZN(new_n1355_));
  INV_X1     g0713(.I(\in0[77] ), .ZN(new_n1356_));
  INV_X1     g0714(.I(\in1[77] ), .ZN(new_n1357_));
  NAND2_X1   g0715(.A1(\in0[76] ), .A2(\in1[76] ), .ZN(new_n1358_));
  AOI21_X1   g0716(.A1(new_n1356_), .A2(new_n1357_), .B(new_n1358_), .ZN(new_n1359_));
  AOI22_X1   g0717(.A1(\in0[78] ), .A2(\in1[79] ), .B1(\in0[79] ), .B2(\in1[78] ), .ZN(new_n1360_));
  NOR2_X1    g0718(.A1(new_n1356_), .A2(new_n1357_), .ZN(new_n1361_));
  NOR3_X1    g0719(.A1(new_n1359_), .A2(new_n1360_), .A3(new_n1361_), .ZN(new_n1362_));
  NOR2_X1    g0720(.A1(\in0[79] ), .A2(\in1[79] ), .ZN(new_n1363_));
  NAND2_X1   g0721(.A1(\in0[78] ), .A2(\in1[78] ), .ZN(new_n1364_));
  NOR2_X1    g0722(.A1(new_n1363_), .A2(new_n1364_), .ZN(new_n1365_));
  AOI21_X1   g0723(.A1(\in0[79] ), .A2(\in1[79] ), .B(new_n1365_), .ZN(new_n1366_));
  AOI22_X1   g0724(.A1(\in0[76] ), .A2(\in1[77] ), .B1(\in0[77] ), .B2(\in1[76] ), .ZN(new_n1367_));
  OR3_X2     g0725(.A1(new_n1366_), .A2(new_n1360_), .A3(new_n1367_), .Z(new_n1368_));
  AOI22_X1   g0726(.A1(\in0[74] ), .A2(\in1[75] ), .B1(\in0[75] ), .B2(\in1[74] ), .ZN(new_n1369_));
  INV_X1     g0727(.I(new_n1369_), .ZN(new_n1370_));
  INV_X1     g0728(.I(\in0[72] ), .ZN(new_n1371_));
  INV_X1     g0729(.I(\in1[72] ), .ZN(new_n1372_));
  NAND2_X1   g0730(.A1(\in0[74] ), .A2(\in1[73] ), .ZN(new_n1373_));
  NAND2_X1   g0731(.A1(\in0[73] ), .A2(\in1[74] ), .ZN(new_n1374_));
  NAND4_X1   g0732(.A1(new_n1373_), .A2(new_n1374_), .A3(new_n1371_), .A4(new_n1372_), .ZN(new_n1375_));
  INV_X1     g0733(.I(\in0[75] ), .ZN(new_n1376_));
  INV_X1     g0734(.I(\in1[73] ), .ZN(new_n1377_));
  NOR3_X1    g0735(.A1(new_n1376_), .A2(new_n1377_), .A3(\in0[73] ), .ZN(new_n1378_));
  AOI22_X1   g0736(.A1(new_n1375_), .A2(new_n1378_), .B1(new_n1370_), .B2(\in1[75] ), .ZN(new_n1379_));
  OAI21_X1   g0737(.A1(new_n1368_), .A2(new_n1362_), .B(new_n1379_), .ZN(new_n1380_));
  INV_X1     g0738(.I(\in0[101] ), .ZN(new_n1381_));
  INV_X1     g0739(.I(\in1[101] ), .ZN(new_n1382_));
  NAND2_X1   g0740(.A1(\in0[100] ), .A2(\in1[100] ), .ZN(new_n1383_));
  AOI21_X1   g0741(.A1(new_n1381_), .A2(new_n1382_), .B(new_n1383_), .ZN(new_n1384_));
  AOI22_X1   g0742(.A1(\in0[102] ), .A2(\in1[103] ), .B1(\in0[103] ), .B2(\in1[102] ), .ZN(new_n1385_));
  NOR2_X1    g0743(.A1(new_n1381_), .A2(new_n1382_), .ZN(new_n1386_));
  NOR3_X1    g0744(.A1(new_n1384_), .A2(new_n1385_), .A3(new_n1386_), .ZN(new_n1387_));
  NOR2_X1    g0745(.A1(\in0[103] ), .A2(\in1[103] ), .ZN(new_n1388_));
  NAND2_X1   g0746(.A1(\in0[102] ), .A2(\in1[102] ), .ZN(new_n1389_));
  NOR2_X1    g0747(.A1(new_n1388_), .A2(new_n1389_), .ZN(new_n1390_));
  AOI21_X1   g0748(.A1(\in0[103] ), .A2(\in1[103] ), .B(new_n1390_), .ZN(new_n1391_));
  AOI22_X1   g0749(.A1(\in0[100] ), .A2(\in1[101] ), .B1(\in0[101] ), .B2(\in1[100] ), .ZN(new_n1392_));
  OR3_X2     g0750(.A1(new_n1391_), .A2(new_n1385_), .A3(new_n1392_), .Z(new_n1393_));
  INV_X1     g0751(.I(new_n1267_), .ZN(new_n1394_));
  INV_X1     g0752(.I(\in0[96] ), .ZN(new_n1395_));
  INV_X1     g0753(.I(\in1[96] ), .ZN(new_n1396_));
  NAND2_X1   g0754(.A1(\in0[98] ), .A2(\in1[97] ), .ZN(new_n1397_));
  NAND2_X1   g0755(.A1(\in0[97] ), .A2(\in1[98] ), .ZN(new_n1398_));
  NAND4_X1   g0756(.A1(new_n1397_), .A2(new_n1398_), .A3(new_n1395_), .A4(new_n1396_), .ZN(new_n1399_));
  INV_X1     g0757(.I(\in0[99] ), .ZN(new_n1400_));
  NOR3_X1    g0758(.A1(new_n1400_), .A2(new_n1266_), .A3(\in0[97] ), .ZN(new_n1401_));
  AOI22_X1   g0759(.A1(new_n1399_), .A2(new_n1401_), .B1(new_n1394_), .B2(\in1[99] ), .ZN(new_n1402_));
  OAI21_X1   g0760(.A1(new_n1393_), .A2(new_n1387_), .B(new_n1402_), .ZN(new_n1403_));
  NAND3_X1   g0761(.A1(new_n1380_), .A2(new_n1403_), .A3(new_n1355_), .ZN(new_n1404_));
  AOI22_X1   g0762(.A1(\in0[70] ), .A2(\in1[71] ), .B1(\in0[71] ), .B2(\in1[70] ), .ZN(new_n1405_));
  AOI22_X1   g0763(.A1(\in0[68] ), .A2(\in1[69] ), .B1(\in0[69] ), .B2(\in1[68] ), .ZN(new_n1406_));
  INV_X1     g0764(.I(\in0[69] ), .ZN(new_n1407_));
  INV_X1     g0765(.I(\in1[69] ), .ZN(new_n1408_));
  NAND2_X1   g0766(.A1(\in0[68] ), .A2(\in1[68] ), .ZN(new_n1409_));
  AOI21_X1   g0767(.A1(new_n1407_), .A2(new_n1408_), .B(new_n1409_), .ZN(new_n1410_));
  NOR2_X1    g0768(.A1(new_n1407_), .A2(new_n1408_), .ZN(new_n1411_));
  NOR3_X1    g0769(.A1(new_n1410_), .A2(new_n1405_), .A3(new_n1411_), .ZN(new_n1412_));
  OAI21_X1   g0770(.A1(\in0[73] ), .A2(new_n1377_), .B(new_n1369_), .ZN(new_n1413_));
  NAND2_X1   g0771(.A1(\in0[71] ), .A2(\in1[71] ), .ZN(new_n1414_));
  NOR2_X1    g0772(.A1(\in0[71] ), .A2(\in1[71] ), .ZN(new_n1415_));
  NAND2_X1   g0773(.A1(\in0[70] ), .A2(\in1[70] ), .ZN(new_n1416_));
  OAI21_X1   g0774(.A1(new_n1415_), .A2(new_n1416_), .B(new_n1414_), .ZN(new_n1417_));
  NAND4_X1   g0775(.A1(new_n1413_), .A2(\in0[72] ), .A3(\in1[72] ), .A4(new_n1417_), .ZN(new_n1418_));
  OAI22_X1   g0776(.A1(new_n1418_), .A2(new_n1412_), .B1(new_n1405_), .B2(new_n1406_), .ZN(new_n1419_));
  INV_X1     g0777(.I(\in0[31] ), .ZN(new_n1420_));
  AOI22_X1   g0778(.A1(\in0[38] ), .A2(\in1[39] ), .B1(\in0[39] ), .B2(\in1[38] ), .ZN(new_n1421_));
  NAND2_X1   g0779(.A1(\in0[37] ), .A2(\in1[36] ), .ZN(new_n1422_));
  NAND2_X1   g0780(.A1(\in0[36] ), .A2(\in1[37] ), .ZN(new_n1423_));
  AOI21_X1   g0781(.A1(new_n1422_), .A2(new_n1423_), .B(new_n1421_), .ZN(new_n1424_));
  INV_X1     g0782(.I(\in0[32] ), .ZN(new_n1425_));
  INV_X1     g0783(.I(\in0[33] ), .ZN(new_n1426_));
  INV_X1     g0784(.I(\in1[32] ), .ZN(new_n1427_));
  INV_X1     g0785(.I(\in1[33] ), .ZN(new_n1428_));
  OAI22_X1   g0786(.A1(new_n1425_), .A2(new_n1428_), .B1(new_n1426_), .B2(new_n1427_), .ZN(new_n1429_));
  NAND2_X1   g0787(.A1(\in0[35] ), .A2(\in1[34] ), .ZN(new_n1430_));
  NAND2_X1   g0788(.A1(\in0[34] ), .A2(\in1[35] ), .ZN(new_n1431_));
  NAND2_X1   g0789(.A1(new_n1430_), .A2(new_n1431_), .ZN(new_n1432_));
  NAND3_X1   g0790(.A1(new_n1424_), .A2(new_n1429_), .A3(new_n1432_), .ZN(new_n1433_));
  NAND2_X1   g0791(.A1(new_n1433_), .A2(new_n1420_), .ZN(new_n1434_));
  INV_X1     g0792(.I(\in1[31] ), .ZN(new_n1435_));
  OAI21_X1   g0793(.A1(new_n1433_), .A2(new_n1420_), .B(new_n1435_), .ZN(new_n1436_));
  NAND3_X1   g0794(.A1(new_n1419_), .A2(new_n1434_), .A3(new_n1436_), .ZN(new_n1437_));
  INV_X1     g0795(.I(\in0[81] ), .ZN(new_n1438_));
  NAND2_X1   g0796(.A1(\in0[83] ), .A2(\in1[82] ), .ZN(new_n1439_));
  NAND2_X1   g0797(.A1(\in0[82] ), .A2(\in1[83] ), .ZN(new_n1440_));
  NAND2_X1   g0798(.A1(new_n1439_), .A2(new_n1440_), .ZN(new_n1441_));
  AOI21_X1   g0799(.A1(new_n1438_), .A2(\in1[81] ), .B(new_n1441_), .ZN(new_n1442_));
  NAND2_X1   g0800(.A1(\in0[80] ), .A2(\in1[80] ), .ZN(new_n1443_));
  INV_X1     g0801(.I(\in0[80] ), .ZN(new_n1444_));
  INV_X1     g0802(.I(\in1[80] ), .ZN(new_n1445_));
  NAND2_X1   g0803(.A1(\in0[82] ), .A2(\in1[81] ), .ZN(new_n1446_));
  NAND2_X1   g0804(.A1(\in0[81] ), .A2(\in1[82] ), .ZN(new_n1447_));
  NAND4_X1   g0805(.A1(new_n1446_), .A2(new_n1447_), .A3(new_n1444_), .A4(new_n1445_), .ZN(new_n1448_));
  AND3_X2    g0806(.A1(new_n1438_), .A2(\in0[83] ), .A3(\in1[81] ), .Z(new_n1449_));
  AOI22_X1   g0807(.A1(new_n1449_), .A2(new_n1448_), .B1(\in1[83] ), .B2(new_n1441_), .ZN(new_n1450_));
  AOI22_X1   g0808(.A1(\in0[86] ), .A2(\in1[87] ), .B1(\in0[87] ), .B2(\in1[86] ), .ZN(new_n1451_));
  AOI22_X1   g0809(.A1(\in0[84] ), .A2(\in1[85] ), .B1(\in0[85] ), .B2(\in1[84] ), .ZN(new_n1452_));
  OR2_X2     g0810(.A1(new_n1451_), .A2(new_n1452_), .Z(new_n1453_));
  OAI22_X1   g0811(.A1(new_n1450_), .A2(new_n1453_), .B1(new_n1442_), .B2(new_n1443_), .ZN(new_n1454_));
  INV_X1     g0812(.I(\in0[87] ), .ZN(new_n1455_));
  INV_X1     g0813(.I(\in1[87] ), .ZN(new_n1456_));
  NOR2_X1    g0814(.A1(new_n1455_), .A2(new_n1456_), .ZN(new_n1457_));
  NAND2_X1   g0815(.A1(new_n1455_), .A2(new_n1456_), .ZN(new_n1458_));
  AND2_X2    g0816(.A1(\in0[86] ), .A2(\in1[86] ), .Z(new_n1459_));
  AOI21_X1   g0817(.A1(new_n1458_), .A2(new_n1459_), .B(new_n1457_), .ZN(new_n1460_));
  INV_X1     g0818(.I(\in0[85] ), .ZN(new_n1461_));
  INV_X1     g0819(.I(\in1[85] ), .ZN(new_n1462_));
  NAND2_X1   g0820(.A1(\in0[84] ), .A2(\in1[84] ), .ZN(new_n1463_));
  AOI21_X1   g0821(.A1(new_n1461_), .A2(new_n1462_), .B(new_n1463_), .ZN(new_n1464_));
  NOR2_X1    g0822(.A1(new_n1461_), .A2(new_n1462_), .ZN(new_n1465_));
  NOR3_X1    g0823(.A1(new_n1464_), .A2(new_n1451_), .A3(new_n1465_), .ZN(new_n1466_));
  NAND2_X1   g0824(.A1(\in0[91] ), .A2(\in1[90] ), .ZN(new_n1467_));
  NAND2_X1   g0825(.A1(\in0[90] ), .A2(\in1[91] ), .ZN(new_n1468_));
  NAND2_X1   g0826(.A1(new_n1467_), .A2(new_n1468_), .ZN(new_n1469_));
  INV_X1     g0827(.I(\in0[88] ), .ZN(new_n1470_));
  INV_X1     g0828(.I(\in1[88] ), .ZN(new_n1471_));
  NAND2_X1   g0829(.A1(\in0[90] ), .A2(\in1[89] ), .ZN(new_n1472_));
  NAND2_X1   g0830(.A1(\in0[89] ), .A2(\in1[90] ), .ZN(new_n1473_));
  NAND4_X1   g0831(.A1(new_n1472_), .A2(new_n1473_), .A3(new_n1470_), .A4(new_n1471_), .ZN(new_n1474_));
  INV_X1     g0832(.I(\in0[91] ), .ZN(new_n1475_));
  INV_X1     g0833(.I(\in1[89] ), .ZN(new_n1476_));
  NOR3_X1    g0834(.A1(new_n1475_), .A2(new_n1476_), .A3(\in0[89] ), .ZN(new_n1477_));
  AOI22_X1   g0835(.A1(new_n1474_), .A2(new_n1477_), .B1(new_n1469_), .B2(\in1[91] ), .ZN(new_n1478_));
  NOR2_X1    g0836(.A1(new_n1476_), .A2(\in0[89] ), .ZN(new_n1479_));
  NOR2_X1    g0837(.A1(new_n1470_), .A2(new_n1471_), .ZN(new_n1480_));
  OAI21_X1   g0838(.A1(new_n1469_), .A2(new_n1479_), .B(new_n1480_), .ZN(new_n1481_));
  OAI22_X1   g0839(.A1(new_n1478_), .A2(new_n1481_), .B1(new_n1466_), .B2(new_n1460_), .ZN(new_n1482_));
  NAND2_X1   g0840(.A1(new_n1454_), .A2(new_n1482_), .ZN(new_n1483_));
  NOR4_X1    g0841(.A1(new_n1404_), .A2(new_n1337_), .A3(new_n1437_), .A4(new_n1483_), .ZN(new_n1484_));
  INV_X1     g0842(.I(\in0[59] ), .ZN(new_n1485_));
  AOI22_X1   g0843(.A1(\in0[57] ), .A2(\in1[58] ), .B1(\in0[58] ), .B2(\in1[57] ), .ZN(new_n1486_));
  OR2_X2     g0844(.A1(\in0[56] ), .A2(\in1[56] ), .Z(new_n1487_));
  AND2_X2    g0845(.A1(\in0[57] ), .A2(\in1[57] ), .Z(new_n1488_));
  AOI21_X1   g0846(.A1(new_n1488_), .A2(new_n1487_), .B(new_n1486_), .ZN(new_n1489_));
  NAND2_X1   g0847(.A1(\in0[63] ), .A2(\in1[62] ), .ZN(new_n1490_));
  NAND2_X1   g0848(.A1(\in0[62] ), .A2(\in1[63] ), .ZN(new_n1491_));
  NAND2_X1   g0849(.A1(new_n1490_), .A2(new_n1491_), .ZN(new_n1492_));
  NAND2_X1   g0850(.A1(\in0[61] ), .A2(\in1[60] ), .ZN(new_n1493_));
  NAND2_X1   g0851(.A1(\in0[60] ), .A2(\in1[61] ), .ZN(new_n1494_));
  NAND2_X1   g0852(.A1(new_n1493_), .A2(new_n1494_), .ZN(new_n1495_));
  NAND2_X1   g0853(.A1(\in0[59] ), .A2(\in1[58] ), .ZN(new_n1496_));
  NAND2_X1   g0854(.A1(\in0[58] ), .A2(\in1[59] ), .ZN(new_n1497_));
  NAND2_X1   g0855(.A1(new_n1496_), .A2(new_n1497_), .ZN(new_n1498_));
  NAND3_X1   g0856(.A1(new_n1492_), .A2(new_n1495_), .A3(new_n1498_), .ZN(new_n1499_));
  OAI21_X1   g0857(.A1(new_n1499_), .A2(new_n1489_), .B(new_n1485_), .ZN(new_n1500_));
  NAND2_X1   g0858(.A1(\in0[63] ), .A2(\in1[63] ), .ZN(new_n1501_));
  NOR2_X1    g0859(.A1(\in0[63] ), .A2(\in1[63] ), .ZN(new_n1502_));
  NAND2_X1   g0860(.A1(\in0[62] ), .A2(\in1[62] ), .ZN(new_n1503_));
  OAI21_X1   g0861(.A1(new_n1502_), .A2(new_n1503_), .B(new_n1501_), .ZN(new_n1504_));
  AOI21_X1   g0862(.A1(new_n1500_), .A2(\in1[59] ), .B(new_n1504_), .ZN(new_n1505_));
  NAND2_X1   g0863(.A1(\in0[61] ), .A2(\in1[61] ), .ZN(new_n1506_));
  NOR2_X1    g0864(.A1(\in0[61] ), .A2(\in1[61] ), .ZN(new_n1507_));
  NAND2_X1   g0865(.A1(\in0[60] ), .A2(\in1[60] ), .ZN(new_n1508_));
  OAI21_X1   g0866(.A1(new_n1507_), .A2(new_n1508_), .B(new_n1506_), .ZN(new_n1509_));
  NAND2_X1   g0867(.A1(new_n1509_), .A2(new_n1492_), .ZN(new_n1510_));
  INV_X1     g0868(.I(\in1[67] ), .ZN(new_n1511_));
  AOI22_X1   g0869(.A1(\in0[66] ), .A2(\in1[67] ), .B1(\in0[67] ), .B2(\in1[66] ), .ZN(new_n1512_));
  NOR2_X1    g0870(.A1(new_n1512_), .A2(new_n1511_), .ZN(new_n1513_));
  NAND2_X1   g0871(.A1(\in0[66] ), .A2(\in1[65] ), .ZN(new_n1514_));
  AND2_X2    g0872(.A1(\in0[65] ), .A2(\in1[66] ), .Z(new_n1515_));
  NOR3_X1    g0873(.A1(new_n1515_), .A2(\in0[64] ), .A3(\in1[64] ), .ZN(new_n1516_));
  NAND2_X1   g0874(.A1(new_n1516_), .A2(new_n1514_), .ZN(new_n1517_));
  INV_X1     g0875(.I(\in0[67] ), .ZN(new_n1518_));
  INV_X1     g0876(.I(\in0[65] ), .ZN(new_n1519_));
  NAND2_X1   g0877(.A1(new_n1519_), .A2(\in1[65] ), .ZN(new_n1520_));
  NOR2_X1    g0878(.A1(new_n1520_), .A2(new_n1518_), .ZN(new_n1521_));
  AOI21_X1   g0879(.A1(new_n1517_), .A2(new_n1521_), .B(new_n1513_), .ZN(new_n1522_));
  NAND2_X1   g0880(.A1(new_n1512_), .A2(new_n1520_), .ZN(new_n1523_));
  NAND3_X1   g0881(.A1(new_n1523_), .A2(\in0[64] ), .A3(\in1[64] ), .ZN(new_n1524_));
  OAI22_X1   g0882(.A1(new_n1505_), .A2(new_n1510_), .B1(new_n1522_), .B2(new_n1524_), .ZN(new_n1525_));
  INV_X1     g0883(.I(\in0[35] ), .ZN(new_n1526_));
  AOI22_X1   g0884(.A1(\in0[33] ), .A2(\in1[34] ), .B1(\in0[34] ), .B2(\in1[33] ), .ZN(new_n1527_));
  NAND2_X1   g0885(.A1(new_n1425_), .A2(new_n1427_), .ZN(new_n1528_));
  NOR2_X1    g0886(.A1(new_n1426_), .A2(new_n1428_), .ZN(new_n1529_));
  AOI21_X1   g0887(.A1(new_n1529_), .A2(new_n1528_), .B(new_n1527_), .ZN(new_n1530_));
  NAND2_X1   g0888(.A1(new_n1424_), .A2(new_n1432_), .ZN(new_n1531_));
  OAI21_X1   g0889(.A1(new_n1531_), .A2(new_n1530_), .B(new_n1526_), .ZN(new_n1532_));
  NAND2_X1   g0890(.A1(\in0[39] ), .A2(\in1[39] ), .ZN(new_n1533_));
  NOR2_X1    g0891(.A1(\in0[39] ), .A2(\in1[39] ), .ZN(new_n1534_));
  NAND2_X1   g0892(.A1(\in0[38] ), .A2(\in1[38] ), .ZN(new_n1535_));
  OAI21_X1   g0893(.A1(new_n1534_), .A2(new_n1535_), .B(new_n1533_), .ZN(new_n1536_));
  AOI21_X1   g0894(.A1(new_n1532_), .A2(\in1[35] ), .B(new_n1536_), .ZN(new_n1537_));
  INV_X1     g0895(.I(new_n1421_), .ZN(new_n1538_));
  NAND2_X1   g0896(.A1(\in0[37] ), .A2(\in1[37] ), .ZN(new_n1539_));
  NOR2_X1    g0897(.A1(\in0[37] ), .A2(\in1[37] ), .ZN(new_n1540_));
  NAND2_X1   g0898(.A1(\in0[36] ), .A2(\in1[36] ), .ZN(new_n1541_));
  OAI21_X1   g0899(.A1(new_n1540_), .A2(new_n1541_), .B(new_n1539_), .ZN(new_n1542_));
  NAND2_X1   g0900(.A1(new_n1542_), .A2(new_n1538_), .ZN(new_n1543_));
  INV_X1     g0901(.I(\in0[43] ), .ZN(new_n1544_));
  AOI22_X1   g0902(.A1(\in0[41] ), .A2(\in1[42] ), .B1(\in0[42] ), .B2(\in1[41] ), .ZN(new_n1545_));
  INV_X1     g0903(.I(\in0[40] ), .ZN(new_n1546_));
  INV_X1     g0904(.I(\in1[40] ), .ZN(new_n1547_));
  NAND2_X1   g0905(.A1(new_n1546_), .A2(new_n1547_), .ZN(new_n1548_));
  INV_X1     g0906(.I(\in0[41] ), .ZN(new_n1549_));
  INV_X1     g0907(.I(\in1[41] ), .ZN(new_n1550_));
  NOR2_X1    g0908(.A1(new_n1549_), .A2(new_n1550_), .ZN(new_n1551_));
  AOI21_X1   g0909(.A1(new_n1551_), .A2(new_n1548_), .B(new_n1545_), .ZN(new_n1552_));
  AOI22_X1   g0910(.A1(\in0[46] ), .A2(\in1[47] ), .B1(\in0[47] ), .B2(\in1[46] ), .ZN(new_n1553_));
  AOI22_X1   g0911(.A1(\in0[44] ), .A2(\in1[45] ), .B1(\in0[45] ), .B2(\in1[44] ), .ZN(new_n1554_));
  AOI22_X1   g0912(.A1(\in0[42] ), .A2(\in1[43] ), .B1(\in0[43] ), .B2(\in1[42] ), .ZN(new_n1555_));
  NOR3_X1    g0913(.A1(new_n1553_), .A2(new_n1554_), .A3(new_n1555_), .ZN(new_n1556_));
  INV_X1     g0914(.I(new_n1556_), .ZN(new_n1557_));
  OAI21_X1   g0915(.A1(new_n1557_), .A2(new_n1552_), .B(new_n1544_), .ZN(new_n1558_));
  NAND2_X1   g0916(.A1(\in0[47] ), .A2(\in1[47] ), .ZN(new_n1559_));
  NOR2_X1    g0917(.A1(\in0[47] ), .A2(\in1[47] ), .ZN(new_n1560_));
  NAND2_X1   g0918(.A1(\in0[46] ), .A2(\in1[46] ), .ZN(new_n1561_));
  OAI21_X1   g0919(.A1(new_n1560_), .A2(new_n1561_), .B(new_n1559_), .ZN(new_n1562_));
  AOI21_X1   g0920(.A1(new_n1558_), .A2(\in1[43] ), .B(new_n1562_), .ZN(new_n1563_));
  INV_X1     g0921(.I(new_n1553_), .ZN(new_n1564_));
  NAND2_X1   g0922(.A1(\in0[45] ), .A2(\in1[45] ), .ZN(new_n1565_));
  NOR2_X1    g0923(.A1(\in0[45] ), .A2(\in1[45] ), .ZN(new_n1566_));
  NAND2_X1   g0924(.A1(\in0[44] ), .A2(\in1[44] ), .ZN(new_n1567_));
  OAI21_X1   g0925(.A1(new_n1566_), .A2(new_n1567_), .B(new_n1565_), .ZN(new_n1568_));
  OAI22_X1   g0926(.A1(new_n1546_), .A2(new_n1550_), .B1(new_n1549_), .B2(new_n1547_), .ZN(new_n1569_));
  NAND4_X1   g0927(.A1(new_n1556_), .A2(new_n1564_), .A3(new_n1568_), .A4(new_n1569_), .ZN(new_n1570_));
  OAI22_X1   g0928(.A1(new_n1537_), .A2(new_n1543_), .B1(new_n1563_), .B2(new_n1570_), .ZN(new_n1571_));
  INV_X1     g0929(.I(\in1[53] ), .ZN(new_n1572_));
  NOR2_X1    g0930(.A1(new_n1572_), .A2(\in0[53] ), .ZN(new_n1573_));
  INV_X1     g0931(.I(new_n1573_), .ZN(new_n1574_));
  AOI22_X1   g0932(.A1(\in0[54] ), .A2(\in1[55] ), .B1(\in0[55] ), .B2(\in1[54] ), .ZN(new_n1575_));
  NAND2_X1   g0933(.A1(new_n1574_), .A2(new_n1575_), .ZN(new_n1576_));
  AND3_X2    g0934(.A1(new_n1576_), .A2(\in0[52] ), .A3(\in1[52] ), .Z(new_n1577_));
  INV_X1     g0935(.I(new_n1577_), .ZN(new_n1578_));
  INV_X1     g0936(.I(\in0[48] ), .ZN(new_n1579_));
  INV_X1     g0937(.I(\in0[49] ), .ZN(new_n1580_));
  INV_X1     g0938(.I(\in1[48] ), .ZN(new_n1581_));
  INV_X1     g0939(.I(\in1[49] ), .ZN(new_n1582_));
  OAI22_X1   g0940(.A1(new_n1579_), .A2(new_n1582_), .B1(new_n1580_), .B2(new_n1581_), .ZN(new_n1583_));
  NAND2_X1   g0941(.A1(\in0[51] ), .A2(\in1[50] ), .ZN(new_n1584_));
  NAND2_X1   g0942(.A1(\in0[50] ), .A2(\in1[51] ), .ZN(new_n1585_));
  NAND2_X1   g0943(.A1(new_n1584_), .A2(new_n1585_), .ZN(new_n1586_));
  NAND2_X1   g0944(.A1(new_n1583_), .A2(new_n1586_), .ZN(new_n1587_));
  INV_X1     g0945(.I(\in0[51] ), .ZN(new_n1588_));
  AOI22_X1   g0946(.A1(\in0[49] ), .A2(\in1[50] ), .B1(\in0[50] ), .B2(\in1[49] ), .ZN(new_n1589_));
  NOR2_X1    g0947(.A1(\in0[48] ), .A2(\in1[48] ), .ZN(new_n1590_));
  NOR3_X1    g0948(.A1(new_n1590_), .A2(new_n1580_), .A3(new_n1582_), .ZN(new_n1591_));
  OAI21_X1   g0949(.A1(new_n1589_), .A2(new_n1591_), .B(new_n1586_), .ZN(new_n1592_));
  OAI21_X1   g0950(.A1(new_n1578_), .A2(new_n1592_), .B(new_n1588_), .ZN(new_n1593_));
  INV_X1     g0951(.I(\in0[53] ), .ZN(new_n1594_));
  INV_X1     g0952(.I(\in0[54] ), .ZN(new_n1595_));
  INV_X1     g0953(.I(\in1[54] ), .ZN(new_n1596_));
  OAI22_X1   g0954(.A1(new_n1594_), .A2(new_n1596_), .B1(new_n1595_), .B2(new_n1572_), .ZN(new_n1597_));
  INV_X1     g0955(.I(\in0[52] ), .ZN(new_n1598_));
  OR3_X2     g0956(.A1(new_n1573_), .A2(new_n1598_), .A3(\in1[52] ), .Z(new_n1599_));
  AOI21_X1   g0957(.A1(new_n1599_), .A2(new_n1597_), .B(new_n1575_), .ZN(new_n1600_));
  AOI21_X1   g0958(.A1(new_n1593_), .A2(\in1[51] ), .B(new_n1600_), .ZN(new_n1601_));
  AOI22_X1   g0959(.A1(\in0[56] ), .A2(\in1[57] ), .B1(\in0[57] ), .B2(\in1[56] ), .ZN(new_n1602_));
  NAND2_X1   g0960(.A1(\in0[55] ), .A2(\in1[55] ), .ZN(new_n1603_));
  NOR2_X1    g0961(.A1(new_n1602_), .A2(new_n1603_), .ZN(new_n1604_));
  NAND4_X1   g0962(.A1(new_n1604_), .A2(new_n1492_), .A3(new_n1495_), .A4(new_n1498_), .ZN(new_n1605_));
  OAI22_X1   g0963(.A1(new_n1601_), .A2(new_n1605_), .B1(new_n1578_), .B2(new_n1587_), .ZN(new_n1606_));
  NAND4_X1   g0964(.A1(new_n1606_), .A2(new_n1484_), .A3(new_n1525_), .A4(new_n1571_), .ZN(new_n1607_));
  AOI21_X1   g0965(.A1(new_n1257_), .A2(new_n1139_), .B(new_n1607_), .ZN(new_n1608_));
  AOI21_X1   g0966(.A1(new_n1608_), .A2(new_n1135_), .B(new_n1134_), .ZN(new_n1609_));
  AOI21_X1   g0967(.A1(new_n1129_), .A2(new_n643_), .B(new_n854_), .ZN(new_n1610_));
  INV_X1     g0968(.I(new_n1610_), .ZN(new_n1611_));
  NOR2_X1    g0969(.A1(new_n1611_), .A2(new_n1609_), .ZN(new_n1612_));
  NOR2_X1    g0970(.A1(new_n1135_), .A2(\in0[127] ), .ZN(new_n1613_));
  INV_X1     g0971(.I(new_n1613_), .ZN(new_n1614_));
  NAND2_X1   g0972(.A1(new_n1608_), .A2(new_n1614_), .ZN(new_n1615_));
  NOR2_X1    g0973(.A1(new_n1615_), .A2(\in1[30] ), .ZN(new_n1616_));
  AOI21_X1   g0974(.A1(new_n1137_), .A2(new_n1615_), .B(new_n1616_), .ZN(new_n1617_));
  INV_X1     g0975(.I(new_n1617_), .ZN(new_n1618_));
  INV_X1     g0976(.I(\in3[30] ), .ZN(new_n1619_));
  INV_X1     g0977(.I(new_n651_), .ZN(new_n1620_));
  INV_X1     g0978(.I(new_n656_), .ZN(new_n1621_));
  INV_X1     g0979(.I(new_n663_), .ZN(new_n1622_));
  INV_X1     g0980(.I(new_n668_), .ZN(new_n1623_));
  INV_X1     g0981(.I(new_n675_), .ZN(new_n1624_));
  INV_X1     g0982(.I(new_n681_), .ZN(new_n1625_));
  NOR3_X1    g0983(.A1(\in2[0] ), .A2(\in2[1] ), .A3(\in3[1] ), .ZN(new_n1626_));
  NOR2_X1    g0984(.A1(new_n1131_), .A2(\in3[0] ), .ZN(new_n1627_));
  INV_X1     g0985(.I(\in2[1] ), .ZN(new_n1628_));
  NAND2_X1   g0986(.A1(new_n1628_), .A2(\in3[0] ), .ZN(new_n1629_));
  NOR4_X1    g0987(.A1(new_n1627_), .A2(new_n1629_), .A3(new_n1626_), .A4(new_n693_), .ZN(new_n1630_));
  OAI22_X1   g0988(.A1(new_n1630_), .A2(new_n690_), .B1(new_n685_), .B2(\in3[3] ), .ZN(new_n1631_));
  AOI22_X1   g0989(.A1(new_n1631_), .A2(new_n686_), .B1(\in2[4] ), .B2(new_n682_), .ZN(new_n1632_));
  OAI21_X1   g0990(.A1(new_n1632_), .A2(new_n683_), .B(new_n708_), .ZN(new_n1633_));
  AOI22_X1   g0991(.A1(new_n1633_), .A2(new_n1625_), .B1(\in2[8] ), .B2(new_n676_), .ZN(new_n1634_));
  OAI21_X1   g0992(.A1(new_n1634_), .A2(new_n677_), .B(new_n718_), .ZN(new_n1635_));
  INV_X1     g0993(.I(new_n726_), .ZN(new_n1636_));
  AOI21_X1   g0994(.A1(new_n1635_), .A2(new_n1624_), .B(new_n1636_), .ZN(new_n1637_));
  OAI21_X1   g0995(.A1(new_n1637_), .A2(new_n671_), .B(new_n728_), .ZN(new_n1638_));
  INV_X1     g0996(.I(new_n731_), .ZN(new_n1639_));
  AOI21_X1   g0997(.A1(new_n1638_), .A2(new_n1623_), .B(new_n1639_), .ZN(new_n1640_));
  OAI21_X1   g0998(.A1(new_n1640_), .A2(new_n665_), .B(new_n738_), .ZN(new_n1641_));
  INV_X1     g0999(.I(new_n746_), .ZN(new_n1642_));
  AOI21_X1   g1000(.A1(new_n1641_), .A2(new_n1622_), .B(new_n1642_), .ZN(new_n1643_));
  OAI21_X1   g1001(.A1(new_n1643_), .A2(new_n659_), .B(new_n748_), .ZN(new_n1644_));
  INV_X1     g1002(.I(new_n751_), .ZN(new_n1645_));
  AOI21_X1   g1003(.A1(new_n1644_), .A2(new_n1621_), .B(new_n1645_), .ZN(new_n1646_));
  OAI21_X1   g1004(.A1(new_n1646_), .A2(new_n653_), .B(new_n758_), .ZN(new_n1647_));
  INV_X1     g1005(.I(new_n766_), .ZN(new_n1648_));
  AOI21_X1   g1006(.A1(new_n1647_), .A2(new_n1620_), .B(new_n1648_), .ZN(new_n1649_));
  INV_X1     g1007(.I(new_n1128_), .ZN(new_n1650_));
  OAI21_X1   g1008(.A1(new_n1649_), .A2(new_n647_), .B(new_n1650_), .ZN(new_n1651_));
  NOR2_X1    g1009(.A1(new_n1651_), .A2(new_n644_), .ZN(new_n1652_));
  NOR2_X1    g1010(.A1(new_n1652_), .A2(\in2[30] ), .ZN(new_n1653_));
  AOI21_X1   g1011(.A1(new_n1619_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n1654_));
  INV_X1     g1012(.I(new_n1654_), .ZN(new_n1655_));
  NAND2_X1   g1013(.A1(new_n1618_), .A2(new_n1655_), .ZN(new_n1656_));
  NOR2_X1    g1014(.A1(new_n1615_), .A2(\in1[27] ), .ZN(new_n1657_));
  AOI21_X1   g1015(.A1(new_n1141_), .A2(new_n1615_), .B(new_n1657_), .ZN(new_n1658_));
  INV_X1     g1016(.I(\in3[27] ), .ZN(new_n1659_));
  NOR2_X1    g1017(.A1(new_n1652_), .A2(\in2[27] ), .ZN(new_n1660_));
  AOI21_X1   g1018(.A1(new_n1659_), .A2(new_n1652_), .B(new_n1660_), .ZN(new_n1661_));
  NOR2_X1    g1019(.A1(new_n1658_), .A2(new_n1661_), .ZN(new_n1662_));
  NOR2_X1    g1020(.A1(new_n1652_), .A2(\in2[24] ), .ZN(new_n1663_));
  AOI21_X1   g1021(.A1(new_n652_), .A2(new_n1652_), .B(new_n1663_), .ZN(new_n1664_));
  NOR2_X1    g1022(.A1(new_n1615_), .A2(\in1[24] ), .ZN(new_n1665_));
  AOI21_X1   g1023(.A1(new_n1239_), .A2(new_n1615_), .B(new_n1665_), .ZN(new_n1666_));
  INV_X1     g1024(.I(new_n1666_), .ZN(new_n1667_));
  NAND2_X1   g1025(.A1(new_n1667_), .A2(new_n1664_), .ZN(new_n1668_));
  NOR2_X1    g1026(.A1(new_n1652_), .A2(\in2[23] ), .ZN(new_n1669_));
  AOI21_X1   g1027(.A1(new_n655_), .A2(new_n1652_), .B(new_n1669_), .ZN(new_n1670_));
  INV_X1     g1028(.I(new_n1670_), .ZN(new_n1671_));
  NOR2_X1    g1029(.A1(new_n1615_), .A2(\in1[23] ), .ZN(new_n1672_));
  AOI21_X1   g1030(.A1(new_n1146_), .A2(new_n1615_), .B(new_n1672_), .ZN(new_n1673_));
  NOR2_X1    g1031(.A1(new_n1671_), .A2(new_n1673_), .ZN(new_n1674_));
  NOR2_X1    g1032(.A1(new_n1615_), .A2(\in1[22] ), .ZN(new_n1675_));
  AOI21_X1   g1033(.A1(new_n1150_), .A2(new_n1615_), .B(new_n1675_), .ZN(new_n1676_));
  INV_X1     g1034(.I(new_n1676_), .ZN(new_n1677_));
  INV_X1     g1035(.I(\in3[22] ), .ZN(new_n1678_));
  NOR2_X1    g1036(.A1(new_n1652_), .A2(\in2[22] ), .ZN(new_n1679_));
  AOI21_X1   g1037(.A1(new_n1678_), .A2(new_n1652_), .B(new_n1679_), .ZN(new_n1680_));
  INV_X1     g1038(.I(new_n1680_), .ZN(new_n1681_));
  NAND2_X1   g1039(.A1(new_n1677_), .A2(new_n1681_), .ZN(new_n1682_));
  NOR2_X1    g1040(.A1(new_n1615_), .A2(\in1[19] ), .ZN(new_n1683_));
  AOI21_X1   g1041(.A1(new_n1154_), .A2(new_n1615_), .B(new_n1683_), .ZN(new_n1684_));
  INV_X1     g1042(.I(\in3[19] ), .ZN(new_n1685_));
  NOR2_X1    g1043(.A1(new_n1652_), .A2(\in2[19] ), .ZN(new_n1686_));
  AOI21_X1   g1044(.A1(new_n1685_), .A2(new_n1652_), .B(new_n1686_), .ZN(new_n1687_));
  NOR2_X1    g1045(.A1(new_n1684_), .A2(new_n1687_), .ZN(new_n1688_));
  NOR2_X1    g1046(.A1(new_n1652_), .A2(\in2[16] ), .ZN(new_n1689_));
  AOI21_X1   g1047(.A1(new_n664_), .A2(new_n1652_), .B(new_n1689_), .ZN(new_n1690_));
  NOR2_X1    g1048(.A1(new_n1615_), .A2(\in1[16] ), .ZN(new_n1691_));
  AOI21_X1   g1049(.A1(new_n1218_), .A2(new_n1615_), .B(new_n1691_), .ZN(new_n1692_));
  INV_X1     g1050(.I(new_n1692_), .ZN(new_n1693_));
  NAND2_X1   g1051(.A1(new_n1693_), .A2(new_n1690_), .ZN(new_n1694_));
  NOR2_X1    g1052(.A1(new_n1652_), .A2(\in2[15] ), .ZN(new_n1695_));
  AOI21_X1   g1053(.A1(new_n667_), .A2(new_n1652_), .B(new_n1695_), .ZN(new_n1696_));
  INV_X1     g1054(.I(new_n1696_), .ZN(new_n1697_));
  NOR2_X1    g1055(.A1(new_n1615_), .A2(\in1[15] ), .ZN(new_n1698_));
  AOI21_X1   g1056(.A1(new_n1159_), .A2(new_n1615_), .B(new_n1698_), .ZN(new_n1699_));
  NOR2_X1    g1057(.A1(new_n1697_), .A2(new_n1699_), .ZN(new_n1700_));
  NOR2_X1    g1058(.A1(new_n1615_), .A2(\in1[14] ), .ZN(new_n1701_));
  AOI21_X1   g1059(.A1(new_n1163_), .A2(new_n1615_), .B(new_n1701_), .ZN(new_n1702_));
  INV_X1     g1060(.I(new_n1702_), .ZN(new_n1703_));
  INV_X1     g1061(.I(\in3[14] ), .ZN(new_n1704_));
  NOR2_X1    g1062(.A1(new_n1652_), .A2(\in2[14] ), .ZN(new_n1705_));
  AOI21_X1   g1063(.A1(new_n1704_), .A2(new_n1652_), .B(new_n1705_), .ZN(new_n1706_));
  INV_X1     g1064(.I(new_n1706_), .ZN(new_n1707_));
  NAND2_X1   g1065(.A1(new_n1703_), .A2(new_n1707_), .ZN(new_n1708_));
  NAND2_X1   g1066(.A1(new_n1615_), .A2(new_n1167_), .ZN(new_n1709_));
  OAI21_X1   g1067(.A1(\in1[11] ), .A2(new_n1615_), .B(new_n1709_), .ZN(new_n1710_));
  INV_X1     g1068(.I(new_n1710_), .ZN(new_n1711_));
  INV_X1     g1069(.I(\in3[11] ), .ZN(new_n1712_));
  NOR2_X1    g1070(.A1(new_n1652_), .A2(\in2[11] ), .ZN(new_n1713_));
  AOI21_X1   g1071(.A1(new_n1712_), .A2(new_n1652_), .B(new_n1713_), .ZN(new_n1714_));
  NOR2_X1    g1072(.A1(new_n1711_), .A2(new_n1714_), .ZN(new_n1715_));
  NAND2_X1   g1073(.A1(new_n1652_), .A2(new_n676_), .ZN(new_n1716_));
  OAI21_X1   g1074(.A1(\in2[8] ), .A2(new_n1652_), .B(new_n1716_), .ZN(new_n1717_));
  NOR2_X1    g1075(.A1(new_n1615_), .A2(\in1[7] ), .ZN(new_n1718_));
  AOI21_X1   g1076(.A1(new_n1173_), .A2(new_n1615_), .B(new_n1718_), .ZN(new_n1719_));
  INV_X1     g1077(.I(new_n1719_), .ZN(new_n1720_));
  INV_X1     g1078(.I(\in3[7] ), .ZN(new_n1721_));
  NOR2_X1    g1079(.A1(new_n1652_), .A2(\in2[7] ), .ZN(new_n1722_));
  AOI21_X1   g1080(.A1(new_n1721_), .A2(new_n1652_), .B(new_n1722_), .ZN(new_n1723_));
  NOR2_X1    g1081(.A1(new_n1720_), .A2(new_n1723_), .ZN(new_n1724_));
  NAND2_X1   g1082(.A1(new_n1724_), .A2(new_n1717_), .ZN(new_n1725_));
  INV_X1     g1083(.I(\in3[5] ), .ZN(new_n1726_));
  NOR2_X1    g1084(.A1(new_n1652_), .A2(\in2[5] ), .ZN(new_n1727_));
  AOI21_X1   g1085(.A1(new_n1726_), .A2(new_n1652_), .B(new_n1727_), .ZN(new_n1728_));
  INV_X1     g1086(.I(\in0[5] ), .ZN(new_n1729_));
  NOR2_X1    g1087(.A1(new_n1615_), .A2(\in1[5] ), .ZN(new_n1730_));
  AOI21_X1   g1088(.A1(new_n1729_), .A2(new_n1615_), .B(new_n1730_), .ZN(new_n1731_));
  INV_X1     g1089(.I(new_n1731_), .ZN(new_n1732_));
  NAND2_X1   g1090(.A1(new_n1732_), .A2(new_n1728_), .ZN(new_n1733_));
  NAND2_X1   g1091(.A1(new_n1652_), .A2(new_n682_), .ZN(new_n1734_));
  OAI21_X1   g1092(.A1(\in2[4] ), .A2(new_n1652_), .B(new_n1734_), .ZN(new_n1735_));
  INV_X1     g1093(.I(\in0[4] ), .ZN(new_n1736_));
  NOR2_X1    g1094(.A1(new_n1615_), .A2(\in1[4] ), .ZN(new_n1737_));
  AOI21_X1   g1095(.A1(new_n1736_), .A2(new_n1615_), .B(new_n1737_), .ZN(new_n1738_));
  NOR2_X1    g1096(.A1(new_n1738_), .A2(new_n1735_), .ZN(new_n1739_));
  AOI21_X1   g1097(.A1(new_n1608_), .A2(new_n1614_), .B(\in0[3] ), .ZN(new_n1740_));
  INV_X1     g1098(.I(new_n1142_), .ZN(new_n1741_));
  INV_X1     g1099(.I(new_n1155_), .ZN(new_n1742_));
  INV_X1     g1100(.I(new_n1168_), .ZN(new_n1743_));
  INV_X1     g1101(.I(new_n1174_), .ZN(new_n1744_));
  AOI22_X1   g1102(.A1(new_n1187_), .A2(new_n1179_), .B1(\in0[4] ), .B2(new_n1175_), .ZN(new_n1745_));
  OAI21_X1   g1103(.A1(new_n1745_), .A2(new_n1176_), .B(new_n1196_), .ZN(new_n1746_));
  AOI22_X1   g1104(.A1(new_n1746_), .A2(new_n1744_), .B1(\in0[8] ), .B2(new_n1169_), .ZN(new_n1747_));
  OAI21_X1   g1105(.A1(new_n1747_), .A2(new_n1170_), .B(new_n1206_), .ZN(new_n1748_));
  INV_X1     g1106(.I(new_n1214_), .ZN(new_n1749_));
  AOI21_X1   g1107(.A1(new_n1748_), .A2(new_n1743_), .B(new_n1749_), .ZN(new_n1750_));
  NOR2_X1    g1108(.A1(new_n1750_), .A2(new_n1164_), .ZN(new_n1751_));
  OAI21_X1   g1109(.A1(new_n1751_), .A2(new_n1216_), .B(new_n1160_), .ZN(new_n1752_));
  AOI21_X1   g1110(.A1(new_n1752_), .A2(new_n1220_), .B(new_n1157_), .ZN(new_n1753_));
  OAI21_X1   g1111(.A1(new_n1753_), .A2(new_n1228_), .B(new_n1742_), .ZN(new_n1754_));
  AOI21_X1   g1112(.A1(new_n1754_), .A2(new_n1235_), .B(new_n1151_), .ZN(new_n1755_));
  OAI21_X1   g1113(.A1(new_n1755_), .A2(new_n1237_), .B(new_n1147_), .ZN(new_n1756_));
  AOI21_X1   g1114(.A1(new_n1756_), .A2(new_n1241_), .B(new_n1144_), .ZN(new_n1757_));
  OAI21_X1   g1115(.A1(new_n1757_), .A2(new_n1249_), .B(new_n1741_), .ZN(new_n1758_));
  AOI21_X1   g1116(.A1(new_n1758_), .A2(new_n1256_), .B(new_n1138_), .ZN(new_n1759_));
  NOR4_X1    g1117(.A1(new_n1759_), .A2(\in1[3] ), .A3(new_n1607_), .A4(new_n1613_), .ZN(new_n1760_));
  OR2_X2     g1118(.A1(new_n1740_), .A2(new_n1760_), .Z(new_n1761_));
  INV_X1     g1119(.I(new_n644_), .ZN(new_n1762_));
  AOI21_X1   g1120(.A1(new_n1129_), .A2(new_n1762_), .B(\in2[3] ), .ZN(new_n1763_));
  NOR3_X1    g1121(.A1(new_n1651_), .A2(\in3[3] ), .A3(new_n644_), .ZN(new_n1764_));
  OR2_X2     g1122(.A1(new_n1764_), .A2(new_n1763_), .Z(new_n1765_));
  NAND2_X1   g1123(.A1(new_n1761_), .A2(new_n1765_), .ZN(new_n1766_));
  INV_X1     g1124(.I(\in0[1] ), .ZN(new_n1767_));
  NAND2_X1   g1125(.A1(new_n1615_), .A2(new_n1767_), .ZN(new_n1768_));
  OAI21_X1   g1126(.A1(\in1[1] ), .A2(new_n1615_), .B(new_n1768_), .ZN(new_n1769_));
  INV_X1     g1127(.I(\in0[0] ), .ZN(new_n1770_));
  OAI22_X1   g1128(.A1(new_n1750_), .A2(new_n1164_), .B1(new_n1159_), .B2(\in1[15] ), .ZN(new_n1771_));
  AOI21_X1   g1129(.A1(new_n1771_), .A2(new_n1160_), .B(new_n1219_), .ZN(new_n1772_));
  OAI21_X1   g1130(.A1(new_n1772_), .A2(new_n1157_), .B(new_n1227_), .ZN(new_n1773_));
  INV_X1     g1131(.I(new_n1235_), .ZN(new_n1774_));
  AOI21_X1   g1132(.A1(new_n1773_), .A2(new_n1742_), .B(new_n1774_), .ZN(new_n1775_));
  OAI22_X1   g1133(.A1(new_n1775_), .A2(new_n1151_), .B1(new_n1146_), .B2(\in1[23] ), .ZN(new_n1776_));
  AOI21_X1   g1134(.A1(new_n1776_), .A2(new_n1147_), .B(new_n1240_), .ZN(new_n1777_));
  OAI21_X1   g1135(.A1(new_n1777_), .A2(new_n1144_), .B(new_n1248_), .ZN(new_n1778_));
  INV_X1     g1136(.I(new_n1256_), .ZN(new_n1779_));
  AOI21_X1   g1137(.A1(new_n1778_), .A2(new_n1741_), .B(new_n1779_), .ZN(new_n1780_));
  INV_X1     g1138(.I(new_n1607_), .ZN(new_n1781_));
  OAI21_X1   g1139(.A1(new_n1780_), .A2(new_n1138_), .B(new_n1781_), .ZN(new_n1782_));
  NOR2_X1    g1140(.A1(new_n1782_), .A2(new_n1613_), .ZN(new_n1783_));
  NAND3_X1   g1141(.A1(new_n1133_), .A2(\in1[0] ), .A3(new_n1783_), .ZN(new_n1784_));
  INV_X1     g1142(.I(\in1[0] ), .ZN(new_n1785_));
  NAND3_X1   g1143(.A1(new_n1133_), .A2(new_n1785_), .A3(new_n1615_), .ZN(new_n1786_));
  AOI21_X1   g1144(.A1(new_n1784_), .A2(new_n1786_), .B(new_n1770_), .ZN(new_n1787_));
  NAND4_X1   g1145(.A1(new_n1129_), .A2(\in2[2] ), .A3(\in3[2] ), .A4(new_n644_), .ZN(new_n1788_));
  NAND4_X1   g1146(.A1(new_n1129_), .A2(new_n688_), .A3(new_n689_), .A4(new_n644_), .ZN(new_n1789_));
  NAND2_X1   g1147(.A1(new_n1788_), .A2(new_n1789_), .ZN(new_n1790_));
  NAND3_X1   g1148(.A1(new_n1790_), .A2(\in1[2] ), .A3(new_n1783_), .ZN(new_n1791_));
  NAND4_X1   g1149(.A1(new_n1783_), .A2(new_n1788_), .A3(new_n1789_), .A4(new_n1181_), .ZN(new_n1792_));
  AOI21_X1   g1150(.A1(new_n1791_), .A2(new_n1792_), .B(new_n1180_), .ZN(new_n1793_));
  AOI21_X1   g1151(.A1(new_n1787_), .A2(new_n1793_), .B(new_n1769_), .ZN(new_n1794_));
  AND2_X2    g1152(.A1(new_n1788_), .A2(new_n1789_), .Z(new_n1795_));
  NOR4_X1    g1153(.A1(new_n1740_), .A2(new_n1764_), .A3(new_n1760_), .A4(new_n1763_), .ZN(new_n1796_));
  INV_X1     g1154(.I(\in3[1] ), .ZN(new_n1797_));
  AOI21_X1   g1155(.A1(new_n1129_), .A2(new_n1762_), .B(\in2[1] ), .ZN(new_n1798_));
  AOI21_X1   g1156(.A1(new_n1652_), .A2(new_n1797_), .B(new_n1798_), .ZN(new_n1799_));
  NAND3_X1   g1157(.A1(new_n1608_), .A2(new_n1181_), .A3(new_n1614_), .ZN(new_n1800_));
  OAI21_X1   g1158(.A1(new_n1782_), .A2(new_n1613_), .B(new_n1180_), .ZN(new_n1801_));
  NAND2_X1   g1159(.A1(new_n1801_), .A2(new_n1800_), .ZN(new_n1802_));
  NOR4_X1    g1160(.A1(new_n1796_), .A2(new_n1795_), .A3(new_n1802_), .A4(new_n1799_), .ZN(new_n1803_));
  OAI21_X1   g1161(.A1(new_n1787_), .A2(new_n1793_), .B(new_n1803_), .ZN(new_n1804_));
  OAI21_X1   g1162(.A1(new_n1794_), .A2(new_n1804_), .B(new_n1766_), .ZN(new_n1805_));
  NAND2_X1   g1163(.A1(new_n1738_), .A2(new_n1735_), .ZN(new_n1806_));
  AOI21_X1   g1164(.A1(new_n1805_), .A2(new_n1806_), .B(new_n1739_), .ZN(new_n1807_));
  NOR2_X1    g1165(.A1(new_n1732_), .A2(new_n1728_), .ZN(new_n1808_));
  OAI21_X1   g1166(.A1(new_n1807_), .A2(new_n1808_), .B(new_n1733_), .ZN(new_n1809_));
  NAND2_X1   g1167(.A1(new_n1615_), .A2(new_n1172_), .ZN(new_n1810_));
  OAI21_X1   g1168(.A1(\in1[6] ), .A2(new_n1615_), .B(new_n1810_), .ZN(new_n1811_));
  NAND2_X1   g1169(.A1(new_n1652_), .A2(new_n703_), .ZN(new_n1812_));
  OAI21_X1   g1170(.A1(\in2[6] ), .A2(new_n1652_), .B(new_n1812_), .ZN(new_n1813_));
  INV_X1     g1171(.I(new_n1723_), .ZN(new_n1814_));
  NOR2_X1    g1172(.A1(new_n1814_), .A2(new_n1719_), .ZN(new_n1815_));
  AOI21_X1   g1173(.A1(new_n1815_), .A2(new_n1813_), .B(new_n1811_), .ZN(new_n1816_));
  NOR2_X1    g1174(.A1(new_n1724_), .A2(new_n1717_), .ZN(new_n1817_));
  NOR2_X1    g1175(.A1(new_n1815_), .A2(new_n1813_), .ZN(new_n1818_));
  INV_X1     g1176(.I(\in0[8] ), .ZN(new_n1819_));
  NAND2_X1   g1177(.A1(new_n1615_), .A2(new_n1819_), .ZN(new_n1820_));
  OAI21_X1   g1178(.A1(\in1[8] ), .A2(new_n1615_), .B(new_n1820_), .ZN(new_n1821_));
  INV_X1     g1179(.I(new_n1821_), .ZN(new_n1822_));
  NOR4_X1    g1180(.A1(new_n1816_), .A2(new_n1817_), .A3(new_n1818_), .A4(new_n1822_), .ZN(new_n1823_));
  NAND2_X1   g1181(.A1(new_n1809_), .A2(new_n1823_), .ZN(new_n1824_));
  INV_X1     g1182(.I(\in0[9] ), .ZN(new_n1825_));
  NOR2_X1    g1183(.A1(new_n1615_), .A2(\in1[9] ), .ZN(new_n1826_));
  AOI21_X1   g1184(.A1(new_n1825_), .A2(new_n1615_), .B(new_n1826_), .ZN(new_n1827_));
  INV_X1     g1185(.I(\in3[9] ), .ZN(new_n1828_));
  NOR2_X1    g1186(.A1(new_n1652_), .A2(\in2[9] ), .ZN(new_n1829_));
  AOI21_X1   g1187(.A1(new_n1828_), .A2(new_n1652_), .B(new_n1829_), .ZN(new_n1830_));
  NOR2_X1    g1188(.A1(new_n1652_), .A2(\in2[10] ), .ZN(new_n1831_));
  AOI21_X1   g1189(.A1(new_n713_), .A2(new_n1652_), .B(new_n1831_), .ZN(new_n1832_));
  NAND2_X1   g1190(.A1(new_n1615_), .A2(new_n1166_), .ZN(new_n1833_));
  OAI21_X1   g1191(.A1(\in1[10] ), .A2(new_n1615_), .B(new_n1833_), .ZN(new_n1834_));
  NAND2_X1   g1192(.A1(new_n1834_), .A2(new_n1832_), .ZN(new_n1835_));
  OAI21_X1   g1193(.A1(new_n1835_), .A2(new_n1830_), .B(new_n1827_), .ZN(new_n1836_));
  INV_X1     g1194(.I(new_n1714_), .ZN(new_n1837_));
  NOR2_X1    g1195(.A1(new_n1837_), .A2(new_n1710_), .ZN(new_n1838_));
  NOR4_X1    g1196(.A1(new_n1838_), .A2(new_n1830_), .A3(new_n1832_), .A4(new_n1834_), .ZN(new_n1839_));
  NAND2_X1   g1197(.A1(new_n1839_), .A2(new_n1836_), .ZN(new_n1840_));
  AOI21_X1   g1198(.A1(new_n1824_), .A2(new_n1725_), .B(new_n1840_), .ZN(new_n1841_));
  INV_X1     g1199(.I(\in0[12] ), .ZN(new_n1842_));
  NOR2_X1    g1200(.A1(new_n1615_), .A2(\in1[12] ), .ZN(new_n1843_));
  AOI21_X1   g1201(.A1(new_n1842_), .A2(new_n1615_), .B(new_n1843_), .ZN(new_n1844_));
  INV_X1     g1202(.I(\in3[12] ), .ZN(new_n1845_));
  NOR2_X1    g1203(.A1(new_n1652_), .A2(\in2[12] ), .ZN(new_n1846_));
  AOI21_X1   g1204(.A1(new_n1845_), .A2(new_n1652_), .B(new_n1846_), .ZN(new_n1847_));
  INV_X1     g1205(.I(new_n1847_), .ZN(new_n1848_));
  NOR2_X1    g1206(.A1(new_n1652_), .A2(\in2[13] ), .ZN(new_n1849_));
  AOI21_X1   g1207(.A1(new_n721_), .A2(new_n1652_), .B(new_n1849_), .ZN(new_n1850_));
  NOR2_X1    g1208(.A1(new_n1615_), .A2(\in1[13] ), .ZN(new_n1851_));
  AOI21_X1   g1209(.A1(new_n1162_), .A2(new_n1615_), .B(new_n1851_), .ZN(new_n1852_));
  INV_X1     g1210(.I(new_n1852_), .ZN(new_n1853_));
  NAND3_X1   g1211(.A1(new_n1853_), .A2(new_n1848_), .A3(new_n1850_), .ZN(new_n1854_));
  INV_X1     g1212(.I(new_n1850_), .ZN(new_n1855_));
  NAND2_X1   g1213(.A1(new_n1702_), .A2(new_n1706_), .ZN(new_n1856_));
  NAND4_X1   g1214(.A1(new_n1856_), .A2(new_n1848_), .A3(new_n1855_), .A4(new_n1852_), .ZN(new_n1857_));
  AOI21_X1   g1215(.A1(new_n1854_), .A2(new_n1844_), .B(new_n1857_), .ZN(new_n1858_));
  OAI21_X1   g1216(.A1(new_n1841_), .A2(new_n1715_), .B(new_n1858_), .ZN(new_n1859_));
  INV_X1     g1217(.I(new_n1699_), .ZN(new_n1860_));
  NOR2_X1    g1218(.A1(new_n1860_), .A2(new_n1696_), .ZN(new_n1861_));
  AOI21_X1   g1219(.A1(new_n1859_), .A2(new_n1708_), .B(new_n1861_), .ZN(new_n1862_));
  INV_X1     g1220(.I(new_n1690_), .ZN(new_n1863_));
  NAND2_X1   g1221(.A1(new_n1863_), .A2(new_n1692_), .ZN(new_n1864_));
  OAI21_X1   g1222(.A1(new_n1862_), .A2(new_n1700_), .B(new_n1864_), .ZN(new_n1865_));
  INV_X1     g1223(.I(\in0[17] ), .ZN(new_n1866_));
  NOR2_X1    g1224(.A1(new_n1615_), .A2(\in1[17] ), .ZN(new_n1867_));
  AOI21_X1   g1225(.A1(new_n1866_), .A2(new_n1615_), .B(new_n1867_), .ZN(new_n1868_));
  INV_X1     g1226(.I(new_n1868_), .ZN(new_n1869_));
  INV_X1     g1227(.I(\in3[17] ), .ZN(new_n1870_));
  NOR2_X1    g1228(.A1(new_n1652_), .A2(\in2[17] ), .ZN(new_n1871_));
  AOI21_X1   g1229(.A1(new_n1870_), .A2(new_n1652_), .B(new_n1871_), .ZN(new_n1872_));
  NOR2_X1    g1230(.A1(new_n1652_), .A2(\in2[18] ), .ZN(new_n1873_));
  AOI21_X1   g1231(.A1(new_n733_), .A2(new_n1652_), .B(new_n1873_), .ZN(new_n1874_));
  INV_X1     g1232(.I(new_n1874_), .ZN(new_n1875_));
  NOR2_X1    g1233(.A1(new_n1615_), .A2(\in1[18] ), .ZN(new_n1876_));
  AOI21_X1   g1234(.A1(new_n1153_), .A2(new_n1615_), .B(new_n1876_), .ZN(new_n1877_));
  NOR3_X1    g1235(.A1(new_n1875_), .A2(new_n1872_), .A3(new_n1877_), .ZN(new_n1878_));
  INV_X1     g1236(.I(new_n1877_), .ZN(new_n1879_));
  INV_X1     g1237(.I(new_n1684_), .ZN(new_n1880_));
  INV_X1     g1238(.I(new_n1687_), .ZN(new_n1881_));
  NOR2_X1    g1239(.A1(new_n1880_), .A2(new_n1881_), .ZN(new_n1882_));
  NOR4_X1    g1240(.A1(new_n1882_), .A2(new_n1872_), .A3(new_n1874_), .A4(new_n1879_), .ZN(new_n1883_));
  OAI21_X1   g1241(.A1(new_n1869_), .A2(new_n1878_), .B(new_n1883_), .ZN(new_n1884_));
  AOI21_X1   g1242(.A1(new_n1865_), .A2(new_n1694_), .B(new_n1884_), .ZN(new_n1885_));
  INV_X1     g1243(.I(\in0[20] ), .ZN(new_n1886_));
  NOR2_X1    g1244(.A1(new_n1615_), .A2(\in1[20] ), .ZN(new_n1887_));
  AOI21_X1   g1245(.A1(new_n1886_), .A2(new_n1615_), .B(new_n1887_), .ZN(new_n1888_));
  INV_X1     g1246(.I(\in3[20] ), .ZN(new_n1889_));
  NOR2_X1    g1247(.A1(new_n1652_), .A2(\in2[20] ), .ZN(new_n1890_));
  AOI21_X1   g1248(.A1(new_n1889_), .A2(new_n1652_), .B(new_n1890_), .ZN(new_n1891_));
  INV_X1     g1249(.I(new_n1891_), .ZN(new_n1892_));
  NOR2_X1    g1250(.A1(new_n1652_), .A2(\in2[21] ), .ZN(new_n1893_));
  AOI21_X1   g1251(.A1(new_n741_), .A2(new_n1652_), .B(new_n1893_), .ZN(new_n1894_));
  NOR2_X1    g1252(.A1(new_n1615_), .A2(\in1[21] ), .ZN(new_n1895_));
  AOI21_X1   g1253(.A1(new_n1149_), .A2(new_n1615_), .B(new_n1895_), .ZN(new_n1896_));
  INV_X1     g1254(.I(new_n1896_), .ZN(new_n1897_));
  NAND3_X1   g1255(.A1(new_n1897_), .A2(new_n1892_), .A3(new_n1894_), .ZN(new_n1898_));
  INV_X1     g1256(.I(new_n1894_), .ZN(new_n1899_));
  NAND2_X1   g1257(.A1(new_n1676_), .A2(new_n1680_), .ZN(new_n1900_));
  NAND4_X1   g1258(.A1(new_n1900_), .A2(new_n1892_), .A3(new_n1899_), .A4(new_n1896_), .ZN(new_n1901_));
  AOI21_X1   g1259(.A1(new_n1898_), .A2(new_n1888_), .B(new_n1901_), .ZN(new_n1902_));
  OAI21_X1   g1260(.A1(new_n1885_), .A2(new_n1688_), .B(new_n1902_), .ZN(new_n1903_));
  INV_X1     g1261(.I(new_n1673_), .ZN(new_n1904_));
  NOR2_X1    g1262(.A1(new_n1904_), .A2(new_n1670_), .ZN(new_n1905_));
  AOI21_X1   g1263(.A1(new_n1903_), .A2(new_n1682_), .B(new_n1905_), .ZN(new_n1906_));
  INV_X1     g1264(.I(new_n1664_), .ZN(new_n1907_));
  NAND2_X1   g1265(.A1(new_n1907_), .A2(new_n1666_), .ZN(new_n1908_));
  OAI21_X1   g1266(.A1(new_n1906_), .A2(new_n1674_), .B(new_n1908_), .ZN(new_n1909_));
  INV_X1     g1267(.I(\in0[25] ), .ZN(new_n1910_));
  NOR2_X1    g1268(.A1(new_n1615_), .A2(\in1[25] ), .ZN(new_n1911_));
  AOI21_X1   g1269(.A1(new_n1910_), .A2(new_n1615_), .B(new_n1911_), .ZN(new_n1912_));
  INV_X1     g1270(.I(new_n1912_), .ZN(new_n1913_));
  INV_X1     g1271(.I(\in3[25] ), .ZN(new_n1914_));
  NOR2_X1    g1272(.A1(new_n1652_), .A2(\in2[25] ), .ZN(new_n1915_));
  AOI21_X1   g1273(.A1(new_n1914_), .A2(new_n1652_), .B(new_n1915_), .ZN(new_n1916_));
  NOR2_X1    g1274(.A1(new_n1652_), .A2(\in2[26] ), .ZN(new_n1917_));
  AOI21_X1   g1275(.A1(new_n753_), .A2(new_n1652_), .B(new_n1917_), .ZN(new_n1918_));
  INV_X1     g1276(.I(new_n1918_), .ZN(new_n1919_));
  NOR2_X1    g1277(.A1(new_n1615_), .A2(\in1[26] ), .ZN(new_n1920_));
  AOI21_X1   g1278(.A1(new_n1140_), .A2(new_n1615_), .B(new_n1920_), .ZN(new_n1921_));
  NOR3_X1    g1279(.A1(new_n1919_), .A2(new_n1916_), .A3(new_n1921_), .ZN(new_n1922_));
  INV_X1     g1280(.I(new_n1921_), .ZN(new_n1923_));
  INV_X1     g1281(.I(new_n1658_), .ZN(new_n1924_));
  INV_X1     g1282(.I(new_n1661_), .ZN(new_n1925_));
  NOR2_X1    g1283(.A1(new_n1924_), .A2(new_n1925_), .ZN(new_n1926_));
  NOR4_X1    g1284(.A1(new_n1926_), .A2(new_n1916_), .A3(new_n1918_), .A4(new_n1923_), .ZN(new_n1927_));
  OAI21_X1   g1285(.A1(new_n1913_), .A2(new_n1922_), .B(new_n1927_), .ZN(new_n1928_));
  AOI21_X1   g1286(.A1(new_n1909_), .A2(new_n1668_), .B(new_n1928_), .ZN(new_n1929_));
  INV_X1     g1287(.I(\in0[28] ), .ZN(new_n1930_));
  NOR2_X1    g1288(.A1(new_n1615_), .A2(\in1[28] ), .ZN(new_n1931_));
  AOI21_X1   g1289(.A1(new_n1930_), .A2(new_n1615_), .B(new_n1931_), .ZN(new_n1932_));
  INV_X1     g1290(.I(\in3[28] ), .ZN(new_n1933_));
  NOR2_X1    g1291(.A1(new_n1652_), .A2(\in2[28] ), .ZN(new_n1934_));
  AOI21_X1   g1292(.A1(new_n1933_), .A2(new_n1652_), .B(new_n1934_), .ZN(new_n1935_));
  INV_X1     g1293(.I(new_n1935_), .ZN(new_n1936_));
  NOR2_X1    g1294(.A1(new_n1652_), .A2(\in2[29] ), .ZN(new_n1937_));
  AOI21_X1   g1295(.A1(new_n761_), .A2(new_n1652_), .B(new_n1937_), .ZN(new_n1938_));
  NOR2_X1    g1296(.A1(new_n1615_), .A2(\in1[29] ), .ZN(new_n1939_));
  AOI21_X1   g1297(.A1(new_n1136_), .A2(new_n1615_), .B(new_n1939_), .ZN(new_n1940_));
  INV_X1     g1298(.I(new_n1940_), .ZN(new_n1941_));
  NAND3_X1   g1299(.A1(new_n1941_), .A2(new_n1936_), .A3(new_n1938_), .ZN(new_n1942_));
  INV_X1     g1300(.I(new_n1938_), .ZN(new_n1943_));
  NAND2_X1   g1301(.A1(new_n1617_), .A2(new_n1654_), .ZN(new_n1944_));
  NAND4_X1   g1302(.A1(new_n1944_), .A2(new_n1936_), .A3(new_n1943_), .A4(new_n1940_), .ZN(new_n1945_));
  AOI21_X1   g1303(.A1(new_n1942_), .A2(new_n1932_), .B(new_n1945_), .ZN(new_n1946_));
  OAI21_X1   g1304(.A1(new_n1929_), .A2(new_n1662_), .B(new_n1946_), .ZN(new_n1947_));
  NOR2_X1    g1305(.A1(new_n1652_), .A2(\in2[51] ), .ZN(new_n1948_));
  AOI21_X1   g1306(.A1(new_n1108_), .A2(new_n1652_), .B(new_n1948_), .ZN(new_n1949_));
  NOR2_X1    g1307(.A1(new_n1615_), .A2(\in1[49] ), .ZN(new_n1950_));
  AOI21_X1   g1308(.A1(new_n1580_), .A2(new_n1615_), .B(new_n1950_), .ZN(new_n1951_));
  NOR2_X1    g1309(.A1(new_n1615_), .A2(\in1[51] ), .ZN(new_n1952_));
  AOI21_X1   g1310(.A1(new_n1588_), .A2(new_n1615_), .B(new_n1952_), .ZN(new_n1953_));
  NOR2_X1    g1311(.A1(new_n1652_), .A2(\in2[49] ), .ZN(new_n1954_));
  AOI21_X1   g1312(.A1(new_n1103_), .A2(new_n1652_), .B(new_n1954_), .ZN(new_n1955_));
  OAI22_X1   g1313(.A1(new_n1949_), .A2(new_n1951_), .B1(new_n1953_), .B2(new_n1955_), .ZN(new_n1956_));
  INV_X1     g1314(.I(\in0[50] ), .ZN(new_n1957_));
  NOR2_X1    g1315(.A1(new_n1615_), .A2(\in1[50] ), .ZN(new_n1958_));
  AOI21_X1   g1316(.A1(new_n1957_), .A2(new_n1615_), .B(new_n1958_), .ZN(new_n1959_));
  NOR2_X1    g1317(.A1(new_n1652_), .A2(\in2[50] ), .ZN(new_n1960_));
  AOI21_X1   g1318(.A1(new_n1107_), .A2(new_n1652_), .B(new_n1960_), .ZN(new_n1961_));
  INV_X1     g1319(.I(new_n1961_), .ZN(new_n1962_));
  OAI21_X1   g1320(.A1(new_n1959_), .A2(new_n1962_), .B(new_n1956_), .ZN(new_n1963_));
  NOR2_X1    g1321(.A1(new_n1652_), .A2(\in2[52] ), .ZN(new_n1964_));
  AOI21_X1   g1322(.A1(new_n1119_), .A2(new_n1652_), .B(new_n1964_), .ZN(new_n1965_));
  INV_X1     g1323(.I(new_n1965_), .ZN(new_n1966_));
  NOR2_X1    g1324(.A1(new_n1615_), .A2(\in1[52] ), .ZN(new_n1967_));
  AOI21_X1   g1325(.A1(new_n1598_), .A2(new_n1615_), .B(new_n1967_), .ZN(new_n1968_));
  NOR2_X1    g1326(.A1(new_n1966_), .A2(new_n1968_), .ZN(new_n1969_));
  INV_X1     g1327(.I(\in3[54] ), .ZN(new_n1970_));
  NOR2_X1    g1328(.A1(new_n1652_), .A2(\in2[54] ), .ZN(new_n1971_));
  AOI21_X1   g1329(.A1(new_n1970_), .A2(new_n1652_), .B(new_n1971_), .ZN(new_n1972_));
  INV_X1     g1330(.I(\in0[55] ), .ZN(new_n1973_));
  NOR2_X1    g1331(.A1(new_n1615_), .A2(\in1[55] ), .ZN(new_n1974_));
  AOI21_X1   g1332(.A1(new_n1973_), .A2(new_n1615_), .B(new_n1974_), .ZN(new_n1975_));
  NOR2_X1    g1333(.A1(new_n1615_), .A2(\in1[54] ), .ZN(new_n1976_));
  AOI21_X1   g1334(.A1(new_n1595_), .A2(new_n1615_), .B(new_n1976_), .ZN(new_n1977_));
  INV_X1     g1335(.I(\in3[55] ), .ZN(new_n1978_));
  NOR2_X1    g1336(.A1(new_n1652_), .A2(\in2[55] ), .ZN(new_n1979_));
  AOI21_X1   g1337(.A1(new_n1978_), .A2(new_n1652_), .B(new_n1979_), .ZN(new_n1980_));
  OAI22_X1   g1338(.A1(new_n1972_), .A2(new_n1975_), .B1(new_n1977_), .B2(new_n1980_), .ZN(new_n1981_));
  NOR2_X1    g1339(.A1(new_n1652_), .A2(\in2[53] ), .ZN(new_n1982_));
  AOI21_X1   g1340(.A1(new_n1093_), .A2(new_n1652_), .B(new_n1982_), .ZN(new_n1983_));
  NOR2_X1    g1341(.A1(new_n1615_), .A2(\in1[53] ), .ZN(new_n1984_));
  AOI21_X1   g1342(.A1(new_n1594_), .A2(new_n1615_), .B(new_n1984_), .ZN(new_n1985_));
  NOR2_X1    g1343(.A1(new_n1985_), .A2(new_n1983_), .ZN(new_n1986_));
  OAI21_X1   g1344(.A1(new_n1981_), .A2(new_n1969_), .B(new_n1986_), .ZN(new_n1987_));
  NAND2_X1   g1345(.A1(new_n1963_), .A2(new_n1987_), .ZN(new_n1988_));
  NOR2_X1    g1346(.A1(new_n1615_), .A2(\in1[48] ), .ZN(new_n1989_));
  AOI21_X1   g1347(.A1(new_n1579_), .A2(new_n1615_), .B(new_n1989_), .ZN(new_n1990_));
  NOR2_X1    g1348(.A1(new_n1652_), .A2(\in2[48] ), .ZN(new_n1991_));
  AOI21_X1   g1349(.A1(new_n1102_), .A2(new_n1652_), .B(new_n1991_), .ZN(new_n1992_));
  NOR2_X1    g1350(.A1(new_n1990_), .A2(new_n1992_), .ZN(new_n1993_));
  INV_X1     g1351(.I(new_n1975_), .ZN(new_n1994_));
  INV_X1     g1352(.I(new_n1985_), .ZN(new_n1995_));
  INV_X1     g1353(.I(new_n1977_), .ZN(new_n1996_));
  NOR2_X1    g1354(.A1(new_n1996_), .A2(new_n1972_), .ZN(new_n1997_));
  NAND2_X1   g1355(.A1(new_n1997_), .A2(new_n1995_), .ZN(new_n1998_));
  NAND2_X1   g1356(.A1(new_n1998_), .A2(new_n1983_), .ZN(new_n1999_));
  INV_X1     g1357(.I(new_n1968_), .ZN(new_n2000_));
  NOR2_X1    g1358(.A1(new_n1997_), .A2(new_n1995_), .ZN(new_n2001_));
  NOR4_X1    g1359(.A1(new_n2001_), .A2(new_n1965_), .A3(new_n2000_), .A4(new_n1980_), .ZN(new_n2002_));
  AOI22_X1   g1360(.A1(new_n2002_), .A2(new_n1999_), .B1(new_n1994_), .B2(new_n1981_), .ZN(new_n2003_));
  NOR2_X1    g1361(.A1(new_n1953_), .A2(new_n1959_), .ZN(new_n2004_));
  NAND2_X1   g1362(.A1(new_n1953_), .A2(new_n1959_), .ZN(new_n2005_));
  NOR2_X1    g1363(.A1(new_n1949_), .A2(new_n1961_), .ZN(new_n2006_));
  AOI21_X1   g1364(.A1(new_n2005_), .A2(new_n2006_), .B(new_n2004_), .ZN(new_n2007_));
  OAI21_X1   g1365(.A1(new_n2003_), .A2(new_n1987_), .B(new_n2007_), .ZN(new_n2008_));
  INV_X1     g1366(.I(new_n1992_), .ZN(new_n2009_));
  INV_X1     g1367(.I(new_n1951_), .ZN(new_n2010_));
  NOR3_X1    g1368(.A1(new_n1963_), .A2(new_n2010_), .A3(new_n1955_), .ZN(new_n2011_));
  NOR2_X1    g1369(.A1(new_n2011_), .A2(new_n2009_), .ZN(new_n2012_));
  INV_X1     g1370(.I(\in3[61] ), .ZN(new_n2013_));
  NOR2_X1    g1371(.A1(new_n1652_), .A2(\in2[61] ), .ZN(new_n2014_));
  AOI21_X1   g1372(.A1(new_n2013_), .A2(new_n1652_), .B(new_n2014_), .ZN(new_n2015_));
  INV_X1     g1373(.I(new_n2015_), .ZN(new_n2016_));
  INV_X1     g1374(.I(\in0[61] ), .ZN(new_n2017_));
  NOR2_X1    g1375(.A1(new_n1615_), .A2(\in1[61] ), .ZN(new_n2018_));
  AOI21_X1   g1376(.A1(new_n2017_), .A2(new_n1615_), .B(new_n2018_), .ZN(new_n2019_));
  INV_X1     g1377(.I(\in3[62] ), .ZN(new_n2020_));
  NOR2_X1    g1378(.A1(new_n1652_), .A2(\in2[62] ), .ZN(new_n2021_));
  AOI21_X1   g1379(.A1(new_n2020_), .A2(new_n1652_), .B(new_n2021_), .ZN(new_n2022_));
  INV_X1     g1380(.I(new_n2022_), .ZN(new_n2023_));
  INV_X1     g1381(.I(\in0[63] ), .ZN(new_n2024_));
  NOR2_X1    g1382(.A1(new_n1615_), .A2(\in1[63] ), .ZN(new_n2025_));
  AOI21_X1   g1383(.A1(new_n2024_), .A2(new_n1615_), .B(new_n2025_), .ZN(new_n2026_));
  INV_X1     g1384(.I(new_n2026_), .ZN(new_n2027_));
  INV_X1     g1385(.I(\in0[62] ), .ZN(new_n2028_));
  NOR2_X1    g1386(.A1(new_n1615_), .A2(\in1[62] ), .ZN(new_n2029_));
  AOI21_X1   g1387(.A1(new_n2028_), .A2(new_n1615_), .B(new_n2029_), .ZN(new_n2030_));
  INV_X1     g1388(.I(new_n2030_), .ZN(new_n2031_));
  INV_X1     g1389(.I(\in3[63] ), .ZN(new_n2032_));
  NOR2_X1    g1390(.A1(new_n1652_), .A2(\in2[63] ), .ZN(new_n2033_));
  AOI21_X1   g1391(.A1(new_n2032_), .A2(new_n1652_), .B(new_n2033_), .ZN(new_n2034_));
  INV_X1     g1392(.I(new_n2034_), .ZN(new_n2035_));
  AOI22_X1   g1393(.A1(new_n2023_), .A2(new_n2027_), .B1(new_n2031_), .B2(new_n2035_), .ZN(new_n2036_));
  OAI21_X1   g1394(.A1(new_n2016_), .A2(new_n2019_), .B(new_n2036_), .ZN(new_n2037_));
  INV_X1     g1395(.I(\in3[60] ), .ZN(new_n2038_));
  NOR2_X1    g1396(.A1(new_n1652_), .A2(\in2[60] ), .ZN(new_n2039_));
  AOI21_X1   g1397(.A1(new_n2038_), .A2(new_n1652_), .B(new_n2039_), .ZN(new_n2040_));
  INV_X1     g1398(.I(new_n2040_), .ZN(new_n2041_));
  INV_X1     g1399(.I(\in0[60] ), .ZN(new_n2042_));
  NOR2_X1    g1400(.A1(new_n1615_), .A2(\in1[60] ), .ZN(new_n2043_));
  AOI21_X1   g1401(.A1(new_n2042_), .A2(new_n1615_), .B(new_n2043_), .ZN(new_n2044_));
  INV_X1     g1402(.I(new_n2044_), .ZN(new_n2045_));
  NAND3_X1   g1403(.A1(new_n2037_), .A2(new_n2041_), .A3(new_n2045_), .ZN(new_n2046_));
  INV_X1     g1404(.I(new_n1990_), .ZN(new_n2047_));
  NOR2_X1    g1405(.A1(new_n1652_), .A2(\in2[58] ), .ZN(new_n2048_));
  AOI21_X1   g1406(.A1(new_n1018_), .A2(new_n1652_), .B(new_n2048_), .ZN(new_n2049_));
  NOR2_X1    g1407(.A1(new_n1615_), .A2(\in1[59] ), .ZN(new_n2050_));
  AOI21_X1   g1408(.A1(new_n1485_), .A2(new_n1615_), .B(new_n2050_), .ZN(new_n2051_));
  INV_X1     g1409(.I(\in0[58] ), .ZN(new_n2052_));
  NOR2_X1    g1410(.A1(new_n1615_), .A2(\in1[58] ), .ZN(new_n2053_));
  AOI21_X1   g1411(.A1(new_n2052_), .A2(new_n1615_), .B(new_n2053_), .ZN(new_n2054_));
  NOR2_X1    g1412(.A1(new_n1652_), .A2(\in2[59] ), .ZN(new_n2055_));
  AOI21_X1   g1413(.A1(new_n1019_), .A2(new_n1652_), .B(new_n2055_), .ZN(new_n2056_));
  OAI22_X1   g1414(.A1(new_n2049_), .A2(new_n2051_), .B1(new_n2054_), .B2(new_n2056_), .ZN(new_n2057_));
  INV_X1     g1415(.I(\in3[56] ), .ZN(new_n2058_));
  NOR2_X1    g1416(.A1(new_n1652_), .A2(\in2[56] ), .ZN(new_n2059_));
  AOI21_X1   g1417(.A1(new_n2058_), .A2(new_n1652_), .B(new_n2059_), .ZN(new_n2060_));
  INV_X1     g1418(.I(\in0[57] ), .ZN(new_n2061_));
  NOR2_X1    g1419(.A1(new_n1615_), .A2(\in1[57] ), .ZN(new_n2062_));
  AOI21_X1   g1420(.A1(new_n2061_), .A2(new_n1615_), .B(new_n2062_), .ZN(new_n2063_));
  INV_X1     g1421(.I(\in0[56] ), .ZN(new_n2064_));
  NOR2_X1    g1422(.A1(new_n1615_), .A2(\in1[56] ), .ZN(new_n2065_));
  AOI21_X1   g1423(.A1(new_n2064_), .A2(new_n1615_), .B(new_n2065_), .ZN(new_n2066_));
  INV_X1     g1424(.I(\in3[57] ), .ZN(new_n2067_));
  NOR2_X1    g1425(.A1(new_n1652_), .A2(\in2[57] ), .ZN(new_n2068_));
  AOI21_X1   g1426(.A1(new_n2067_), .A2(new_n1652_), .B(new_n2068_), .ZN(new_n2069_));
  OAI22_X1   g1427(.A1(new_n2060_), .A2(new_n2063_), .B1(new_n2066_), .B2(new_n2069_), .ZN(new_n2070_));
  NAND3_X1   g1428(.A1(new_n2057_), .A2(new_n2070_), .A3(new_n2047_), .ZN(new_n2071_));
  NOR3_X1    g1429(.A1(new_n2012_), .A2(new_n2046_), .A3(new_n2071_), .ZN(new_n2072_));
  AOI22_X1   g1430(.A1(new_n2008_), .A2(new_n2072_), .B1(new_n1988_), .B2(new_n1993_), .ZN(new_n2073_));
  NOR2_X1    g1431(.A1(new_n1652_), .A2(\in2[117] ), .ZN(new_n2074_));
  AOI21_X1   g1432(.A1(new_n837_), .A2(new_n1652_), .B(new_n2074_), .ZN(new_n2075_));
  INV_X1     g1433(.I(new_n2075_), .ZN(new_n2076_));
  NOR2_X1    g1434(.A1(new_n1615_), .A2(\in1[117] ), .ZN(new_n2077_));
  AOI21_X1   g1435(.A1(new_n1322_), .A2(new_n1615_), .B(new_n2077_), .ZN(new_n2078_));
  INV_X1     g1436(.I(\in3[118] ), .ZN(new_n2079_));
  NOR2_X1    g1437(.A1(new_n1652_), .A2(\in2[118] ), .ZN(new_n2080_));
  AOI21_X1   g1438(.A1(new_n2079_), .A2(new_n1652_), .B(new_n2080_), .ZN(new_n2081_));
  INV_X1     g1439(.I(new_n2081_), .ZN(new_n2082_));
  INV_X1     g1440(.I(\in0[119] ), .ZN(new_n2083_));
  NOR2_X1    g1441(.A1(new_n1615_), .A2(\in1[119] ), .ZN(new_n2084_));
  AOI21_X1   g1442(.A1(new_n2083_), .A2(new_n1615_), .B(new_n2084_), .ZN(new_n2085_));
  INV_X1     g1443(.I(new_n2085_), .ZN(new_n2086_));
  INV_X1     g1444(.I(\in0[118] ), .ZN(new_n2087_));
  NOR2_X1    g1445(.A1(new_n1615_), .A2(\in1[118] ), .ZN(new_n2088_));
  AOI21_X1   g1446(.A1(new_n2087_), .A2(new_n1615_), .B(new_n2088_), .ZN(new_n2089_));
  INV_X1     g1447(.I(new_n2089_), .ZN(new_n2090_));
  INV_X1     g1448(.I(\in3[119] ), .ZN(new_n2091_));
  NOR2_X1    g1449(.A1(new_n1652_), .A2(\in2[119] ), .ZN(new_n2092_));
  AOI21_X1   g1450(.A1(new_n2091_), .A2(new_n1652_), .B(new_n2092_), .ZN(new_n2093_));
  INV_X1     g1451(.I(new_n2093_), .ZN(new_n2094_));
  AOI22_X1   g1452(.A1(new_n2082_), .A2(new_n2086_), .B1(new_n2090_), .B2(new_n2094_), .ZN(new_n2095_));
  OAI21_X1   g1453(.A1(new_n2076_), .A2(new_n2078_), .B(new_n2095_), .ZN(new_n2096_));
  INV_X1     g1454(.I(\in3[116] ), .ZN(new_n2097_));
  NOR2_X1    g1455(.A1(new_n1652_), .A2(\in2[116] ), .ZN(new_n2098_));
  AOI21_X1   g1456(.A1(new_n2097_), .A2(new_n1652_), .B(new_n2098_), .ZN(new_n2099_));
  INV_X1     g1457(.I(new_n2099_), .ZN(new_n2100_));
  INV_X1     g1458(.I(\in0[116] ), .ZN(new_n2101_));
  NOR2_X1    g1459(.A1(new_n1615_), .A2(\in1[116] ), .ZN(new_n2102_));
  AOI21_X1   g1460(.A1(new_n2101_), .A2(new_n1615_), .B(new_n2102_), .ZN(new_n2103_));
  INV_X1     g1461(.I(new_n2103_), .ZN(new_n2104_));
  NAND3_X1   g1462(.A1(new_n2096_), .A2(new_n2100_), .A3(new_n2104_), .ZN(new_n2105_));
  INV_X1     g1463(.I(new_n2078_), .ZN(new_n2106_));
  NOR2_X1    g1464(.A1(new_n2106_), .A2(new_n2104_), .ZN(new_n2107_));
  NOR3_X1    g1465(.A1(new_n2107_), .A2(new_n2075_), .A3(new_n2099_), .ZN(new_n2108_));
  NOR2_X1    g1466(.A1(new_n2078_), .A2(new_n2103_), .ZN(new_n2109_));
  NOR3_X1    g1467(.A1(new_n2108_), .A2(new_n2095_), .A3(new_n2109_), .ZN(new_n2110_));
  NOR2_X1    g1468(.A1(new_n1652_), .A2(\in2[120] ), .ZN(new_n2111_));
  AOI21_X1   g1469(.A1(new_n863_), .A2(new_n1652_), .B(new_n2111_), .ZN(new_n2112_));
  INV_X1     g1470(.I(new_n2112_), .ZN(new_n2113_));
  NOR2_X1    g1471(.A1(new_n1615_), .A2(\in1[120] ), .ZN(new_n2114_));
  AOI21_X1   g1472(.A1(new_n1347_), .A2(new_n1615_), .B(new_n2114_), .ZN(new_n2115_));
  INV_X1     g1473(.I(\in3[122] ), .ZN(new_n2116_));
  NOR2_X1    g1474(.A1(new_n1652_), .A2(\in2[122] ), .ZN(new_n2117_));
  AOI21_X1   g1475(.A1(new_n2116_), .A2(new_n1652_), .B(new_n2117_), .ZN(new_n2118_));
  INV_X1     g1476(.I(new_n2118_), .ZN(new_n2119_));
  NOR2_X1    g1477(.A1(new_n1615_), .A2(\in1[123] ), .ZN(new_n2120_));
  AOI21_X1   g1478(.A1(new_n1352_), .A2(new_n1615_), .B(new_n2120_), .ZN(new_n2121_));
  INV_X1     g1479(.I(new_n2121_), .ZN(new_n2122_));
  INV_X1     g1480(.I(\in0[122] ), .ZN(new_n2123_));
  NOR2_X1    g1481(.A1(new_n1615_), .A2(\in1[122] ), .ZN(new_n2124_));
  AOI21_X1   g1482(.A1(new_n2123_), .A2(new_n1615_), .B(new_n2124_), .ZN(new_n2125_));
  INV_X1     g1483(.I(new_n2125_), .ZN(new_n2126_));
  INV_X1     g1484(.I(\in3[123] ), .ZN(new_n2127_));
  NOR2_X1    g1485(.A1(new_n1652_), .A2(\in2[123] ), .ZN(new_n2128_));
  AOI21_X1   g1486(.A1(new_n2127_), .A2(new_n1652_), .B(new_n2128_), .ZN(new_n2129_));
  INV_X1     g1487(.I(new_n2129_), .ZN(new_n2130_));
  AOI22_X1   g1488(.A1(new_n2119_), .A2(new_n2122_), .B1(new_n2126_), .B2(new_n2130_), .ZN(new_n2131_));
  OAI21_X1   g1489(.A1(new_n2113_), .A2(new_n2115_), .B(new_n2131_), .ZN(new_n2132_));
  NAND2_X1   g1490(.A1(new_n2086_), .A2(new_n2090_), .ZN(new_n2133_));
  NOR2_X1    g1491(.A1(new_n2086_), .A2(new_n2090_), .ZN(new_n2134_));
  NAND2_X1   g1492(.A1(new_n2082_), .A2(new_n2094_), .ZN(new_n2135_));
  OAI21_X1   g1493(.A1(new_n2134_), .A2(new_n2135_), .B(new_n2133_), .ZN(new_n2136_));
  NOR2_X1    g1494(.A1(new_n1652_), .A2(\in2[121] ), .ZN(new_n2137_));
  AOI21_X1   g1495(.A1(new_n842_), .A2(new_n1652_), .B(new_n2137_), .ZN(new_n2138_));
  INV_X1     g1496(.I(new_n2138_), .ZN(new_n2139_));
  INV_X1     g1497(.I(\in0[121] ), .ZN(new_n2140_));
  NOR2_X1    g1498(.A1(new_n1615_), .A2(\in1[121] ), .ZN(new_n2141_));
  AOI21_X1   g1499(.A1(new_n2140_), .A2(new_n1615_), .B(new_n2141_), .ZN(new_n2142_));
  INV_X1     g1500(.I(new_n2142_), .ZN(new_n2143_));
  NAND4_X1   g1501(.A1(new_n2132_), .A2(new_n2136_), .A3(new_n2139_), .A4(new_n2143_), .ZN(new_n2144_));
  OAI21_X1   g1502(.A1(new_n2144_), .A2(new_n2110_), .B(new_n2105_), .ZN(new_n2145_));
  NOR2_X1    g1503(.A1(new_n1652_), .A2(\in2[104] ), .ZN(new_n2146_));
  AOI21_X1   g1504(.A1(new_n795_), .A2(new_n1652_), .B(new_n2146_), .ZN(new_n2147_));
  NOR2_X1    g1505(.A1(new_n1615_), .A2(\in1[104] ), .ZN(new_n2148_));
  AOI21_X1   g1506(.A1(new_n1281_), .A2(new_n1615_), .B(new_n2148_), .ZN(new_n2149_));
  INV_X1     g1507(.I(new_n2149_), .ZN(new_n2150_));
  NOR2_X1    g1508(.A1(new_n1652_), .A2(\in2[106] ), .ZN(new_n2151_));
  AOI21_X1   g1509(.A1(new_n789_), .A2(new_n1652_), .B(new_n2151_), .ZN(new_n2152_));
  INV_X1     g1510(.I(\in0[107] ), .ZN(new_n2153_));
  NOR2_X1    g1511(.A1(new_n1615_), .A2(\in1[107] ), .ZN(new_n2154_));
  AOI21_X1   g1512(.A1(new_n2153_), .A2(new_n1615_), .B(new_n2154_), .ZN(new_n2155_));
  INV_X1     g1513(.I(\in0[106] ), .ZN(new_n2156_));
  NOR2_X1    g1514(.A1(new_n1615_), .A2(\in1[106] ), .ZN(new_n2157_));
  AOI21_X1   g1515(.A1(new_n2156_), .A2(new_n1615_), .B(new_n2157_), .ZN(new_n2158_));
  NOR2_X1    g1516(.A1(new_n1652_), .A2(\in2[107] ), .ZN(new_n2159_));
  AOI21_X1   g1517(.A1(new_n790_), .A2(new_n1652_), .B(new_n2159_), .ZN(new_n2160_));
  OAI22_X1   g1518(.A1(new_n2152_), .A2(new_n2155_), .B1(new_n2158_), .B2(new_n2160_), .ZN(new_n2161_));
  AOI21_X1   g1519(.A1(new_n2147_), .A2(new_n2150_), .B(new_n2161_), .ZN(new_n2162_));
  NOR2_X1    g1520(.A1(new_n1652_), .A2(\in2[105] ), .ZN(new_n2163_));
  AOI21_X1   g1521(.A1(new_n785_), .A2(new_n1652_), .B(new_n2163_), .ZN(new_n2164_));
  INV_X1     g1522(.I(new_n2164_), .ZN(new_n2165_));
  NOR2_X1    g1523(.A1(new_n1615_), .A2(\in1[105] ), .ZN(new_n2166_));
  AOI21_X1   g1524(.A1(new_n1275_), .A2(new_n1615_), .B(new_n2166_), .ZN(new_n2167_));
  INV_X1     g1525(.I(new_n2167_), .ZN(new_n2168_));
  NAND2_X1   g1526(.A1(new_n2168_), .A2(new_n2165_), .ZN(new_n2169_));
  INV_X1     g1527(.I(new_n2155_), .ZN(new_n2170_));
  INV_X1     g1528(.I(new_n2158_), .ZN(new_n2171_));
  NOR2_X1    g1529(.A1(new_n2171_), .A2(new_n2152_), .ZN(new_n2172_));
  NAND2_X1   g1530(.A1(new_n2172_), .A2(new_n2168_), .ZN(new_n2173_));
  NAND2_X1   g1531(.A1(new_n2173_), .A2(new_n2164_), .ZN(new_n2174_));
  NOR2_X1    g1532(.A1(new_n2172_), .A2(new_n2168_), .ZN(new_n2175_));
  NOR4_X1    g1533(.A1(new_n2175_), .A2(new_n2147_), .A3(new_n2150_), .A4(new_n2160_), .ZN(new_n2176_));
  AOI22_X1   g1534(.A1(new_n2176_), .A2(new_n2174_), .B1(new_n2170_), .B2(new_n2161_), .ZN(new_n2177_));
  NOR2_X1    g1535(.A1(new_n1652_), .A2(\in2[109] ), .ZN(new_n2178_));
  AOI21_X1   g1536(.A1(new_n812_), .A2(new_n1652_), .B(new_n2178_), .ZN(new_n2179_));
  INV_X1     g1537(.I(new_n2179_), .ZN(new_n2180_));
  NOR2_X1    g1538(.A1(new_n1615_), .A2(\in1[109] ), .ZN(new_n2181_));
  AOI21_X1   g1539(.A1(new_n1298_), .A2(new_n1615_), .B(new_n2181_), .ZN(new_n2182_));
  NOR2_X1    g1540(.A1(new_n2180_), .A2(new_n2182_), .ZN(new_n2183_));
  INV_X1     g1541(.I(\in3[110] ), .ZN(new_n2184_));
  NOR2_X1    g1542(.A1(new_n1652_), .A2(\in2[110] ), .ZN(new_n2185_));
  AOI21_X1   g1543(.A1(new_n2184_), .A2(new_n1652_), .B(new_n2185_), .ZN(new_n2186_));
  NOR2_X1    g1544(.A1(new_n1615_), .A2(\in1[111] ), .ZN(new_n2187_));
  AOI21_X1   g1545(.A1(new_n1292_), .A2(new_n1615_), .B(new_n2187_), .ZN(new_n2188_));
  INV_X1     g1546(.I(\in0[110] ), .ZN(new_n2189_));
  NOR2_X1    g1547(.A1(new_n1615_), .A2(\in1[110] ), .ZN(new_n2190_));
  AOI21_X1   g1548(.A1(new_n2189_), .A2(new_n1615_), .B(new_n2190_), .ZN(new_n2191_));
  NOR2_X1    g1549(.A1(new_n1652_), .A2(\in2[111] ), .ZN(new_n2192_));
  AOI21_X1   g1550(.A1(new_n806_), .A2(new_n1652_), .B(new_n2192_), .ZN(new_n2193_));
  OAI22_X1   g1551(.A1(new_n2186_), .A2(new_n2188_), .B1(new_n2191_), .B2(new_n2193_), .ZN(new_n2194_));
  INV_X1     g1552(.I(\in3[108] ), .ZN(new_n2195_));
  NOR2_X1    g1553(.A1(new_n1652_), .A2(\in2[108] ), .ZN(new_n2196_));
  AOI21_X1   g1554(.A1(new_n2195_), .A2(new_n1652_), .B(new_n2196_), .ZN(new_n2197_));
  INV_X1     g1555(.I(\in0[108] ), .ZN(new_n2198_));
  NOR2_X1    g1556(.A1(new_n1615_), .A2(\in1[108] ), .ZN(new_n2199_));
  AOI21_X1   g1557(.A1(new_n2198_), .A2(new_n1615_), .B(new_n2199_), .ZN(new_n2200_));
  NOR2_X1    g1558(.A1(new_n2200_), .A2(new_n2197_), .ZN(new_n2201_));
  OAI21_X1   g1559(.A1(new_n2194_), .A2(new_n2183_), .B(new_n2201_), .ZN(new_n2202_));
  OAI22_X1   g1560(.A1(new_n2177_), .A2(new_n2202_), .B1(new_n2162_), .B2(new_n2169_), .ZN(new_n2203_));
  NOR2_X1    g1561(.A1(new_n2188_), .A2(new_n2191_), .ZN(new_n2204_));
  INV_X1     g1562(.I(new_n2188_), .ZN(new_n2205_));
  INV_X1     g1563(.I(new_n2191_), .ZN(new_n2206_));
  NOR2_X1    g1564(.A1(new_n2205_), .A2(new_n2206_), .ZN(new_n2207_));
  NOR3_X1    g1565(.A1(new_n2207_), .A2(new_n2186_), .A3(new_n2193_), .ZN(new_n2208_));
  INV_X1     g1566(.I(new_n2182_), .ZN(new_n2209_));
  INV_X1     g1567(.I(new_n2200_), .ZN(new_n2210_));
  NOR2_X1    g1568(.A1(new_n2209_), .A2(new_n2210_), .ZN(new_n2211_));
  NOR3_X1    g1569(.A1(new_n2211_), .A2(new_n2179_), .A3(new_n2197_), .ZN(new_n2212_));
  OAI21_X1   g1570(.A1(new_n2182_), .A2(new_n2200_), .B(new_n2194_), .ZN(new_n2213_));
  OAI22_X1   g1571(.A1(new_n2212_), .A2(new_n2213_), .B1(new_n2208_), .B2(new_n2204_), .ZN(new_n2214_));
  NOR2_X1    g1572(.A1(new_n1615_), .A2(\in1[115] ), .ZN(new_n2215_));
  AOI21_X1   g1573(.A1(new_n1312_), .A2(new_n1615_), .B(new_n2215_), .ZN(new_n2216_));
  INV_X1     g1574(.I(new_n2216_), .ZN(new_n2217_));
  NOR2_X1    g1575(.A1(new_n1652_), .A2(\in2[114] ), .ZN(new_n2218_));
  AOI21_X1   g1576(.A1(new_n819_), .A2(new_n1652_), .B(new_n2218_), .ZN(new_n2219_));
  INV_X1     g1577(.I(\in0[114] ), .ZN(new_n2220_));
  NOR2_X1    g1578(.A1(new_n1615_), .A2(\in1[114] ), .ZN(new_n2221_));
  AOI21_X1   g1579(.A1(new_n2220_), .A2(new_n1615_), .B(new_n2221_), .ZN(new_n2222_));
  NOR2_X1    g1580(.A1(new_n1652_), .A2(\in2[115] ), .ZN(new_n2223_));
  AOI21_X1   g1581(.A1(new_n820_), .A2(new_n1652_), .B(new_n2223_), .ZN(new_n2224_));
  OAI22_X1   g1582(.A1(new_n2216_), .A2(new_n2219_), .B1(new_n2222_), .B2(new_n2224_), .ZN(new_n2225_));
  NOR2_X1    g1583(.A1(new_n1652_), .A2(\in2[113] ), .ZN(new_n2226_));
  AOI21_X1   g1584(.A1(new_n827_), .A2(new_n1652_), .B(new_n2226_), .ZN(new_n2227_));
  INV_X1     g1585(.I(\in0[113] ), .ZN(new_n2228_));
  NOR2_X1    g1586(.A1(new_n1615_), .A2(\in1[113] ), .ZN(new_n2229_));
  AOI21_X1   g1587(.A1(new_n2228_), .A2(new_n1615_), .B(new_n2229_), .ZN(new_n2230_));
  INV_X1     g1588(.I(new_n2230_), .ZN(new_n2231_));
  INV_X1     g1589(.I(new_n2222_), .ZN(new_n2232_));
  NOR2_X1    g1590(.A1(new_n2232_), .A2(new_n2219_), .ZN(new_n2233_));
  NAND2_X1   g1591(.A1(new_n2233_), .A2(new_n2231_), .ZN(new_n2234_));
  NAND2_X1   g1592(.A1(new_n2234_), .A2(new_n2227_), .ZN(new_n2235_));
  NOR2_X1    g1593(.A1(new_n2233_), .A2(new_n2231_), .ZN(new_n2236_));
  NOR2_X1    g1594(.A1(new_n1652_), .A2(\in2[112] ), .ZN(new_n2237_));
  AOI21_X1   g1595(.A1(new_n823_), .A2(new_n1652_), .B(new_n2237_), .ZN(new_n2238_));
  NOR2_X1    g1596(.A1(new_n1615_), .A2(\in1[112] ), .ZN(new_n2239_));
  AOI21_X1   g1597(.A1(new_n1307_), .A2(new_n1615_), .B(new_n2239_), .ZN(new_n2240_));
  INV_X1     g1598(.I(new_n2240_), .ZN(new_n2241_));
  NOR4_X1    g1599(.A1(new_n2236_), .A2(new_n2224_), .A3(new_n2238_), .A4(new_n2241_), .ZN(new_n2242_));
  AOI22_X1   g1600(.A1(new_n2242_), .A2(new_n2235_), .B1(new_n2217_), .B2(new_n2225_), .ZN(new_n2243_));
  INV_X1     g1601(.I(new_n2238_), .ZN(new_n2244_));
  NOR2_X1    g1602(.A1(new_n2244_), .A2(new_n2240_), .ZN(new_n2245_));
  NOR2_X1    g1603(.A1(new_n2230_), .A2(new_n2227_), .ZN(new_n2246_));
  OAI21_X1   g1604(.A1(new_n2225_), .A2(new_n2245_), .B(new_n2246_), .ZN(new_n2247_));
  OAI21_X1   g1605(.A1(new_n2243_), .A2(new_n2247_), .B(new_n2214_), .ZN(new_n2248_));
  NAND3_X1   g1606(.A1(new_n2203_), .A2(new_n2248_), .A3(new_n2145_), .ZN(new_n2249_));
  NOR2_X1    g1607(.A1(new_n1652_), .A2(\in2[80] ), .ZN(new_n2250_));
  AOI21_X1   g1608(.A1(new_n965_), .A2(new_n1652_), .B(new_n2250_), .ZN(new_n2251_));
  NOR2_X1    g1609(.A1(new_n1615_), .A2(\in1[80] ), .ZN(new_n2252_));
  AOI21_X1   g1610(.A1(new_n1444_), .A2(new_n1615_), .B(new_n2252_), .ZN(new_n2253_));
  INV_X1     g1611(.I(new_n2253_), .ZN(new_n2254_));
  NOR2_X1    g1612(.A1(new_n1652_), .A2(\in2[82] ), .ZN(new_n2255_));
  AOI21_X1   g1613(.A1(new_n959_), .A2(new_n1652_), .B(new_n2255_), .ZN(new_n2256_));
  INV_X1     g1614(.I(\in0[83] ), .ZN(new_n2257_));
  NOR2_X1    g1615(.A1(new_n1615_), .A2(\in1[83] ), .ZN(new_n2258_));
  AOI21_X1   g1616(.A1(new_n2257_), .A2(new_n1615_), .B(new_n2258_), .ZN(new_n2259_));
  INV_X1     g1617(.I(\in0[82] ), .ZN(new_n2260_));
  NOR2_X1    g1618(.A1(new_n1615_), .A2(\in1[82] ), .ZN(new_n2261_));
  AOI21_X1   g1619(.A1(new_n2260_), .A2(new_n1615_), .B(new_n2261_), .ZN(new_n2262_));
  NOR2_X1    g1620(.A1(new_n1652_), .A2(\in2[83] ), .ZN(new_n2263_));
  AOI21_X1   g1621(.A1(new_n960_), .A2(new_n1652_), .B(new_n2263_), .ZN(new_n2264_));
  OAI22_X1   g1622(.A1(new_n2256_), .A2(new_n2259_), .B1(new_n2262_), .B2(new_n2264_), .ZN(new_n2265_));
  AOI21_X1   g1623(.A1(new_n2251_), .A2(new_n2254_), .B(new_n2265_), .ZN(new_n2266_));
  NOR2_X1    g1624(.A1(new_n1652_), .A2(\in2[81] ), .ZN(new_n2267_));
  AOI21_X1   g1625(.A1(new_n955_), .A2(new_n1652_), .B(new_n2267_), .ZN(new_n2268_));
  INV_X1     g1626(.I(new_n2268_), .ZN(new_n2269_));
  NOR2_X1    g1627(.A1(new_n1615_), .A2(\in1[81] ), .ZN(new_n2270_));
  AOI21_X1   g1628(.A1(new_n1438_), .A2(new_n1615_), .B(new_n2270_), .ZN(new_n2271_));
  INV_X1     g1629(.I(new_n2271_), .ZN(new_n2272_));
  NAND2_X1   g1630(.A1(new_n2272_), .A2(new_n2269_), .ZN(new_n2273_));
  INV_X1     g1631(.I(new_n2259_), .ZN(new_n2274_));
  INV_X1     g1632(.I(new_n2262_), .ZN(new_n2275_));
  NOR2_X1    g1633(.A1(new_n2275_), .A2(new_n2256_), .ZN(new_n2276_));
  NAND2_X1   g1634(.A1(new_n2276_), .A2(new_n2272_), .ZN(new_n2277_));
  NAND2_X1   g1635(.A1(new_n2277_), .A2(new_n2268_), .ZN(new_n2278_));
  NOR2_X1    g1636(.A1(new_n2276_), .A2(new_n2272_), .ZN(new_n2279_));
  NOR4_X1    g1637(.A1(new_n2279_), .A2(new_n2251_), .A3(new_n2254_), .A4(new_n2264_), .ZN(new_n2280_));
  AOI22_X1   g1638(.A1(new_n2280_), .A2(new_n2278_), .B1(new_n2274_), .B2(new_n2265_), .ZN(new_n2281_));
  NOR2_X1    g1639(.A1(new_n1652_), .A2(\in2[85] ), .ZN(new_n2282_));
  AOI21_X1   g1640(.A1(new_n982_), .A2(new_n1652_), .B(new_n2282_), .ZN(new_n2283_));
  INV_X1     g1641(.I(new_n2283_), .ZN(new_n2284_));
  NOR2_X1    g1642(.A1(new_n1615_), .A2(\in1[85] ), .ZN(new_n2285_));
  AOI21_X1   g1643(.A1(new_n1461_), .A2(new_n1615_), .B(new_n2285_), .ZN(new_n2286_));
  NOR2_X1    g1644(.A1(new_n2284_), .A2(new_n2286_), .ZN(new_n2287_));
  INV_X1     g1645(.I(\in3[86] ), .ZN(new_n2288_));
  NOR2_X1    g1646(.A1(new_n1652_), .A2(\in2[86] ), .ZN(new_n2289_));
  AOI21_X1   g1647(.A1(new_n2288_), .A2(new_n1652_), .B(new_n2289_), .ZN(new_n2290_));
  NOR2_X1    g1648(.A1(new_n1615_), .A2(\in1[87] ), .ZN(new_n2291_));
  AOI21_X1   g1649(.A1(new_n1455_), .A2(new_n1615_), .B(new_n2291_), .ZN(new_n2292_));
  INV_X1     g1650(.I(\in0[86] ), .ZN(new_n2293_));
  NOR2_X1    g1651(.A1(new_n1615_), .A2(\in1[86] ), .ZN(new_n2294_));
  AOI21_X1   g1652(.A1(new_n2293_), .A2(new_n1615_), .B(new_n2294_), .ZN(new_n2295_));
  NOR2_X1    g1653(.A1(new_n1652_), .A2(\in2[87] ), .ZN(new_n2296_));
  AOI21_X1   g1654(.A1(new_n976_), .A2(new_n1652_), .B(new_n2296_), .ZN(new_n2297_));
  OAI22_X1   g1655(.A1(new_n2290_), .A2(new_n2292_), .B1(new_n2295_), .B2(new_n2297_), .ZN(new_n2298_));
  INV_X1     g1656(.I(\in3[84] ), .ZN(new_n2299_));
  NOR2_X1    g1657(.A1(new_n1652_), .A2(\in2[84] ), .ZN(new_n2300_));
  AOI21_X1   g1658(.A1(new_n2299_), .A2(new_n1652_), .B(new_n2300_), .ZN(new_n2301_));
  INV_X1     g1659(.I(\in0[84] ), .ZN(new_n2302_));
  NOR2_X1    g1660(.A1(new_n1615_), .A2(\in1[84] ), .ZN(new_n2303_));
  AOI21_X1   g1661(.A1(new_n2302_), .A2(new_n1615_), .B(new_n2303_), .ZN(new_n2304_));
  NOR2_X1    g1662(.A1(new_n2304_), .A2(new_n2301_), .ZN(new_n2305_));
  OAI21_X1   g1663(.A1(new_n2298_), .A2(new_n2287_), .B(new_n2305_), .ZN(new_n2306_));
  OAI22_X1   g1664(.A1(new_n2281_), .A2(new_n2306_), .B1(new_n2266_), .B2(new_n2273_), .ZN(new_n2307_));
  NOR2_X1    g1665(.A1(new_n2292_), .A2(new_n2295_), .ZN(new_n2308_));
  INV_X1     g1666(.I(new_n2292_), .ZN(new_n2309_));
  INV_X1     g1667(.I(new_n2295_), .ZN(new_n2310_));
  NOR2_X1    g1668(.A1(new_n2309_), .A2(new_n2310_), .ZN(new_n2311_));
  NOR3_X1    g1669(.A1(new_n2311_), .A2(new_n2290_), .A3(new_n2297_), .ZN(new_n2312_));
  INV_X1     g1670(.I(new_n2286_), .ZN(new_n2313_));
  INV_X1     g1671(.I(new_n2304_), .ZN(new_n2314_));
  NOR2_X1    g1672(.A1(new_n2313_), .A2(new_n2314_), .ZN(new_n2315_));
  NOR3_X1    g1673(.A1(new_n2315_), .A2(new_n2283_), .A3(new_n2301_), .ZN(new_n2316_));
  OAI21_X1   g1674(.A1(new_n2286_), .A2(new_n2304_), .B(new_n2298_), .ZN(new_n2317_));
  OAI22_X1   g1675(.A1(new_n2316_), .A2(new_n2317_), .B1(new_n2312_), .B2(new_n2308_), .ZN(new_n2318_));
  NOR2_X1    g1676(.A1(new_n1615_), .A2(\in1[91] ), .ZN(new_n2319_));
  AOI21_X1   g1677(.A1(new_n1475_), .A2(new_n1615_), .B(new_n2319_), .ZN(new_n2320_));
  INV_X1     g1678(.I(new_n2320_), .ZN(new_n2321_));
  NOR2_X1    g1679(.A1(new_n1652_), .A2(\in2[90] ), .ZN(new_n2322_));
  AOI21_X1   g1680(.A1(new_n989_), .A2(new_n1652_), .B(new_n2322_), .ZN(new_n2323_));
  INV_X1     g1681(.I(\in0[90] ), .ZN(new_n2324_));
  NOR2_X1    g1682(.A1(new_n1615_), .A2(\in1[90] ), .ZN(new_n2325_));
  AOI21_X1   g1683(.A1(new_n2324_), .A2(new_n1615_), .B(new_n2325_), .ZN(new_n2326_));
  NOR2_X1    g1684(.A1(new_n1652_), .A2(\in2[91] ), .ZN(new_n2327_));
  AOI21_X1   g1685(.A1(new_n990_), .A2(new_n1652_), .B(new_n2327_), .ZN(new_n2328_));
  OAI22_X1   g1686(.A1(new_n2320_), .A2(new_n2323_), .B1(new_n2326_), .B2(new_n2328_), .ZN(new_n2329_));
  NOR2_X1    g1687(.A1(new_n1652_), .A2(\in2[89] ), .ZN(new_n2330_));
  AOI21_X1   g1688(.A1(new_n997_), .A2(new_n1652_), .B(new_n2330_), .ZN(new_n2331_));
  INV_X1     g1689(.I(\in0[89] ), .ZN(new_n2332_));
  NOR2_X1    g1690(.A1(new_n1615_), .A2(\in1[89] ), .ZN(new_n2333_));
  AOI21_X1   g1691(.A1(new_n2332_), .A2(new_n1615_), .B(new_n2333_), .ZN(new_n2334_));
  INV_X1     g1692(.I(new_n2334_), .ZN(new_n2335_));
  INV_X1     g1693(.I(new_n2326_), .ZN(new_n2336_));
  NOR2_X1    g1694(.A1(new_n2336_), .A2(new_n2323_), .ZN(new_n2337_));
  NAND2_X1   g1695(.A1(new_n2337_), .A2(new_n2335_), .ZN(new_n2338_));
  NAND2_X1   g1696(.A1(new_n2338_), .A2(new_n2331_), .ZN(new_n2339_));
  NOR2_X1    g1697(.A1(new_n2337_), .A2(new_n2335_), .ZN(new_n2340_));
  NOR2_X1    g1698(.A1(new_n1652_), .A2(\in2[88] ), .ZN(new_n2341_));
  AOI21_X1   g1699(.A1(new_n993_), .A2(new_n1652_), .B(new_n2341_), .ZN(new_n2342_));
  NOR2_X1    g1700(.A1(new_n1615_), .A2(\in1[88] ), .ZN(new_n2343_));
  AOI21_X1   g1701(.A1(new_n1470_), .A2(new_n1615_), .B(new_n2343_), .ZN(new_n2344_));
  INV_X1     g1702(.I(new_n2344_), .ZN(new_n2345_));
  NOR4_X1    g1703(.A1(new_n2340_), .A2(new_n2328_), .A3(new_n2342_), .A4(new_n2345_), .ZN(new_n2346_));
  AOI22_X1   g1704(.A1(new_n2346_), .A2(new_n2339_), .B1(new_n2321_), .B2(new_n2329_), .ZN(new_n2347_));
  INV_X1     g1705(.I(new_n2342_), .ZN(new_n2348_));
  NOR2_X1    g1706(.A1(new_n2348_), .A2(new_n2344_), .ZN(new_n2349_));
  NOR2_X1    g1707(.A1(new_n2334_), .A2(new_n2331_), .ZN(new_n2350_));
  OAI21_X1   g1708(.A1(new_n2329_), .A2(new_n2349_), .B(new_n2350_), .ZN(new_n2351_));
  OAI21_X1   g1709(.A1(new_n2347_), .A2(new_n2351_), .B(new_n2318_), .ZN(new_n2352_));
  NOR2_X1    g1710(.A1(new_n1652_), .A2(\in2[93] ), .ZN(new_n2353_));
  AOI21_X1   g1711(.A1(new_n771_), .A2(new_n1652_), .B(new_n2353_), .ZN(new_n2354_));
  INV_X1     g1712(.I(new_n2354_), .ZN(new_n2355_));
  NOR2_X1    g1713(.A1(new_n1615_), .A2(\in1[93] ), .ZN(new_n2356_));
  AOI21_X1   g1714(.A1(new_n1260_), .A2(new_n1615_), .B(new_n2356_), .ZN(new_n2357_));
  INV_X1     g1715(.I(\in3[94] ), .ZN(new_n2358_));
  NOR2_X1    g1716(.A1(new_n1652_), .A2(\in2[94] ), .ZN(new_n2359_));
  AOI21_X1   g1717(.A1(new_n2358_), .A2(new_n1652_), .B(new_n2359_), .ZN(new_n2360_));
  INV_X1     g1718(.I(new_n2360_), .ZN(new_n2361_));
  INV_X1     g1719(.I(\in0[95] ), .ZN(new_n2362_));
  NOR2_X1    g1720(.A1(new_n1615_), .A2(\in1[95] ), .ZN(new_n2363_));
  AOI21_X1   g1721(.A1(new_n2362_), .A2(new_n1615_), .B(new_n2363_), .ZN(new_n2364_));
  INV_X1     g1722(.I(new_n2364_), .ZN(new_n2365_));
  INV_X1     g1723(.I(\in0[94] ), .ZN(new_n2366_));
  NOR2_X1    g1724(.A1(new_n1615_), .A2(\in1[94] ), .ZN(new_n2367_));
  AOI21_X1   g1725(.A1(new_n2366_), .A2(new_n1615_), .B(new_n2367_), .ZN(new_n2368_));
  INV_X1     g1726(.I(new_n2368_), .ZN(new_n2369_));
  INV_X1     g1727(.I(\in3[95] ), .ZN(new_n2370_));
  NOR2_X1    g1728(.A1(new_n1652_), .A2(\in2[95] ), .ZN(new_n2371_));
  AOI21_X1   g1729(.A1(new_n2370_), .A2(new_n1652_), .B(new_n2371_), .ZN(new_n2372_));
  INV_X1     g1730(.I(new_n2372_), .ZN(new_n2373_));
  AOI22_X1   g1731(.A1(new_n2361_), .A2(new_n2365_), .B1(new_n2369_), .B2(new_n2373_), .ZN(new_n2374_));
  OAI21_X1   g1732(.A1(new_n2355_), .A2(new_n2357_), .B(new_n2374_), .ZN(new_n2375_));
  INV_X1     g1733(.I(\in3[92] ), .ZN(new_n2376_));
  NOR2_X1    g1734(.A1(new_n1652_), .A2(\in2[92] ), .ZN(new_n2377_));
  AOI21_X1   g1735(.A1(new_n2376_), .A2(new_n1652_), .B(new_n2377_), .ZN(new_n2378_));
  INV_X1     g1736(.I(new_n2378_), .ZN(new_n2379_));
  INV_X1     g1737(.I(\in0[92] ), .ZN(new_n2380_));
  NOR2_X1    g1738(.A1(new_n1615_), .A2(\in1[92] ), .ZN(new_n2381_));
  AOI21_X1   g1739(.A1(new_n2380_), .A2(new_n1615_), .B(new_n2381_), .ZN(new_n2382_));
  INV_X1     g1740(.I(new_n2382_), .ZN(new_n2383_));
  NAND3_X1   g1741(.A1(new_n2375_), .A2(new_n2379_), .A3(new_n2383_), .ZN(new_n2384_));
  INV_X1     g1742(.I(new_n2357_), .ZN(new_n2385_));
  NOR2_X1    g1743(.A1(new_n2385_), .A2(new_n2383_), .ZN(new_n2386_));
  NOR3_X1    g1744(.A1(new_n2386_), .A2(new_n2354_), .A3(new_n2378_), .ZN(new_n2387_));
  NOR2_X1    g1745(.A1(new_n2357_), .A2(new_n2382_), .ZN(new_n2388_));
  NOR3_X1    g1746(.A1(new_n2387_), .A2(new_n2374_), .A3(new_n2388_), .ZN(new_n2389_));
  NOR2_X1    g1747(.A1(new_n1652_), .A2(\in2[96] ), .ZN(new_n2390_));
  AOI21_X1   g1748(.A1(new_n911_), .A2(new_n1652_), .B(new_n2390_), .ZN(new_n2391_));
  INV_X1     g1749(.I(new_n2391_), .ZN(new_n2392_));
  NOR2_X1    g1750(.A1(new_n1615_), .A2(\in1[96] ), .ZN(new_n2393_));
  AOI21_X1   g1751(.A1(new_n1395_), .A2(new_n1615_), .B(new_n2393_), .ZN(new_n2394_));
  INV_X1     g1752(.I(\in3[98] ), .ZN(new_n2395_));
  NOR2_X1    g1753(.A1(new_n1652_), .A2(\in2[98] ), .ZN(new_n2396_));
  AOI21_X1   g1754(.A1(new_n2395_), .A2(new_n1652_), .B(new_n2396_), .ZN(new_n2397_));
  INV_X1     g1755(.I(new_n2397_), .ZN(new_n2398_));
  NOR2_X1    g1756(.A1(new_n1615_), .A2(\in1[99] ), .ZN(new_n2399_));
  AOI21_X1   g1757(.A1(new_n1400_), .A2(new_n1615_), .B(new_n2399_), .ZN(new_n2400_));
  INV_X1     g1758(.I(new_n2400_), .ZN(new_n2401_));
  INV_X1     g1759(.I(\in0[98] ), .ZN(new_n2402_));
  NOR2_X1    g1760(.A1(new_n1615_), .A2(\in1[98] ), .ZN(new_n2403_));
  AOI21_X1   g1761(.A1(new_n2402_), .A2(new_n1615_), .B(new_n2403_), .ZN(new_n2404_));
  INV_X1     g1762(.I(new_n2404_), .ZN(new_n2405_));
  INV_X1     g1763(.I(\in3[99] ), .ZN(new_n2406_));
  NOR2_X1    g1764(.A1(new_n1652_), .A2(\in2[99] ), .ZN(new_n2407_));
  AOI21_X1   g1765(.A1(new_n2406_), .A2(new_n1652_), .B(new_n2407_), .ZN(new_n2408_));
  INV_X1     g1766(.I(new_n2408_), .ZN(new_n2409_));
  AOI22_X1   g1767(.A1(new_n2398_), .A2(new_n2401_), .B1(new_n2405_), .B2(new_n2409_), .ZN(new_n2410_));
  OAI21_X1   g1768(.A1(new_n2392_), .A2(new_n2394_), .B(new_n2410_), .ZN(new_n2411_));
  NAND2_X1   g1769(.A1(new_n2365_), .A2(new_n2369_), .ZN(new_n2412_));
  NOR2_X1    g1770(.A1(new_n2365_), .A2(new_n2369_), .ZN(new_n2413_));
  NAND2_X1   g1771(.A1(new_n2361_), .A2(new_n2373_), .ZN(new_n2414_));
  OAI21_X1   g1772(.A1(new_n2413_), .A2(new_n2414_), .B(new_n2412_), .ZN(new_n2415_));
  NOR2_X1    g1773(.A1(new_n1652_), .A2(\in2[97] ), .ZN(new_n2416_));
  AOI21_X1   g1774(.A1(new_n776_), .A2(new_n1652_), .B(new_n2416_), .ZN(new_n2417_));
  INV_X1     g1775(.I(new_n2417_), .ZN(new_n2418_));
  INV_X1     g1776(.I(\in0[97] ), .ZN(new_n2419_));
  NOR2_X1    g1777(.A1(new_n1615_), .A2(\in1[97] ), .ZN(new_n2420_));
  AOI21_X1   g1778(.A1(new_n2419_), .A2(new_n1615_), .B(new_n2420_), .ZN(new_n2421_));
  INV_X1     g1779(.I(new_n2421_), .ZN(new_n2422_));
  NAND4_X1   g1780(.A1(new_n2411_), .A2(new_n2415_), .A3(new_n2418_), .A4(new_n2422_), .ZN(new_n2423_));
  OAI21_X1   g1781(.A1(new_n2423_), .A2(new_n2389_), .B(new_n2384_), .ZN(new_n2424_));
  NOR2_X1    g1782(.A1(new_n1615_), .A2(\in1[101] ), .ZN(new_n2425_));
  AOI21_X1   g1783(.A1(new_n1381_), .A2(new_n1615_), .B(new_n2425_), .ZN(new_n2426_));
  INV_X1     g1784(.I(\in0[100] ), .ZN(new_n2427_));
  NOR2_X1    g1785(.A1(new_n1615_), .A2(\in1[100] ), .ZN(new_n2428_));
  AOI21_X1   g1786(.A1(new_n2427_), .A2(new_n1615_), .B(new_n2428_), .ZN(new_n2429_));
  NAND2_X1   g1787(.A1(new_n2426_), .A2(new_n2429_), .ZN(new_n2430_));
  NOR2_X1    g1788(.A1(new_n1652_), .A2(\in2[101] ), .ZN(new_n2431_));
  AOI21_X1   g1789(.A1(new_n897_), .A2(new_n1652_), .B(new_n2431_), .ZN(new_n2432_));
  INV_X1     g1790(.I(new_n2432_), .ZN(new_n2433_));
  INV_X1     g1791(.I(\in3[100] ), .ZN(new_n2434_));
  NOR2_X1    g1792(.A1(new_n1652_), .A2(\in2[100] ), .ZN(new_n2435_));
  AOI21_X1   g1793(.A1(new_n2434_), .A2(new_n1652_), .B(new_n2435_), .ZN(new_n2436_));
  INV_X1     g1794(.I(new_n2436_), .ZN(new_n2437_));
  NAND3_X1   g1795(.A1(new_n2430_), .A2(new_n2433_), .A3(new_n2437_), .ZN(new_n2438_));
  INV_X1     g1796(.I(new_n2426_), .ZN(new_n2439_));
  INV_X1     g1797(.I(new_n2429_), .ZN(new_n2440_));
  INV_X1     g1798(.I(\in3[102] ), .ZN(new_n2441_));
  NOR2_X1    g1799(.A1(new_n1652_), .A2(\in2[102] ), .ZN(new_n2442_));
  AOI21_X1   g1800(.A1(new_n2441_), .A2(new_n1652_), .B(new_n2442_), .ZN(new_n2443_));
  INV_X1     g1801(.I(new_n2443_), .ZN(new_n2444_));
  INV_X1     g1802(.I(\in0[103] ), .ZN(new_n2445_));
  NOR2_X1    g1803(.A1(new_n1615_), .A2(\in1[103] ), .ZN(new_n2446_));
  AOI21_X1   g1804(.A1(new_n2445_), .A2(new_n1615_), .B(new_n2446_), .ZN(new_n2447_));
  INV_X1     g1805(.I(new_n2447_), .ZN(new_n2448_));
  INV_X1     g1806(.I(\in0[102] ), .ZN(new_n2449_));
  NOR2_X1    g1807(.A1(new_n1615_), .A2(\in1[102] ), .ZN(new_n2450_));
  AOI21_X1   g1808(.A1(new_n2449_), .A2(new_n1615_), .B(new_n2450_), .ZN(new_n2451_));
  INV_X1     g1809(.I(new_n2451_), .ZN(new_n2452_));
  INV_X1     g1810(.I(\in3[103] ), .ZN(new_n2453_));
  NOR2_X1    g1811(.A1(new_n1652_), .A2(\in2[103] ), .ZN(new_n2454_));
  AOI21_X1   g1812(.A1(new_n2453_), .A2(new_n1652_), .B(new_n2454_), .ZN(new_n2455_));
  INV_X1     g1813(.I(new_n2455_), .ZN(new_n2456_));
  AOI22_X1   g1814(.A1(new_n2444_), .A2(new_n2448_), .B1(new_n2452_), .B2(new_n2456_), .ZN(new_n2457_));
  AOI21_X1   g1815(.A1(new_n2439_), .A2(new_n2440_), .B(new_n2457_), .ZN(new_n2458_));
  NAND2_X1   g1816(.A1(new_n2458_), .A2(new_n2438_), .ZN(new_n2459_));
  NAND2_X1   g1817(.A1(new_n2448_), .A2(new_n2452_), .ZN(new_n2460_));
  NOR2_X1    g1818(.A1(new_n2448_), .A2(new_n2452_), .ZN(new_n2461_));
  NAND2_X1   g1819(.A1(new_n2444_), .A2(new_n2456_), .ZN(new_n2462_));
  OAI21_X1   g1820(.A1(new_n2461_), .A2(new_n2462_), .B(new_n2460_), .ZN(new_n2463_));
  OAI21_X1   g1821(.A1(new_n2426_), .A2(new_n2433_), .B(new_n2457_), .ZN(new_n2464_));
  NOR2_X1    g1822(.A1(new_n2429_), .A2(new_n2436_), .ZN(new_n2465_));
  NAND4_X1   g1823(.A1(new_n2459_), .A2(new_n2463_), .A3(new_n2464_), .A4(new_n2465_), .ZN(new_n2466_));
  INV_X1     g1824(.I(new_n2410_), .ZN(new_n2467_));
  NOR2_X1    g1825(.A1(new_n2405_), .A2(new_n2397_), .ZN(new_n2468_));
  NAND2_X1   g1826(.A1(new_n2468_), .A2(new_n2422_), .ZN(new_n2469_));
  NAND2_X1   g1827(.A1(new_n2469_), .A2(new_n2417_), .ZN(new_n2470_));
  INV_X1     g1828(.I(new_n2394_), .ZN(new_n2471_));
  NOR2_X1    g1829(.A1(new_n2468_), .A2(new_n2422_), .ZN(new_n2472_));
  NOR4_X1    g1830(.A1(new_n2472_), .A2(new_n2391_), .A3(new_n2471_), .A4(new_n2408_), .ZN(new_n2473_));
  AOI22_X1   g1831(.A1(new_n2473_), .A2(new_n2470_), .B1(new_n2401_), .B2(new_n2467_), .ZN(new_n2474_));
  NAND2_X1   g1832(.A1(new_n2466_), .A2(new_n2474_), .ZN(new_n2475_));
  NAND4_X1   g1833(.A1(new_n2475_), .A2(new_n2307_), .A3(new_n2352_), .A4(new_n2424_), .ZN(new_n2476_));
  NOR3_X1    g1834(.A1(new_n2476_), .A2(new_n2073_), .A3(new_n2249_), .ZN(new_n2477_));
  NOR2_X1    g1835(.A1(new_n1652_), .A2(\in2[33] ), .ZN(new_n2478_));
  AOI21_X1   g1836(.A1(new_n943_), .A2(new_n1652_), .B(new_n2478_), .ZN(new_n2479_));
  NOR2_X1    g1837(.A1(new_n1615_), .A2(\in1[32] ), .ZN(new_n2480_));
  AOI21_X1   g1838(.A1(new_n1425_), .A2(new_n1615_), .B(new_n2480_), .ZN(new_n2481_));
  NOR2_X1    g1839(.A1(new_n1615_), .A2(\in1[33] ), .ZN(new_n2482_));
  AOI21_X1   g1840(.A1(new_n1426_), .A2(new_n1615_), .B(new_n2482_), .ZN(new_n2483_));
  NOR2_X1    g1841(.A1(new_n1652_), .A2(\in2[32] ), .ZN(new_n2484_));
  AOI21_X1   g1842(.A1(new_n942_), .A2(new_n1652_), .B(new_n2484_), .ZN(new_n2485_));
  OAI22_X1   g1843(.A1(new_n2479_), .A2(new_n2481_), .B1(new_n2483_), .B2(new_n2485_), .ZN(new_n2486_));
  NOR2_X1    g1844(.A1(new_n1652_), .A2(\in2[35] ), .ZN(new_n2487_));
  AOI21_X1   g1845(.A1(new_n948_), .A2(new_n1652_), .B(new_n2487_), .ZN(new_n2488_));
  NOR2_X1    g1846(.A1(new_n1615_), .A2(\in1[35] ), .ZN(new_n2489_));
  AOI21_X1   g1847(.A1(new_n1526_), .A2(new_n1615_), .B(new_n2489_), .ZN(new_n2490_));
  OAI22_X1   g1848(.A1(new_n2479_), .A2(new_n2490_), .B1(new_n2483_), .B2(new_n2488_), .ZN(new_n2491_));
  INV_X1     g1849(.I(\in0[34] ), .ZN(new_n2492_));
  NOR2_X1    g1850(.A1(new_n1615_), .A2(\in1[34] ), .ZN(new_n2493_));
  AOI21_X1   g1851(.A1(new_n2492_), .A2(new_n1615_), .B(new_n2493_), .ZN(new_n2494_));
  NOR2_X1    g1852(.A1(new_n1652_), .A2(\in2[34] ), .ZN(new_n2495_));
  AOI21_X1   g1853(.A1(new_n947_), .A2(new_n1652_), .B(new_n2495_), .ZN(new_n2496_));
  INV_X1     g1854(.I(new_n2496_), .ZN(new_n2497_));
  OAI21_X1   g1855(.A1(new_n2494_), .A2(new_n2497_), .B(new_n2491_), .ZN(new_n2498_));
  INV_X1     g1856(.I(\in3[37] ), .ZN(new_n2499_));
  NOR2_X1    g1857(.A1(new_n1652_), .A2(\in2[37] ), .ZN(new_n2500_));
  AOI21_X1   g1858(.A1(new_n2499_), .A2(new_n1652_), .B(new_n2500_), .ZN(new_n2501_));
  INV_X1     g1859(.I(new_n2501_), .ZN(new_n2502_));
  INV_X1     g1860(.I(\in0[37] ), .ZN(new_n2503_));
  NOR2_X1    g1861(.A1(new_n1615_), .A2(\in1[37] ), .ZN(new_n2504_));
  AOI21_X1   g1862(.A1(new_n2503_), .A2(new_n1615_), .B(new_n2504_), .ZN(new_n2505_));
  NOR2_X1    g1863(.A1(new_n2502_), .A2(new_n2505_), .ZN(new_n2506_));
  INV_X1     g1864(.I(\in3[38] ), .ZN(new_n2507_));
  NOR2_X1    g1865(.A1(new_n1652_), .A2(\in2[38] ), .ZN(new_n2508_));
  AOI21_X1   g1866(.A1(new_n2507_), .A2(new_n1652_), .B(new_n2508_), .ZN(new_n2509_));
  INV_X1     g1867(.I(\in0[39] ), .ZN(new_n2510_));
  NOR2_X1    g1868(.A1(new_n1615_), .A2(\in1[39] ), .ZN(new_n2511_));
  AOI21_X1   g1869(.A1(new_n2510_), .A2(new_n1615_), .B(new_n2511_), .ZN(new_n2512_));
  INV_X1     g1870(.I(\in0[38] ), .ZN(new_n2513_));
  NOR2_X1    g1871(.A1(new_n1615_), .A2(\in1[38] ), .ZN(new_n2514_));
  AOI21_X1   g1872(.A1(new_n2513_), .A2(new_n1615_), .B(new_n2514_), .ZN(new_n2515_));
  INV_X1     g1873(.I(\in3[39] ), .ZN(new_n2516_));
  NOR2_X1    g1874(.A1(new_n1652_), .A2(\in2[39] ), .ZN(new_n2517_));
  AOI21_X1   g1875(.A1(new_n2516_), .A2(new_n1652_), .B(new_n2517_), .ZN(new_n2518_));
  OAI22_X1   g1876(.A1(new_n2509_), .A2(new_n2512_), .B1(new_n2515_), .B2(new_n2518_), .ZN(new_n2519_));
  INV_X1     g1877(.I(\in3[36] ), .ZN(new_n2520_));
  NOR2_X1    g1878(.A1(new_n1652_), .A2(\in2[36] ), .ZN(new_n2521_));
  AOI21_X1   g1879(.A1(new_n2520_), .A2(new_n1652_), .B(new_n2521_), .ZN(new_n2522_));
  INV_X1     g1880(.I(\in0[36] ), .ZN(new_n2523_));
  NOR2_X1    g1881(.A1(new_n1615_), .A2(\in1[36] ), .ZN(new_n2524_));
  AOI21_X1   g1882(.A1(new_n2523_), .A2(new_n1615_), .B(new_n2524_), .ZN(new_n2525_));
  NOR2_X1    g1883(.A1(new_n2525_), .A2(new_n2522_), .ZN(new_n2526_));
  OAI21_X1   g1884(.A1(new_n2519_), .A2(new_n2506_), .B(new_n2526_), .ZN(new_n2527_));
  NOR2_X1    g1885(.A1(new_n2490_), .A2(new_n2494_), .ZN(new_n2528_));
  NAND2_X1   g1886(.A1(new_n2490_), .A2(new_n2494_), .ZN(new_n2529_));
  NOR2_X1    g1887(.A1(new_n2488_), .A2(new_n2496_), .ZN(new_n2530_));
  AOI21_X1   g1888(.A1(new_n2529_), .A2(new_n2530_), .B(new_n2528_), .ZN(new_n2531_));
  OAI21_X1   g1889(.A1(new_n2527_), .A2(new_n2531_), .B(new_n2498_), .ZN(new_n2532_));
  INV_X1     g1890(.I(new_n2512_), .ZN(new_n2533_));
  INV_X1     g1891(.I(new_n2515_), .ZN(new_n2534_));
  NAND2_X1   g1892(.A1(new_n2533_), .A2(new_n2534_), .ZN(new_n2535_));
  NOR2_X1    g1893(.A1(new_n2533_), .A2(new_n2534_), .ZN(new_n2536_));
  INV_X1     g1894(.I(new_n2509_), .ZN(new_n2537_));
  INV_X1     g1895(.I(new_n2518_), .ZN(new_n2538_));
  NAND2_X1   g1896(.A1(new_n2537_), .A2(new_n2538_), .ZN(new_n2539_));
  OAI21_X1   g1897(.A1(new_n2536_), .A2(new_n2539_), .B(new_n2535_), .ZN(new_n2540_));
  AOI21_X1   g1898(.A1(new_n2532_), .A2(new_n2486_), .B(new_n2540_), .ZN(new_n2541_));
  NOR2_X1    g1899(.A1(new_n2505_), .A2(new_n2525_), .ZN(new_n2542_));
  INV_X1     g1900(.I(new_n2505_), .ZN(new_n2543_));
  INV_X1     g1901(.I(new_n2525_), .ZN(new_n2544_));
  NOR2_X1    g1902(.A1(new_n2543_), .A2(new_n2544_), .ZN(new_n2545_));
  NOR3_X1    g1903(.A1(new_n2545_), .A2(new_n2501_), .A3(new_n2522_), .ZN(new_n2546_));
  OAI21_X1   g1904(.A1(new_n2546_), .A2(new_n2542_), .B(new_n2519_), .ZN(new_n2547_));
  INV_X1     g1905(.I(\in0[45] ), .ZN(new_n2548_));
  NOR2_X1    g1906(.A1(new_n1615_), .A2(\in1[45] ), .ZN(new_n2549_));
  AOI21_X1   g1907(.A1(new_n2548_), .A2(new_n1615_), .B(new_n2549_), .ZN(new_n2550_));
  INV_X1     g1908(.I(\in3[45] ), .ZN(new_n2551_));
  NOR2_X1    g1909(.A1(new_n1652_), .A2(\in2[45] ), .ZN(new_n2552_));
  AOI21_X1   g1910(.A1(new_n2551_), .A2(new_n1652_), .B(new_n2552_), .ZN(new_n2553_));
  INV_X1     g1911(.I(\in3[46] ), .ZN(new_n2554_));
  NOR2_X1    g1912(.A1(new_n1652_), .A2(\in2[46] ), .ZN(new_n2555_));
  AOI21_X1   g1913(.A1(new_n2554_), .A2(new_n1652_), .B(new_n2555_), .ZN(new_n2556_));
  INV_X1     g1914(.I(new_n2556_), .ZN(new_n2557_));
  INV_X1     g1915(.I(\in0[47] ), .ZN(new_n2558_));
  NOR2_X1    g1916(.A1(new_n1615_), .A2(\in1[47] ), .ZN(new_n2559_));
  AOI21_X1   g1917(.A1(new_n2558_), .A2(new_n1615_), .B(new_n2559_), .ZN(new_n2560_));
  INV_X1     g1918(.I(new_n2560_), .ZN(new_n2561_));
  INV_X1     g1919(.I(\in0[46] ), .ZN(new_n2562_));
  NOR2_X1    g1920(.A1(new_n1615_), .A2(\in1[46] ), .ZN(new_n2563_));
  AOI21_X1   g1921(.A1(new_n2562_), .A2(new_n1615_), .B(new_n2563_), .ZN(new_n2564_));
  INV_X1     g1922(.I(new_n2564_), .ZN(new_n2565_));
  INV_X1     g1923(.I(\in3[47] ), .ZN(new_n2566_));
  NOR2_X1    g1924(.A1(new_n1652_), .A2(\in2[47] ), .ZN(new_n2567_));
  AOI21_X1   g1925(.A1(new_n2566_), .A2(new_n1652_), .B(new_n2567_), .ZN(new_n2568_));
  INV_X1     g1926(.I(new_n2568_), .ZN(new_n2569_));
  AOI22_X1   g1927(.A1(new_n2557_), .A2(new_n2561_), .B1(new_n2565_), .B2(new_n2569_), .ZN(new_n2570_));
  OAI21_X1   g1928(.A1(new_n2570_), .A2(new_n2553_), .B(new_n2550_), .ZN(new_n2571_));
  INV_X1     g1929(.I(\in3[44] ), .ZN(new_n2572_));
  NOR2_X1    g1930(.A1(new_n1652_), .A2(\in2[44] ), .ZN(new_n2573_));
  AOI21_X1   g1931(.A1(new_n2572_), .A2(new_n1652_), .B(new_n2573_), .ZN(new_n2574_));
  INV_X1     g1932(.I(new_n2574_), .ZN(new_n2575_));
  INV_X1     g1933(.I(\in0[44] ), .ZN(new_n2576_));
  NOR2_X1    g1934(.A1(new_n1615_), .A2(\in1[44] ), .ZN(new_n2577_));
  AOI21_X1   g1935(.A1(new_n2576_), .A2(new_n1615_), .B(new_n2577_), .ZN(new_n2578_));
  NAND2_X1   g1936(.A1(new_n2575_), .A2(new_n2578_), .ZN(new_n2579_));
  AOI21_X1   g1937(.A1(new_n2570_), .A2(new_n2553_), .B(new_n2579_), .ZN(new_n2580_));
  NAND2_X1   g1938(.A1(new_n2561_), .A2(new_n2565_), .ZN(new_n2581_));
  NOR2_X1    g1939(.A1(new_n2561_), .A2(new_n2565_), .ZN(new_n2582_));
  NAND2_X1   g1940(.A1(new_n2557_), .A2(new_n2569_), .ZN(new_n2583_));
  OAI21_X1   g1941(.A1(new_n2582_), .A2(new_n2583_), .B(new_n2581_), .ZN(new_n2584_));
  AOI21_X1   g1942(.A1(new_n2580_), .A2(new_n2571_), .B(new_n2584_), .ZN(new_n2585_));
  NOR2_X1    g1943(.A1(new_n1615_), .A2(\in1[43] ), .ZN(new_n2586_));
  AOI21_X1   g1944(.A1(new_n1544_), .A2(new_n1615_), .B(new_n2586_), .ZN(new_n2587_));
  INV_X1     g1945(.I(new_n2587_), .ZN(new_n2588_));
  INV_X1     g1946(.I(\in3[42] ), .ZN(new_n2589_));
  NOR2_X1    g1947(.A1(new_n1652_), .A2(\in2[42] ), .ZN(new_n2590_));
  AOI21_X1   g1948(.A1(new_n2589_), .A2(new_n1652_), .B(new_n2590_), .ZN(new_n2591_));
  INV_X1     g1949(.I(new_n2591_), .ZN(new_n2592_));
  INV_X1     g1950(.I(\in0[42] ), .ZN(new_n2593_));
  NOR2_X1    g1951(.A1(new_n1615_), .A2(\in1[42] ), .ZN(new_n2594_));
  AOI21_X1   g1952(.A1(new_n2593_), .A2(new_n1615_), .B(new_n2594_), .ZN(new_n2595_));
  INV_X1     g1953(.I(new_n2595_), .ZN(new_n2596_));
  INV_X1     g1954(.I(\in3[43] ), .ZN(new_n2597_));
  NOR2_X1    g1955(.A1(new_n1652_), .A2(\in2[43] ), .ZN(new_n2598_));
  AOI21_X1   g1956(.A1(new_n2597_), .A2(new_n1652_), .B(new_n2598_), .ZN(new_n2599_));
  INV_X1     g1957(.I(new_n2599_), .ZN(new_n2600_));
  AOI22_X1   g1958(.A1(new_n2588_), .A2(new_n2592_), .B1(new_n2596_), .B2(new_n2600_), .ZN(new_n2601_));
  INV_X1     g1959(.I(new_n2601_), .ZN(new_n2602_));
  NOR2_X1    g1960(.A1(new_n1652_), .A2(\in2[41] ), .ZN(new_n2603_));
  AOI21_X1   g1961(.A1(new_n1071_), .A2(new_n1652_), .B(new_n2603_), .ZN(new_n2604_));
  INV_X1     g1962(.I(new_n2604_), .ZN(new_n2605_));
  NOR2_X1    g1963(.A1(new_n1615_), .A2(\in1[41] ), .ZN(new_n2606_));
  AOI21_X1   g1964(.A1(new_n1549_), .A2(new_n1615_), .B(new_n2606_), .ZN(new_n2607_));
  INV_X1     g1965(.I(new_n2607_), .ZN(new_n2608_));
  NOR2_X1    g1966(.A1(new_n2596_), .A2(new_n2591_), .ZN(new_n2609_));
  AOI21_X1   g1967(.A1(new_n2609_), .A2(new_n2608_), .B(new_n2605_), .ZN(new_n2610_));
  NOR2_X1    g1968(.A1(new_n1652_), .A2(\in2[40] ), .ZN(new_n2611_));
  AOI21_X1   g1969(.A1(new_n1068_), .A2(new_n1652_), .B(new_n2611_), .ZN(new_n2612_));
  NOR2_X1    g1970(.A1(new_n1615_), .A2(\in1[40] ), .ZN(new_n2613_));
  AOI21_X1   g1971(.A1(new_n1546_), .A2(new_n1615_), .B(new_n2613_), .ZN(new_n2614_));
  INV_X1     g1972(.I(new_n2614_), .ZN(new_n2615_));
  NOR3_X1    g1973(.A1(new_n2615_), .A2(new_n2599_), .A3(new_n2612_), .ZN(new_n2616_));
  OAI21_X1   g1974(.A1(new_n2608_), .A2(new_n2609_), .B(new_n2616_), .ZN(new_n2617_));
  OAI22_X1   g1975(.A1(new_n2617_), .A2(new_n2610_), .B1(new_n2587_), .B2(new_n2601_), .ZN(new_n2618_));
  INV_X1     g1976(.I(new_n2578_), .ZN(new_n2619_));
  INV_X1     g1977(.I(new_n2553_), .ZN(new_n2620_));
  OAI21_X1   g1978(.A1(new_n2550_), .A2(new_n2620_), .B(new_n2570_), .ZN(new_n2621_));
  AND3_X2    g1979(.A1(new_n2621_), .A2(new_n2575_), .A3(new_n2619_), .Z(new_n2622_));
  OAI22_X1   g1980(.A1(new_n2604_), .A2(new_n2614_), .B1(new_n2607_), .B2(new_n2612_), .ZN(new_n2623_));
  NAND4_X1   g1981(.A1(new_n2622_), .A2(new_n2602_), .A3(new_n2618_), .A4(new_n2623_), .ZN(new_n2624_));
  OAI22_X1   g1982(.A1(new_n2624_), .A2(new_n2585_), .B1(new_n2541_), .B2(new_n2547_), .ZN(new_n2625_));
  NOR2_X1    g1983(.A1(new_n1652_), .A2(\in2[31] ), .ZN(new_n2626_));
  AOI21_X1   g1984(.A1(new_n952_), .A2(new_n1652_), .B(new_n2626_), .ZN(new_n2627_));
  INV_X1     g1985(.I(new_n2627_), .ZN(new_n2628_));
  INV_X1     g1986(.I(new_n2481_), .ZN(new_n2629_));
  INV_X1     g1987(.I(new_n2485_), .ZN(new_n2630_));
  NAND2_X1   g1988(.A1(new_n2629_), .A2(new_n2630_), .ZN(new_n2631_));
  AOI21_X1   g1989(.A1(new_n2498_), .A2(new_n2527_), .B(new_n2631_), .ZN(new_n2632_));
  INV_X1     g1990(.I(\in3[125] ), .ZN(new_n2633_));
  NOR2_X1    g1991(.A1(new_n1652_), .A2(\in2[125] ), .ZN(new_n2634_));
  AOI21_X1   g1992(.A1(new_n2633_), .A2(new_n1652_), .B(new_n2634_), .ZN(new_n2635_));
  NOR2_X1    g1993(.A1(new_n1615_), .A2(\in1[126] ), .ZN(new_n2636_));
  AOI21_X1   g1994(.A1(new_n1342_), .A2(new_n1615_), .B(new_n2636_), .ZN(new_n2637_));
  INV_X1     g1995(.I(\in0[125] ), .ZN(new_n2638_));
  NOR2_X1    g1996(.A1(new_n1615_), .A2(\in1[125] ), .ZN(new_n2639_));
  AOI21_X1   g1997(.A1(new_n2638_), .A2(new_n1615_), .B(new_n2639_), .ZN(new_n2640_));
  NOR2_X1    g1998(.A1(new_n1652_), .A2(\in2[126] ), .ZN(new_n2641_));
  AOI21_X1   g1999(.A1(new_n858_), .A2(new_n1652_), .B(new_n2641_), .ZN(new_n2642_));
  OAI22_X1   g2000(.A1(new_n2635_), .A2(new_n2637_), .B1(new_n2640_), .B2(new_n2642_), .ZN(new_n2643_));
  INV_X1     g2001(.I(new_n1609_), .ZN(new_n2644_));
  INV_X1     g2002(.I(new_n2637_), .ZN(new_n2645_));
  NOR4_X1    g2003(.A1(new_n2645_), .A2(new_n2644_), .A3(new_n1610_), .A4(new_n2642_), .ZN(new_n2646_));
  NOR2_X1    g2004(.A1(new_n2646_), .A2(new_n2643_), .ZN(new_n2647_));
  AOI21_X1   g2005(.A1(new_n1609_), .A2(new_n1611_), .B(new_n2643_), .ZN(new_n2648_));
  INV_X1     g2006(.I(new_n2635_), .ZN(new_n2649_));
  INV_X1     g2007(.I(new_n2640_), .ZN(new_n2650_));
  INV_X1     g2008(.I(\in0[124] ), .ZN(new_n2651_));
  NOR2_X1    g2009(.A1(new_n1615_), .A2(\in1[124] ), .ZN(new_n2652_));
  AOI21_X1   g2010(.A1(new_n2651_), .A2(new_n1615_), .B(new_n2652_), .ZN(new_n2653_));
  INV_X1     g2011(.I(new_n2653_), .ZN(new_n2654_));
  INV_X1     g2012(.I(\in3[124] ), .ZN(new_n2655_));
  NOR2_X1    g2013(.A1(new_n1652_), .A2(\in2[124] ), .ZN(new_n2656_));
  AOI21_X1   g2014(.A1(new_n2655_), .A2(new_n1652_), .B(new_n2656_), .ZN(new_n2657_));
  INV_X1     g2015(.I(new_n2657_), .ZN(new_n2658_));
  AOI22_X1   g2016(.A1(new_n2649_), .A2(new_n2654_), .B1(new_n2650_), .B2(new_n2658_), .ZN(new_n2659_));
  NAND2_X1   g2017(.A1(new_n2654_), .A2(new_n2658_), .ZN(new_n2660_));
  NOR4_X1    g2018(.A1(new_n2647_), .A2(new_n2648_), .A3(new_n2659_), .A4(new_n2660_), .ZN(new_n2661_));
  NOR2_X1    g2019(.A1(new_n2126_), .A2(new_n2118_), .ZN(new_n2662_));
  AOI21_X1   g2020(.A1(new_n2662_), .A2(new_n2143_), .B(new_n2139_), .ZN(new_n2663_));
  INV_X1     g2021(.I(new_n2115_), .ZN(new_n2664_));
  NOR3_X1    g2022(.A1(new_n2664_), .A2(new_n2112_), .A3(new_n2129_), .ZN(new_n2665_));
  OAI21_X1   g2023(.A1(new_n2143_), .A2(new_n2662_), .B(new_n2665_), .ZN(new_n2666_));
  OAI22_X1   g2024(.A1(new_n2666_), .A2(new_n2663_), .B1(new_n2121_), .B2(new_n2131_), .ZN(new_n2667_));
  OAI22_X1   g2025(.A1(new_n2667_), .A2(new_n2661_), .B1(new_n2628_), .B2(new_n2632_), .ZN(new_n2668_));
  NOR2_X1    g2026(.A1(new_n1652_), .A2(\in2[69] ), .ZN(new_n2669_));
  AOI21_X1   g2027(.A1(new_n923_), .A2(new_n1652_), .B(new_n2669_), .ZN(new_n2670_));
  NOR2_X1    g2028(.A1(new_n1615_), .A2(\in1[69] ), .ZN(new_n2671_));
  AOI21_X1   g2029(.A1(new_n1407_), .A2(new_n1615_), .B(new_n2671_), .ZN(new_n2672_));
  INV_X1     g2030(.I(new_n2672_), .ZN(new_n2673_));
  NAND2_X1   g2031(.A1(new_n2673_), .A2(new_n2670_), .ZN(new_n2674_));
  INV_X1     g2032(.I(\in3[70] ), .ZN(new_n2675_));
  NOR2_X1    g2033(.A1(new_n1652_), .A2(\in2[70] ), .ZN(new_n2676_));
  AOI21_X1   g2034(.A1(new_n2675_), .A2(new_n1652_), .B(new_n2676_), .ZN(new_n2677_));
  INV_X1     g2035(.I(new_n2677_), .ZN(new_n2678_));
  INV_X1     g2036(.I(\in0[71] ), .ZN(new_n2679_));
  NOR2_X1    g2037(.A1(new_n1615_), .A2(\in1[71] ), .ZN(new_n2680_));
  AOI21_X1   g2038(.A1(new_n2679_), .A2(new_n1615_), .B(new_n2680_), .ZN(new_n2681_));
  INV_X1     g2039(.I(new_n2681_), .ZN(new_n2682_));
  INV_X1     g2040(.I(\in0[70] ), .ZN(new_n2683_));
  NOR2_X1    g2041(.A1(new_n1615_), .A2(\in1[70] ), .ZN(new_n2684_));
  AOI21_X1   g2042(.A1(new_n2683_), .A2(new_n1615_), .B(new_n2684_), .ZN(new_n2685_));
  INV_X1     g2043(.I(new_n2685_), .ZN(new_n2686_));
  INV_X1     g2044(.I(\in3[71] ), .ZN(new_n2687_));
  NOR2_X1    g2045(.A1(new_n1652_), .A2(\in2[71] ), .ZN(new_n2688_));
  AOI21_X1   g2046(.A1(new_n2687_), .A2(new_n1652_), .B(new_n2688_), .ZN(new_n2689_));
  INV_X1     g2047(.I(new_n2689_), .ZN(new_n2690_));
  AOI22_X1   g2048(.A1(new_n2678_), .A2(new_n2682_), .B1(new_n2686_), .B2(new_n2690_), .ZN(new_n2691_));
  INV_X1     g2049(.I(\in3[68] ), .ZN(new_n2692_));
  NOR2_X1    g2050(.A1(new_n1652_), .A2(\in2[68] ), .ZN(new_n2693_));
  AOI21_X1   g2051(.A1(new_n2692_), .A2(new_n1652_), .B(new_n2693_), .ZN(new_n2694_));
  INV_X1     g2052(.I(new_n2694_), .ZN(new_n2695_));
  INV_X1     g2053(.I(\in0[68] ), .ZN(new_n2696_));
  NOR2_X1    g2054(.A1(new_n1615_), .A2(\in1[68] ), .ZN(new_n2697_));
  AOI21_X1   g2055(.A1(new_n2696_), .A2(new_n1615_), .B(new_n2697_), .ZN(new_n2698_));
  INV_X1     g2056(.I(new_n2698_), .ZN(new_n2699_));
  NAND2_X1   g2057(.A1(new_n2699_), .A2(new_n2695_), .ZN(new_n2700_));
  AOI21_X1   g2058(.A1(new_n2691_), .A2(new_n2674_), .B(new_n2700_), .ZN(new_n2701_));
  NOR2_X1    g2059(.A1(new_n2673_), .A2(new_n2699_), .ZN(new_n2702_));
  NOR3_X1    g2060(.A1(new_n2702_), .A2(new_n2670_), .A3(new_n2694_), .ZN(new_n2703_));
  NOR2_X1    g2061(.A1(new_n2672_), .A2(new_n2698_), .ZN(new_n2704_));
  NOR3_X1    g2062(.A1(new_n2703_), .A2(new_n2691_), .A3(new_n2704_), .ZN(new_n2705_));
  NOR2_X1    g2063(.A1(new_n1652_), .A2(\in2[72] ), .ZN(new_n2706_));
  AOI21_X1   g2064(.A1(new_n887_), .A2(new_n1652_), .B(new_n2706_), .ZN(new_n2707_));
  NOR2_X1    g2065(.A1(new_n1615_), .A2(\in1[72] ), .ZN(new_n2708_));
  AOI21_X1   g2066(.A1(new_n1371_), .A2(new_n1615_), .B(new_n2708_), .ZN(new_n2709_));
  INV_X1     g2067(.I(new_n2709_), .ZN(new_n2710_));
  INV_X1     g2068(.I(\in3[74] ), .ZN(new_n2711_));
  NOR2_X1    g2069(.A1(new_n1652_), .A2(\in2[74] ), .ZN(new_n2712_));
  AOI21_X1   g2070(.A1(new_n2711_), .A2(new_n1652_), .B(new_n2712_), .ZN(new_n2713_));
  INV_X1     g2071(.I(new_n2713_), .ZN(new_n2714_));
  NOR2_X1    g2072(.A1(new_n1615_), .A2(\in1[75] ), .ZN(new_n2715_));
  AOI21_X1   g2073(.A1(new_n1376_), .A2(new_n1615_), .B(new_n2715_), .ZN(new_n2716_));
  INV_X1     g2074(.I(new_n2716_), .ZN(new_n2717_));
  INV_X1     g2075(.I(\in0[74] ), .ZN(new_n2718_));
  NOR2_X1    g2076(.A1(new_n1615_), .A2(\in1[74] ), .ZN(new_n2719_));
  AOI21_X1   g2077(.A1(new_n2718_), .A2(new_n1615_), .B(new_n2719_), .ZN(new_n2720_));
  INV_X1     g2078(.I(new_n2720_), .ZN(new_n2721_));
  INV_X1     g2079(.I(\in3[75] ), .ZN(new_n2722_));
  NOR2_X1    g2080(.A1(new_n1652_), .A2(\in2[75] ), .ZN(new_n2723_));
  AOI21_X1   g2081(.A1(new_n2722_), .A2(new_n1652_), .B(new_n2723_), .ZN(new_n2724_));
  INV_X1     g2082(.I(new_n2724_), .ZN(new_n2725_));
  AOI22_X1   g2083(.A1(new_n2714_), .A2(new_n2717_), .B1(new_n2721_), .B2(new_n2725_), .ZN(new_n2726_));
  INV_X1     g2084(.I(new_n2726_), .ZN(new_n2727_));
  AOI21_X1   g2085(.A1(new_n2707_), .A2(new_n2710_), .B(new_n2727_), .ZN(new_n2728_));
  NOR2_X1    g2086(.A1(new_n2682_), .A2(new_n2686_), .ZN(new_n2729_));
  NOR3_X1    g2087(.A1(new_n2729_), .A2(new_n2677_), .A3(new_n2689_), .ZN(new_n2730_));
  AOI21_X1   g2088(.A1(new_n2682_), .A2(new_n2686_), .B(new_n2730_), .ZN(new_n2731_));
  NOR2_X1    g2089(.A1(new_n1652_), .A2(\in2[73] ), .ZN(new_n2732_));
  AOI21_X1   g2090(.A1(new_n892_), .A2(new_n1652_), .B(new_n2732_), .ZN(new_n2733_));
  INV_X1     g2091(.I(new_n2733_), .ZN(new_n2734_));
  INV_X1     g2092(.I(\in0[73] ), .ZN(new_n2735_));
  NOR2_X1    g2093(.A1(new_n1615_), .A2(\in1[73] ), .ZN(new_n2736_));
  AOI21_X1   g2094(.A1(new_n2735_), .A2(new_n1615_), .B(new_n2736_), .ZN(new_n2737_));
  INV_X1     g2095(.I(new_n2737_), .ZN(new_n2738_));
  NAND2_X1   g2096(.A1(new_n2738_), .A2(new_n2734_), .ZN(new_n2739_));
  NOR4_X1    g2097(.A1(new_n2728_), .A2(new_n2731_), .A3(new_n2705_), .A4(new_n2739_), .ZN(new_n2740_));
  NOR2_X1    g2098(.A1(new_n1615_), .A2(\in1[77] ), .ZN(new_n2741_));
  AOI21_X1   g2099(.A1(new_n1356_), .A2(new_n1615_), .B(new_n2741_), .ZN(new_n2742_));
  INV_X1     g2100(.I(new_n2742_), .ZN(new_n2743_));
  INV_X1     g2101(.I(\in0[76] ), .ZN(new_n2744_));
  NOR2_X1    g2102(.A1(new_n1615_), .A2(\in1[76] ), .ZN(new_n2745_));
  AOI21_X1   g2103(.A1(new_n2744_), .A2(new_n1615_), .B(new_n2745_), .ZN(new_n2746_));
  INV_X1     g2104(.I(new_n2746_), .ZN(new_n2747_));
  NOR2_X1    g2105(.A1(new_n2743_), .A2(new_n2747_), .ZN(new_n2748_));
  NOR2_X1    g2106(.A1(new_n1652_), .A2(\in2[77] ), .ZN(new_n2749_));
  AOI21_X1   g2107(.A1(new_n872_), .A2(new_n1652_), .B(new_n2749_), .ZN(new_n2750_));
  INV_X1     g2108(.I(\in3[76] ), .ZN(new_n2751_));
  NOR2_X1    g2109(.A1(new_n1652_), .A2(\in2[76] ), .ZN(new_n2752_));
  AOI21_X1   g2110(.A1(new_n2751_), .A2(new_n1652_), .B(new_n2752_), .ZN(new_n2753_));
  NOR3_X1    g2111(.A1(new_n2748_), .A2(new_n2750_), .A3(new_n2753_), .ZN(new_n2754_));
  INV_X1     g2112(.I(\in3[78] ), .ZN(new_n2755_));
  NOR2_X1    g2113(.A1(new_n1652_), .A2(\in2[78] ), .ZN(new_n2756_));
  AOI21_X1   g2114(.A1(new_n2755_), .A2(new_n1652_), .B(new_n2756_), .ZN(new_n2757_));
  INV_X1     g2115(.I(new_n2757_), .ZN(new_n2758_));
  INV_X1     g2116(.I(\in0[79] ), .ZN(new_n2759_));
  NOR2_X1    g2117(.A1(new_n1615_), .A2(\in1[79] ), .ZN(new_n2760_));
  AOI21_X1   g2118(.A1(new_n2759_), .A2(new_n1615_), .B(new_n2760_), .ZN(new_n2761_));
  INV_X1     g2119(.I(new_n2761_), .ZN(new_n2762_));
  INV_X1     g2120(.I(\in0[78] ), .ZN(new_n2763_));
  NOR2_X1    g2121(.A1(new_n1615_), .A2(\in1[78] ), .ZN(new_n2764_));
  AOI21_X1   g2122(.A1(new_n2763_), .A2(new_n1615_), .B(new_n2764_), .ZN(new_n2765_));
  INV_X1     g2123(.I(new_n2765_), .ZN(new_n2766_));
  INV_X1     g2124(.I(\in3[79] ), .ZN(new_n2767_));
  NOR2_X1    g2125(.A1(new_n1652_), .A2(\in2[79] ), .ZN(new_n2768_));
  AOI21_X1   g2126(.A1(new_n2767_), .A2(new_n1652_), .B(new_n2768_), .ZN(new_n2769_));
  INV_X1     g2127(.I(new_n2769_), .ZN(new_n2770_));
  AOI22_X1   g2128(.A1(new_n2758_), .A2(new_n2762_), .B1(new_n2766_), .B2(new_n2770_), .ZN(new_n2771_));
  NOR2_X1    g2129(.A1(new_n2742_), .A2(new_n2746_), .ZN(new_n2772_));
  NOR3_X1    g2130(.A1(new_n2754_), .A2(new_n2771_), .A3(new_n2772_), .ZN(new_n2773_));
  NOR2_X1    g2131(.A1(new_n2761_), .A2(new_n2765_), .ZN(new_n2774_));
  NAND2_X1   g2132(.A1(new_n2761_), .A2(new_n2765_), .ZN(new_n2775_));
  NOR2_X1    g2133(.A1(new_n2757_), .A2(new_n2769_), .ZN(new_n2776_));
  AOI21_X1   g2134(.A1(new_n2775_), .A2(new_n2776_), .B(new_n2774_), .ZN(new_n2777_));
  INV_X1     g2135(.I(new_n2753_), .ZN(new_n2778_));
  INV_X1     g2136(.I(new_n2750_), .ZN(new_n2779_));
  OAI21_X1   g2137(.A1(new_n2742_), .A2(new_n2779_), .B(new_n2771_), .ZN(new_n2780_));
  NAND3_X1   g2138(.A1(new_n2780_), .A2(new_n2747_), .A3(new_n2778_), .ZN(new_n2781_));
  NOR3_X1    g2139(.A1(new_n2781_), .A2(new_n2773_), .A3(new_n2777_), .ZN(new_n2782_));
  NOR2_X1    g2140(.A1(new_n2721_), .A2(new_n2713_), .ZN(new_n2783_));
  AOI21_X1   g2141(.A1(new_n2783_), .A2(new_n2738_), .B(new_n2734_), .ZN(new_n2784_));
  NOR3_X1    g2142(.A1(new_n2710_), .A2(new_n2707_), .A3(new_n2724_), .ZN(new_n2785_));
  OAI21_X1   g2143(.A1(new_n2738_), .A2(new_n2783_), .B(new_n2785_), .ZN(new_n2786_));
  OAI22_X1   g2144(.A1(new_n2786_), .A2(new_n2784_), .B1(new_n2716_), .B2(new_n2726_), .ZN(new_n2787_));
  OAI22_X1   g2145(.A1(new_n2782_), .A2(new_n2787_), .B1(new_n2740_), .B2(new_n2701_), .ZN(new_n2788_));
  NOR2_X1    g2146(.A1(new_n1615_), .A2(\in1[31] ), .ZN(new_n2789_));
  AOI21_X1   g2147(.A1(new_n1420_), .A2(new_n1615_), .B(new_n2789_), .ZN(new_n2790_));
  INV_X1     g2148(.I(new_n2790_), .ZN(new_n2791_));
  AOI21_X1   g2149(.A1(new_n2632_), .A2(new_n2628_), .B(new_n2791_), .ZN(new_n2792_));
  INV_X1     g2150(.I(new_n2019_), .ZN(new_n2793_));
  INV_X1     g2151(.I(new_n2036_), .ZN(new_n2794_));
  AOI21_X1   g2152(.A1(new_n2794_), .A2(new_n2016_), .B(new_n2793_), .ZN(new_n2795_));
  NOR2_X1    g2153(.A1(new_n2045_), .A2(new_n2040_), .ZN(new_n2796_));
  OAI21_X1   g2154(.A1(new_n2794_), .A2(new_n2016_), .B(new_n2796_), .ZN(new_n2797_));
  NOR2_X1    g2155(.A1(new_n2026_), .A2(new_n2030_), .ZN(new_n2798_));
  NAND2_X1   g2156(.A1(new_n2026_), .A2(new_n2030_), .ZN(new_n2799_));
  NOR2_X1    g2157(.A1(new_n2022_), .A2(new_n2034_), .ZN(new_n2800_));
  AOI21_X1   g2158(.A1(new_n2799_), .A2(new_n2800_), .B(new_n2798_), .ZN(new_n2801_));
  OAI21_X1   g2159(.A1(new_n2795_), .A2(new_n2797_), .B(new_n2801_), .ZN(new_n2802_));
  INV_X1     g2160(.I(new_n2051_), .ZN(new_n2803_));
  NAND2_X1   g2161(.A1(new_n2057_), .A2(new_n2803_), .ZN(new_n2804_));
  INV_X1     g2162(.I(new_n2056_), .ZN(new_n2805_));
  INV_X1     g2163(.I(new_n2049_), .ZN(new_n2806_));
  NAND2_X1   g2164(.A1(new_n2806_), .A2(new_n2054_), .ZN(new_n2807_));
  OAI21_X1   g2165(.A1(new_n2807_), .A2(new_n2063_), .B(new_n2069_), .ZN(new_n2808_));
  NAND2_X1   g2166(.A1(new_n2807_), .A2(new_n2063_), .ZN(new_n2809_));
  INV_X1     g2167(.I(new_n2066_), .ZN(new_n2810_));
  NOR2_X1    g2168(.A1(new_n2810_), .A2(new_n2060_), .ZN(new_n2811_));
  NAND4_X1   g2169(.A1(new_n2808_), .A2(new_n2809_), .A3(new_n2805_), .A4(new_n2811_), .ZN(new_n2812_));
  AOI21_X1   g2170(.A1(new_n2812_), .A2(new_n2804_), .B(new_n2046_), .ZN(new_n2813_));
  NOR2_X1    g2171(.A1(new_n1615_), .A2(\in1[67] ), .ZN(new_n2814_));
  AOI21_X1   g2172(.A1(new_n1518_), .A2(new_n1615_), .B(new_n2814_), .ZN(new_n2815_));
  INV_X1     g2173(.I(new_n2815_), .ZN(new_n2816_));
  NOR2_X1    g2174(.A1(new_n1652_), .A2(\in2[66] ), .ZN(new_n2817_));
  AOI21_X1   g2175(.A1(new_n1038_), .A2(new_n1652_), .B(new_n2817_), .ZN(new_n2818_));
  INV_X1     g2176(.I(new_n2818_), .ZN(new_n2819_));
  INV_X1     g2177(.I(\in0[66] ), .ZN(new_n2820_));
  NOR2_X1    g2178(.A1(new_n1615_), .A2(\in1[66] ), .ZN(new_n2821_));
  AOI21_X1   g2179(.A1(new_n2820_), .A2(new_n1615_), .B(new_n2821_), .ZN(new_n2822_));
  INV_X1     g2180(.I(new_n2822_), .ZN(new_n2823_));
  NOR2_X1    g2181(.A1(new_n1652_), .A2(\in2[67] ), .ZN(new_n2824_));
  AOI21_X1   g2182(.A1(new_n1033_), .A2(new_n1652_), .B(new_n2824_), .ZN(new_n2825_));
  INV_X1     g2183(.I(new_n2825_), .ZN(new_n2826_));
  AOI22_X1   g2184(.A1(new_n2816_), .A2(new_n2819_), .B1(new_n2823_), .B2(new_n2826_), .ZN(new_n2827_));
  NOR2_X1    g2185(.A1(new_n1652_), .A2(\in2[65] ), .ZN(new_n2828_));
  AOI21_X1   g2186(.A1(new_n1044_), .A2(new_n1652_), .B(new_n2828_), .ZN(new_n2829_));
  INV_X1     g2187(.I(new_n2829_), .ZN(new_n2830_));
  NOR2_X1    g2188(.A1(new_n1615_), .A2(\in1[65] ), .ZN(new_n2831_));
  AOI21_X1   g2189(.A1(new_n1519_), .A2(new_n1615_), .B(new_n2831_), .ZN(new_n2832_));
  INV_X1     g2190(.I(new_n2832_), .ZN(new_n2833_));
  NOR2_X1    g2191(.A1(new_n2823_), .A2(new_n2818_), .ZN(new_n2834_));
  AOI21_X1   g2192(.A1(new_n2834_), .A2(new_n2833_), .B(new_n2830_), .ZN(new_n2835_));
  INV_X1     g2193(.I(\in3[64] ), .ZN(new_n2836_));
  NOR2_X1    g2194(.A1(new_n1652_), .A2(\in2[64] ), .ZN(new_n2837_));
  AOI21_X1   g2195(.A1(new_n2836_), .A2(new_n1652_), .B(new_n2837_), .ZN(new_n2838_));
  INV_X1     g2196(.I(\in0[64] ), .ZN(new_n2839_));
  NOR2_X1    g2197(.A1(new_n1615_), .A2(\in1[64] ), .ZN(new_n2840_));
  AOI21_X1   g2198(.A1(new_n2839_), .A2(new_n1615_), .B(new_n2840_), .ZN(new_n2841_));
  INV_X1     g2199(.I(new_n2841_), .ZN(new_n2842_));
  NOR3_X1    g2200(.A1(new_n2842_), .A2(new_n2825_), .A3(new_n2838_), .ZN(new_n2843_));
  OAI21_X1   g2201(.A1(new_n2833_), .A2(new_n2834_), .B(new_n2843_), .ZN(new_n2844_));
  OAI22_X1   g2202(.A1(new_n2844_), .A2(new_n2835_), .B1(new_n2815_), .B2(new_n2827_), .ZN(new_n2845_));
  NAND2_X1   g2203(.A1(new_n2842_), .A2(new_n2838_), .ZN(new_n2846_));
  NAND2_X1   g2204(.A1(new_n2833_), .A2(new_n2830_), .ZN(new_n2847_));
  AOI21_X1   g2205(.A1(new_n2827_), .A2(new_n2846_), .B(new_n2847_), .ZN(new_n2848_));
  AOI22_X1   g2206(.A1(new_n2813_), .A2(new_n2802_), .B1(new_n2845_), .B2(new_n2848_), .ZN(new_n2849_));
  NOR4_X1    g2207(.A1(new_n2849_), .A2(new_n2788_), .A3(new_n2668_), .A4(new_n2792_), .ZN(new_n2850_));
  NAND3_X1   g2208(.A1(new_n2477_), .A2(new_n2625_), .A3(new_n2850_), .ZN(new_n2851_));
  AOI21_X1   g2209(.A1(new_n1947_), .A2(new_n1656_), .B(new_n2851_), .ZN(new_n2852_));
  NOR2_X1    g2210(.A1(new_n1615_), .A2(\in1[0] ), .ZN(new_n2853_));
  AOI21_X1   g2211(.A1(new_n1770_), .A2(new_n1615_), .B(new_n2853_), .ZN(new_n2854_));
  INV_X1     g2212(.I(new_n2854_), .ZN(new_n2855_));
  NAND4_X1   g2213(.A1(new_n2852_), .A2(new_n1133_), .A3(new_n1612_), .A4(new_n2855_), .ZN(new_n2856_));
  INV_X1     g2214(.I(new_n1133_), .ZN(new_n2857_));
  NAND4_X1   g2215(.A1(new_n2852_), .A2(new_n2857_), .A3(new_n1612_), .A4(new_n2854_), .ZN(new_n2858_));
  NAND2_X1   g2216(.A1(new_n2856_), .A2(new_n2858_), .ZN(\result[0] ));
  INV_X1     g2217(.I(new_n1799_), .ZN(new_n2860_));
  NAND4_X1   g2218(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1769_), .A4(new_n2860_), .ZN(new_n2861_));
  INV_X1     g2219(.I(new_n1769_), .ZN(new_n2862_));
  NAND4_X1   g2220(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2862_), .A4(new_n1799_), .ZN(new_n2863_));
  NAND2_X1   g2221(.A1(new_n2861_), .A2(new_n2863_), .ZN(\result[1] ));
  NAND4_X1   g2222(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1790_), .A4(new_n1802_), .ZN(new_n2865_));
  INV_X1     g2223(.I(new_n1802_), .ZN(new_n2866_));
  NAND4_X1   g2224(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1795_), .A4(new_n2866_), .ZN(new_n2867_));
  NAND2_X1   g2225(.A1(new_n2865_), .A2(new_n2867_), .ZN(\result[2] ));
  NAND4_X1   g2226(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1761_), .A4(new_n1765_), .ZN(new_n2869_));
  INV_X1     g2227(.I(new_n1761_), .ZN(new_n2870_));
  INV_X1     g2228(.I(new_n1765_), .ZN(new_n2871_));
  NAND4_X1   g2229(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2870_), .A4(new_n2871_), .ZN(new_n2872_));
  NAND2_X1   g2230(.A1(new_n2869_), .A2(new_n2872_), .ZN(\result[3] ));
  INV_X1     g2231(.I(new_n1738_), .ZN(new_n2874_));
  NAND4_X1   g2232(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1735_), .A4(new_n2874_), .ZN(new_n2875_));
  INV_X1     g2233(.I(new_n1735_), .ZN(new_n2876_));
  NAND4_X1   g2234(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2876_), .A4(new_n1738_), .ZN(new_n2877_));
  NAND2_X1   g2235(.A1(new_n2875_), .A2(new_n2877_), .ZN(\result[4] ));
  INV_X1     g2236(.I(new_n1728_), .ZN(new_n2879_));
  NAND4_X1   g2237(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2879_), .A4(new_n1732_), .ZN(new_n2880_));
  NAND4_X1   g2238(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1728_), .A4(new_n1731_), .ZN(new_n2881_));
  NAND2_X1   g2239(.A1(new_n2880_), .A2(new_n2881_), .ZN(\result[5] ));
  NAND4_X1   g2240(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1811_), .A4(new_n1813_), .ZN(new_n2883_));
  INV_X1     g2241(.I(new_n1811_), .ZN(new_n2884_));
  INV_X1     g2242(.I(new_n1813_), .ZN(new_n2885_));
  NAND4_X1   g2243(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2884_), .A4(new_n2885_), .ZN(new_n2886_));
  NAND2_X1   g2244(.A1(new_n2883_), .A2(new_n2886_), .ZN(\result[6] ));
  NAND4_X1   g2245(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1720_), .A4(new_n1814_), .ZN(new_n2888_));
  NAND4_X1   g2246(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1719_), .A4(new_n1723_), .ZN(new_n2889_));
  NAND2_X1   g2247(.A1(new_n2888_), .A2(new_n2889_), .ZN(\result[7] ));
  NAND4_X1   g2248(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1717_), .A4(new_n1821_), .ZN(new_n2891_));
  INV_X1     g2249(.I(new_n1717_), .ZN(new_n2892_));
  NAND4_X1   g2250(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2892_), .A4(new_n1822_), .ZN(new_n2893_));
  NAND2_X1   g2251(.A1(new_n2891_), .A2(new_n2893_), .ZN(\result[8] ));
  INV_X1     g2252(.I(new_n1827_), .ZN(new_n2895_));
  INV_X1     g2253(.I(new_n1830_), .ZN(new_n2896_));
  NAND4_X1   g2254(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2895_), .A4(new_n2896_), .ZN(new_n2897_));
  NAND4_X1   g2255(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1827_), .A4(new_n1830_), .ZN(new_n2898_));
  NAND2_X1   g2256(.A1(new_n2897_), .A2(new_n2898_), .ZN(\result[9] ));
  INV_X1     g2257(.I(new_n1832_), .ZN(new_n2900_));
  NAND4_X1   g2258(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2900_), .A4(new_n1834_), .ZN(new_n2901_));
  INV_X1     g2259(.I(new_n1834_), .ZN(new_n2902_));
  NAND4_X1   g2260(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1832_), .A4(new_n2902_), .ZN(new_n2903_));
  NAND2_X1   g2261(.A1(new_n2901_), .A2(new_n2903_), .ZN(\result[10] ));
  NAND4_X1   g2262(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1710_), .A4(new_n1837_), .ZN(new_n2905_));
  NAND4_X1   g2263(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1711_), .A4(new_n1714_), .ZN(new_n2906_));
  NAND2_X1   g2264(.A1(new_n2905_), .A2(new_n2906_), .ZN(\result[11] ));
  INV_X1     g2265(.I(new_n1844_), .ZN(new_n2908_));
  NAND4_X1   g2266(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2908_), .A4(new_n1848_), .ZN(new_n2909_));
  NAND4_X1   g2267(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1844_), .A4(new_n1847_), .ZN(new_n2910_));
  NAND2_X1   g2268(.A1(new_n2909_), .A2(new_n2910_), .ZN(\result[12] ));
  NAND4_X1   g2269(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1855_), .A4(new_n1853_), .ZN(new_n2912_));
  NAND4_X1   g2270(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1850_), .A4(new_n1852_), .ZN(new_n2913_));
  NAND2_X1   g2271(.A1(new_n2912_), .A2(new_n2913_), .ZN(\result[13] ));
  NAND4_X1   g2272(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1703_), .A4(new_n1707_), .ZN(new_n2915_));
  NAND4_X1   g2273(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1702_), .A4(new_n1706_), .ZN(new_n2916_));
  NAND2_X1   g2274(.A1(new_n2915_), .A2(new_n2916_), .ZN(\result[14] ));
  NAND4_X1   g2275(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1697_), .A4(new_n1860_), .ZN(new_n2918_));
  NAND4_X1   g2276(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1696_), .A4(new_n1699_), .ZN(new_n2919_));
  NAND2_X1   g2277(.A1(new_n2918_), .A2(new_n2919_), .ZN(\result[15] ));
  NAND4_X1   g2278(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1863_), .A4(new_n1693_), .ZN(new_n2921_));
  NAND4_X1   g2279(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1690_), .A4(new_n1692_), .ZN(new_n2922_));
  NAND2_X1   g2280(.A1(new_n2921_), .A2(new_n2922_), .ZN(\result[16] ));
  INV_X1     g2281(.I(new_n1872_), .ZN(new_n2924_));
  NAND4_X1   g2282(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1869_), .A4(new_n2924_), .ZN(new_n2925_));
  NAND4_X1   g2283(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1868_), .A4(new_n1872_), .ZN(new_n2926_));
  NAND2_X1   g2284(.A1(new_n2925_), .A2(new_n2926_), .ZN(\result[17] ));
  NAND4_X1   g2285(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1875_), .A4(new_n1879_), .ZN(new_n2928_));
  NAND4_X1   g2286(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1874_), .A4(new_n1877_), .ZN(new_n2929_));
  NAND2_X1   g2287(.A1(new_n2928_), .A2(new_n2929_), .ZN(\result[18] ));
  NAND4_X1   g2288(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1880_), .A4(new_n1881_), .ZN(new_n2931_));
  NAND4_X1   g2289(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1684_), .A4(new_n1687_), .ZN(new_n2932_));
  NAND2_X1   g2290(.A1(new_n2931_), .A2(new_n2932_), .ZN(\result[19] ));
  INV_X1     g2291(.I(new_n1888_), .ZN(new_n2934_));
  NAND4_X1   g2292(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2934_), .A4(new_n1892_), .ZN(new_n2935_));
  NAND4_X1   g2293(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1888_), .A4(new_n1891_), .ZN(new_n2936_));
  NAND2_X1   g2294(.A1(new_n2935_), .A2(new_n2936_), .ZN(\result[20] ));
  NAND4_X1   g2295(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1899_), .A4(new_n1897_), .ZN(new_n2938_));
  NAND4_X1   g2296(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1894_), .A4(new_n1896_), .ZN(new_n2939_));
  NAND2_X1   g2297(.A1(new_n2938_), .A2(new_n2939_), .ZN(\result[21] ));
  NAND4_X1   g2298(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1677_), .A4(new_n1681_), .ZN(new_n2941_));
  NAND4_X1   g2299(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1676_), .A4(new_n1680_), .ZN(new_n2942_));
  NAND2_X1   g2300(.A1(new_n2941_), .A2(new_n2942_), .ZN(\result[22] ));
  NAND4_X1   g2301(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1671_), .A4(new_n1904_), .ZN(new_n2944_));
  NAND4_X1   g2302(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1670_), .A4(new_n1673_), .ZN(new_n2945_));
  NAND2_X1   g2303(.A1(new_n2944_), .A2(new_n2945_), .ZN(\result[23] ));
  NAND4_X1   g2304(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1907_), .A4(new_n1667_), .ZN(new_n2947_));
  NAND4_X1   g2305(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1664_), .A4(new_n1666_), .ZN(new_n2948_));
  NAND2_X1   g2306(.A1(new_n2947_), .A2(new_n2948_), .ZN(\result[24] ));
  INV_X1     g2307(.I(new_n1916_), .ZN(new_n2950_));
  NAND4_X1   g2308(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1913_), .A4(new_n2950_), .ZN(new_n2951_));
  NAND4_X1   g2309(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1912_), .A4(new_n1916_), .ZN(new_n2952_));
  NAND2_X1   g2310(.A1(new_n2951_), .A2(new_n2952_), .ZN(\result[25] ));
  NAND4_X1   g2311(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1919_), .A4(new_n1923_), .ZN(new_n2954_));
  NAND4_X1   g2312(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1918_), .A4(new_n1921_), .ZN(new_n2955_));
  NAND2_X1   g2313(.A1(new_n2954_), .A2(new_n2955_), .ZN(\result[26] ));
  NAND4_X1   g2314(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1924_), .A4(new_n1925_), .ZN(new_n2957_));
  NAND4_X1   g2315(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1658_), .A4(new_n1661_), .ZN(new_n2958_));
  NAND2_X1   g2316(.A1(new_n2957_), .A2(new_n2958_), .ZN(\result[27] ));
  INV_X1     g2317(.I(new_n1932_), .ZN(new_n2960_));
  NAND4_X1   g2318(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2960_), .A4(new_n1936_), .ZN(new_n2961_));
  NAND4_X1   g2319(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1932_), .A4(new_n1935_), .ZN(new_n2962_));
  NAND2_X1   g2320(.A1(new_n2961_), .A2(new_n2962_), .ZN(\result[28] ));
  NAND4_X1   g2321(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1943_), .A4(new_n1941_), .ZN(new_n2964_));
  NAND4_X1   g2322(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1938_), .A4(new_n1940_), .ZN(new_n2965_));
  NAND2_X1   g2323(.A1(new_n2964_), .A2(new_n2965_), .ZN(\result[29] ));
  NAND4_X1   g2324(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1618_), .A4(new_n1655_), .ZN(new_n2967_));
  NAND4_X1   g2325(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1617_), .A4(new_n1654_), .ZN(new_n2968_));
  NAND2_X1   g2326(.A1(new_n2967_), .A2(new_n2968_), .ZN(\result[30] ));
  NAND4_X1   g2327(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2628_), .A4(new_n2791_), .ZN(new_n2970_));
  NAND4_X1   g2328(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2627_), .A4(new_n2790_), .ZN(new_n2971_));
  NAND2_X1   g2329(.A1(new_n2970_), .A2(new_n2971_), .ZN(\result[31] ));
  NAND4_X1   g2330(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2629_), .A4(new_n2630_), .ZN(new_n2973_));
  NAND4_X1   g2331(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2481_), .A4(new_n2485_), .ZN(new_n2974_));
  NAND2_X1   g2332(.A1(new_n2973_), .A2(new_n2974_), .ZN(\result[32] ));
  INV_X1     g2333(.I(new_n2479_), .ZN(new_n2976_));
  INV_X1     g2334(.I(new_n2483_), .ZN(new_n2977_));
  NAND4_X1   g2335(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2976_), .A4(new_n2977_), .ZN(new_n2978_));
  NAND4_X1   g2336(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2479_), .A4(new_n2483_), .ZN(new_n2979_));
  NAND2_X1   g2337(.A1(new_n2978_), .A2(new_n2979_), .ZN(\result[33] ));
  INV_X1     g2338(.I(new_n2494_), .ZN(new_n2981_));
  NAND4_X1   g2339(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2981_), .A4(new_n2497_), .ZN(new_n2982_));
  NAND4_X1   g2340(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2494_), .A4(new_n2496_), .ZN(new_n2983_));
  NAND2_X1   g2341(.A1(new_n2982_), .A2(new_n2983_), .ZN(\result[34] ));
  INV_X1     g2342(.I(new_n2488_), .ZN(new_n2985_));
  INV_X1     g2343(.I(new_n2490_), .ZN(new_n2986_));
  NAND4_X1   g2344(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2985_), .A4(new_n2986_), .ZN(new_n2987_));
  NAND4_X1   g2345(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2488_), .A4(new_n2490_), .ZN(new_n2988_));
  NAND2_X1   g2346(.A1(new_n2987_), .A2(new_n2988_), .ZN(\result[35] ));
  INV_X1     g2347(.I(new_n2522_), .ZN(new_n2990_));
  NAND4_X1   g2348(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2990_), .A4(new_n2544_), .ZN(new_n2991_));
  NAND4_X1   g2349(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2522_), .A4(new_n2525_), .ZN(new_n2992_));
  NAND2_X1   g2350(.A1(new_n2991_), .A2(new_n2992_), .ZN(\result[36] ));
  NAND4_X1   g2351(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2502_), .A4(new_n2543_), .ZN(new_n2994_));
  NAND4_X1   g2352(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2501_), .A4(new_n2505_), .ZN(new_n2995_));
  NAND2_X1   g2353(.A1(new_n2994_), .A2(new_n2995_), .ZN(\result[37] ));
  NAND4_X1   g2354(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2537_), .A4(new_n2534_), .ZN(new_n2997_));
  NAND4_X1   g2355(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2509_), .A4(new_n2515_), .ZN(new_n2998_));
  NAND2_X1   g2356(.A1(new_n2997_), .A2(new_n2998_), .ZN(\result[38] ));
  NAND4_X1   g2357(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2533_), .A4(new_n2538_), .ZN(new_n3000_));
  NAND4_X1   g2358(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2512_), .A4(new_n2518_), .ZN(new_n3001_));
  NAND2_X1   g2359(.A1(new_n3000_), .A2(new_n3001_), .ZN(\result[39] ));
  INV_X1     g2360(.I(new_n2612_), .ZN(new_n3003_));
  NAND4_X1   g2361(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3003_), .A4(new_n2615_), .ZN(new_n3004_));
  NAND4_X1   g2362(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2612_), .A4(new_n2614_), .ZN(new_n3005_));
  NAND2_X1   g2363(.A1(new_n3004_), .A2(new_n3005_), .ZN(\result[40] ));
  NAND4_X1   g2364(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2605_), .A4(new_n2608_), .ZN(new_n3007_));
  NAND4_X1   g2365(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2604_), .A4(new_n2607_), .ZN(new_n3008_));
  NAND2_X1   g2366(.A1(new_n3007_), .A2(new_n3008_), .ZN(\result[41] ));
  NAND4_X1   g2367(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2592_), .A4(new_n2596_), .ZN(new_n3010_));
  NAND4_X1   g2368(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2591_), .A4(new_n2595_), .ZN(new_n3011_));
  NAND2_X1   g2369(.A1(new_n3010_), .A2(new_n3011_), .ZN(\result[42] ));
  NAND4_X1   g2370(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2588_), .A4(new_n2600_), .ZN(new_n3013_));
  NAND4_X1   g2371(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2587_), .A4(new_n2599_), .ZN(new_n3014_));
  NAND2_X1   g2372(.A1(new_n3013_), .A2(new_n3014_), .ZN(\result[43] ));
  NAND4_X1   g2373(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2575_), .A4(new_n2619_), .ZN(new_n3016_));
  NAND4_X1   g2374(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2574_), .A4(new_n2578_), .ZN(new_n3017_));
  NAND2_X1   g2375(.A1(new_n3016_), .A2(new_n3017_), .ZN(\result[44] ));
  INV_X1     g2376(.I(new_n2550_), .ZN(new_n3019_));
  NAND4_X1   g2377(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3019_), .A4(new_n2620_), .ZN(new_n3020_));
  NAND4_X1   g2378(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2550_), .A4(new_n2553_), .ZN(new_n3021_));
  NAND2_X1   g2379(.A1(new_n3020_), .A2(new_n3021_), .ZN(\result[45] ));
  NAND4_X1   g2380(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2557_), .A4(new_n2565_), .ZN(new_n3023_));
  NAND4_X1   g2381(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2556_), .A4(new_n2564_), .ZN(new_n3024_));
  NAND2_X1   g2382(.A1(new_n3023_), .A2(new_n3024_), .ZN(\result[46] ));
  NAND4_X1   g2383(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2561_), .A4(new_n2569_), .ZN(new_n3026_));
  NAND4_X1   g2384(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2560_), .A4(new_n2568_), .ZN(new_n3027_));
  NAND2_X1   g2385(.A1(new_n3026_), .A2(new_n3027_), .ZN(\result[47] ));
  NAND4_X1   g2386(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2047_), .A4(new_n2009_), .ZN(new_n3029_));
  NAND4_X1   g2387(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1990_), .A4(new_n1992_), .ZN(new_n3030_));
  NAND2_X1   g2388(.A1(new_n3029_), .A2(new_n3030_), .ZN(\result[48] ));
  INV_X1     g2389(.I(new_n1955_), .ZN(new_n3032_));
  NAND4_X1   g2390(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2010_), .A4(new_n3032_), .ZN(new_n3033_));
  NAND4_X1   g2391(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1951_), .A4(new_n1955_), .ZN(new_n3034_));
  NAND2_X1   g2392(.A1(new_n3033_), .A2(new_n3034_), .ZN(\result[49] ));
  INV_X1     g2393(.I(new_n1959_), .ZN(new_n3036_));
  NAND4_X1   g2394(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3036_), .A4(new_n1962_), .ZN(new_n3037_));
  NAND4_X1   g2395(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1959_), .A4(new_n1961_), .ZN(new_n3038_));
  NAND2_X1   g2396(.A1(new_n3037_), .A2(new_n3038_), .ZN(\result[50] ));
  INV_X1     g2397(.I(new_n1949_), .ZN(new_n3040_));
  INV_X1     g2398(.I(new_n1953_), .ZN(new_n3041_));
  NAND4_X1   g2399(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3040_), .A4(new_n3041_), .ZN(new_n3042_));
  NAND4_X1   g2400(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1949_), .A4(new_n1953_), .ZN(new_n3043_));
  NAND2_X1   g2401(.A1(new_n3042_), .A2(new_n3043_), .ZN(\result[51] ));
  NAND4_X1   g2402(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1966_), .A4(new_n2000_), .ZN(new_n3045_));
  NAND4_X1   g2403(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1965_), .A4(new_n1968_), .ZN(new_n3046_));
  NAND2_X1   g2404(.A1(new_n3045_), .A2(new_n3046_), .ZN(\result[52] ));
  INV_X1     g2405(.I(new_n1983_), .ZN(new_n3048_));
  NAND4_X1   g2406(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3048_), .A4(new_n1995_), .ZN(new_n3049_));
  NAND4_X1   g2407(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1983_), .A4(new_n1985_), .ZN(new_n3050_));
  NAND2_X1   g2408(.A1(new_n3049_), .A2(new_n3050_), .ZN(\result[53] ));
  INV_X1     g2409(.I(new_n1972_), .ZN(new_n3052_));
  NAND4_X1   g2410(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3052_), .A4(new_n1996_), .ZN(new_n3053_));
  NAND4_X1   g2411(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1972_), .A4(new_n1977_), .ZN(new_n3054_));
  NAND2_X1   g2412(.A1(new_n3053_), .A2(new_n3054_), .ZN(\result[54] ));
  INV_X1     g2413(.I(new_n1980_), .ZN(new_n3056_));
  NAND4_X1   g2414(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1994_), .A4(new_n3056_), .ZN(new_n3057_));
  NAND4_X1   g2415(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1975_), .A4(new_n1980_), .ZN(new_n3058_));
  NAND2_X1   g2416(.A1(new_n3057_), .A2(new_n3058_), .ZN(\result[55] ));
  INV_X1     g2417(.I(new_n2060_), .ZN(new_n3060_));
  NAND4_X1   g2418(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3060_), .A4(new_n2810_), .ZN(new_n3061_));
  NAND4_X1   g2419(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2060_), .A4(new_n2066_), .ZN(new_n3062_));
  NAND2_X1   g2420(.A1(new_n3061_), .A2(new_n3062_), .ZN(\result[56] ));
  INV_X1     g2421(.I(new_n2063_), .ZN(new_n3064_));
  INV_X1     g2422(.I(new_n2069_), .ZN(new_n3065_));
  NAND4_X1   g2423(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3064_), .A4(new_n3065_), .ZN(new_n3066_));
  NAND4_X1   g2424(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2063_), .A4(new_n2069_), .ZN(new_n3067_));
  NAND2_X1   g2425(.A1(new_n3066_), .A2(new_n3067_), .ZN(\result[57] ));
  INV_X1     g2426(.I(new_n2054_), .ZN(new_n3069_));
  NAND4_X1   g2427(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2806_), .A4(new_n3069_), .ZN(new_n3070_));
  NAND4_X1   g2428(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2049_), .A4(new_n2054_), .ZN(new_n3071_));
  NAND2_X1   g2429(.A1(new_n3070_), .A2(new_n3071_), .ZN(\result[58] ));
  NAND4_X1   g2430(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2803_), .A4(new_n2805_), .ZN(new_n3073_));
  NAND4_X1   g2431(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2051_), .A4(new_n2056_), .ZN(new_n3074_));
  NAND2_X1   g2432(.A1(new_n3073_), .A2(new_n3074_), .ZN(\result[59] ));
  NAND4_X1   g2433(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2041_), .A4(new_n2045_), .ZN(new_n3076_));
  NAND4_X1   g2434(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2040_), .A4(new_n2044_), .ZN(new_n3077_));
  NAND2_X1   g2435(.A1(new_n3076_), .A2(new_n3077_), .ZN(\result[60] ));
  NAND4_X1   g2436(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2016_), .A4(new_n2793_), .ZN(new_n3079_));
  NAND4_X1   g2437(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2015_), .A4(new_n2019_), .ZN(new_n3080_));
  NAND2_X1   g2438(.A1(new_n3079_), .A2(new_n3080_), .ZN(\result[61] ));
  NAND4_X1   g2439(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2023_), .A4(new_n2031_), .ZN(new_n3082_));
  NAND4_X1   g2440(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2022_), .A4(new_n2030_), .ZN(new_n3083_));
  NAND2_X1   g2441(.A1(new_n3082_), .A2(new_n3083_), .ZN(\result[62] ));
  NAND4_X1   g2442(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2027_), .A4(new_n2035_), .ZN(new_n3085_));
  NAND4_X1   g2443(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2026_), .A4(new_n2034_), .ZN(new_n3086_));
  NAND2_X1   g2444(.A1(new_n3085_), .A2(new_n3086_), .ZN(\result[63] ));
  INV_X1     g2445(.I(new_n2838_), .ZN(new_n3088_));
  NAND4_X1   g2446(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3088_), .A4(new_n2842_), .ZN(new_n3089_));
  NAND4_X1   g2447(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2838_), .A4(new_n2841_), .ZN(new_n3090_));
  NAND2_X1   g2448(.A1(new_n3089_), .A2(new_n3090_), .ZN(\result[64] ));
  NAND4_X1   g2449(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2830_), .A4(new_n2833_), .ZN(new_n3092_));
  NAND4_X1   g2450(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2829_), .A4(new_n2832_), .ZN(new_n3093_));
  NAND2_X1   g2451(.A1(new_n3092_), .A2(new_n3093_), .ZN(\result[65] ));
  NAND4_X1   g2452(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2819_), .A4(new_n2823_), .ZN(new_n3095_));
  NAND4_X1   g2453(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2818_), .A4(new_n2822_), .ZN(new_n3096_));
  NAND2_X1   g2454(.A1(new_n3095_), .A2(new_n3096_), .ZN(\result[66] ));
  NAND4_X1   g2455(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2816_), .A4(new_n2826_), .ZN(new_n3098_));
  NAND4_X1   g2456(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2815_), .A4(new_n2825_), .ZN(new_n3099_));
  NAND2_X1   g2457(.A1(new_n3098_), .A2(new_n3099_), .ZN(\result[67] ));
  NAND4_X1   g2458(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2695_), .A4(new_n2699_), .ZN(new_n3101_));
  NAND4_X1   g2459(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2694_), .A4(new_n2698_), .ZN(new_n3102_));
  NAND2_X1   g2460(.A1(new_n3101_), .A2(new_n3102_), .ZN(\result[68] ));
  INV_X1     g2461(.I(new_n2670_), .ZN(new_n3104_));
  NAND4_X1   g2462(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3104_), .A4(new_n2673_), .ZN(new_n3105_));
  NAND4_X1   g2463(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2670_), .A4(new_n2672_), .ZN(new_n3106_));
  NAND2_X1   g2464(.A1(new_n3105_), .A2(new_n3106_), .ZN(\result[69] ));
  NAND4_X1   g2465(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2678_), .A4(new_n2686_), .ZN(new_n3108_));
  NAND4_X1   g2466(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2677_), .A4(new_n2685_), .ZN(new_n3109_));
  NAND2_X1   g2467(.A1(new_n3108_), .A2(new_n3109_), .ZN(\result[70] ));
  NAND4_X1   g2468(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2682_), .A4(new_n2690_), .ZN(new_n3111_));
  NAND4_X1   g2469(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2681_), .A4(new_n2689_), .ZN(new_n3112_));
  NAND2_X1   g2470(.A1(new_n3111_), .A2(new_n3112_), .ZN(\result[71] ));
  INV_X1     g2471(.I(new_n2707_), .ZN(new_n3114_));
  NAND4_X1   g2472(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3114_), .A4(new_n2710_), .ZN(new_n3115_));
  NAND4_X1   g2473(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2707_), .A4(new_n2709_), .ZN(new_n3116_));
  NAND2_X1   g2474(.A1(new_n3115_), .A2(new_n3116_), .ZN(\result[72] ));
  NAND4_X1   g2475(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2734_), .A4(new_n2738_), .ZN(new_n3118_));
  NAND4_X1   g2476(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2733_), .A4(new_n2737_), .ZN(new_n3119_));
  NAND2_X1   g2477(.A1(new_n3118_), .A2(new_n3119_), .ZN(\result[73] ));
  NAND4_X1   g2478(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2714_), .A4(new_n2721_), .ZN(new_n3121_));
  NAND4_X1   g2479(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2713_), .A4(new_n2720_), .ZN(new_n3122_));
  NAND2_X1   g2480(.A1(new_n3121_), .A2(new_n3122_), .ZN(\result[74] ));
  NAND4_X1   g2481(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2717_), .A4(new_n2725_), .ZN(new_n3124_));
  NAND4_X1   g2482(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2716_), .A4(new_n2724_), .ZN(new_n3125_));
  NAND2_X1   g2483(.A1(new_n3124_), .A2(new_n3125_), .ZN(\result[75] ));
  NAND4_X1   g2484(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2747_), .A4(new_n2778_), .ZN(new_n3127_));
  NAND4_X1   g2485(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2746_), .A4(new_n2753_), .ZN(new_n3128_));
  NAND2_X1   g2486(.A1(new_n3127_), .A2(new_n3128_), .ZN(\result[76] ));
  NAND4_X1   g2487(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2743_), .A4(new_n2779_), .ZN(new_n3130_));
  NAND4_X1   g2488(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2742_), .A4(new_n2750_), .ZN(new_n3131_));
  NAND2_X1   g2489(.A1(new_n3130_), .A2(new_n3131_), .ZN(\result[77] ));
  NAND4_X1   g2490(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2758_), .A4(new_n2766_), .ZN(new_n3133_));
  NAND4_X1   g2491(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2757_), .A4(new_n2765_), .ZN(new_n3134_));
  NAND2_X1   g2492(.A1(new_n3133_), .A2(new_n3134_), .ZN(\result[78] ));
  NAND4_X1   g2493(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2762_), .A4(new_n2770_), .ZN(new_n3136_));
  NAND4_X1   g2494(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2761_), .A4(new_n2769_), .ZN(new_n3137_));
  NAND2_X1   g2495(.A1(new_n3136_), .A2(new_n3137_), .ZN(\result[79] ));
  INV_X1     g2496(.I(new_n2251_), .ZN(new_n3139_));
  NAND4_X1   g2497(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3139_), .A4(new_n2254_), .ZN(new_n3140_));
  NAND4_X1   g2498(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2251_), .A4(new_n2253_), .ZN(new_n3141_));
  NAND2_X1   g2499(.A1(new_n3140_), .A2(new_n3141_), .ZN(\result[80] ));
  NAND4_X1   g2500(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2269_), .A4(new_n2272_), .ZN(new_n3143_));
  NAND4_X1   g2501(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2268_), .A4(new_n2271_), .ZN(new_n3144_));
  NAND2_X1   g2502(.A1(new_n3143_), .A2(new_n3144_), .ZN(\result[81] ));
  INV_X1     g2503(.I(new_n2256_), .ZN(new_n3146_));
  NAND4_X1   g2504(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3146_), .A4(new_n2275_), .ZN(new_n3147_));
  NAND4_X1   g2505(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2256_), .A4(new_n2262_), .ZN(new_n3148_));
  NAND2_X1   g2506(.A1(new_n3147_), .A2(new_n3148_), .ZN(\result[82] ));
  INV_X1     g2507(.I(new_n2264_), .ZN(new_n3150_));
  NAND4_X1   g2508(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2274_), .A4(new_n3150_), .ZN(new_n3151_));
  NAND4_X1   g2509(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2259_), .A4(new_n2264_), .ZN(new_n3152_));
  NAND2_X1   g2510(.A1(new_n3151_), .A2(new_n3152_), .ZN(\result[83] ));
  INV_X1     g2511(.I(new_n2301_), .ZN(new_n3154_));
  NAND4_X1   g2512(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3154_), .A4(new_n2314_), .ZN(new_n3155_));
  NAND4_X1   g2513(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2301_), .A4(new_n2304_), .ZN(new_n3156_));
  NAND2_X1   g2514(.A1(new_n3155_), .A2(new_n3156_), .ZN(\result[84] ));
  NAND4_X1   g2515(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2284_), .A4(new_n2313_), .ZN(new_n3158_));
  NAND4_X1   g2516(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2283_), .A4(new_n2286_), .ZN(new_n3159_));
  NAND2_X1   g2517(.A1(new_n3158_), .A2(new_n3159_), .ZN(\result[85] ));
  INV_X1     g2518(.I(new_n2290_), .ZN(new_n3161_));
  NAND4_X1   g2519(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3161_), .A4(new_n2310_), .ZN(new_n3162_));
  NAND4_X1   g2520(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2290_), .A4(new_n2295_), .ZN(new_n3163_));
  NAND2_X1   g2521(.A1(new_n3162_), .A2(new_n3163_), .ZN(\result[86] ));
  INV_X1     g2522(.I(new_n2297_), .ZN(new_n3165_));
  NAND4_X1   g2523(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2309_), .A4(new_n3165_), .ZN(new_n3166_));
  NAND4_X1   g2524(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2292_), .A4(new_n2297_), .ZN(new_n3167_));
  NAND2_X1   g2525(.A1(new_n3166_), .A2(new_n3167_), .ZN(\result[87] ));
  NAND4_X1   g2526(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2348_), .A4(new_n2345_), .ZN(new_n3169_));
  NAND4_X1   g2527(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2342_), .A4(new_n2344_), .ZN(new_n3170_));
  NAND2_X1   g2528(.A1(new_n3169_), .A2(new_n3170_), .ZN(\result[88] ));
  INV_X1     g2529(.I(new_n2331_), .ZN(new_n3172_));
  NAND4_X1   g2530(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3172_), .A4(new_n2335_), .ZN(new_n3173_));
  NAND4_X1   g2531(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2331_), .A4(new_n2334_), .ZN(new_n3174_));
  NAND2_X1   g2532(.A1(new_n3173_), .A2(new_n3174_), .ZN(\result[89] ));
  INV_X1     g2533(.I(new_n2323_), .ZN(new_n3176_));
  NAND4_X1   g2534(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3176_), .A4(new_n2336_), .ZN(new_n3177_));
  NAND4_X1   g2535(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2323_), .A4(new_n2326_), .ZN(new_n3178_));
  NAND2_X1   g2536(.A1(new_n3177_), .A2(new_n3178_), .ZN(\result[90] ));
  INV_X1     g2537(.I(new_n2328_), .ZN(new_n3180_));
  NAND4_X1   g2538(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2321_), .A4(new_n3180_), .ZN(new_n3181_));
  NAND4_X1   g2539(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2320_), .A4(new_n2328_), .ZN(new_n3182_));
  NAND2_X1   g2540(.A1(new_n3181_), .A2(new_n3182_), .ZN(\result[91] ));
  NAND4_X1   g2541(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2379_), .A4(new_n2383_), .ZN(new_n3184_));
  NAND4_X1   g2542(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2378_), .A4(new_n2382_), .ZN(new_n3185_));
  NAND2_X1   g2543(.A1(new_n3184_), .A2(new_n3185_), .ZN(\result[92] ));
  NAND4_X1   g2544(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2355_), .A4(new_n2385_), .ZN(new_n3187_));
  NAND4_X1   g2545(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2354_), .A4(new_n2357_), .ZN(new_n3188_));
  NAND2_X1   g2546(.A1(new_n3187_), .A2(new_n3188_), .ZN(\result[93] ));
  NAND4_X1   g2547(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2361_), .A4(new_n2369_), .ZN(new_n3190_));
  NAND4_X1   g2548(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2360_), .A4(new_n2368_), .ZN(new_n3191_));
  NAND2_X1   g2549(.A1(new_n3190_), .A2(new_n3191_), .ZN(\result[94] ));
  NAND4_X1   g2550(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2365_), .A4(new_n2373_), .ZN(new_n3193_));
  NAND4_X1   g2551(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2364_), .A4(new_n2372_), .ZN(new_n3194_));
  NAND2_X1   g2552(.A1(new_n3193_), .A2(new_n3194_), .ZN(\result[95] ));
  NAND4_X1   g2553(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2392_), .A4(new_n2471_), .ZN(new_n3196_));
  NAND4_X1   g2554(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2391_), .A4(new_n2394_), .ZN(new_n3197_));
  NAND2_X1   g2555(.A1(new_n3196_), .A2(new_n3197_), .ZN(\result[96] ));
  NAND4_X1   g2556(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2418_), .A4(new_n2422_), .ZN(new_n3199_));
  NAND4_X1   g2557(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2417_), .A4(new_n2421_), .ZN(new_n3200_));
  NAND2_X1   g2558(.A1(new_n3199_), .A2(new_n3200_), .ZN(\result[97] ));
  NAND4_X1   g2559(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2398_), .A4(new_n2405_), .ZN(new_n3202_));
  NAND4_X1   g2560(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2397_), .A4(new_n2404_), .ZN(new_n3203_));
  NAND2_X1   g2561(.A1(new_n3202_), .A2(new_n3203_), .ZN(\result[98] ));
  NAND4_X1   g2562(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2401_), .A4(new_n2409_), .ZN(new_n3205_));
  NAND4_X1   g2563(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2400_), .A4(new_n2408_), .ZN(new_n3206_));
  NAND2_X1   g2564(.A1(new_n3205_), .A2(new_n3206_), .ZN(\result[99] ));
  NAND4_X1   g2565(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2440_), .A4(new_n2437_), .ZN(new_n3208_));
  NAND4_X1   g2566(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2429_), .A4(new_n2436_), .ZN(new_n3209_));
  NAND2_X1   g2567(.A1(new_n3208_), .A2(new_n3209_), .ZN(\result[100] ));
  NAND4_X1   g2568(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2439_), .A4(new_n2433_), .ZN(new_n3211_));
  NAND4_X1   g2569(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2426_), .A4(new_n2432_), .ZN(new_n3212_));
  NAND2_X1   g2570(.A1(new_n3211_), .A2(new_n3212_), .ZN(\result[101] ));
  NAND4_X1   g2571(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2444_), .A4(new_n2452_), .ZN(new_n3214_));
  NAND4_X1   g2572(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2443_), .A4(new_n2451_), .ZN(new_n3215_));
  NAND2_X1   g2573(.A1(new_n3214_), .A2(new_n3215_), .ZN(\result[102] ));
  NAND4_X1   g2574(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2448_), .A4(new_n2456_), .ZN(new_n3217_));
  NAND4_X1   g2575(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2447_), .A4(new_n2455_), .ZN(new_n3218_));
  NAND2_X1   g2576(.A1(new_n3217_), .A2(new_n3218_), .ZN(\result[103] ));
  INV_X1     g2577(.I(new_n2147_), .ZN(new_n3220_));
  NAND4_X1   g2578(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3220_), .A4(new_n2150_), .ZN(new_n3221_));
  NAND4_X1   g2579(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2147_), .A4(new_n2149_), .ZN(new_n3222_));
  NAND2_X1   g2580(.A1(new_n3221_), .A2(new_n3222_), .ZN(\result[104] ));
  NAND4_X1   g2581(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2165_), .A4(new_n2168_), .ZN(new_n3224_));
  NAND4_X1   g2582(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2164_), .A4(new_n2167_), .ZN(new_n3225_));
  NAND2_X1   g2583(.A1(new_n3224_), .A2(new_n3225_), .ZN(\result[105] ));
  INV_X1     g2584(.I(new_n2152_), .ZN(new_n3227_));
  NAND4_X1   g2585(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3227_), .A4(new_n2171_), .ZN(new_n3228_));
  NAND4_X1   g2586(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2152_), .A4(new_n2158_), .ZN(new_n3229_));
  NAND2_X1   g2587(.A1(new_n3228_), .A2(new_n3229_), .ZN(\result[106] ));
  INV_X1     g2588(.I(new_n2160_), .ZN(new_n3231_));
  NAND4_X1   g2589(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2170_), .A4(new_n3231_), .ZN(new_n3232_));
  NAND4_X1   g2590(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2155_), .A4(new_n2160_), .ZN(new_n3233_));
  NAND2_X1   g2591(.A1(new_n3232_), .A2(new_n3233_), .ZN(\result[107] ));
  INV_X1     g2592(.I(new_n2197_), .ZN(new_n3235_));
  NAND4_X1   g2593(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3235_), .A4(new_n2210_), .ZN(new_n3236_));
  NAND4_X1   g2594(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2197_), .A4(new_n2200_), .ZN(new_n3237_));
  NAND2_X1   g2595(.A1(new_n3236_), .A2(new_n3237_), .ZN(\result[108] ));
  NAND4_X1   g2596(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2180_), .A4(new_n2209_), .ZN(new_n3239_));
  NAND4_X1   g2597(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2179_), .A4(new_n2182_), .ZN(new_n3240_));
  NAND2_X1   g2598(.A1(new_n3239_), .A2(new_n3240_), .ZN(\result[109] ));
  INV_X1     g2599(.I(new_n2186_), .ZN(new_n3242_));
  NAND4_X1   g2600(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3242_), .A4(new_n2206_), .ZN(new_n3243_));
  NAND4_X1   g2601(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2186_), .A4(new_n2191_), .ZN(new_n3244_));
  NAND2_X1   g2602(.A1(new_n3243_), .A2(new_n3244_), .ZN(\result[110] ));
  INV_X1     g2603(.I(new_n2193_), .ZN(new_n3246_));
  NAND4_X1   g2604(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2205_), .A4(new_n3246_), .ZN(new_n3247_));
  NAND4_X1   g2605(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2188_), .A4(new_n2193_), .ZN(new_n3248_));
  NAND2_X1   g2606(.A1(new_n3247_), .A2(new_n3248_), .ZN(\result[111] ));
  NAND4_X1   g2607(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2244_), .A4(new_n2241_), .ZN(new_n3250_));
  NAND4_X1   g2608(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2238_), .A4(new_n2240_), .ZN(new_n3251_));
  NAND2_X1   g2609(.A1(new_n3250_), .A2(new_n3251_), .ZN(\result[112] ));
  INV_X1     g2610(.I(new_n2227_), .ZN(new_n3253_));
  NAND4_X1   g2611(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3253_), .A4(new_n2231_), .ZN(new_n3254_));
  NAND4_X1   g2612(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2227_), .A4(new_n2230_), .ZN(new_n3255_));
  NAND2_X1   g2613(.A1(new_n3254_), .A2(new_n3255_), .ZN(\result[113] ));
  INV_X1     g2614(.I(new_n2219_), .ZN(new_n3257_));
  NAND4_X1   g2615(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n3257_), .A4(new_n2232_), .ZN(new_n3258_));
  NAND4_X1   g2616(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2219_), .A4(new_n2222_), .ZN(new_n3259_));
  NAND2_X1   g2617(.A1(new_n3258_), .A2(new_n3259_), .ZN(\result[114] ));
  INV_X1     g2618(.I(new_n2224_), .ZN(new_n3261_));
  NAND4_X1   g2619(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2217_), .A4(new_n3261_), .ZN(new_n3262_));
  NAND4_X1   g2620(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2216_), .A4(new_n2224_), .ZN(new_n3263_));
  NAND2_X1   g2621(.A1(new_n3262_), .A2(new_n3263_), .ZN(\result[115] ));
  NAND4_X1   g2622(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2100_), .A4(new_n2104_), .ZN(new_n3265_));
  NAND4_X1   g2623(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2099_), .A4(new_n2103_), .ZN(new_n3266_));
  NAND2_X1   g2624(.A1(new_n3265_), .A2(new_n3266_), .ZN(\result[116] ));
  NAND4_X1   g2625(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2076_), .A4(new_n2106_), .ZN(new_n3268_));
  NAND4_X1   g2626(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2075_), .A4(new_n2078_), .ZN(new_n3269_));
  NAND2_X1   g2627(.A1(new_n3268_), .A2(new_n3269_), .ZN(\result[117] ));
  NAND4_X1   g2628(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2082_), .A4(new_n2090_), .ZN(new_n3271_));
  NAND4_X1   g2629(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2081_), .A4(new_n2089_), .ZN(new_n3272_));
  NAND2_X1   g2630(.A1(new_n3271_), .A2(new_n3272_), .ZN(\result[118] ));
  NAND4_X1   g2631(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2086_), .A4(new_n2094_), .ZN(new_n3274_));
  NAND4_X1   g2632(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2085_), .A4(new_n2093_), .ZN(new_n3275_));
  NAND2_X1   g2633(.A1(new_n3274_), .A2(new_n3275_), .ZN(\result[119] ));
  NAND4_X1   g2634(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2113_), .A4(new_n2664_), .ZN(new_n3277_));
  NAND4_X1   g2635(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2112_), .A4(new_n2115_), .ZN(new_n3278_));
  NAND2_X1   g2636(.A1(new_n3277_), .A2(new_n3278_), .ZN(\result[120] ));
  NAND4_X1   g2637(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2139_), .A4(new_n2143_), .ZN(new_n3280_));
  NAND4_X1   g2638(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2138_), .A4(new_n2142_), .ZN(new_n3281_));
  NAND2_X1   g2639(.A1(new_n3280_), .A2(new_n3281_), .ZN(\result[121] ));
  NAND4_X1   g2640(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2119_), .A4(new_n2126_), .ZN(new_n3283_));
  NAND4_X1   g2641(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2118_), .A4(new_n2125_), .ZN(new_n3284_));
  NAND2_X1   g2642(.A1(new_n3283_), .A2(new_n3284_), .ZN(\result[122] ));
  NAND4_X1   g2643(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2122_), .A4(new_n2130_), .ZN(new_n3286_));
  NAND4_X1   g2644(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2121_), .A4(new_n2129_), .ZN(new_n3287_));
  NAND2_X1   g2645(.A1(new_n3286_), .A2(new_n3287_), .ZN(\result[123] ));
  NAND4_X1   g2646(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2654_), .A4(new_n2658_), .ZN(new_n3289_));
  NAND4_X1   g2647(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2653_), .A4(new_n2657_), .ZN(new_n3290_));
  NAND2_X1   g2648(.A1(new_n3289_), .A2(new_n3290_), .ZN(\result[124] ));
  NAND4_X1   g2649(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2649_), .A4(new_n2650_), .ZN(new_n3292_));
  NAND4_X1   g2650(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2635_), .A4(new_n2640_), .ZN(new_n3293_));
  NAND2_X1   g2651(.A1(new_n3292_), .A2(new_n3293_), .ZN(\result[125] ));
  INV_X1     g2652(.I(new_n2642_), .ZN(new_n3295_));
  NAND4_X1   g2653(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2645_), .A4(new_n3295_), .ZN(new_n3296_));
  NAND4_X1   g2654(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n2637_), .A4(new_n2642_), .ZN(new_n3297_));
  NAND2_X1   g2655(.A1(new_n3296_), .A2(new_n3297_), .ZN(\result[126] ));
  AOI21_X1   g2656(.A1(new_n2852_), .A2(new_n1611_), .B(new_n2644_), .ZN(\result[127] ));
  NAND4_X1   g2657(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1783_), .A4(new_n1652_), .ZN(new_n3300_));
  INV_X1     g2658(.I(new_n1652_), .ZN(new_n3301_));
  NAND4_X1   g2659(.A1(new_n2852_), .A2(new_n1612_), .A3(new_n1615_), .A4(new_n3301_), .ZN(new_n3302_));
  NAND2_X1   g2660(.A1(new_n3300_), .A2(new_n3302_), .ZN(\address[0] ));
  INV_X1     g2661(.I(new_n1612_), .ZN(new_n3304_));
  AND2_X2    g2662(.A1(new_n2852_), .A2(new_n3304_), .Z(\address[1] ));
endmodule


